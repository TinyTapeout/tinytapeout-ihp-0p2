module tt_um_vc32_cpu (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire _15022_;
 wire _15023_;
 wire _15024_;
 wire _15025_;
 wire _15026_;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire _15031_;
 wire _15032_;
 wire _15033_;
 wire _15034_;
 wire _15035_;
 wire _15036_;
 wire _15037_;
 wire _15038_;
 wire _15039_;
 wire _15040_;
 wire _15041_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire _15045_;
 wire _15046_;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire _15051_;
 wire _15052_;
 wire _15053_;
 wire _15054_;
 wire _15055_;
 wire _15056_;
 wire _15057_;
 wire _15058_;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire _15062_;
 wire _15063_;
 wire _15064_;
 wire _15065_;
 wire _15066_;
 wire _15067_;
 wire _15068_;
 wire _15069_;
 wire _15070_;
 wire _15071_;
 wire _15072_;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire _15078_;
 wire _15079_;
 wire _15080_;
 wire _15081_;
 wire _15082_;
 wire _15083_;
 wire _15084_;
 wire _15085_;
 wire _15086_;
 wire _15087_;
 wire _15088_;
 wire _15089_;
 wire _15090_;
 wire _15091_;
 wire _15092_;
 wire _15093_;
 wire _15094_;
 wire _15095_;
 wire _15096_;
 wire _15097_;
 wire _15098_;
 wire _15099_;
 wire _15100_;
 wire _15101_;
 wire _15102_;
 wire clknet_leaf_0_clk;
 wire \cpu.addr[10] ;
 wire \cpu.addr[11] ;
 wire \cpu.addr[12] ;
 wire \cpu.addr[13] ;
 wire \cpu.addr[14] ;
 wire \cpu.addr[15] ;
 wire \cpu.addr[1] ;
 wire \cpu.addr[2] ;
 wire \cpu.addr[3] ;
 wire \cpu.addr[4] ;
 wire \cpu.addr[5] ;
 wire \cpu.addr[6] ;
 wire \cpu.addr[7] ;
 wire \cpu.addr[8] ;
 wire \cpu.addr[9] ;
 wire \cpu.br ;
 wire \cpu.cond[0] ;
 wire \cpu.cond[1] ;
 wire \cpu.cond[2] ;
 wire \cpu.d_flush_all ;
 wire \cpu.d_rstrobe_d ;
 wire \cpu.d_wstrobe_d ;
 wire \cpu.dcache.flush_write ;
 wire \cpu.dcache.r_data[0][0] ;
 wire \cpu.dcache.r_data[0][10] ;
 wire \cpu.dcache.r_data[0][11] ;
 wire \cpu.dcache.r_data[0][12] ;
 wire \cpu.dcache.r_data[0][13] ;
 wire \cpu.dcache.r_data[0][14] ;
 wire \cpu.dcache.r_data[0][15] ;
 wire \cpu.dcache.r_data[0][16] ;
 wire \cpu.dcache.r_data[0][17] ;
 wire \cpu.dcache.r_data[0][18] ;
 wire \cpu.dcache.r_data[0][19] ;
 wire \cpu.dcache.r_data[0][1] ;
 wire \cpu.dcache.r_data[0][20] ;
 wire \cpu.dcache.r_data[0][21] ;
 wire \cpu.dcache.r_data[0][22] ;
 wire \cpu.dcache.r_data[0][23] ;
 wire \cpu.dcache.r_data[0][24] ;
 wire \cpu.dcache.r_data[0][25] ;
 wire \cpu.dcache.r_data[0][26] ;
 wire \cpu.dcache.r_data[0][27] ;
 wire \cpu.dcache.r_data[0][28] ;
 wire \cpu.dcache.r_data[0][29] ;
 wire \cpu.dcache.r_data[0][2] ;
 wire \cpu.dcache.r_data[0][30] ;
 wire \cpu.dcache.r_data[0][31] ;
 wire \cpu.dcache.r_data[0][3] ;
 wire \cpu.dcache.r_data[0][4] ;
 wire \cpu.dcache.r_data[0][5] ;
 wire \cpu.dcache.r_data[0][6] ;
 wire \cpu.dcache.r_data[0][7] ;
 wire \cpu.dcache.r_data[0][8] ;
 wire \cpu.dcache.r_data[0][9] ;
 wire \cpu.dcache.r_data[1][0] ;
 wire \cpu.dcache.r_data[1][10] ;
 wire \cpu.dcache.r_data[1][11] ;
 wire \cpu.dcache.r_data[1][12] ;
 wire \cpu.dcache.r_data[1][13] ;
 wire \cpu.dcache.r_data[1][14] ;
 wire \cpu.dcache.r_data[1][15] ;
 wire \cpu.dcache.r_data[1][16] ;
 wire \cpu.dcache.r_data[1][17] ;
 wire \cpu.dcache.r_data[1][18] ;
 wire \cpu.dcache.r_data[1][19] ;
 wire \cpu.dcache.r_data[1][1] ;
 wire \cpu.dcache.r_data[1][20] ;
 wire \cpu.dcache.r_data[1][21] ;
 wire \cpu.dcache.r_data[1][22] ;
 wire \cpu.dcache.r_data[1][23] ;
 wire \cpu.dcache.r_data[1][24] ;
 wire \cpu.dcache.r_data[1][25] ;
 wire \cpu.dcache.r_data[1][26] ;
 wire \cpu.dcache.r_data[1][27] ;
 wire \cpu.dcache.r_data[1][28] ;
 wire \cpu.dcache.r_data[1][29] ;
 wire \cpu.dcache.r_data[1][2] ;
 wire \cpu.dcache.r_data[1][30] ;
 wire \cpu.dcache.r_data[1][31] ;
 wire \cpu.dcache.r_data[1][3] ;
 wire \cpu.dcache.r_data[1][4] ;
 wire \cpu.dcache.r_data[1][5] ;
 wire \cpu.dcache.r_data[1][6] ;
 wire \cpu.dcache.r_data[1][7] ;
 wire \cpu.dcache.r_data[1][8] ;
 wire \cpu.dcache.r_data[1][9] ;
 wire \cpu.dcache.r_data[2][0] ;
 wire \cpu.dcache.r_data[2][10] ;
 wire \cpu.dcache.r_data[2][11] ;
 wire \cpu.dcache.r_data[2][12] ;
 wire \cpu.dcache.r_data[2][13] ;
 wire \cpu.dcache.r_data[2][14] ;
 wire \cpu.dcache.r_data[2][15] ;
 wire \cpu.dcache.r_data[2][16] ;
 wire \cpu.dcache.r_data[2][17] ;
 wire \cpu.dcache.r_data[2][18] ;
 wire \cpu.dcache.r_data[2][19] ;
 wire \cpu.dcache.r_data[2][1] ;
 wire \cpu.dcache.r_data[2][20] ;
 wire \cpu.dcache.r_data[2][21] ;
 wire \cpu.dcache.r_data[2][22] ;
 wire \cpu.dcache.r_data[2][23] ;
 wire \cpu.dcache.r_data[2][24] ;
 wire \cpu.dcache.r_data[2][25] ;
 wire \cpu.dcache.r_data[2][26] ;
 wire \cpu.dcache.r_data[2][27] ;
 wire \cpu.dcache.r_data[2][28] ;
 wire \cpu.dcache.r_data[2][29] ;
 wire \cpu.dcache.r_data[2][2] ;
 wire \cpu.dcache.r_data[2][30] ;
 wire \cpu.dcache.r_data[2][31] ;
 wire \cpu.dcache.r_data[2][3] ;
 wire \cpu.dcache.r_data[2][4] ;
 wire \cpu.dcache.r_data[2][5] ;
 wire \cpu.dcache.r_data[2][6] ;
 wire \cpu.dcache.r_data[2][7] ;
 wire \cpu.dcache.r_data[2][8] ;
 wire \cpu.dcache.r_data[2][9] ;
 wire \cpu.dcache.r_data[3][0] ;
 wire \cpu.dcache.r_data[3][10] ;
 wire \cpu.dcache.r_data[3][11] ;
 wire \cpu.dcache.r_data[3][12] ;
 wire \cpu.dcache.r_data[3][13] ;
 wire \cpu.dcache.r_data[3][14] ;
 wire \cpu.dcache.r_data[3][15] ;
 wire \cpu.dcache.r_data[3][16] ;
 wire \cpu.dcache.r_data[3][17] ;
 wire \cpu.dcache.r_data[3][18] ;
 wire \cpu.dcache.r_data[3][19] ;
 wire \cpu.dcache.r_data[3][1] ;
 wire \cpu.dcache.r_data[3][20] ;
 wire \cpu.dcache.r_data[3][21] ;
 wire \cpu.dcache.r_data[3][22] ;
 wire \cpu.dcache.r_data[3][23] ;
 wire \cpu.dcache.r_data[3][24] ;
 wire \cpu.dcache.r_data[3][25] ;
 wire \cpu.dcache.r_data[3][26] ;
 wire \cpu.dcache.r_data[3][27] ;
 wire \cpu.dcache.r_data[3][28] ;
 wire \cpu.dcache.r_data[3][29] ;
 wire \cpu.dcache.r_data[3][2] ;
 wire \cpu.dcache.r_data[3][30] ;
 wire \cpu.dcache.r_data[3][31] ;
 wire \cpu.dcache.r_data[3][3] ;
 wire \cpu.dcache.r_data[3][4] ;
 wire \cpu.dcache.r_data[3][5] ;
 wire \cpu.dcache.r_data[3][6] ;
 wire \cpu.dcache.r_data[3][7] ;
 wire \cpu.dcache.r_data[3][8] ;
 wire \cpu.dcache.r_data[3][9] ;
 wire \cpu.dcache.r_data[4][0] ;
 wire \cpu.dcache.r_data[4][10] ;
 wire \cpu.dcache.r_data[4][11] ;
 wire \cpu.dcache.r_data[4][12] ;
 wire \cpu.dcache.r_data[4][13] ;
 wire \cpu.dcache.r_data[4][14] ;
 wire \cpu.dcache.r_data[4][15] ;
 wire \cpu.dcache.r_data[4][16] ;
 wire \cpu.dcache.r_data[4][17] ;
 wire \cpu.dcache.r_data[4][18] ;
 wire \cpu.dcache.r_data[4][19] ;
 wire \cpu.dcache.r_data[4][1] ;
 wire \cpu.dcache.r_data[4][20] ;
 wire \cpu.dcache.r_data[4][21] ;
 wire \cpu.dcache.r_data[4][22] ;
 wire \cpu.dcache.r_data[4][23] ;
 wire \cpu.dcache.r_data[4][24] ;
 wire \cpu.dcache.r_data[4][25] ;
 wire \cpu.dcache.r_data[4][26] ;
 wire \cpu.dcache.r_data[4][27] ;
 wire \cpu.dcache.r_data[4][28] ;
 wire \cpu.dcache.r_data[4][29] ;
 wire \cpu.dcache.r_data[4][2] ;
 wire \cpu.dcache.r_data[4][30] ;
 wire \cpu.dcache.r_data[4][31] ;
 wire \cpu.dcache.r_data[4][3] ;
 wire \cpu.dcache.r_data[4][4] ;
 wire \cpu.dcache.r_data[4][5] ;
 wire \cpu.dcache.r_data[4][6] ;
 wire \cpu.dcache.r_data[4][7] ;
 wire \cpu.dcache.r_data[4][8] ;
 wire \cpu.dcache.r_data[4][9] ;
 wire \cpu.dcache.r_data[5][0] ;
 wire \cpu.dcache.r_data[5][10] ;
 wire \cpu.dcache.r_data[5][11] ;
 wire \cpu.dcache.r_data[5][12] ;
 wire \cpu.dcache.r_data[5][13] ;
 wire \cpu.dcache.r_data[5][14] ;
 wire \cpu.dcache.r_data[5][15] ;
 wire \cpu.dcache.r_data[5][16] ;
 wire \cpu.dcache.r_data[5][17] ;
 wire \cpu.dcache.r_data[5][18] ;
 wire \cpu.dcache.r_data[5][19] ;
 wire \cpu.dcache.r_data[5][1] ;
 wire \cpu.dcache.r_data[5][20] ;
 wire \cpu.dcache.r_data[5][21] ;
 wire \cpu.dcache.r_data[5][22] ;
 wire \cpu.dcache.r_data[5][23] ;
 wire \cpu.dcache.r_data[5][24] ;
 wire \cpu.dcache.r_data[5][25] ;
 wire \cpu.dcache.r_data[5][26] ;
 wire \cpu.dcache.r_data[5][27] ;
 wire \cpu.dcache.r_data[5][28] ;
 wire \cpu.dcache.r_data[5][29] ;
 wire \cpu.dcache.r_data[5][2] ;
 wire \cpu.dcache.r_data[5][30] ;
 wire \cpu.dcache.r_data[5][31] ;
 wire \cpu.dcache.r_data[5][3] ;
 wire \cpu.dcache.r_data[5][4] ;
 wire \cpu.dcache.r_data[5][5] ;
 wire \cpu.dcache.r_data[5][6] ;
 wire \cpu.dcache.r_data[5][7] ;
 wire \cpu.dcache.r_data[5][8] ;
 wire \cpu.dcache.r_data[5][9] ;
 wire \cpu.dcache.r_data[6][0] ;
 wire \cpu.dcache.r_data[6][10] ;
 wire \cpu.dcache.r_data[6][11] ;
 wire \cpu.dcache.r_data[6][12] ;
 wire \cpu.dcache.r_data[6][13] ;
 wire \cpu.dcache.r_data[6][14] ;
 wire \cpu.dcache.r_data[6][15] ;
 wire \cpu.dcache.r_data[6][16] ;
 wire \cpu.dcache.r_data[6][17] ;
 wire \cpu.dcache.r_data[6][18] ;
 wire \cpu.dcache.r_data[6][19] ;
 wire \cpu.dcache.r_data[6][1] ;
 wire \cpu.dcache.r_data[6][20] ;
 wire \cpu.dcache.r_data[6][21] ;
 wire \cpu.dcache.r_data[6][22] ;
 wire \cpu.dcache.r_data[6][23] ;
 wire \cpu.dcache.r_data[6][24] ;
 wire \cpu.dcache.r_data[6][25] ;
 wire \cpu.dcache.r_data[6][26] ;
 wire \cpu.dcache.r_data[6][27] ;
 wire \cpu.dcache.r_data[6][28] ;
 wire \cpu.dcache.r_data[6][29] ;
 wire \cpu.dcache.r_data[6][2] ;
 wire \cpu.dcache.r_data[6][30] ;
 wire \cpu.dcache.r_data[6][31] ;
 wire \cpu.dcache.r_data[6][3] ;
 wire \cpu.dcache.r_data[6][4] ;
 wire \cpu.dcache.r_data[6][5] ;
 wire \cpu.dcache.r_data[6][6] ;
 wire \cpu.dcache.r_data[6][7] ;
 wire \cpu.dcache.r_data[6][8] ;
 wire \cpu.dcache.r_data[6][9] ;
 wire \cpu.dcache.r_data[7][0] ;
 wire \cpu.dcache.r_data[7][10] ;
 wire \cpu.dcache.r_data[7][11] ;
 wire \cpu.dcache.r_data[7][12] ;
 wire \cpu.dcache.r_data[7][13] ;
 wire \cpu.dcache.r_data[7][14] ;
 wire \cpu.dcache.r_data[7][15] ;
 wire \cpu.dcache.r_data[7][16] ;
 wire \cpu.dcache.r_data[7][17] ;
 wire \cpu.dcache.r_data[7][18] ;
 wire \cpu.dcache.r_data[7][19] ;
 wire \cpu.dcache.r_data[7][1] ;
 wire \cpu.dcache.r_data[7][20] ;
 wire \cpu.dcache.r_data[7][21] ;
 wire \cpu.dcache.r_data[7][22] ;
 wire \cpu.dcache.r_data[7][23] ;
 wire \cpu.dcache.r_data[7][24] ;
 wire \cpu.dcache.r_data[7][25] ;
 wire \cpu.dcache.r_data[7][26] ;
 wire \cpu.dcache.r_data[7][27] ;
 wire \cpu.dcache.r_data[7][28] ;
 wire \cpu.dcache.r_data[7][29] ;
 wire \cpu.dcache.r_data[7][2] ;
 wire \cpu.dcache.r_data[7][30] ;
 wire \cpu.dcache.r_data[7][31] ;
 wire \cpu.dcache.r_data[7][3] ;
 wire \cpu.dcache.r_data[7][4] ;
 wire \cpu.dcache.r_data[7][5] ;
 wire \cpu.dcache.r_data[7][6] ;
 wire \cpu.dcache.r_data[7][7] ;
 wire \cpu.dcache.r_data[7][8] ;
 wire \cpu.dcache.r_data[7][9] ;
 wire \cpu.dcache.r_dirty[0] ;
 wire \cpu.dcache.r_dirty[1] ;
 wire \cpu.dcache.r_dirty[2] ;
 wire \cpu.dcache.r_dirty[3] ;
 wire \cpu.dcache.r_dirty[4] ;
 wire \cpu.dcache.r_dirty[5] ;
 wire \cpu.dcache.r_dirty[6] ;
 wire \cpu.dcache.r_dirty[7] ;
 wire \cpu.dcache.r_offset[0] ;
 wire \cpu.dcache.r_offset[1] ;
 wire \cpu.dcache.r_offset[2] ;
 wire \cpu.dcache.r_tag[0][10] ;
 wire \cpu.dcache.r_tag[0][11] ;
 wire \cpu.dcache.r_tag[0][12] ;
 wire \cpu.dcache.r_tag[0][13] ;
 wire \cpu.dcache.r_tag[0][14] ;
 wire \cpu.dcache.r_tag[0][15] ;
 wire \cpu.dcache.r_tag[0][16] ;
 wire \cpu.dcache.r_tag[0][17] ;
 wire \cpu.dcache.r_tag[0][18] ;
 wire \cpu.dcache.r_tag[0][19] ;
 wire \cpu.dcache.r_tag[0][20] ;
 wire \cpu.dcache.r_tag[0][21] ;
 wire \cpu.dcache.r_tag[0][22] ;
 wire \cpu.dcache.r_tag[0][23] ;
 wire \cpu.dcache.r_tag[0][5] ;
 wire \cpu.dcache.r_tag[0][6] ;
 wire \cpu.dcache.r_tag[0][7] ;
 wire \cpu.dcache.r_tag[0][8] ;
 wire \cpu.dcache.r_tag[0][9] ;
 wire \cpu.dcache.r_tag[1][10] ;
 wire \cpu.dcache.r_tag[1][11] ;
 wire \cpu.dcache.r_tag[1][12] ;
 wire \cpu.dcache.r_tag[1][13] ;
 wire \cpu.dcache.r_tag[1][14] ;
 wire \cpu.dcache.r_tag[1][15] ;
 wire \cpu.dcache.r_tag[1][16] ;
 wire \cpu.dcache.r_tag[1][17] ;
 wire \cpu.dcache.r_tag[1][18] ;
 wire \cpu.dcache.r_tag[1][19] ;
 wire \cpu.dcache.r_tag[1][20] ;
 wire \cpu.dcache.r_tag[1][21] ;
 wire \cpu.dcache.r_tag[1][22] ;
 wire \cpu.dcache.r_tag[1][23] ;
 wire \cpu.dcache.r_tag[1][5] ;
 wire \cpu.dcache.r_tag[1][6] ;
 wire \cpu.dcache.r_tag[1][7] ;
 wire \cpu.dcache.r_tag[1][8] ;
 wire \cpu.dcache.r_tag[1][9] ;
 wire \cpu.dcache.r_tag[2][10] ;
 wire \cpu.dcache.r_tag[2][11] ;
 wire \cpu.dcache.r_tag[2][12] ;
 wire \cpu.dcache.r_tag[2][13] ;
 wire \cpu.dcache.r_tag[2][14] ;
 wire \cpu.dcache.r_tag[2][15] ;
 wire \cpu.dcache.r_tag[2][16] ;
 wire \cpu.dcache.r_tag[2][17] ;
 wire \cpu.dcache.r_tag[2][18] ;
 wire \cpu.dcache.r_tag[2][19] ;
 wire \cpu.dcache.r_tag[2][20] ;
 wire \cpu.dcache.r_tag[2][21] ;
 wire \cpu.dcache.r_tag[2][22] ;
 wire \cpu.dcache.r_tag[2][23] ;
 wire \cpu.dcache.r_tag[2][5] ;
 wire \cpu.dcache.r_tag[2][6] ;
 wire \cpu.dcache.r_tag[2][7] ;
 wire \cpu.dcache.r_tag[2][8] ;
 wire \cpu.dcache.r_tag[2][9] ;
 wire \cpu.dcache.r_tag[3][10] ;
 wire \cpu.dcache.r_tag[3][11] ;
 wire \cpu.dcache.r_tag[3][12] ;
 wire \cpu.dcache.r_tag[3][13] ;
 wire \cpu.dcache.r_tag[3][14] ;
 wire \cpu.dcache.r_tag[3][15] ;
 wire \cpu.dcache.r_tag[3][16] ;
 wire \cpu.dcache.r_tag[3][17] ;
 wire \cpu.dcache.r_tag[3][18] ;
 wire \cpu.dcache.r_tag[3][19] ;
 wire \cpu.dcache.r_tag[3][20] ;
 wire \cpu.dcache.r_tag[3][21] ;
 wire \cpu.dcache.r_tag[3][22] ;
 wire \cpu.dcache.r_tag[3][23] ;
 wire \cpu.dcache.r_tag[3][5] ;
 wire \cpu.dcache.r_tag[3][6] ;
 wire \cpu.dcache.r_tag[3][7] ;
 wire \cpu.dcache.r_tag[3][8] ;
 wire \cpu.dcache.r_tag[3][9] ;
 wire \cpu.dcache.r_tag[4][10] ;
 wire \cpu.dcache.r_tag[4][11] ;
 wire \cpu.dcache.r_tag[4][12] ;
 wire \cpu.dcache.r_tag[4][13] ;
 wire \cpu.dcache.r_tag[4][14] ;
 wire \cpu.dcache.r_tag[4][15] ;
 wire \cpu.dcache.r_tag[4][16] ;
 wire \cpu.dcache.r_tag[4][17] ;
 wire \cpu.dcache.r_tag[4][18] ;
 wire \cpu.dcache.r_tag[4][19] ;
 wire \cpu.dcache.r_tag[4][20] ;
 wire \cpu.dcache.r_tag[4][21] ;
 wire \cpu.dcache.r_tag[4][22] ;
 wire \cpu.dcache.r_tag[4][23] ;
 wire \cpu.dcache.r_tag[4][5] ;
 wire \cpu.dcache.r_tag[4][6] ;
 wire \cpu.dcache.r_tag[4][7] ;
 wire \cpu.dcache.r_tag[4][8] ;
 wire \cpu.dcache.r_tag[4][9] ;
 wire \cpu.dcache.r_tag[5][10] ;
 wire \cpu.dcache.r_tag[5][11] ;
 wire \cpu.dcache.r_tag[5][12] ;
 wire \cpu.dcache.r_tag[5][13] ;
 wire \cpu.dcache.r_tag[5][14] ;
 wire \cpu.dcache.r_tag[5][15] ;
 wire \cpu.dcache.r_tag[5][16] ;
 wire \cpu.dcache.r_tag[5][17] ;
 wire \cpu.dcache.r_tag[5][18] ;
 wire \cpu.dcache.r_tag[5][19] ;
 wire \cpu.dcache.r_tag[5][20] ;
 wire \cpu.dcache.r_tag[5][21] ;
 wire \cpu.dcache.r_tag[5][22] ;
 wire \cpu.dcache.r_tag[5][23] ;
 wire \cpu.dcache.r_tag[5][5] ;
 wire \cpu.dcache.r_tag[5][6] ;
 wire \cpu.dcache.r_tag[5][7] ;
 wire \cpu.dcache.r_tag[5][8] ;
 wire \cpu.dcache.r_tag[5][9] ;
 wire \cpu.dcache.r_tag[6][10] ;
 wire \cpu.dcache.r_tag[6][11] ;
 wire \cpu.dcache.r_tag[6][12] ;
 wire \cpu.dcache.r_tag[6][13] ;
 wire \cpu.dcache.r_tag[6][14] ;
 wire \cpu.dcache.r_tag[6][15] ;
 wire \cpu.dcache.r_tag[6][16] ;
 wire \cpu.dcache.r_tag[6][17] ;
 wire \cpu.dcache.r_tag[6][18] ;
 wire \cpu.dcache.r_tag[6][19] ;
 wire \cpu.dcache.r_tag[6][20] ;
 wire \cpu.dcache.r_tag[6][21] ;
 wire \cpu.dcache.r_tag[6][22] ;
 wire \cpu.dcache.r_tag[6][23] ;
 wire \cpu.dcache.r_tag[6][5] ;
 wire \cpu.dcache.r_tag[6][6] ;
 wire \cpu.dcache.r_tag[6][7] ;
 wire \cpu.dcache.r_tag[6][8] ;
 wire \cpu.dcache.r_tag[6][9] ;
 wire \cpu.dcache.r_tag[7][10] ;
 wire \cpu.dcache.r_tag[7][11] ;
 wire \cpu.dcache.r_tag[7][12] ;
 wire \cpu.dcache.r_tag[7][13] ;
 wire \cpu.dcache.r_tag[7][14] ;
 wire \cpu.dcache.r_tag[7][15] ;
 wire \cpu.dcache.r_tag[7][16] ;
 wire \cpu.dcache.r_tag[7][17] ;
 wire \cpu.dcache.r_tag[7][18] ;
 wire \cpu.dcache.r_tag[7][19] ;
 wire \cpu.dcache.r_tag[7][20] ;
 wire \cpu.dcache.r_tag[7][21] ;
 wire \cpu.dcache.r_tag[7][22] ;
 wire \cpu.dcache.r_tag[7][23] ;
 wire \cpu.dcache.r_tag[7][5] ;
 wire \cpu.dcache.r_tag[7][6] ;
 wire \cpu.dcache.r_tag[7][7] ;
 wire \cpu.dcache.r_tag[7][8] ;
 wire \cpu.dcache.r_tag[7][9] ;
 wire \cpu.dcache.r_valid[0] ;
 wire \cpu.dcache.r_valid[1] ;
 wire \cpu.dcache.r_valid[2] ;
 wire \cpu.dcache.r_valid[3] ;
 wire \cpu.dcache.r_valid[4] ;
 wire \cpu.dcache.r_valid[5] ;
 wire \cpu.dcache.r_valid[6] ;
 wire \cpu.dcache.r_valid[7] ;
 wire \cpu.dcache.wdata[0] ;
 wire \cpu.dcache.wdata[10] ;
 wire \cpu.dcache.wdata[11] ;
 wire \cpu.dcache.wdata[12] ;
 wire \cpu.dcache.wdata[13] ;
 wire \cpu.dcache.wdata[14] ;
 wire \cpu.dcache.wdata[15] ;
 wire \cpu.dcache.wdata[1] ;
 wire \cpu.dcache.wdata[2] ;
 wire \cpu.dcache.wdata[3] ;
 wire \cpu.dcache.wdata[4] ;
 wire \cpu.dcache.wdata[5] ;
 wire \cpu.dcache.wdata[6] ;
 wire \cpu.dcache.wdata[7] ;
 wire \cpu.dcache.wdata[8] ;
 wire \cpu.dcache.wdata[9] ;
 wire \cpu.dec.div ;
 wire \cpu.dec.do_flush_all ;
 wire \cpu.dec.do_flush_write ;
 wire \cpu.dec.do_inv_mmu ;
 wire \cpu.dec.imm[0] ;
 wire \cpu.dec.imm[10] ;
 wire \cpu.dec.imm[11] ;
 wire \cpu.dec.imm[12] ;
 wire \cpu.dec.imm[13] ;
 wire \cpu.dec.imm[14] ;
 wire \cpu.dec.imm[15] ;
 wire \cpu.dec.imm[1] ;
 wire \cpu.dec.imm[2] ;
 wire \cpu.dec.imm[3] ;
 wire \cpu.dec.imm[4] ;
 wire \cpu.dec.imm[5] ;
 wire \cpu.dec.imm[6] ;
 wire \cpu.dec.imm[7] ;
 wire \cpu.dec.imm[8] ;
 wire \cpu.dec.imm[9] ;
 wire \cpu.dec.io ;
 wire \cpu.dec.iready ;
 wire \cpu.dec.jmp ;
 wire \cpu.dec.load ;
 wire \cpu.dec.mult ;
 wire \cpu.dec.needs_rs2 ;
 wire \cpu.dec.r_op[10] ;
 wire \cpu.dec.r_op[1] ;
 wire \cpu.dec.r_op[2] ;
 wire \cpu.dec.r_op[3] ;
 wire \cpu.dec.r_op[4] ;
 wire \cpu.dec.r_op[5] ;
 wire \cpu.dec.r_op[6] ;
 wire \cpu.dec.r_op[7] ;
 wire \cpu.dec.r_op[8] ;
 wire \cpu.dec.r_op[9] ;
 wire \cpu.dec.r_rd[0] ;
 wire \cpu.dec.r_rd[1] ;
 wire \cpu.dec.r_rd[2] ;
 wire \cpu.dec.r_rd[3] ;
 wire \cpu.dec.r_rs1[0] ;
 wire \cpu.dec.r_rs1[1] ;
 wire \cpu.dec.r_rs1[2] ;
 wire \cpu.dec.r_rs1[3] ;
 wire \cpu.dec.r_rs2[0] ;
 wire \cpu.dec.r_rs2[1] ;
 wire \cpu.dec.r_rs2[2] ;
 wire \cpu.dec.r_rs2[3] ;
 wire \cpu.dec.r_rs2_inv ;
 wire \cpu.dec.r_rs2_pc ;
 wire \cpu.dec.r_set_cc ;
 wire \cpu.dec.r_store ;
 wire \cpu.dec.r_swapsp ;
 wire \cpu.dec.r_sys_call ;
 wire \cpu.dec.r_trap ;
 wire \cpu.dec.supmode ;
 wire \cpu.dec.user_io ;
 wire \cpu.ex.c_div_running ;
 wire \cpu.ex.c_mult[0] ;
 wire \cpu.ex.c_mult[10] ;
 wire \cpu.ex.c_mult[11] ;
 wire \cpu.ex.c_mult[12] ;
 wire \cpu.ex.c_mult[13] ;
 wire \cpu.ex.c_mult[14] ;
 wire \cpu.ex.c_mult[15] ;
 wire \cpu.ex.c_mult[1] ;
 wire \cpu.ex.c_mult[2] ;
 wire \cpu.ex.c_mult[3] ;
 wire \cpu.ex.c_mult[4] ;
 wire \cpu.ex.c_mult[5] ;
 wire \cpu.ex.c_mult[6] ;
 wire \cpu.ex.c_mult[7] ;
 wire \cpu.ex.c_mult[8] ;
 wire \cpu.ex.c_mult[9] ;
 wire \cpu.ex.c_mult_off[0] ;
 wire \cpu.ex.c_mult_off[1] ;
 wire \cpu.ex.c_mult_off[2] ;
 wire \cpu.ex.c_mult_off[3] ;
 wire \cpu.ex.c_mult_running ;
 wire \cpu.ex.genblk3.c_supmode ;
 wire \cpu.ex.genblk3.r_mmu_d_proxy ;
 wire \cpu.ex.genblk3.r_mmu_enable ;
 wire \cpu.ex.genblk3.r_prev_supmode ;
 wire \cpu.ex.i_flush_all ;
 wire \cpu.ex.ifetch ;
 wire \cpu.ex.io_access ;
 wire \cpu.ex.mmu_read[12] ;
 wire \cpu.ex.mmu_read[13] ;
 wire \cpu.ex.mmu_read[14] ;
 wire \cpu.ex.mmu_read[15] ;
 wire \cpu.ex.mmu_read[1] ;
 wire \cpu.ex.mmu_read[2] ;
 wire \cpu.ex.mmu_read[3] ;
 wire \cpu.ex.mmu_reg_data[0] ;
 wire \cpu.ex.pc[10] ;
 wire \cpu.ex.pc[11] ;
 wire \cpu.ex.pc[12] ;
 wire \cpu.ex.pc[13] ;
 wire \cpu.ex.pc[14] ;
 wire \cpu.ex.pc[15] ;
 wire \cpu.ex.pc[1] ;
 wire \cpu.ex.pc[2] ;
 wire \cpu.ex.pc[3] ;
 wire \cpu.ex.pc[4] ;
 wire \cpu.ex.pc[5] ;
 wire \cpu.ex.pc[6] ;
 wire \cpu.ex.pc[7] ;
 wire \cpu.ex.pc[8] ;
 wire \cpu.ex.pc[9] ;
 wire \cpu.ex.r_10[0] ;
 wire \cpu.ex.r_10[10] ;
 wire \cpu.ex.r_10[11] ;
 wire \cpu.ex.r_10[12] ;
 wire \cpu.ex.r_10[13] ;
 wire \cpu.ex.r_10[14] ;
 wire \cpu.ex.r_10[15] ;
 wire \cpu.ex.r_10[1] ;
 wire \cpu.ex.r_10[2] ;
 wire \cpu.ex.r_10[3] ;
 wire \cpu.ex.r_10[4] ;
 wire \cpu.ex.r_10[5] ;
 wire \cpu.ex.r_10[6] ;
 wire \cpu.ex.r_10[7] ;
 wire \cpu.ex.r_10[8] ;
 wire \cpu.ex.r_10[9] ;
 wire \cpu.ex.r_11[0] ;
 wire \cpu.ex.r_11[10] ;
 wire \cpu.ex.r_11[11] ;
 wire \cpu.ex.r_11[12] ;
 wire \cpu.ex.r_11[13] ;
 wire \cpu.ex.r_11[14] ;
 wire \cpu.ex.r_11[15] ;
 wire \cpu.ex.r_11[1] ;
 wire \cpu.ex.r_11[2] ;
 wire \cpu.ex.r_11[3] ;
 wire \cpu.ex.r_11[4] ;
 wire \cpu.ex.r_11[5] ;
 wire \cpu.ex.r_11[6] ;
 wire \cpu.ex.r_11[7] ;
 wire \cpu.ex.r_11[8] ;
 wire \cpu.ex.r_11[9] ;
 wire \cpu.ex.r_12[0] ;
 wire \cpu.ex.r_12[10] ;
 wire \cpu.ex.r_12[11] ;
 wire \cpu.ex.r_12[12] ;
 wire \cpu.ex.r_12[13] ;
 wire \cpu.ex.r_12[14] ;
 wire \cpu.ex.r_12[15] ;
 wire \cpu.ex.r_12[1] ;
 wire \cpu.ex.r_12[2] ;
 wire \cpu.ex.r_12[3] ;
 wire \cpu.ex.r_12[4] ;
 wire \cpu.ex.r_12[5] ;
 wire \cpu.ex.r_12[6] ;
 wire \cpu.ex.r_12[7] ;
 wire \cpu.ex.r_12[8] ;
 wire \cpu.ex.r_12[9] ;
 wire \cpu.ex.r_13[0] ;
 wire \cpu.ex.r_13[10] ;
 wire \cpu.ex.r_13[11] ;
 wire \cpu.ex.r_13[12] ;
 wire \cpu.ex.r_13[13] ;
 wire \cpu.ex.r_13[14] ;
 wire \cpu.ex.r_13[15] ;
 wire \cpu.ex.r_13[1] ;
 wire \cpu.ex.r_13[2] ;
 wire \cpu.ex.r_13[3] ;
 wire \cpu.ex.r_13[4] ;
 wire \cpu.ex.r_13[5] ;
 wire \cpu.ex.r_13[6] ;
 wire \cpu.ex.r_13[7] ;
 wire \cpu.ex.r_13[8] ;
 wire \cpu.ex.r_13[9] ;
 wire \cpu.ex.r_14[0] ;
 wire \cpu.ex.r_14[10] ;
 wire \cpu.ex.r_14[11] ;
 wire \cpu.ex.r_14[12] ;
 wire \cpu.ex.r_14[13] ;
 wire \cpu.ex.r_14[14] ;
 wire \cpu.ex.r_14[15] ;
 wire \cpu.ex.r_14[1] ;
 wire \cpu.ex.r_14[2] ;
 wire \cpu.ex.r_14[3] ;
 wire \cpu.ex.r_14[4] ;
 wire \cpu.ex.r_14[5] ;
 wire \cpu.ex.r_14[6] ;
 wire \cpu.ex.r_14[7] ;
 wire \cpu.ex.r_14[8] ;
 wire \cpu.ex.r_14[9] ;
 wire \cpu.ex.r_15[0] ;
 wire \cpu.ex.r_15[10] ;
 wire \cpu.ex.r_15[11] ;
 wire \cpu.ex.r_15[12] ;
 wire \cpu.ex.r_15[13] ;
 wire \cpu.ex.r_15[14] ;
 wire \cpu.ex.r_15[15] ;
 wire \cpu.ex.r_15[1] ;
 wire \cpu.ex.r_15[2] ;
 wire \cpu.ex.r_15[3] ;
 wire \cpu.ex.r_15[4] ;
 wire \cpu.ex.r_15[5] ;
 wire \cpu.ex.r_15[6] ;
 wire \cpu.ex.r_15[7] ;
 wire \cpu.ex.r_15[8] ;
 wire \cpu.ex.r_15[9] ;
 wire \cpu.ex.r_8[0] ;
 wire \cpu.ex.r_8[10] ;
 wire \cpu.ex.r_8[11] ;
 wire \cpu.ex.r_8[12] ;
 wire \cpu.ex.r_8[13] ;
 wire \cpu.ex.r_8[14] ;
 wire \cpu.ex.r_8[15] ;
 wire \cpu.ex.r_8[1] ;
 wire \cpu.ex.r_8[2] ;
 wire \cpu.ex.r_8[3] ;
 wire \cpu.ex.r_8[4] ;
 wire \cpu.ex.r_8[5] ;
 wire \cpu.ex.r_8[6] ;
 wire \cpu.ex.r_8[7] ;
 wire \cpu.ex.r_8[8] ;
 wire \cpu.ex.r_8[9] ;
 wire \cpu.ex.r_9[0] ;
 wire \cpu.ex.r_9[10] ;
 wire \cpu.ex.r_9[11] ;
 wire \cpu.ex.r_9[12] ;
 wire \cpu.ex.r_9[13] ;
 wire \cpu.ex.r_9[14] ;
 wire \cpu.ex.r_9[15] ;
 wire \cpu.ex.r_9[1] ;
 wire \cpu.ex.r_9[2] ;
 wire \cpu.ex.r_9[3] ;
 wire \cpu.ex.r_9[4] ;
 wire \cpu.ex.r_9[5] ;
 wire \cpu.ex.r_9[6] ;
 wire \cpu.ex.r_9[7] ;
 wire \cpu.ex.r_9[8] ;
 wire \cpu.ex.r_9[9] ;
 wire \cpu.ex.r_branch_stall ;
 wire \cpu.ex.r_cc ;
 wire \cpu.ex.r_div_running ;
 wire \cpu.ex.r_epc[10] ;
 wire \cpu.ex.r_epc[11] ;
 wire \cpu.ex.r_epc[12] ;
 wire \cpu.ex.r_epc[13] ;
 wire \cpu.ex.r_epc[14] ;
 wire \cpu.ex.r_epc[15] ;
 wire \cpu.ex.r_epc[1] ;
 wire \cpu.ex.r_epc[2] ;
 wire \cpu.ex.r_epc[3] ;
 wire \cpu.ex.r_epc[4] ;
 wire \cpu.ex.r_epc[5] ;
 wire \cpu.ex.r_epc[6] ;
 wire \cpu.ex.r_epc[7] ;
 wire \cpu.ex.r_epc[8] ;
 wire \cpu.ex.r_epc[9] ;
 wire \cpu.ex.r_ie ;
 wire \cpu.ex.r_lr[10] ;
 wire \cpu.ex.r_lr[11] ;
 wire \cpu.ex.r_lr[12] ;
 wire \cpu.ex.r_lr[13] ;
 wire \cpu.ex.r_lr[14] ;
 wire \cpu.ex.r_lr[15] ;
 wire \cpu.ex.r_lr[1] ;
 wire \cpu.ex.r_lr[2] ;
 wire \cpu.ex.r_lr[3] ;
 wire \cpu.ex.r_lr[4] ;
 wire \cpu.ex.r_lr[5] ;
 wire \cpu.ex.r_lr[6] ;
 wire \cpu.ex.r_lr[7] ;
 wire \cpu.ex.r_lr[8] ;
 wire \cpu.ex.r_lr[9] ;
 wire \cpu.ex.r_mult[0] ;
 wire \cpu.ex.r_mult[10] ;
 wire \cpu.ex.r_mult[11] ;
 wire \cpu.ex.r_mult[12] ;
 wire \cpu.ex.r_mult[13] ;
 wire \cpu.ex.r_mult[14] ;
 wire \cpu.ex.r_mult[15] ;
 wire \cpu.ex.r_mult[16] ;
 wire \cpu.ex.r_mult[17] ;
 wire \cpu.ex.r_mult[18] ;
 wire \cpu.ex.r_mult[19] ;
 wire \cpu.ex.r_mult[1] ;
 wire \cpu.ex.r_mult[20] ;
 wire \cpu.ex.r_mult[21] ;
 wire \cpu.ex.r_mult[22] ;
 wire \cpu.ex.r_mult[23] ;
 wire \cpu.ex.r_mult[24] ;
 wire \cpu.ex.r_mult[25] ;
 wire \cpu.ex.r_mult[26] ;
 wire \cpu.ex.r_mult[27] ;
 wire \cpu.ex.r_mult[28] ;
 wire \cpu.ex.r_mult[29] ;
 wire \cpu.ex.r_mult[2] ;
 wire \cpu.ex.r_mult[30] ;
 wire \cpu.ex.r_mult[31] ;
 wire \cpu.ex.r_mult[3] ;
 wire \cpu.ex.r_mult[4] ;
 wire \cpu.ex.r_mult[5] ;
 wire \cpu.ex.r_mult[6] ;
 wire \cpu.ex.r_mult[7] ;
 wire \cpu.ex.r_mult[8] ;
 wire \cpu.ex.r_mult[9] ;
 wire \cpu.ex.r_mult_off[0] ;
 wire \cpu.ex.r_mult_off[1] ;
 wire \cpu.ex.r_mult_off[2] ;
 wire \cpu.ex.r_mult_off[3] ;
 wire \cpu.ex.r_mult_running ;
 wire \cpu.ex.r_prev_ie ;
 wire \cpu.ex.r_read_stall ;
 wire \cpu.ex.r_set_cc ;
 wire \cpu.ex.r_sp[10] ;
 wire \cpu.ex.r_sp[11] ;
 wire \cpu.ex.r_sp[12] ;
 wire \cpu.ex.r_sp[13] ;
 wire \cpu.ex.r_sp[14] ;
 wire \cpu.ex.r_sp[15] ;
 wire \cpu.ex.r_sp[1] ;
 wire \cpu.ex.r_sp[2] ;
 wire \cpu.ex.r_sp[3] ;
 wire \cpu.ex.r_sp[4] ;
 wire \cpu.ex.r_sp[5] ;
 wire \cpu.ex.r_sp[6] ;
 wire \cpu.ex.r_sp[7] ;
 wire \cpu.ex.r_sp[8] ;
 wire \cpu.ex.r_sp[9] ;
 wire \cpu.ex.r_stmp[0] ;
 wire \cpu.ex.r_stmp[10] ;
 wire \cpu.ex.r_stmp[11] ;
 wire \cpu.ex.r_stmp[12] ;
 wire \cpu.ex.r_stmp[13] ;
 wire \cpu.ex.r_stmp[14] ;
 wire \cpu.ex.r_stmp[15] ;
 wire \cpu.ex.r_stmp[1] ;
 wire \cpu.ex.r_stmp[2] ;
 wire \cpu.ex.r_stmp[3] ;
 wire \cpu.ex.r_stmp[4] ;
 wire \cpu.ex.r_stmp[5] ;
 wire \cpu.ex.r_stmp[6] ;
 wire \cpu.ex.r_stmp[7] ;
 wire \cpu.ex.r_stmp[8] ;
 wire \cpu.ex.r_stmp[9] ;
 wire \cpu.ex.r_wb_addr[0] ;
 wire \cpu.ex.r_wb_addr[1] ;
 wire \cpu.ex.r_wb_addr[2] ;
 wire \cpu.ex.r_wb_addr[3] ;
 wire \cpu.ex.r_wb_swapsp ;
 wire \cpu.ex.r_wb_valid ;
 wire \cpu.ex.r_wmask[0] ;
 wire \cpu.ex.r_wmask[1] ;
 wire \cpu.genblk1.mmu.r_valid_d[0] ;
 wire \cpu.genblk1.mmu.r_valid_d[10] ;
 wire \cpu.genblk1.mmu.r_valid_d[11] ;
 wire \cpu.genblk1.mmu.r_valid_d[12] ;
 wire \cpu.genblk1.mmu.r_valid_d[13] ;
 wire \cpu.genblk1.mmu.r_valid_d[14] ;
 wire \cpu.genblk1.mmu.r_valid_d[15] ;
 wire \cpu.genblk1.mmu.r_valid_d[16] ;
 wire \cpu.genblk1.mmu.r_valid_d[17] ;
 wire \cpu.genblk1.mmu.r_valid_d[18] ;
 wire \cpu.genblk1.mmu.r_valid_d[19] ;
 wire \cpu.genblk1.mmu.r_valid_d[1] ;
 wire \cpu.genblk1.mmu.r_valid_d[20] ;
 wire \cpu.genblk1.mmu.r_valid_d[21] ;
 wire \cpu.genblk1.mmu.r_valid_d[22] ;
 wire \cpu.genblk1.mmu.r_valid_d[23] ;
 wire \cpu.genblk1.mmu.r_valid_d[24] ;
 wire \cpu.genblk1.mmu.r_valid_d[25] ;
 wire \cpu.genblk1.mmu.r_valid_d[26] ;
 wire \cpu.genblk1.mmu.r_valid_d[27] ;
 wire \cpu.genblk1.mmu.r_valid_d[28] ;
 wire \cpu.genblk1.mmu.r_valid_d[29] ;
 wire \cpu.genblk1.mmu.r_valid_d[2] ;
 wire \cpu.genblk1.mmu.r_valid_d[30] ;
 wire \cpu.genblk1.mmu.r_valid_d[31] ;
 wire \cpu.genblk1.mmu.r_valid_d[3] ;
 wire \cpu.genblk1.mmu.r_valid_d[4] ;
 wire \cpu.genblk1.mmu.r_valid_d[5] ;
 wire \cpu.genblk1.mmu.r_valid_d[6] ;
 wire \cpu.genblk1.mmu.r_valid_d[7] ;
 wire \cpu.genblk1.mmu.r_valid_d[8] ;
 wire \cpu.genblk1.mmu.r_valid_d[9] ;
 wire \cpu.genblk1.mmu.r_valid_i[0] ;
 wire \cpu.genblk1.mmu.r_valid_i[10] ;
 wire \cpu.genblk1.mmu.r_valid_i[11] ;
 wire \cpu.genblk1.mmu.r_valid_i[12] ;
 wire \cpu.genblk1.mmu.r_valid_i[13] ;
 wire \cpu.genblk1.mmu.r_valid_i[14] ;
 wire \cpu.genblk1.mmu.r_valid_i[15] ;
 wire \cpu.genblk1.mmu.r_valid_i[16] ;
 wire \cpu.genblk1.mmu.r_valid_i[17] ;
 wire \cpu.genblk1.mmu.r_valid_i[18] ;
 wire \cpu.genblk1.mmu.r_valid_i[19] ;
 wire \cpu.genblk1.mmu.r_valid_i[1] ;
 wire \cpu.genblk1.mmu.r_valid_i[20] ;
 wire \cpu.genblk1.mmu.r_valid_i[21] ;
 wire \cpu.genblk1.mmu.r_valid_i[22] ;
 wire \cpu.genblk1.mmu.r_valid_i[23] ;
 wire \cpu.genblk1.mmu.r_valid_i[24] ;
 wire \cpu.genblk1.mmu.r_valid_i[25] ;
 wire \cpu.genblk1.mmu.r_valid_i[26] ;
 wire \cpu.genblk1.mmu.r_valid_i[27] ;
 wire \cpu.genblk1.mmu.r_valid_i[28] ;
 wire \cpu.genblk1.mmu.r_valid_i[29] ;
 wire \cpu.genblk1.mmu.r_valid_i[2] ;
 wire \cpu.genblk1.mmu.r_valid_i[30] ;
 wire \cpu.genblk1.mmu.r_valid_i[31] ;
 wire \cpu.genblk1.mmu.r_valid_i[3] ;
 wire \cpu.genblk1.mmu.r_valid_i[4] ;
 wire \cpu.genblk1.mmu.r_valid_i[5] ;
 wire \cpu.genblk1.mmu.r_valid_i[6] ;
 wire \cpu.genblk1.mmu.r_valid_i[7] ;
 wire \cpu.genblk1.mmu.r_valid_i[8] ;
 wire \cpu.genblk1.mmu.r_valid_i[9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][9] ;
 wire \cpu.genblk1.mmu.r_writeable_d[0] ;
 wire \cpu.genblk1.mmu.r_writeable_d[10] ;
 wire \cpu.genblk1.mmu.r_writeable_d[11] ;
 wire \cpu.genblk1.mmu.r_writeable_d[12] ;
 wire \cpu.genblk1.mmu.r_writeable_d[13] ;
 wire \cpu.genblk1.mmu.r_writeable_d[14] ;
 wire \cpu.genblk1.mmu.r_writeable_d[15] ;
 wire \cpu.genblk1.mmu.r_writeable_d[16] ;
 wire \cpu.genblk1.mmu.r_writeable_d[17] ;
 wire \cpu.genblk1.mmu.r_writeable_d[18] ;
 wire \cpu.genblk1.mmu.r_writeable_d[19] ;
 wire \cpu.genblk1.mmu.r_writeable_d[1] ;
 wire \cpu.genblk1.mmu.r_writeable_d[20] ;
 wire \cpu.genblk1.mmu.r_writeable_d[21] ;
 wire \cpu.genblk1.mmu.r_writeable_d[22] ;
 wire \cpu.genblk1.mmu.r_writeable_d[23] ;
 wire \cpu.genblk1.mmu.r_writeable_d[24] ;
 wire \cpu.genblk1.mmu.r_writeable_d[25] ;
 wire \cpu.genblk1.mmu.r_writeable_d[26] ;
 wire \cpu.genblk1.mmu.r_writeable_d[27] ;
 wire \cpu.genblk1.mmu.r_writeable_d[28] ;
 wire \cpu.genblk1.mmu.r_writeable_d[29] ;
 wire \cpu.genblk1.mmu.r_writeable_d[2] ;
 wire \cpu.genblk1.mmu.r_writeable_d[30] ;
 wire \cpu.genblk1.mmu.r_writeable_d[31] ;
 wire \cpu.genblk1.mmu.r_writeable_d[3] ;
 wire \cpu.genblk1.mmu.r_writeable_d[4] ;
 wire \cpu.genblk1.mmu.r_writeable_d[5] ;
 wire \cpu.genblk1.mmu.r_writeable_d[6] ;
 wire \cpu.genblk1.mmu.r_writeable_d[7] ;
 wire \cpu.genblk1.mmu.r_writeable_d[8] ;
 wire \cpu.genblk1.mmu.r_writeable_d[9] ;
 wire \cpu.gpio.genblk1[3].srcs_o[0] ;
 wire \cpu.gpio.genblk1[3].srcs_o[11] ;
 wire \cpu.gpio.genblk1[3].srcs_o[1] ;
 wire \cpu.gpio.genblk1[3].srcs_o[2] ;
 wire \cpu.gpio.genblk1[3].srcs_o[3] ;
 wire \cpu.gpio.genblk1[3].srcs_o[4] ;
 wire \cpu.gpio.genblk1[3].srcs_o[5] ;
 wire \cpu.gpio.genblk1[3].srcs_o[6] ;
 wire \cpu.gpio.genblk1[3].srcs_o[7] ;
 wire \cpu.gpio.genblk1[3].srcs_o[8] ;
 wire \cpu.gpio.genblk1[4].srcs_o[0] ;
 wire \cpu.gpio.genblk1[5].srcs_o[0] ;
 wire \cpu.gpio.genblk1[6].srcs_o[0] ;
 wire \cpu.gpio.genblk1[7].srcs_o[0] ;
 wire \cpu.gpio.genblk2[4].srcs_io[0] ;
 wire \cpu.gpio.genblk2[5].srcs_io[0] ;
 wire \cpu.gpio.genblk2[6].srcs_io[0] ;
 wire \cpu.gpio.genblk2[7].srcs_io[0] ;
 wire \cpu.gpio.r_enable_in[0] ;
 wire \cpu.gpio.r_enable_in[1] ;
 wire \cpu.gpio.r_enable_in[2] ;
 wire \cpu.gpio.r_enable_in[3] ;
 wire \cpu.gpio.r_enable_in[4] ;
 wire \cpu.gpio.r_enable_in[5] ;
 wire \cpu.gpio.r_enable_in[6] ;
 wire \cpu.gpio.r_enable_in[7] ;
 wire \cpu.gpio.r_enable_io[4] ;
 wire \cpu.gpio.r_enable_io[5] ;
 wire \cpu.gpio.r_enable_io[6] ;
 wire \cpu.gpio.r_enable_io[7] ;
 wire \cpu.gpio.r_spi_miso_src[0][0] ;
 wire \cpu.gpio.r_spi_miso_src[0][1] ;
 wire \cpu.gpio.r_spi_miso_src[0][2] ;
 wire \cpu.gpio.r_spi_miso_src[0][3] ;
 wire \cpu.gpio.r_spi_miso_src[1][0] ;
 wire \cpu.gpio.r_spi_miso_src[1][1] ;
 wire \cpu.gpio.r_spi_miso_src[1][2] ;
 wire \cpu.gpio.r_spi_miso_src[1][3] ;
 wire \cpu.gpio.r_src_io[4][0] ;
 wire \cpu.gpio.r_src_io[4][1] ;
 wire \cpu.gpio.r_src_io[4][2] ;
 wire \cpu.gpio.r_src_io[4][3] ;
 wire \cpu.gpio.r_src_io[5][0] ;
 wire \cpu.gpio.r_src_io[5][1] ;
 wire \cpu.gpio.r_src_io[5][2] ;
 wire \cpu.gpio.r_src_io[5][3] ;
 wire \cpu.gpio.r_src_io[6][0] ;
 wire \cpu.gpio.r_src_io[6][1] ;
 wire \cpu.gpio.r_src_io[6][2] ;
 wire \cpu.gpio.r_src_io[6][3] ;
 wire \cpu.gpio.r_src_io[7][0] ;
 wire \cpu.gpio.r_src_io[7][1] ;
 wire \cpu.gpio.r_src_io[7][2] ;
 wire \cpu.gpio.r_src_io[7][3] ;
 wire \cpu.gpio.r_src_o[3][0] ;
 wire \cpu.gpio.r_src_o[3][1] ;
 wire \cpu.gpio.r_src_o[3][2] ;
 wire \cpu.gpio.r_src_o[3][3] ;
 wire \cpu.gpio.r_src_o[4][0] ;
 wire \cpu.gpio.r_src_o[4][1] ;
 wire \cpu.gpio.r_src_o[4][2] ;
 wire \cpu.gpio.r_src_o[4][3] ;
 wire \cpu.gpio.r_src_o[5][0] ;
 wire \cpu.gpio.r_src_o[5][1] ;
 wire \cpu.gpio.r_src_o[5][2] ;
 wire \cpu.gpio.r_src_o[5][3] ;
 wire \cpu.gpio.r_src_o[6][0] ;
 wire \cpu.gpio.r_src_o[6][1] ;
 wire \cpu.gpio.r_src_o[6][2] ;
 wire \cpu.gpio.r_src_o[6][3] ;
 wire \cpu.gpio.r_src_o[7][0] ;
 wire \cpu.gpio.r_src_o[7][1] ;
 wire \cpu.gpio.r_src_o[7][2] ;
 wire \cpu.gpio.r_src_o[7][3] ;
 wire \cpu.gpio.r_uart_rx_src[0] ;
 wire \cpu.gpio.r_uart_rx_src[1] ;
 wire \cpu.gpio.r_uart_rx_src[2] ;
 wire \cpu.gpio.uart_rx ;
 wire \cpu.i_wstrobe_d ;
 wire \cpu.icache.r_data[0][0] ;
 wire \cpu.icache.r_data[0][10] ;
 wire \cpu.icache.r_data[0][11] ;
 wire \cpu.icache.r_data[0][12] ;
 wire \cpu.icache.r_data[0][13] ;
 wire \cpu.icache.r_data[0][14] ;
 wire \cpu.icache.r_data[0][15] ;
 wire \cpu.icache.r_data[0][16] ;
 wire \cpu.icache.r_data[0][17] ;
 wire \cpu.icache.r_data[0][18] ;
 wire \cpu.icache.r_data[0][19] ;
 wire \cpu.icache.r_data[0][1] ;
 wire \cpu.icache.r_data[0][20] ;
 wire \cpu.icache.r_data[0][21] ;
 wire \cpu.icache.r_data[0][22] ;
 wire \cpu.icache.r_data[0][23] ;
 wire \cpu.icache.r_data[0][24] ;
 wire \cpu.icache.r_data[0][25] ;
 wire \cpu.icache.r_data[0][26] ;
 wire \cpu.icache.r_data[0][27] ;
 wire \cpu.icache.r_data[0][28] ;
 wire \cpu.icache.r_data[0][29] ;
 wire \cpu.icache.r_data[0][2] ;
 wire \cpu.icache.r_data[0][30] ;
 wire \cpu.icache.r_data[0][31] ;
 wire \cpu.icache.r_data[0][3] ;
 wire \cpu.icache.r_data[0][4] ;
 wire \cpu.icache.r_data[0][5] ;
 wire \cpu.icache.r_data[0][6] ;
 wire \cpu.icache.r_data[0][7] ;
 wire \cpu.icache.r_data[0][8] ;
 wire \cpu.icache.r_data[0][9] ;
 wire \cpu.icache.r_data[1][0] ;
 wire \cpu.icache.r_data[1][10] ;
 wire \cpu.icache.r_data[1][11] ;
 wire \cpu.icache.r_data[1][12] ;
 wire \cpu.icache.r_data[1][13] ;
 wire \cpu.icache.r_data[1][14] ;
 wire \cpu.icache.r_data[1][15] ;
 wire \cpu.icache.r_data[1][16] ;
 wire \cpu.icache.r_data[1][17] ;
 wire \cpu.icache.r_data[1][18] ;
 wire \cpu.icache.r_data[1][19] ;
 wire \cpu.icache.r_data[1][1] ;
 wire \cpu.icache.r_data[1][20] ;
 wire \cpu.icache.r_data[1][21] ;
 wire \cpu.icache.r_data[1][22] ;
 wire \cpu.icache.r_data[1][23] ;
 wire \cpu.icache.r_data[1][24] ;
 wire \cpu.icache.r_data[1][25] ;
 wire \cpu.icache.r_data[1][26] ;
 wire \cpu.icache.r_data[1][27] ;
 wire \cpu.icache.r_data[1][28] ;
 wire \cpu.icache.r_data[1][29] ;
 wire \cpu.icache.r_data[1][2] ;
 wire \cpu.icache.r_data[1][30] ;
 wire \cpu.icache.r_data[1][31] ;
 wire \cpu.icache.r_data[1][3] ;
 wire \cpu.icache.r_data[1][4] ;
 wire \cpu.icache.r_data[1][5] ;
 wire \cpu.icache.r_data[1][6] ;
 wire \cpu.icache.r_data[1][7] ;
 wire \cpu.icache.r_data[1][8] ;
 wire \cpu.icache.r_data[1][9] ;
 wire \cpu.icache.r_data[2][0] ;
 wire \cpu.icache.r_data[2][10] ;
 wire \cpu.icache.r_data[2][11] ;
 wire \cpu.icache.r_data[2][12] ;
 wire \cpu.icache.r_data[2][13] ;
 wire \cpu.icache.r_data[2][14] ;
 wire \cpu.icache.r_data[2][15] ;
 wire \cpu.icache.r_data[2][16] ;
 wire \cpu.icache.r_data[2][17] ;
 wire \cpu.icache.r_data[2][18] ;
 wire \cpu.icache.r_data[2][19] ;
 wire \cpu.icache.r_data[2][1] ;
 wire \cpu.icache.r_data[2][20] ;
 wire \cpu.icache.r_data[2][21] ;
 wire \cpu.icache.r_data[2][22] ;
 wire \cpu.icache.r_data[2][23] ;
 wire \cpu.icache.r_data[2][24] ;
 wire \cpu.icache.r_data[2][25] ;
 wire \cpu.icache.r_data[2][26] ;
 wire \cpu.icache.r_data[2][27] ;
 wire \cpu.icache.r_data[2][28] ;
 wire \cpu.icache.r_data[2][29] ;
 wire \cpu.icache.r_data[2][2] ;
 wire \cpu.icache.r_data[2][30] ;
 wire \cpu.icache.r_data[2][31] ;
 wire \cpu.icache.r_data[2][3] ;
 wire \cpu.icache.r_data[2][4] ;
 wire \cpu.icache.r_data[2][5] ;
 wire \cpu.icache.r_data[2][6] ;
 wire \cpu.icache.r_data[2][7] ;
 wire \cpu.icache.r_data[2][8] ;
 wire \cpu.icache.r_data[2][9] ;
 wire \cpu.icache.r_data[3][0] ;
 wire \cpu.icache.r_data[3][10] ;
 wire \cpu.icache.r_data[3][11] ;
 wire \cpu.icache.r_data[3][12] ;
 wire \cpu.icache.r_data[3][13] ;
 wire \cpu.icache.r_data[3][14] ;
 wire \cpu.icache.r_data[3][15] ;
 wire \cpu.icache.r_data[3][16] ;
 wire \cpu.icache.r_data[3][17] ;
 wire \cpu.icache.r_data[3][18] ;
 wire \cpu.icache.r_data[3][19] ;
 wire \cpu.icache.r_data[3][1] ;
 wire \cpu.icache.r_data[3][20] ;
 wire \cpu.icache.r_data[3][21] ;
 wire \cpu.icache.r_data[3][22] ;
 wire \cpu.icache.r_data[3][23] ;
 wire \cpu.icache.r_data[3][24] ;
 wire \cpu.icache.r_data[3][25] ;
 wire \cpu.icache.r_data[3][26] ;
 wire \cpu.icache.r_data[3][27] ;
 wire \cpu.icache.r_data[3][28] ;
 wire \cpu.icache.r_data[3][29] ;
 wire \cpu.icache.r_data[3][2] ;
 wire \cpu.icache.r_data[3][30] ;
 wire \cpu.icache.r_data[3][31] ;
 wire \cpu.icache.r_data[3][3] ;
 wire \cpu.icache.r_data[3][4] ;
 wire \cpu.icache.r_data[3][5] ;
 wire \cpu.icache.r_data[3][6] ;
 wire \cpu.icache.r_data[3][7] ;
 wire \cpu.icache.r_data[3][8] ;
 wire \cpu.icache.r_data[3][9] ;
 wire \cpu.icache.r_data[4][0] ;
 wire \cpu.icache.r_data[4][10] ;
 wire \cpu.icache.r_data[4][11] ;
 wire \cpu.icache.r_data[4][12] ;
 wire \cpu.icache.r_data[4][13] ;
 wire \cpu.icache.r_data[4][14] ;
 wire \cpu.icache.r_data[4][15] ;
 wire \cpu.icache.r_data[4][16] ;
 wire \cpu.icache.r_data[4][17] ;
 wire \cpu.icache.r_data[4][18] ;
 wire \cpu.icache.r_data[4][19] ;
 wire \cpu.icache.r_data[4][1] ;
 wire \cpu.icache.r_data[4][20] ;
 wire \cpu.icache.r_data[4][21] ;
 wire \cpu.icache.r_data[4][22] ;
 wire \cpu.icache.r_data[4][23] ;
 wire \cpu.icache.r_data[4][24] ;
 wire \cpu.icache.r_data[4][25] ;
 wire \cpu.icache.r_data[4][26] ;
 wire \cpu.icache.r_data[4][27] ;
 wire \cpu.icache.r_data[4][28] ;
 wire \cpu.icache.r_data[4][29] ;
 wire \cpu.icache.r_data[4][2] ;
 wire \cpu.icache.r_data[4][30] ;
 wire \cpu.icache.r_data[4][31] ;
 wire \cpu.icache.r_data[4][3] ;
 wire \cpu.icache.r_data[4][4] ;
 wire \cpu.icache.r_data[4][5] ;
 wire \cpu.icache.r_data[4][6] ;
 wire \cpu.icache.r_data[4][7] ;
 wire \cpu.icache.r_data[4][8] ;
 wire \cpu.icache.r_data[4][9] ;
 wire \cpu.icache.r_data[5][0] ;
 wire \cpu.icache.r_data[5][10] ;
 wire \cpu.icache.r_data[5][11] ;
 wire \cpu.icache.r_data[5][12] ;
 wire \cpu.icache.r_data[5][13] ;
 wire \cpu.icache.r_data[5][14] ;
 wire \cpu.icache.r_data[5][15] ;
 wire \cpu.icache.r_data[5][16] ;
 wire \cpu.icache.r_data[5][17] ;
 wire \cpu.icache.r_data[5][18] ;
 wire \cpu.icache.r_data[5][19] ;
 wire \cpu.icache.r_data[5][1] ;
 wire \cpu.icache.r_data[5][20] ;
 wire \cpu.icache.r_data[5][21] ;
 wire \cpu.icache.r_data[5][22] ;
 wire \cpu.icache.r_data[5][23] ;
 wire \cpu.icache.r_data[5][24] ;
 wire \cpu.icache.r_data[5][25] ;
 wire \cpu.icache.r_data[5][26] ;
 wire \cpu.icache.r_data[5][27] ;
 wire \cpu.icache.r_data[5][28] ;
 wire \cpu.icache.r_data[5][29] ;
 wire \cpu.icache.r_data[5][2] ;
 wire \cpu.icache.r_data[5][30] ;
 wire \cpu.icache.r_data[5][31] ;
 wire \cpu.icache.r_data[5][3] ;
 wire \cpu.icache.r_data[5][4] ;
 wire \cpu.icache.r_data[5][5] ;
 wire \cpu.icache.r_data[5][6] ;
 wire \cpu.icache.r_data[5][7] ;
 wire \cpu.icache.r_data[5][8] ;
 wire \cpu.icache.r_data[5][9] ;
 wire \cpu.icache.r_data[6][0] ;
 wire \cpu.icache.r_data[6][10] ;
 wire \cpu.icache.r_data[6][11] ;
 wire \cpu.icache.r_data[6][12] ;
 wire \cpu.icache.r_data[6][13] ;
 wire \cpu.icache.r_data[6][14] ;
 wire \cpu.icache.r_data[6][15] ;
 wire \cpu.icache.r_data[6][16] ;
 wire \cpu.icache.r_data[6][17] ;
 wire \cpu.icache.r_data[6][18] ;
 wire \cpu.icache.r_data[6][19] ;
 wire \cpu.icache.r_data[6][1] ;
 wire \cpu.icache.r_data[6][20] ;
 wire \cpu.icache.r_data[6][21] ;
 wire \cpu.icache.r_data[6][22] ;
 wire \cpu.icache.r_data[6][23] ;
 wire \cpu.icache.r_data[6][24] ;
 wire \cpu.icache.r_data[6][25] ;
 wire \cpu.icache.r_data[6][26] ;
 wire \cpu.icache.r_data[6][27] ;
 wire \cpu.icache.r_data[6][28] ;
 wire \cpu.icache.r_data[6][29] ;
 wire \cpu.icache.r_data[6][2] ;
 wire \cpu.icache.r_data[6][30] ;
 wire \cpu.icache.r_data[6][31] ;
 wire \cpu.icache.r_data[6][3] ;
 wire \cpu.icache.r_data[6][4] ;
 wire \cpu.icache.r_data[6][5] ;
 wire \cpu.icache.r_data[6][6] ;
 wire \cpu.icache.r_data[6][7] ;
 wire \cpu.icache.r_data[6][8] ;
 wire \cpu.icache.r_data[6][9] ;
 wire \cpu.icache.r_data[7][0] ;
 wire \cpu.icache.r_data[7][10] ;
 wire \cpu.icache.r_data[7][11] ;
 wire \cpu.icache.r_data[7][12] ;
 wire \cpu.icache.r_data[7][13] ;
 wire \cpu.icache.r_data[7][14] ;
 wire \cpu.icache.r_data[7][15] ;
 wire \cpu.icache.r_data[7][16] ;
 wire \cpu.icache.r_data[7][17] ;
 wire \cpu.icache.r_data[7][18] ;
 wire \cpu.icache.r_data[7][19] ;
 wire \cpu.icache.r_data[7][1] ;
 wire \cpu.icache.r_data[7][20] ;
 wire \cpu.icache.r_data[7][21] ;
 wire \cpu.icache.r_data[7][22] ;
 wire \cpu.icache.r_data[7][23] ;
 wire \cpu.icache.r_data[7][24] ;
 wire \cpu.icache.r_data[7][25] ;
 wire \cpu.icache.r_data[7][26] ;
 wire \cpu.icache.r_data[7][27] ;
 wire \cpu.icache.r_data[7][28] ;
 wire \cpu.icache.r_data[7][29] ;
 wire \cpu.icache.r_data[7][2] ;
 wire \cpu.icache.r_data[7][30] ;
 wire \cpu.icache.r_data[7][31] ;
 wire \cpu.icache.r_data[7][3] ;
 wire \cpu.icache.r_data[7][4] ;
 wire \cpu.icache.r_data[7][5] ;
 wire \cpu.icache.r_data[7][6] ;
 wire \cpu.icache.r_data[7][7] ;
 wire \cpu.icache.r_data[7][8] ;
 wire \cpu.icache.r_data[7][9] ;
 wire \cpu.icache.r_offset[0] ;
 wire \cpu.icache.r_offset[1] ;
 wire \cpu.icache.r_offset[2] ;
 wire \cpu.icache.r_tag[0][10] ;
 wire \cpu.icache.r_tag[0][11] ;
 wire \cpu.icache.r_tag[0][12] ;
 wire \cpu.icache.r_tag[0][13] ;
 wire \cpu.icache.r_tag[0][14] ;
 wire \cpu.icache.r_tag[0][15] ;
 wire \cpu.icache.r_tag[0][16] ;
 wire \cpu.icache.r_tag[0][17] ;
 wire \cpu.icache.r_tag[0][18] ;
 wire \cpu.icache.r_tag[0][19] ;
 wire \cpu.icache.r_tag[0][20] ;
 wire \cpu.icache.r_tag[0][21] ;
 wire \cpu.icache.r_tag[0][22] ;
 wire \cpu.icache.r_tag[0][23] ;
 wire \cpu.icache.r_tag[0][5] ;
 wire \cpu.icache.r_tag[0][6] ;
 wire \cpu.icache.r_tag[0][7] ;
 wire \cpu.icache.r_tag[0][8] ;
 wire \cpu.icache.r_tag[0][9] ;
 wire \cpu.icache.r_tag[1][10] ;
 wire \cpu.icache.r_tag[1][11] ;
 wire \cpu.icache.r_tag[1][12] ;
 wire \cpu.icache.r_tag[1][13] ;
 wire \cpu.icache.r_tag[1][14] ;
 wire \cpu.icache.r_tag[1][15] ;
 wire \cpu.icache.r_tag[1][16] ;
 wire \cpu.icache.r_tag[1][17] ;
 wire \cpu.icache.r_tag[1][18] ;
 wire \cpu.icache.r_tag[1][19] ;
 wire \cpu.icache.r_tag[1][20] ;
 wire \cpu.icache.r_tag[1][21] ;
 wire \cpu.icache.r_tag[1][22] ;
 wire \cpu.icache.r_tag[1][23] ;
 wire \cpu.icache.r_tag[1][5] ;
 wire \cpu.icache.r_tag[1][6] ;
 wire \cpu.icache.r_tag[1][7] ;
 wire \cpu.icache.r_tag[1][8] ;
 wire \cpu.icache.r_tag[1][9] ;
 wire \cpu.icache.r_tag[2][10] ;
 wire \cpu.icache.r_tag[2][11] ;
 wire \cpu.icache.r_tag[2][12] ;
 wire \cpu.icache.r_tag[2][13] ;
 wire \cpu.icache.r_tag[2][14] ;
 wire \cpu.icache.r_tag[2][15] ;
 wire \cpu.icache.r_tag[2][16] ;
 wire \cpu.icache.r_tag[2][17] ;
 wire \cpu.icache.r_tag[2][18] ;
 wire \cpu.icache.r_tag[2][19] ;
 wire \cpu.icache.r_tag[2][20] ;
 wire \cpu.icache.r_tag[2][21] ;
 wire \cpu.icache.r_tag[2][22] ;
 wire \cpu.icache.r_tag[2][23] ;
 wire \cpu.icache.r_tag[2][5] ;
 wire \cpu.icache.r_tag[2][6] ;
 wire \cpu.icache.r_tag[2][7] ;
 wire \cpu.icache.r_tag[2][8] ;
 wire \cpu.icache.r_tag[2][9] ;
 wire \cpu.icache.r_tag[3][10] ;
 wire \cpu.icache.r_tag[3][11] ;
 wire \cpu.icache.r_tag[3][12] ;
 wire \cpu.icache.r_tag[3][13] ;
 wire \cpu.icache.r_tag[3][14] ;
 wire \cpu.icache.r_tag[3][15] ;
 wire \cpu.icache.r_tag[3][16] ;
 wire \cpu.icache.r_tag[3][17] ;
 wire \cpu.icache.r_tag[3][18] ;
 wire \cpu.icache.r_tag[3][19] ;
 wire \cpu.icache.r_tag[3][20] ;
 wire \cpu.icache.r_tag[3][21] ;
 wire \cpu.icache.r_tag[3][22] ;
 wire \cpu.icache.r_tag[3][23] ;
 wire \cpu.icache.r_tag[3][5] ;
 wire \cpu.icache.r_tag[3][6] ;
 wire \cpu.icache.r_tag[3][7] ;
 wire \cpu.icache.r_tag[3][8] ;
 wire \cpu.icache.r_tag[3][9] ;
 wire \cpu.icache.r_tag[4][10] ;
 wire \cpu.icache.r_tag[4][11] ;
 wire \cpu.icache.r_tag[4][12] ;
 wire \cpu.icache.r_tag[4][13] ;
 wire \cpu.icache.r_tag[4][14] ;
 wire \cpu.icache.r_tag[4][15] ;
 wire \cpu.icache.r_tag[4][16] ;
 wire \cpu.icache.r_tag[4][17] ;
 wire \cpu.icache.r_tag[4][18] ;
 wire \cpu.icache.r_tag[4][19] ;
 wire \cpu.icache.r_tag[4][20] ;
 wire \cpu.icache.r_tag[4][21] ;
 wire \cpu.icache.r_tag[4][22] ;
 wire \cpu.icache.r_tag[4][23] ;
 wire \cpu.icache.r_tag[4][5] ;
 wire \cpu.icache.r_tag[4][6] ;
 wire \cpu.icache.r_tag[4][7] ;
 wire \cpu.icache.r_tag[4][8] ;
 wire \cpu.icache.r_tag[4][9] ;
 wire \cpu.icache.r_tag[5][10] ;
 wire \cpu.icache.r_tag[5][11] ;
 wire \cpu.icache.r_tag[5][12] ;
 wire \cpu.icache.r_tag[5][13] ;
 wire \cpu.icache.r_tag[5][14] ;
 wire \cpu.icache.r_tag[5][15] ;
 wire \cpu.icache.r_tag[5][16] ;
 wire \cpu.icache.r_tag[5][17] ;
 wire \cpu.icache.r_tag[5][18] ;
 wire \cpu.icache.r_tag[5][19] ;
 wire \cpu.icache.r_tag[5][20] ;
 wire \cpu.icache.r_tag[5][21] ;
 wire \cpu.icache.r_tag[5][22] ;
 wire \cpu.icache.r_tag[5][23] ;
 wire \cpu.icache.r_tag[5][5] ;
 wire \cpu.icache.r_tag[5][6] ;
 wire \cpu.icache.r_tag[5][7] ;
 wire \cpu.icache.r_tag[5][8] ;
 wire \cpu.icache.r_tag[5][9] ;
 wire \cpu.icache.r_tag[6][10] ;
 wire \cpu.icache.r_tag[6][11] ;
 wire \cpu.icache.r_tag[6][12] ;
 wire \cpu.icache.r_tag[6][13] ;
 wire \cpu.icache.r_tag[6][14] ;
 wire \cpu.icache.r_tag[6][15] ;
 wire \cpu.icache.r_tag[6][16] ;
 wire \cpu.icache.r_tag[6][17] ;
 wire \cpu.icache.r_tag[6][18] ;
 wire \cpu.icache.r_tag[6][19] ;
 wire \cpu.icache.r_tag[6][20] ;
 wire \cpu.icache.r_tag[6][21] ;
 wire \cpu.icache.r_tag[6][22] ;
 wire \cpu.icache.r_tag[6][23] ;
 wire \cpu.icache.r_tag[6][5] ;
 wire \cpu.icache.r_tag[6][6] ;
 wire \cpu.icache.r_tag[6][7] ;
 wire \cpu.icache.r_tag[6][8] ;
 wire \cpu.icache.r_tag[6][9] ;
 wire \cpu.icache.r_tag[7][10] ;
 wire \cpu.icache.r_tag[7][11] ;
 wire \cpu.icache.r_tag[7][12] ;
 wire \cpu.icache.r_tag[7][13] ;
 wire \cpu.icache.r_tag[7][14] ;
 wire \cpu.icache.r_tag[7][15] ;
 wire \cpu.icache.r_tag[7][16] ;
 wire \cpu.icache.r_tag[7][17] ;
 wire \cpu.icache.r_tag[7][18] ;
 wire \cpu.icache.r_tag[7][19] ;
 wire \cpu.icache.r_tag[7][20] ;
 wire \cpu.icache.r_tag[7][21] ;
 wire \cpu.icache.r_tag[7][22] ;
 wire \cpu.icache.r_tag[7][23] ;
 wire \cpu.icache.r_tag[7][5] ;
 wire \cpu.icache.r_tag[7][6] ;
 wire \cpu.icache.r_tag[7][7] ;
 wire \cpu.icache.r_tag[7][8] ;
 wire \cpu.icache.r_tag[7][9] ;
 wire \cpu.icache.r_valid[0] ;
 wire \cpu.icache.r_valid[1] ;
 wire \cpu.icache.r_valid[2] ;
 wire \cpu.icache.r_valid[3] ;
 wire \cpu.icache.r_valid[4] ;
 wire \cpu.icache.r_valid[5] ;
 wire \cpu.icache.r_valid[6] ;
 wire \cpu.icache.r_valid[7] ;
 wire \cpu.intr.r_clock ;
 wire \cpu.intr.r_clock_cmp[0] ;
 wire \cpu.intr.r_clock_cmp[10] ;
 wire \cpu.intr.r_clock_cmp[11] ;
 wire \cpu.intr.r_clock_cmp[12] ;
 wire \cpu.intr.r_clock_cmp[13] ;
 wire \cpu.intr.r_clock_cmp[14] ;
 wire \cpu.intr.r_clock_cmp[15] ;
 wire \cpu.intr.r_clock_cmp[16] ;
 wire \cpu.intr.r_clock_cmp[17] ;
 wire \cpu.intr.r_clock_cmp[18] ;
 wire \cpu.intr.r_clock_cmp[19] ;
 wire \cpu.intr.r_clock_cmp[1] ;
 wire \cpu.intr.r_clock_cmp[20] ;
 wire \cpu.intr.r_clock_cmp[21] ;
 wire \cpu.intr.r_clock_cmp[22] ;
 wire \cpu.intr.r_clock_cmp[23] ;
 wire \cpu.intr.r_clock_cmp[24] ;
 wire \cpu.intr.r_clock_cmp[25] ;
 wire \cpu.intr.r_clock_cmp[26] ;
 wire \cpu.intr.r_clock_cmp[27] ;
 wire \cpu.intr.r_clock_cmp[28] ;
 wire \cpu.intr.r_clock_cmp[29] ;
 wire \cpu.intr.r_clock_cmp[2] ;
 wire \cpu.intr.r_clock_cmp[30] ;
 wire \cpu.intr.r_clock_cmp[31] ;
 wire \cpu.intr.r_clock_cmp[3] ;
 wire \cpu.intr.r_clock_cmp[4] ;
 wire \cpu.intr.r_clock_cmp[5] ;
 wire \cpu.intr.r_clock_cmp[6] ;
 wire \cpu.intr.r_clock_cmp[7] ;
 wire \cpu.intr.r_clock_cmp[8] ;
 wire \cpu.intr.r_clock_cmp[9] ;
 wire \cpu.intr.r_clock_count[0] ;
 wire \cpu.intr.r_clock_count[10] ;
 wire \cpu.intr.r_clock_count[11] ;
 wire \cpu.intr.r_clock_count[12] ;
 wire \cpu.intr.r_clock_count[13] ;
 wire \cpu.intr.r_clock_count[14] ;
 wire \cpu.intr.r_clock_count[15] ;
 wire \cpu.intr.r_clock_count[16] ;
 wire \cpu.intr.r_clock_count[17] ;
 wire \cpu.intr.r_clock_count[18] ;
 wire \cpu.intr.r_clock_count[19] ;
 wire \cpu.intr.r_clock_count[1] ;
 wire \cpu.intr.r_clock_count[20] ;
 wire \cpu.intr.r_clock_count[21] ;
 wire \cpu.intr.r_clock_count[22] ;
 wire \cpu.intr.r_clock_count[23] ;
 wire \cpu.intr.r_clock_count[24] ;
 wire \cpu.intr.r_clock_count[25] ;
 wire \cpu.intr.r_clock_count[26] ;
 wire \cpu.intr.r_clock_count[27] ;
 wire \cpu.intr.r_clock_count[28] ;
 wire \cpu.intr.r_clock_count[29] ;
 wire \cpu.intr.r_clock_count[2] ;
 wire \cpu.intr.r_clock_count[30] ;
 wire \cpu.intr.r_clock_count[31] ;
 wire \cpu.intr.r_clock_count[3] ;
 wire \cpu.intr.r_clock_count[4] ;
 wire \cpu.intr.r_clock_count[5] ;
 wire \cpu.intr.r_clock_count[6] ;
 wire \cpu.intr.r_clock_count[7] ;
 wire \cpu.intr.r_clock_count[8] ;
 wire \cpu.intr.r_clock_count[9] ;
 wire \cpu.intr.r_enable[0] ;
 wire \cpu.intr.r_enable[1] ;
 wire \cpu.intr.r_enable[2] ;
 wire \cpu.intr.r_enable[3] ;
 wire \cpu.intr.r_enable[4] ;
 wire \cpu.intr.r_enable[5] ;
 wire \cpu.intr.r_swi ;
 wire \cpu.intr.r_timer ;
 wire \cpu.intr.r_timer_count[0] ;
 wire \cpu.intr.r_timer_count[10] ;
 wire \cpu.intr.r_timer_count[11] ;
 wire \cpu.intr.r_timer_count[12] ;
 wire \cpu.intr.r_timer_count[13] ;
 wire \cpu.intr.r_timer_count[14] ;
 wire \cpu.intr.r_timer_count[15] ;
 wire \cpu.intr.r_timer_count[16] ;
 wire \cpu.intr.r_timer_count[17] ;
 wire \cpu.intr.r_timer_count[18] ;
 wire \cpu.intr.r_timer_count[19] ;
 wire \cpu.intr.r_timer_count[1] ;
 wire \cpu.intr.r_timer_count[20] ;
 wire \cpu.intr.r_timer_count[21] ;
 wire \cpu.intr.r_timer_count[22] ;
 wire \cpu.intr.r_timer_count[23] ;
 wire \cpu.intr.r_timer_count[2] ;
 wire \cpu.intr.r_timer_count[3] ;
 wire \cpu.intr.r_timer_count[4] ;
 wire \cpu.intr.r_timer_count[5] ;
 wire \cpu.intr.r_timer_count[6] ;
 wire \cpu.intr.r_timer_count[7] ;
 wire \cpu.intr.r_timer_count[8] ;
 wire \cpu.intr.r_timer_count[9] ;
 wire \cpu.intr.r_timer_reload[0] ;
 wire \cpu.intr.r_timer_reload[10] ;
 wire \cpu.intr.r_timer_reload[11] ;
 wire \cpu.intr.r_timer_reload[12] ;
 wire \cpu.intr.r_timer_reload[13] ;
 wire \cpu.intr.r_timer_reload[14] ;
 wire \cpu.intr.r_timer_reload[15] ;
 wire \cpu.intr.r_timer_reload[16] ;
 wire \cpu.intr.r_timer_reload[17] ;
 wire \cpu.intr.r_timer_reload[18] ;
 wire \cpu.intr.r_timer_reload[19] ;
 wire \cpu.intr.r_timer_reload[1] ;
 wire \cpu.intr.r_timer_reload[20] ;
 wire \cpu.intr.r_timer_reload[21] ;
 wire \cpu.intr.r_timer_reload[22] ;
 wire \cpu.intr.r_timer_reload[23] ;
 wire \cpu.intr.r_timer_reload[2] ;
 wire \cpu.intr.r_timer_reload[3] ;
 wire \cpu.intr.r_timer_reload[4] ;
 wire \cpu.intr.r_timer_reload[5] ;
 wire \cpu.intr.r_timer_reload[6] ;
 wire \cpu.intr.r_timer_reload[7] ;
 wire \cpu.intr.r_timer_reload[8] ;
 wire \cpu.intr.r_timer_reload[9] ;
 wire \cpu.intr.spi_intr ;
 wire \cpu.qspi.c_rstrobe_d ;
 wire \cpu.qspi.c_wstrobe_d ;
 wire \cpu.qspi.c_wstrobe_i ;
 wire \cpu.qspi.r_count[0] ;
 wire \cpu.qspi.r_count[1] ;
 wire \cpu.qspi.r_count[2] ;
 wire \cpu.qspi.r_count[3] ;
 wire \cpu.qspi.r_count[4] ;
 wire \cpu.qspi.r_ind ;
 wire \cpu.qspi.r_mask[0] ;
 wire \cpu.qspi.r_mask[1] ;
 wire \cpu.qspi.r_mask[2] ;
 wire \cpu.qspi.r_quad[0] ;
 wire \cpu.qspi.r_quad[1] ;
 wire \cpu.qspi.r_quad[2] ;
 wire \cpu.qspi.r_read_delay[0][0] ;
 wire \cpu.qspi.r_read_delay[0][1] ;
 wire \cpu.qspi.r_read_delay[0][2] ;
 wire \cpu.qspi.r_read_delay[0][3] ;
 wire \cpu.qspi.r_read_delay[1][0] ;
 wire \cpu.qspi.r_read_delay[1][1] ;
 wire \cpu.qspi.r_read_delay[1][2] ;
 wire \cpu.qspi.r_read_delay[1][3] ;
 wire \cpu.qspi.r_read_delay[2][0] ;
 wire \cpu.qspi.r_read_delay[2][1] ;
 wire \cpu.qspi.r_read_delay[2][2] ;
 wire \cpu.qspi.r_read_delay[2][3] ;
 wire \cpu.qspi.r_rom_mode[0] ;
 wire \cpu.qspi.r_rom_mode[1] ;
 wire \cpu.qspi.r_state[0] ;
 wire \cpu.qspi.r_state[10] ;
 wire \cpu.qspi.r_state[11] ;
 wire \cpu.qspi.r_state[12] ;
 wire \cpu.qspi.r_state[13] ;
 wire \cpu.qspi.r_state[14] ;
 wire \cpu.qspi.r_state[15] ;
 wire \cpu.qspi.r_state[16] ;
 wire \cpu.qspi.r_state[17] ;
 wire \cpu.qspi.r_state[1] ;
 wire \cpu.qspi.r_state[2] ;
 wire \cpu.qspi.r_state[3] ;
 wire \cpu.qspi.r_state[4] ;
 wire \cpu.qspi.r_state[5] ;
 wire \cpu.qspi.r_state[6] ;
 wire \cpu.qspi.r_state[7] ;
 wire \cpu.qspi.r_state[8] ;
 wire \cpu.qspi.r_state[9] ;
 wire \cpu.r_clk_invert ;
 wire \cpu.spi.r_bits[0] ;
 wire \cpu.spi.r_bits[1] ;
 wire \cpu.spi.r_bits[2] ;
 wire \cpu.spi.r_clk_count[0][0] ;
 wire \cpu.spi.r_clk_count[0][1] ;
 wire \cpu.spi.r_clk_count[0][2] ;
 wire \cpu.spi.r_clk_count[0][3] ;
 wire \cpu.spi.r_clk_count[0][4] ;
 wire \cpu.spi.r_clk_count[0][5] ;
 wire \cpu.spi.r_clk_count[0][6] ;
 wire \cpu.spi.r_clk_count[0][7] ;
 wire \cpu.spi.r_clk_count[1][0] ;
 wire \cpu.spi.r_clk_count[1][1] ;
 wire \cpu.spi.r_clk_count[1][2] ;
 wire \cpu.spi.r_clk_count[1][3] ;
 wire \cpu.spi.r_clk_count[1][4] ;
 wire \cpu.spi.r_clk_count[1][5] ;
 wire \cpu.spi.r_clk_count[1][6] ;
 wire \cpu.spi.r_clk_count[1][7] ;
 wire \cpu.spi.r_clk_count[2][0] ;
 wire \cpu.spi.r_clk_count[2][1] ;
 wire \cpu.spi.r_clk_count[2][2] ;
 wire \cpu.spi.r_clk_count[2][3] ;
 wire \cpu.spi.r_clk_count[2][4] ;
 wire \cpu.spi.r_clk_count[2][5] ;
 wire \cpu.spi.r_clk_count[2][6] ;
 wire \cpu.spi.r_clk_count[2][7] ;
 wire \cpu.spi.r_count[0] ;
 wire \cpu.spi.r_count[1] ;
 wire \cpu.spi.r_count[2] ;
 wire \cpu.spi.r_count[3] ;
 wire \cpu.spi.r_count[4] ;
 wire \cpu.spi.r_count[5] ;
 wire \cpu.spi.r_count[6] ;
 wire \cpu.spi.r_count[7] ;
 wire \cpu.spi.r_in[0] ;
 wire \cpu.spi.r_in[1] ;
 wire \cpu.spi.r_in[2] ;
 wire \cpu.spi.r_in[3] ;
 wire \cpu.spi.r_in[4] ;
 wire \cpu.spi.r_in[5] ;
 wire \cpu.spi.r_in[6] ;
 wire \cpu.spi.r_in[7] ;
 wire \cpu.spi.r_mode[0][0] ;
 wire \cpu.spi.r_mode[0][1] ;
 wire \cpu.spi.r_mode[1][0] ;
 wire \cpu.spi.r_mode[1][1] ;
 wire \cpu.spi.r_mode[2][0] ;
 wire \cpu.spi.r_mode[2][1] ;
 wire \cpu.spi.r_out[0] ;
 wire \cpu.spi.r_out[1] ;
 wire \cpu.spi.r_out[2] ;
 wire \cpu.spi.r_out[3] ;
 wire \cpu.spi.r_out[4] ;
 wire \cpu.spi.r_out[5] ;
 wire \cpu.spi.r_out[6] ;
 wire \cpu.spi.r_out[7] ;
 wire \cpu.spi.r_ready ;
 wire \cpu.spi.r_searching ;
 wire \cpu.spi.r_sel[0] ;
 wire \cpu.spi.r_sel[1] ;
 wire \cpu.spi.r_src[0] ;
 wire \cpu.spi.r_src[1] ;
 wire \cpu.spi.r_src[2] ;
 wire \cpu.spi.r_state[0] ;
 wire \cpu.spi.r_state[1] ;
 wire \cpu.spi.r_state[2] ;
 wire \cpu.spi.r_state[3] ;
 wire \cpu.spi.r_state[4] ;
 wire \cpu.spi.r_state[5] ;
 wire \cpu.spi.r_state[6] ;
 wire \cpu.spi.r_timeout[0] ;
 wire \cpu.spi.r_timeout[1] ;
 wire \cpu.spi.r_timeout[2] ;
 wire \cpu.spi.r_timeout[3] ;
 wire \cpu.spi.r_timeout[4] ;
 wire \cpu.spi.r_timeout[5] ;
 wire \cpu.spi.r_timeout[6] ;
 wire \cpu.spi.r_timeout[7] ;
 wire \cpu.spi.r_timeout_count[0] ;
 wire \cpu.spi.r_timeout_count[1] ;
 wire \cpu.spi.r_timeout_count[2] ;
 wire \cpu.spi.r_timeout_count[3] ;
 wire \cpu.spi.r_timeout_count[4] ;
 wire \cpu.spi.r_timeout_count[5] ;
 wire \cpu.spi.r_timeout_count[6] ;
 wire \cpu.spi.r_timeout_count[7] ;
 wire \cpu.uart.r_div[0] ;
 wire \cpu.uart.r_div[10] ;
 wire \cpu.uart.r_div[11] ;
 wire \cpu.uart.r_div[1] ;
 wire \cpu.uart.r_div[2] ;
 wire \cpu.uart.r_div[3] ;
 wire \cpu.uart.r_div[4] ;
 wire \cpu.uart.r_div[5] ;
 wire \cpu.uart.r_div[6] ;
 wire \cpu.uart.r_div[7] ;
 wire \cpu.uart.r_div[8] ;
 wire \cpu.uart.r_div[9] ;
 wire \cpu.uart.r_div_value[0] ;
 wire \cpu.uart.r_div_value[10] ;
 wire \cpu.uart.r_div_value[11] ;
 wire \cpu.uart.r_div_value[1] ;
 wire \cpu.uart.r_div_value[2] ;
 wire \cpu.uart.r_div_value[3] ;
 wire \cpu.uart.r_div_value[4] ;
 wire \cpu.uart.r_div_value[5] ;
 wire \cpu.uart.r_div_value[6] ;
 wire \cpu.uart.r_div_value[7] ;
 wire \cpu.uart.r_div_value[8] ;
 wire \cpu.uart.r_div_value[9] ;
 wire \cpu.uart.r_ib[0] ;
 wire \cpu.uart.r_ib[1] ;
 wire \cpu.uart.r_ib[2] ;
 wire \cpu.uart.r_ib[3] ;
 wire \cpu.uart.r_ib[4] ;
 wire \cpu.uart.r_ib[5] ;
 wire \cpu.uart.r_ib[6] ;
 wire \cpu.uart.r_in[0] ;
 wire \cpu.uart.r_in[1] ;
 wire \cpu.uart.r_in[2] ;
 wire \cpu.uart.r_in[3] ;
 wire \cpu.uart.r_in[4] ;
 wire \cpu.uart.r_in[5] ;
 wire \cpu.uart.r_in[6] ;
 wire \cpu.uart.r_in[7] ;
 wire \cpu.uart.r_out[0] ;
 wire \cpu.uart.r_out[1] ;
 wire \cpu.uart.r_out[2] ;
 wire \cpu.uart.r_out[3] ;
 wire \cpu.uart.r_out[4] ;
 wire \cpu.uart.r_out[5] ;
 wire \cpu.uart.r_out[6] ;
 wire \cpu.uart.r_out[7] ;
 wire \cpu.uart.r_r ;
 wire \cpu.uart.r_r_int ;
 wire \cpu.uart.r_r_invert ;
 wire \cpu.uart.r_rcnt[0] ;
 wire \cpu.uart.r_rcnt[1] ;
 wire \cpu.uart.r_rstate[0] ;
 wire \cpu.uart.r_rstate[1] ;
 wire \cpu.uart.r_rstate[2] ;
 wire \cpu.uart.r_rstate[3] ;
 wire \cpu.uart.r_x_int ;
 wire \cpu.uart.r_x_invert ;
 wire \cpu.uart.r_xcnt[0] ;
 wire \cpu.uart.r_xcnt[1] ;
 wire \cpu.uart.r_xstate[0] ;
 wire \cpu.uart.r_xstate[1] ;
 wire \cpu.uart.r_xstate[2] ;
 wire \cpu.uart.r_xstate[3] ;
 wire r_reset;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_253_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_257_clk;
 wire clknet_leaf_258_clk;
 wire clknet_leaf_259_clk;
 wire clknet_leaf_260_clk;
 wire clknet_leaf_261_clk;
 wire clknet_leaf_262_clk;
 wire clknet_leaf_263_clk;
 wire clknet_leaf_264_clk;
 wire clknet_leaf_265_clk;
 wire clknet_leaf_266_clk;
 wire clknet_leaf_267_clk;
 wire clknet_leaf_268_clk;
 wire clknet_leaf_269_clk;
 wire clknet_leaf_270_clk;
 wire clknet_leaf_271_clk;
 wire clknet_leaf_272_clk;
 wire clknet_leaf_273_clk;
 wire clknet_leaf_274_clk;
 wire clknet_leaf_275_clk;
 wire clknet_leaf_276_clk;
 wire clknet_leaf_277_clk;
 wire clknet_leaf_278_clk;
 wire clknet_leaf_279_clk;
 wire clknet_leaf_280_clk;
 wire clknet_leaf_281_clk;
 wire clknet_leaf_282_clk;
 wire clknet_leaf_283_clk;
 wire clknet_leaf_284_clk;
 wire clknet_leaf_285_clk;
 wire clknet_leaf_286_clk;
 wire clknet_leaf_287_clk;
 wire clknet_leaf_288_clk;
 wire clknet_leaf_289_clk;
 wire clknet_leaf_290_clk;
 wire clknet_leaf_291_clk;
 wire clknet_leaf_292_clk;
 wire clknet_leaf_293_clk;
 wire clknet_leaf_294_clk;
 wire clknet_leaf_295_clk;
 wire clknet_leaf_296_clk;
 wire clknet_leaf_297_clk;
 wire clknet_leaf_298_clk;
 wire clknet_leaf_299_clk;
 wire clknet_leaf_300_clk;
 wire clknet_leaf_301_clk;
 wire clknet_leaf_302_clk;
 wire clknet_leaf_303_clk;
 wire clknet_leaf_304_clk;
 wire clknet_leaf_305_clk;
 wire clknet_leaf_306_clk;
 wire clknet_leaf_307_clk;
 wire clknet_leaf_308_clk;
 wire clknet_leaf_309_clk;
 wire clknet_leaf_310_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_6_0__leaf_clk;
 wire clknet_6_1__leaf_clk;
 wire clknet_6_2__leaf_clk;
 wire clknet_6_3__leaf_clk;
 wire clknet_6_4__leaf_clk;
 wire clknet_6_5__leaf_clk;
 wire clknet_6_6__leaf_clk;
 wire clknet_6_7__leaf_clk;
 wire clknet_6_8__leaf_clk;
 wire clknet_6_9__leaf_clk;
 wire clknet_6_10__leaf_clk;
 wire clknet_6_11__leaf_clk;
 wire clknet_6_12__leaf_clk;
 wire clknet_6_13__leaf_clk;
 wire clknet_6_14__leaf_clk;
 wire clknet_6_15__leaf_clk;
 wire clknet_6_16__leaf_clk;
 wire clknet_6_17__leaf_clk;
 wire clknet_6_18__leaf_clk;
 wire clknet_6_19__leaf_clk;
 wire clknet_6_20__leaf_clk;
 wire clknet_6_21__leaf_clk;
 wire clknet_6_22__leaf_clk;
 wire clknet_6_23__leaf_clk;
 wire clknet_6_24__leaf_clk;
 wire clknet_6_25__leaf_clk;
 wire clknet_6_26__leaf_clk;
 wire clknet_6_27__leaf_clk;
 wire clknet_6_28__leaf_clk;
 wire clknet_6_29__leaf_clk;
 wire clknet_6_30__leaf_clk;
 wire clknet_6_31__leaf_clk;
 wire clknet_6_32__leaf_clk;
 wire clknet_6_33__leaf_clk;
 wire clknet_6_34__leaf_clk;
 wire clknet_6_35__leaf_clk;
 wire clknet_6_36__leaf_clk;
 wire clknet_6_37__leaf_clk;
 wire clknet_6_38__leaf_clk;
 wire clknet_6_39__leaf_clk;
 wire clknet_6_40__leaf_clk;
 wire clknet_6_41__leaf_clk;
 wire clknet_6_42__leaf_clk;
 wire clknet_6_43__leaf_clk;
 wire clknet_6_44__leaf_clk;
 wire clknet_6_45__leaf_clk;
 wire clknet_6_46__leaf_clk;
 wire clknet_6_47__leaf_clk;
 wire clknet_6_48__leaf_clk;
 wire clknet_6_49__leaf_clk;
 wire clknet_6_50__leaf_clk;
 wire clknet_6_51__leaf_clk;
 wire clknet_6_52__leaf_clk;
 wire clknet_6_53__leaf_clk;
 wire clknet_6_54__leaf_clk;
 wire clknet_6_55__leaf_clk;
 wire clknet_6_56__leaf_clk;
 wire clknet_6_57__leaf_clk;
 wire clknet_6_58__leaf_clk;
 wire clknet_6_59__leaf_clk;
 wire clknet_6_60__leaf_clk;
 wire clknet_6_61__leaf_clk;
 wire clknet_6_62__leaf_clk;
 wire clknet_6_63__leaf_clk;

 sg13g2_buf_1 _15104_ (.A(\cpu.dec.r_op[5] ),
    .X(_08372_));
 sg13g2_inv_2 _15105_ (.Y(_08373_),
    .A(net1135));
 sg13g2_inv_1 _15106_ (.Y(_08374_),
    .A(_00189_));
 sg13g2_buf_8 _15107_ (.A(\cpu.addr[13] ),
    .X(_08375_));
 sg13g2_buf_1 _15108_ (.A(\cpu.addr[15] ),
    .X(_08376_));
 sg13g2_buf_8 _15109_ (.A(_08376_),
    .X(_08377_));
 sg13g2_nor2_1 _15110_ (.A(net1134),
    .B(net1075),
    .Y(_08378_));
 sg13g2_buf_8 _15111_ (.A(\cpu.addr[12] ),
    .X(_08379_));
 sg13g2_buf_8 _15112_ (.A(\cpu.addr[14] ),
    .X(_08380_));
 sg13g2_buf_8 _15113_ (.A(_08380_),
    .X(_08381_));
 sg13g2_mux4_1 _15114_ (.S0(net1133),
    .A0(\cpu.genblk1.mmu.r_writeable_d[16] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[17] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[20] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[21] ),
    .S1(net1074),
    .X(_08382_));
 sg13g2_nand2_1 _15115_ (.Y(_08383_),
    .A(_08378_),
    .B(_08382_));
 sg13g2_buf_8 _15116_ (.A(net1133),
    .X(_08384_));
 sg13g2_nor2b_1 _15117_ (.A(_08376_),
    .B_N(net1134),
    .Y(_08385_));
 sg13g2_mux2_1 _15118_ (.A0(\cpu.genblk1.mmu.r_writeable_d[19] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[23] ),
    .S(_08380_),
    .X(_08386_));
 sg13g2_nand3_1 _15119_ (.B(_08385_),
    .C(_08386_),
    .A(net1073),
    .Y(_08387_));
 sg13g2_buf_8 _15120_ (.A(_00193_),
    .X(_08388_));
 sg13g2_buf_2 _15121_ (.A(\cpu.ex.r_wmask[1] ),
    .X(_08389_));
 sg13g2_buf_8 _15122_ (.A(\cpu.ex.r_wmask[0] ),
    .X(_08390_));
 sg13g2_nor2_1 _15123_ (.A(_08389_),
    .B(_08390_),
    .Y(_08391_));
 sg13g2_buf_8 _15124_ (.A(_08391_),
    .X(_08392_));
 sg13g2_buf_8 _15125_ (.A(\cpu.ex.io_access ),
    .X(_08393_));
 sg13g2_buf_8 _15126_ (.A(\cpu.ex.genblk3.r_mmu_enable ),
    .X(_08394_));
 sg13g2_nand2b_1 _15127_ (.Y(_08395_),
    .B(net1132),
    .A_N(_08393_));
 sg13g2_buf_2 _15128_ (.A(\cpu.ex.ifetch ),
    .X(_08396_));
 sg13g2_buf_8 _15129_ (.A(\cpu.ex.genblk3.r_mmu_d_proxy ),
    .X(_08397_));
 sg13g2_nor2b_1 _15130_ (.A(_08396_),
    .B_N(_08397_),
    .Y(_08398_));
 sg13g2_nor4_1 _15131_ (.A(_08388_),
    .B(net957),
    .C(_08395_),
    .D(_08398_),
    .Y(_08399_));
 sg13g2_inv_1 _15132_ (.Y(_08400_),
    .A(net1133));
 sg13g2_mux2_1 _15133_ (.A0(\cpu.genblk1.mmu.r_writeable_d[18] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[22] ),
    .S(_08380_),
    .X(_08401_));
 sg13g2_nand3_1 _15134_ (.B(_08385_),
    .C(_08401_),
    .A(_08400_),
    .Y(_08402_));
 sg13g2_and4_1 _15135_ (.A(_08383_),
    .B(_08387_),
    .C(_08399_),
    .D(_08402_),
    .X(_08403_));
 sg13g2_inv_2 _15136_ (.Y(_08404_),
    .A(net1134));
 sg13g2_buf_2 _15137_ (.A(net1074),
    .X(_08405_));
 sg13g2_mux4_1 _15138_ (.S0(_08384_),
    .A0(\cpu.genblk1.mmu.r_writeable_d[24] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[25] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[28] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[29] ),
    .S1(net956),
    .X(_08406_));
 sg13g2_mux4_1 _15139_ (.S0(net1133),
    .A0(\cpu.genblk1.mmu.r_writeable_d[26] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[27] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[30] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[31] ),
    .S1(net1074),
    .X(_08407_));
 sg13g2_and2_1 _15140_ (.A(net1134),
    .B(_08407_),
    .X(_08408_));
 sg13g2_a21oi_1 _15141_ (.A1(_08404_),
    .A2(_08406_),
    .Y(_08409_),
    .B1(_08408_));
 sg13g2_mux4_1 _15142_ (.S0(net1133),
    .A0(\cpu.genblk1.mmu.r_writeable_d[0] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[1] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[4] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[5] ),
    .S1(net1074),
    .X(_08410_));
 sg13g2_nand2_1 _15143_ (.Y(_08411_),
    .A(_08378_),
    .B(_08410_));
 sg13g2_mux2_1 _15144_ (.A0(\cpu.genblk1.mmu.r_writeable_d[3] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[7] ),
    .S(_08381_),
    .X(_08412_));
 sg13g2_nand3_1 _15145_ (.B(_08385_),
    .C(_08412_),
    .A(net1073),
    .Y(_08413_));
 sg13g2_mux2_1 _15146_ (.A0(\cpu.genblk1.mmu.r_writeable_d[2] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[6] ),
    .S(_08380_),
    .X(_08414_));
 sg13g2_nand3_1 _15147_ (.B(_08385_),
    .C(_08414_),
    .A(_08400_),
    .Y(_08415_));
 sg13g2_inv_1 _15148_ (.Y(_08416_),
    .A(_08389_));
 sg13g2_inv_2 _15149_ (.Y(_08417_),
    .A(_08390_));
 sg13g2_inv_1 _15150_ (.Y(_08418_),
    .A(_08388_));
 sg13g2_nand2b_1 _15151_ (.Y(_08419_),
    .B(_08397_),
    .A_N(_08396_));
 sg13g2_a221oi_1 _15152_ (.B2(_08419_),
    .C1(_08395_),
    .B1(_08418_),
    .A1(_08416_),
    .Y(_08420_),
    .A2(_08417_));
 sg13g2_and4_1 _15153_ (.A(_08411_),
    .B(_08413_),
    .C(_08415_),
    .D(_08420_),
    .X(_08421_));
 sg13g2_buf_2 _15154_ (.A(net1134),
    .X(_08422_));
 sg13g2_mux4_1 _15155_ (.S0(_08384_),
    .A0(\cpu.genblk1.mmu.r_writeable_d[8] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[9] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[12] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[13] ),
    .S1(net956),
    .X(_08423_));
 sg13g2_mux4_1 _15156_ (.S0(_08379_),
    .A0(\cpu.genblk1.mmu.r_writeable_d[10] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[11] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[14] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[15] ),
    .S1(_08381_),
    .X(_08424_));
 sg13g2_nand2b_1 _15157_ (.Y(_08425_),
    .B(net1072),
    .A_N(_08424_));
 sg13g2_o21ai_1 _15158_ (.B1(_08425_),
    .Y(_08426_),
    .A1(net1072),
    .A2(_08423_));
 sg13g2_a22oi_1 _15159_ (.Y(_08427_),
    .B1(_08421_),
    .B2(_08426_),
    .A2(_08409_),
    .A1(_08403_));
 sg13g2_inv_4 _15160_ (.A(net1075),
    .Y(_08428_));
 sg13g2_o21ai_1 _15161_ (.B1(_08428_),
    .Y(_08429_),
    .A1(_08403_),
    .A2(_08421_));
 sg13g2_nand2_1 _15162_ (.Y(_08430_),
    .A(_08427_),
    .B(_08429_));
 sg13g2_buf_2 _15163_ (.A(_08430_),
    .X(_08431_));
 sg13g2_buf_1 _15164_ (.A(\cpu.ex.r_read_stall ),
    .X(_08432_));
 sg13g2_nor4_1 _15165_ (.A(_08374_),
    .B(_08432_),
    .C(_08389_),
    .D(_08390_),
    .Y(_08433_));
 sg13g2_buf_2 _15166_ (.A(_08433_),
    .X(_08434_));
 sg13g2_buf_8 _15167_ (.A(\cpu.ex.pc[12] ),
    .X(_08435_));
 sg13g2_nand2b_1 _15168_ (.Y(_08436_),
    .B(_08435_),
    .A_N(\cpu.ex.pc[13] ));
 sg13g2_buf_2 _15169_ (.A(_08436_),
    .X(_08437_));
 sg13g2_buf_8 _15170_ (.A(\cpu.ex.pc[14] ),
    .X(_08438_));
 sg13g2_buf_8 _15171_ (.A(net1131),
    .X(_08439_));
 sg13g2_mux2_1 _15172_ (.A0(\cpu.genblk1.mmu.r_valid_i[9] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[13] ),
    .S(net1071),
    .X(_08440_));
 sg13g2_buf_8 _15173_ (.A(\cpu.ex.pc[13] ),
    .X(_08441_));
 sg13g2_nand2_1 _15174_ (.Y(_08442_),
    .A(_08435_),
    .B(net1130));
 sg13g2_mux2_1 _15175_ (.A0(\cpu.genblk1.mmu.r_valid_i[11] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[15] ),
    .S(net1071),
    .X(_08443_));
 sg13g2_nor2_1 _15176_ (.A(_08442_),
    .B(_08443_),
    .Y(_08444_));
 sg13g2_nand2b_1 _15177_ (.Y(_08445_),
    .B(net1130),
    .A_N(_08435_));
 sg13g2_buf_1 _15178_ (.A(_08445_),
    .X(_08446_));
 sg13g2_mux2_1 _15179_ (.A0(\cpu.genblk1.mmu.r_valid_i[10] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[14] ),
    .S(net1071),
    .X(_08447_));
 sg13g2_nor2_1 _15180_ (.A(_08446_),
    .B(_08447_),
    .Y(_08448_));
 sg13g2_buf_1 _15181_ (.A(_08435_),
    .X(_08449_));
 sg13g2_mux2_1 _15182_ (.A0(\cpu.genblk1.mmu.r_valid_i[8] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[12] ),
    .S(net1071),
    .X(_08450_));
 sg13g2_nor3_1 _15183_ (.A(_08449_),
    .B(net1130),
    .C(_08450_),
    .Y(_08451_));
 sg13g2_buf_8 _15184_ (.A(\cpu.dec.supmode ),
    .X(_08452_));
 sg13g2_buf_2 _15185_ (.A(\cpu.ex.pc[15] ),
    .X(_08453_));
 sg13g2_nand2b_1 _15186_ (.Y(_08454_),
    .B(_08453_),
    .A_N(net1129));
 sg13g2_nor4_1 _15187_ (.A(_08444_),
    .B(_08448_),
    .C(_08451_),
    .D(_08454_),
    .Y(_08455_));
 sg13g2_o21ai_1 _15188_ (.B1(_08455_),
    .Y(_08456_),
    .A1(_08437_),
    .A2(_08440_));
 sg13g2_buf_2 _15189_ (.A(_08396_),
    .X(_08457_));
 sg13g2_nand2_1 _15190_ (.Y(_08458_),
    .A(net1132),
    .B(_08457_));
 sg13g2_mux2_1 _15191_ (.A0(\cpu.genblk1.mmu.r_valid_i[19] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[23] ),
    .S(net1131),
    .X(_08459_));
 sg13g2_nor2_1 _15192_ (.A(_08442_),
    .B(_08459_),
    .Y(_08460_));
 sg13g2_mux2_1 _15193_ (.A0(\cpu.genblk1.mmu.r_valid_i[18] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[22] ),
    .S(net1131),
    .X(_08461_));
 sg13g2_nor2_1 _15194_ (.A(_08446_),
    .B(_08461_),
    .Y(_08462_));
 sg13g2_mux2_1 _15195_ (.A0(\cpu.genblk1.mmu.r_valid_i[16] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[20] ),
    .S(net1131),
    .X(_08463_));
 sg13g2_nor3_1 _15196_ (.A(_08435_),
    .B(net1130),
    .C(_08463_),
    .Y(_08464_));
 sg13g2_mux2_1 _15197_ (.A0(\cpu.genblk1.mmu.r_valid_i[17] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[21] ),
    .S(net1131),
    .X(_08465_));
 sg13g2_nor2b_1 _15198_ (.A(_08453_),
    .B_N(net1129),
    .Y(_08466_));
 sg13g2_o21ai_1 _15199_ (.B1(_08466_),
    .Y(_08467_),
    .A1(_08437_),
    .A2(_08465_));
 sg13g2_nor4_1 _15200_ (.A(_08460_),
    .B(_08462_),
    .C(_08464_),
    .D(_08467_),
    .Y(_08468_));
 sg13g2_mux2_1 _15201_ (.A0(\cpu.genblk1.mmu.r_valid_i[0] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[4] ),
    .S(_08438_),
    .X(_08469_));
 sg13g2_nor3_1 _15202_ (.A(_08435_),
    .B(_08441_),
    .C(_08469_),
    .Y(_08470_));
 sg13g2_mux2_1 _15203_ (.A0(\cpu.genblk1.mmu.r_valid_i[1] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[5] ),
    .S(_08438_),
    .X(_08471_));
 sg13g2_nor2_1 _15204_ (.A(_08437_),
    .B(_08471_),
    .Y(_08472_));
 sg13g2_mux2_1 _15205_ (.A0(\cpu.genblk1.mmu.r_valid_i[3] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[7] ),
    .S(net1071),
    .X(_08473_));
 sg13g2_nor2_1 _15206_ (.A(_08442_),
    .B(_08473_),
    .Y(_08474_));
 sg13g2_mux2_1 _15207_ (.A0(\cpu.genblk1.mmu.r_valid_i[2] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[6] ),
    .S(net1131),
    .X(_08475_));
 sg13g2_nor2_1 _15208_ (.A(_08453_),
    .B(net1129),
    .Y(_08476_));
 sg13g2_o21ai_1 _15209_ (.B1(_08476_),
    .Y(_08477_),
    .A1(_08446_),
    .A2(_08475_));
 sg13g2_nor4_1 _15210_ (.A(_08470_),
    .B(_08472_),
    .C(_08474_),
    .D(_08477_),
    .Y(_08478_));
 sg13g2_mux2_1 _15211_ (.A0(\cpu.genblk1.mmu.r_valid_i[24] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[28] ),
    .S(net1131),
    .X(_08479_));
 sg13g2_nor3_1 _15212_ (.A(_08449_),
    .B(_08441_),
    .C(_08479_),
    .Y(_08480_));
 sg13g2_mux2_1 _15213_ (.A0(\cpu.genblk1.mmu.r_valid_i[25] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[29] ),
    .S(_08439_),
    .X(_08481_));
 sg13g2_nor2_1 _15214_ (.A(_08437_),
    .B(_08481_),
    .Y(_08482_));
 sg13g2_mux2_1 _15215_ (.A0(\cpu.genblk1.mmu.r_valid_i[27] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[31] ),
    .S(_08439_),
    .X(_08483_));
 sg13g2_nor2_1 _15216_ (.A(_08442_),
    .B(_08483_),
    .Y(_08484_));
 sg13g2_mux2_1 _15217_ (.A0(\cpu.genblk1.mmu.r_valid_i[26] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[30] ),
    .S(net1131),
    .X(_08485_));
 sg13g2_and2_1 _15218_ (.A(_08453_),
    .B(net1129),
    .X(_08486_));
 sg13g2_o21ai_1 _15219_ (.B1(_08486_),
    .Y(_08487_),
    .A1(_08446_),
    .A2(_08485_));
 sg13g2_nor4_1 _15220_ (.A(_08480_),
    .B(_08482_),
    .C(_08484_),
    .D(_08487_),
    .Y(_08488_));
 sg13g2_nor4_1 _15221_ (.A(_08458_),
    .B(_08468_),
    .C(_08478_),
    .D(_08488_),
    .Y(_08489_));
 sg13g2_mux4_1 _15222_ (.S0(net1073),
    .A0(\cpu.genblk1.mmu.r_valid_d[18] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[19] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[22] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[23] ),
    .S1(net1074),
    .X(_08490_));
 sg13g2_mux4_1 _15223_ (.S0(net1073),
    .A0(\cpu.genblk1.mmu.r_valid_d[26] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[27] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[30] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[31] ),
    .S1(net956),
    .X(_08491_));
 sg13g2_mux4_1 _15224_ (.S0(net1073),
    .A0(\cpu.genblk1.mmu.r_valid_d[16] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[17] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[20] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[21] ),
    .S1(net1074),
    .X(_08492_));
 sg13g2_mux4_1 _15225_ (.S0(net1073),
    .A0(\cpu.genblk1.mmu.r_valid_d[24] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[25] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[28] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[29] ),
    .S1(net1074),
    .X(_08493_));
 sg13g2_mux4_1 _15226_ (.S0(net1075),
    .A0(_08490_),
    .A1(_08491_),
    .A2(_08492_),
    .A3(_08493_),
    .S1(_08404_),
    .X(_08494_));
 sg13g2_inv_1 _15227_ (.Y(_08495_),
    .A(_08494_));
 sg13g2_nand2_1 _15228_ (.Y(_08496_),
    .A(_08418_),
    .B(_08419_));
 sg13g2_buf_4 _15229_ (.X(_08497_),
    .A(_08496_));
 sg13g2_buf_1 _15230_ (.A(\cpu.ex.mmu_reg_data[0] ),
    .X(_08498_));
 sg13g2_buf_8 _15231_ (.A(\cpu.cond[0] ),
    .X(_08499_));
 sg13g2_buf_1 _15232_ (.A(_00198_),
    .X(_08500_));
 sg13g2_a21oi_1 _15233_ (.A1(_08498_),
    .A2(_08499_),
    .Y(_08501_),
    .B1(_08500_));
 sg13g2_buf_2 _15234_ (.A(_08501_),
    .X(_08502_));
 sg13g2_or2_1 _15235_ (.X(_08503_),
    .B(_08502_),
    .A(_08432_));
 sg13g2_nor2b_2 _15236_ (.A(_08498_),
    .B_N(_08499_),
    .Y(_08504_));
 sg13g2_nand2_1 _15237_ (.Y(_08505_),
    .A(net1132),
    .B(_00197_));
 sg13g2_a21oi_1 _15238_ (.A1(_08500_),
    .A2(_08504_),
    .Y(_08506_),
    .B1(_08505_));
 sg13g2_nor2_1 _15239_ (.A(net957),
    .B(_08395_),
    .Y(_08507_));
 sg13g2_a21oi_1 _15240_ (.A1(_08503_),
    .A2(_08506_),
    .Y(_08508_),
    .B1(_08507_));
 sg13g2_nor2_1 _15241_ (.A(_08497_),
    .B(_08508_),
    .Y(_08509_));
 sg13g2_mux4_1 _15242_ (.S0(net1073),
    .A0(\cpu.genblk1.mmu.r_valid_d[12] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[13] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[14] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[15] ),
    .S1(net1134),
    .X(_08510_));
 sg13g2_and3_1 _15243_ (.X(_08511_),
    .A(net956),
    .B(net1075),
    .C(_08510_));
 sg13g2_inv_1 _15244_ (.Y(_08512_),
    .A(net1074));
 sg13g2_mux4_1 _15245_ (.S0(net1133),
    .A0(\cpu.genblk1.mmu.r_valid_d[8] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[9] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[10] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[11] ),
    .S1(net1134),
    .X(_08513_));
 sg13g2_nand3_1 _15246_ (.B(net1075),
    .C(_08513_),
    .A(_08512_),
    .Y(_08514_));
 sg13g2_nand2_1 _15247_ (.Y(_08515_),
    .A(_08497_),
    .B(_08514_));
 sg13g2_mux4_1 _15248_ (.S0(net1133),
    .A0(\cpu.genblk1.mmu.r_valid_d[4] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[5] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[6] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[7] ),
    .S1(_08375_),
    .X(_08516_));
 sg13g2_nand2_1 _15249_ (.Y(_08517_),
    .A(net956),
    .B(_08516_));
 sg13g2_mux4_1 _15250_ (.S0(net1133),
    .A0(\cpu.genblk1.mmu.r_valid_d[0] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[1] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[2] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[3] ),
    .S1(net1134),
    .X(_08518_));
 sg13g2_nand2_1 _15251_ (.Y(_08519_),
    .A(_08512_),
    .B(_08518_));
 sg13g2_a21oi_1 _15252_ (.A1(_08517_),
    .A2(_08519_),
    .Y(_08520_),
    .B1(net1075));
 sg13g2_nor4_1 _15253_ (.A(_08508_),
    .B(_08511_),
    .C(_08515_),
    .D(_08520_),
    .Y(_08521_));
 sg13g2_a221oi_1 _15254_ (.B2(_08509_),
    .C1(_08521_),
    .B1(_08495_),
    .A1(_08456_),
    .Y(_08522_),
    .A2(_08489_));
 sg13g2_buf_8 _15255_ (.A(_08522_),
    .X(_08523_));
 sg13g2_nor2_1 _15256_ (.A(_08434_),
    .B(net505),
    .Y(_08524_));
 sg13g2_buf_2 _15257_ (.A(_08524_),
    .X(_08525_));
 sg13g2_nor2_1 _15258_ (.A(_08431_),
    .B(_08525_),
    .Y(_08526_));
 sg13g2_buf_1 _15259_ (.A(_08526_),
    .X(_08527_));
 sg13g2_buf_4 _15260_ (.X(_08528_),
    .A(net1070));
 sg13g2_buf_2 _15261_ (.A(_08528_),
    .X(_08529_));
 sg13g2_buf_2 _15262_ (.A(net827),
    .X(_08530_));
 sg13g2_buf_1 _15263_ (.A(net1132),
    .X(_08531_));
 sg13g2_buf_1 _15264_ (.A(net1129),
    .X(_08532_));
 sg13g2_buf_1 _15265_ (.A(_08532_),
    .X(_08533_));
 sg13g2_buf_2 _15266_ (.A(_08528_),
    .X(_08534_));
 sg13g2_buf_2 _15267_ (.A(net826),
    .X(_08535_));
 sg13g2_buf_1 _15268_ (.A(net1130),
    .X(_08536_));
 sg13g2_buf_2 _15269_ (.A(net1066),
    .X(_08537_));
 sg13g2_buf_1 _15270_ (.A(net954),
    .X(_08538_));
 sg13g2_mux4_1 _15271_ (.S0(net718),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][0] ),
    .S1(net825),
    .X(_08539_));
 sg13g2_mux4_1 _15272_ (.S0(net718),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][0] ),
    .S1(net825),
    .X(_08540_));
 sg13g2_mux4_1 _15273_ (.S0(net827),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][0] ),
    .S1(net825),
    .X(_08541_));
 sg13g2_mux4_1 _15274_ (.S0(net718),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][0] ),
    .S1(net825),
    .X(_08542_));
 sg13g2_buf_1 _15275_ (.A(net1071),
    .X(_08543_));
 sg13g2_buf_2 _15276_ (.A(net953),
    .X(_08544_));
 sg13g2_buf_1 _15277_ (.A(_08453_),
    .X(_08545_));
 sg13g2_buf_1 _15278_ (.A(net1065),
    .X(_08546_));
 sg13g2_mux4_1 _15279_ (.S0(net824),
    .A0(_08539_),
    .A1(_08540_),
    .A2(_08541_),
    .A3(_08542_),
    .S1(net952),
    .X(_08547_));
 sg13g2_nand2_1 _15280_ (.Y(_08548_),
    .A(net955),
    .B(_08547_));
 sg13g2_mux4_1 _15281_ (.S0(net718),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][0] ),
    .S1(net825),
    .X(_08549_));
 sg13g2_mux4_1 _15282_ (.S0(_08535_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][0] ),
    .S1(net825),
    .X(_08550_));
 sg13g2_buf_1 _15283_ (.A(net1066),
    .X(_08551_));
 sg13g2_mux4_1 _15284_ (.S0(net827),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][0] ),
    .S1(net951),
    .X(_08552_));
 sg13g2_mux4_1 _15285_ (.S0(net827),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][0] ),
    .S1(_08538_),
    .X(_08553_));
 sg13g2_mux4_1 _15286_ (.S0(net824),
    .A0(_08549_),
    .A1(_08550_),
    .A2(_08552_),
    .A3(_08553_),
    .S1(net952),
    .X(_08554_));
 sg13g2_nand2b_1 _15287_ (.Y(_08555_),
    .B(_08554_),
    .A_N(net1067));
 sg13g2_nand3_1 _15288_ (.B(_08548_),
    .C(_08555_),
    .A(net1068),
    .Y(_08556_));
 sg13g2_o21ai_1 _15289_ (.B1(_08556_),
    .Y(_08557_),
    .A1(net719),
    .A2(net1068));
 sg13g2_buf_2 _15290_ (.A(_08557_),
    .X(_08558_));
 sg13g2_buf_1 _15291_ (.A(_00190_),
    .X(_08559_));
 sg13g2_buf_2 _15292_ (.A(\cpu.ex.pc[3] ),
    .X(_08560_));
 sg13g2_buf_1 _15293_ (.A(\cpu.ex.pc[4] ),
    .X(_08561_));
 sg13g2_inv_2 _15294_ (.Y(_08562_),
    .A(net1127));
 sg13g2_inv_1 _15295_ (.Y(_08563_),
    .A(_08560_));
 sg13g2_buf_2 _15296_ (.A(\cpu.ex.pc[2] ),
    .X(_08564_));
 sg13g2_inv_1 _15297_ (.Y(_08565_),
    .A(net1126));
 sg13g2_buf_1 _15298_ (.A(_08565_),
    .X(_08566_));
 sg13g2_o21ai_1 _15299_ (.B1(net950),
    .Y(_08567_),
    .A1(_08563_),
    .A2(net1127));
 sg13g2_o21ai_1 _15300_ (.B1(_08567_),
    .Y(_08568_),
    .A1(_08560_),
    .A2(_08562_));
 sg13g2_nand2_1 _15301_ (.Y(_08569_),
    .A(net1128),
    .B(_08568_));
 sg13g2_buf_1 _15302_ (.A(_08569_),
    .X(_08570_));
 sg13g2_buf_1 _15303_ (.A(net560),
    .X(_08571_));
 sg13g2_buf_1 _15304_ (.A(net504),
    .X(_08572_));
 sg13g2_buf_1 _15305_ (.A(net453),
    .X(_08573_));
 sg13g2_buf_1 _15306_ (.A(net560),
    .X(_08574_));
 sg13g2_buf_2 _15307_ (.A(net503),
    .X(_08575_));
 sg13g2_nor3_1 _15308_ (.A(net1126),
    .B(_08563_),
    .C(net1127),
    .Y(_08576_));
 sg13g2_buf_2 _15309_ (.A(_08576_),
    .X(_08577_));
 sg13g2_buf_1 _15310_ (.A(_08577_),
    .X(_08578_));
 sg13g2_buf_1 _15311_ (.A(_08578_),
    .X(_08579_));
 sg13g2_buf_1 _15312_ (.A(net641),
    .X(_08580_));
 sg13g2_nor2_1 _15313_ (.A(_08560_),
    .B(net1128),
    .Y(_08581_));
 sg13g2_buf_1 _15314_ (.A(_08581_),
    .X(_08582_));
 sg13g2_and2_1 _15315_ (.A(_08564_),
    .B(net949),
    .X(_08583_));
 sg13g2_buf_2 _15316_ (.A(_08583_),
    .X(_08584_));
 sg13g2_buf_1 _15317_ (.A(_08584_),
    .X(_08585_));
 sg13g2_a22oi_1 _15318_ (.Y(_08586_),
    .B1(net640),
    .B2(\cpu.icache.r_tag[5][12] ),
    .A2(net559),
    .A1(\cpu.icache.r_tag[2][12] ));
 sg13g2_nor3_1 _15319_ (.A(net950),
    .B(_08560_),
    .C(_08561_),
    .Y(_08587_));
 sg13g2_buf_2 _15320_ (.A(_08587_),
    .X(_08588_));
 sg13g2_buf_1 _15321_ (.A(_08588_),
    .X(_08589_));
 sg13g2_buf_1 _15322_ (.A(_08589_),
    .X(_08590_));
 sg13g2_buf_1 _15323_ (.A(net558),
    .X(_08591_));
 sg13g2_buf_1 _15324_ (.A(_08563_),
    .X(_08592_));
 sg13g2_inv_1 _15325_ (.Y(_08593_),
    .A(net1128));
 sg13g2_nor3_1 _15326_ (.A(net950),
    .B(net948),
    .C(_08593_),
    .Y(_08594_));
 sg13g2_buf_2 _15327_ (.A(_08594_),
    .X(_08595_));
 sg13g2_buf_1 _15328_ (.A(_08595_),
    .X(_08596_));
 sg13g2_buf_1 _15329_ (.A(net638),
    .X(_08597_));
 sg13g2_a22oi_1 _15330_ (.Y(_08598_),
    .B1(net557),
    .B2(\cpu.icache.r_tag[3][12] ),
    .A2(_08591_),
    .A1(\cpu.icache.r_tag[1][12] ));
 sg13g2_buf_1 _15331_ (.A(net1128),
    .X(_08599_));
 sg13g2_buf_1 _15332_ (.A(_08599_),
    .X(_08600_));
 sg13g2_buf_1 _15333_ (.A(net947),
    .X(_08601_));
 sg13g2_nor2_1 _15334_ (.A(net950),
    .B(net948),
    .Y(_08602_));
 sg13g2_buf_2 _15335_ (.A(_08602_),
    .X(_08603_));
 sg13g2_buf_1 _15336_ (.A(_08603_),
    .X(_08604_));
 sg13g2_buf_2 _15337_ (.A(_08560_),
    .X(_08605_));
 sg13g2_buf_1 _15338_ (.A(net1063),
    .X(_08606_));
 sg13g2_mux2_1 _15339_ (.A0(\cpu.icache.r_tag[4][12] ),
    .A1(\cpu.icache.r_tag[6][12] ),
    .S(net946),
    .X(_08607_));
 sg13g2_buf_1 _15340_ (.A(net950),
    .X(_08608_));
 sg13g2_a22oi_1 _15341_ (.Y(_08609_),
    .B1(_08607_),
    .B2(net822),
    .A2(net637),
    .A1(\cpu.icache.r_tag[7][12] ));
 sg13g2_or2_1 _15342_ (.X(_08610_),
    .B(_08609_),
    .A(net823));
 sg13g2_nand4_1 _15343_ (.B(_08586_),
    .C(_08598_),
    .A(net452),
    .Y(_08611_),
    .D(_08610_));
 sg13g2_o21ai_1 _15344_ (.B1(_08611_),
    .Y(_08612_),
    .A1(\cpu.icache.r_tag[0][12] ),
    .A2(net416));
 sg13g2_xnor2_1 _15345_ (.Y(_08613_),
    .A(net349),
    .B(_08612_));
 sg13g2_buf_2 _15346_ (.A(_08528_),
    .X(_08614_));
 sg13g2_buf_2 _15347_ (.A(net821),
    .X(_08615_));
 sg13g2_buf_1 _15348_ (.A(net1066),
    .X(_08616_));
 sg13g2_buf_1 _15349_ (.A(net945),
    .X(_08617_));
 sg13g2_mux4_1 _15350_ (.S0(_08615_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][1] ),
    .S1(net820),
    .X(_08618_));
 sg13g2_buf_2 _15351_ (.A(net821),
    .X(_08619_));
 sg13g2_mux4_1 _15352_ (.S0(net715),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][1] ),
    .S1(net820),
    .X(_08620_));
 sg13g2_mux4_1 _15353_ (.S0(_08535_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][1] ),
    .S1(_08538_),
    .X(_08621_));
 sg13g2_buf_1 _15354_ (.A(net945),
    .X(_08622_));
 sg13g2_mux4_1 _15355_ (.S0(net718),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][1] ),
    .S1(_08622_),
    .X(_08623_));
 sg13g2_mux4_1 _15356_ (.S0(net824),
    .A0(_08618_),
    .A1(_08620_),
    .A2(_08621_),
    .A3(_08623_),
    .S1(net952),
    .X(_08624_));
 sg13g2_mux4_1 _15357_ (.S0(net716),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][1] ),
    .S1(net819),
    .X(_08625_));
 sg13g2_mux4_1 _15358_ (.S0(net716),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][1] ),
    .S1(net819),
    .X(_08626_));
 sg13g2_mux4_1 _15359_ (.S0(net718),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][1] ),
    .S1(net825),
    .X(_08627_));
 sg13g2_mux4_1 _15360_ (.S0(net718),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][1] ),
    .S1(net825),
    .X(_08628_));
 sg13g2_mux4_1 _15361_ (.S0(net824),
    .A0(_08625_),
    .A1(_08626_),
    .A2(_08627_),
    .A3(_08628_),
    .S1(net952),
    .X(_08629_));
 sg13g2_mux2_1 _15362_ (.A0(_08624_),
    .A1(_08629_),
    .S(net1067),
    .X(_08630_));
 sg13g2_inv_1 _15363_ (.Y(_08631_),
    .A(net951));
 sg13g2_nor2_1 _15364_ (.A(_08631_),
    .B(net1068),
    .Y(_08632_));
 sg13g2_a21oi_1 _15365_ (.A1(net1068),
    .A2(_08630_),
    .Y(_08633_),
    .B1(_08632_));
 sg13g2_buf_2 _15366_ (.A(_08633_),
    .X(_08634_));
 sg13g2_a22oi_1 _15367_ (.Y(_08635_),
    .B1(net640),
    .B2(\cpu.icache.r_tag[5][13] ),
    .A2(net559),
    .A1(\cpu.icache.r_tag[2][13] ));
 sg13g2_a22oi_1 _15368_ (.Y(_08636_),
    .B1(net557),
    .B2(\cpu.icache.r_tag[3][13] ),
    .A2(net502),
    .A1(\cpu.icache.r_tag[1][13] ));
 sg13g2_mux2_1 _15369_ (.A0(\cpu.icache.r_tag[4][13] ),
    .A1(\cpu.icache.r_tag[6][13] ),
    .S(net946),
    .X(_08637_));
 sg13g2_a22oi_1 _15370_ (.Y(_08638_),
    .B1(_08637_),
    .B2(net822),
    .A2(net637),
    .A1(\cpu.icache.r_tag[7][13] ));
 sg13g2_or2_1 _15371_ (.X(_08639_),
    .B(_08638_),
    .A(net823));
 sg13g2_nand4_1 _15372_ (.B(_08635_),
    .C(_08636_),
    .A(net452),
    .Y(_08640_),
    .D(_08639_));
 sg13g2_o21ai_1 _15373_ (.B1(_08640_),
    .Y(_08641_),
    .A1(\cpu.icache.r_tag[0][13] ),
    .A2(net416));
 sg13g2_xnor2_1 _15374_ (.Y(_08642_),
    .A(net415),
    .B(_08641_));
 sg13g2_nand2_1 _15375_ (.Y(_08643_),
    .A(_08613_),
    .B(_08642_));
 sg13g2_buf_2 _15376_ (.A(_00192_),
    .X(_08644_));
 sg13g2_buf_1 _15377_ (.A(_08644_),
    .X(_08645_));
 sg13g2_mux4_1 _15378_ (.S0(net827),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][4] ),
    .S1(net951),
    .X(_08646_));
 sg13g2_mux4_1 _15379_ (.S0(net827),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][4] ),
    .S1(_08551_),
    .X(_08647_));
 sg13g2_buf_2 _15380_ (.A(_08528_),
    .X(_08648_));
 sg13g2_buf_2 _15381_ (.A(net1066),
    .X(_08649_));
 sg13g2_mux4_1 _15382_ (.S0(net818),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][4] ),
    .S1(net944),
    .X(_08650_));
 sg13g2_mux4_1 _15383_ (.S0(net818),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][4] ),
    .S1(net944),
    .X(_08651_));
 sg13g2_mux4_1 _15384_ (.S0(net953),
    .A0(_08646_),
    .A1(_08647_),
    .A2(_08650_),
    .A3(_08651_),
    .S1(net1065),
    .X(_08652_));
 sg13g2_mux4_1 _15385_ (.S0(net818),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][4] ),
    .S1(net951),
    .X(_08653_));
 sg13g2_mux4_1 _15386_ (.S0(net818),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][4] ),
    .S1(net951),
    .X(_08654_));
 sg13g2_mux4_1 _15387_ (.S0(net818),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][4] ),
    .S1(net944),
    .X(_08655_));
 sg13g2_mux4_1 _15388_ (.S0(net818),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][4] ),
    .S1(net944),
    .X(_08656_));
 sg13g2_mux4_1 _15389_ (.S0(net953),
    .A0(_08653_),
    .A1(_08654_),
    .A2(_08655_),
    .A3(_08656_),
    .S1(net1065),
    .X(_08657_));
 sg13g2_mux2_1 _15390_ (.A0(_08652_),
    .A1(_08657_),
    .S(net1067),
    .X(_08658_));
 sg13g2_nand2b_1 _15391_ (.Y(_08659_),
    .B(_08658_),
    .A_N(net1062));
 sg13g2_buf_2 _15392_ (.A(_08659_),
    .X(_08660_));
 sg13g2_buf_1 _15393_ (.A(net560),
    .X(_08661_));
 sg13g2_buf_1 _15394_ (.A(net717),
    .X(_08662_));
 sg13g2_a22oi_1 _15395_ (.Y(_08663_),
    .B1(net558),
    .B2(\cpu.icache.r_tag[1][16] ),
    .A2(net636),
    .A1(\cpu.icache.r_tag[2][16] ));
 sg13g2_nor3_1 _15396_ (.A(net1126),
    .B(net948),
    .C(net1128),
    .Y(_08664_));
 sg13g2_buf_1 _15397_ (.A(_08664_),
    .X(_08665_));
 sg13g2_buf_1 _15398_ (.A(_08665_),
    .X(_08666_));
 sg13g2_buf_2 _15399_ (.A(net635),
    .X(_08667_));
 sg13g2_a22oi_1 _15400_ (.Y(_08668_),
    .B1(net556),
    .B2(\cpu.icache.r_tag[6][16] ),
    .A2(net557),
    .A1(\cpu.icache.r_tag[3][16] ));
 sg13g2_buf_1 _15401_ (.A(net1126),
    .X(_08669_));
 sg13g2_buf_2 _15402_ (.A(_08669_),
    .X(_08670_));
 sg13g2_buf_1 _15403_ (.A(net1063),
    .X(_08671_));
 sg13g2_mux2_1 _15404_ (.A0(\cpu.icache.r_tag[5][16] ),
    .A1(\cpu.icache.r_tag[7][16] ),
    .S(net942),
    .X(_08672_));
 sg13g2_nor2_2 _15405_ (.A(net1061),
    .B(_08671_),
    .Y(_08673_));
 sg13g2_a22oi_1 _15406_ (.Y(_08674_),
    .B1(_08673_),
    .B2(\cpu.icache.r_tag[4][16] ),
    .A2(_08672_),
    .A1(net943));
 sg13g2_or2_1 _15407_ (.X(_08675_),
    .B(_08674_),
    .A(net947));
 sg13g2_nand4_1 _15408_ (.B(_08663_),
    .C(_08668_),
    .A(net501),
    .Y(_08676_),
    .D(_08675_));
 sg13g2_o21ai_1 _15409_ (.B1(_08676_),
    .Y(_08677_),
    .A1(\cpu.icache.r_tag[0][16] ),
    .A2(net452));
 sg13g2_xnor2_1 _15410_ (.Y(_08678_),
    .A(_08660_),
    .B(_08677_));
 sg13g2_buf_1 _15411_ (.A(_08545_),
    .X(_08679_));
 sg13g2_mux4_1 _15412_ (.S0(_08648_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][3] ),
    .S1(_08649_),
    .X(_08680_));
 sg13g2_mux4_1 _15413_ (.S0(_08648_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][3] ),
    .S1(_08649_),
    .X(_08681_));
 sg13g2_mux4_1 _15414_ (.S0(net818),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][3] ),
    .S1(net944),
    .X(_08682_));
 sg13g2_mux4_1 _15415_ (.S0(net818),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][3] ),
    .S1(net944),
    .X(_08683_));
 sg13g2_mux4_1 _15416_ (.S0(_08543_),
    .A0(_08680_),
    .A1(_08681_),
    .A2(_08682_),
    .A3(_08683_),
    .S1(net1129),
    .X(_08684_));
 sg13g2_nand2b_1 _15417_ (.Y(_08685_),
    .B(net1068),
    .A_N(_08684_));
 sg13g2_buf_2 _15418_ (.A(net821),
    .X(_08686_));
 sg13g2_buf_1 _15419_ (.A(net944),
    .X(_08687_));
 sg13g2_mux4_1 _15420_ (.S0(net714),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][3] ),
    .S1(net817),
    .X(_08688_));
 sg13g2_buf_1 _15421_ (.A(net944),
    .X(_08689_));
 sg13g2_mux4_1 _15422_ (.S0(net714),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][3] ),
    .S1(net816),
    .X(_08690_));
 sg13g2_mux4_1 _15423_ (.S0(net714),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][3] ),
    .S1(net817),
    .X(_08691_));
 sg13g2_mux4_1 _15424_ (.S0(net714),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][3] ),
    .S1(net817),
    .X(_08692_));
 sg13g2_buf_2 _15425_ (.A(net953),
    .X(_08693_));
 sg13g2_mux4_1 _15426_ (.S0(net815),
    .A0(_08688_),
    .A1(_08690_),
    .A2(_08691_),
    .A3(_08692_),
    .S1(net1067),
    .X(_08694_));
 sg13g2_inv_1 _15427_ (.Y(_08695_),
    .A(net1132));
 sg13g2_nor2_1 _15428_ (.A(net941),
    .B(_08695_),
    .Y(_08696_));
 sg13g2_a22oi_1 _15429_ (.Y(_08697_),
    .B1(_08694_),
    .B2(_08696_),
    .A2(_08685_),
    .A1(net941));
 sg13g2_buf_2 _15430_ (.A(_08697_),
    .X(_08698_));
 sg13g2_nor3_1 _15431_ (.A(net950),
    .B(net948),
    .C(_08559_),
    .Y(_08699_));
 sg13g2_buf_2 _15432_ (.A(_08699_),
    .X(_08700_));
 sg13g2_and2_1 _15433_ (.A(\cpu.icache.r_tag[5][15] ),
    .B(_08584_),
    .X(_08701_));
 sg13g2_a221oi_1 _15434_ (.B2(\cpu.icache.r_tag[7][15] ),
    .C1(_08701_),
    .B1(_08700_),
    .A1(\cpu.icache.r_tag[2][15] ),
    .Y(_08702_),
    .A2(net641));
 sg13g2_buf_1 _15435_ (.A(net639),
    .X(_08703_));
 sg13g2_nor3_1 _15436_ (.A(net1126),
    .B(_08560_),
    .C(net1128),
    .Y(_08704_));
 sg13g2_buf_2 _15437_ (.A(_08704_),
    .X(_08705_));
 sg13g2_buf_1 _15438_ (.A(_08705_),
    .X(_08706_));
 sg13g2_a22oi_1 _15439_ (.Y(_08707_),
    .B1(net814),
    .B2(\cpu.icache.r_tag[4][15] ),
    .A2(net555),
    .A1(\cpu.icache.r_tag[1][15] ));
 sg13g2_buf_1 _15440_ (.A(net638),
    .X(_08708_));
 sg13g2_a22oi_1 _15441_ (.Y(_08709_),
    .B1(net556),
    .B2(\cpu.icache.r_tag[6][15] ),
    .A2(net554),
    .A1(\cpu.icache.r_tag[3][15] ));
 sg13g2_nand4_1 _15442_ (.B(_08702_),
    .C(_08707_),
    .A(net501),
    .Y(_08710_),
    .D(_08709_));
 sg13g2_o21ai_1 _15443_ (.B1(_08710_),
    .Y(_08711_),
    .A1(\cpu.icache.r_tag[0][15] ),
    .A2(net453));
 sg13g2_xnor2_1 _15444_ (.Y(_08712_),
    .A(net450),
    .B(_08711_));
 sg13g2_and2_1 _15445_ (.A(_08678_),
    .B(_08712_),
    .X(_08713_));
 sg13g2_buf_2 _15446_ (.A(net821),
    .X(_08714_));
 sg13g2_buf_1 _15447_ (.A(net945),
    .X(_08715_));
 sg13g2_mux4_1 _15448_ (.S0(net713),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][6] ),
    .S1(net813),
    .X(_08716_));
 sg13g2_mux4_1 _15449_ (.S0(net713),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][6] ),
    .S1(net813),
    .X(_08717_));
 sg13g2_mux4_1 _15450_ (.S0(net716),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][6] ),
    .S1(net819),
    .X(_08718_));
 sg13g2_mux4_1 _15451_ (.S0(net716),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][6] ),
    .S1(net820),
    .X(_08719_));
 sg13g2_mux4_1 _15452_ (.S0(net824),
    .A0(_08716_),
    .A1(_08717_),
    .A2(_08718_),
    .A3(_08719_),
    .S1(_08546_),
    .X(_08720_));
 sg13g2_mux4_1 _15453_ (.S0(net715),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][6] ),
    .S1(net820),
    .X(_08721_));
 sg13g2_mux4_1 _15454_ (.S0(net713),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][6] ),
    .S1(net813),
    .X(_08722_));
 sg13g2_mux4_1 _15455_ (.S0(net716),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][6] ),
    .S1(net819),
    .X(_08723_));
 sg13g2_mux4_1 _15456_ (.S0(net716),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][6] ),
    .S1(net819),
    .X(_08724_));
 sg13g2_mux4_1 _15457_ (.S0(_08544_),
    .A0(_08721_),
    .A1(_08722_),
    .A2(_08723_),
    .A3(_08724_),
    .S1(net952),
    .X(_08725_));
 sg13g2_mux2_1 _15458_ (.A0(_08720_),
    .A1(_08725_),
    .S(net955),
    .X(_08726_));
 sg13g2_nand2b_1 _15459_ (.Y(_08727_),
    .B(_08726_),
    .A_N(net1062));
 sg13g2_buf_2 _15460_ (.A(_08727_),
    .X(_08728_));
 sg13g2_a22oi_1 _15461_ (.Y(_08729_),
    .B1(net558),
    .B2(\cpu.icache.r_tag[1][18] ),
    .A2(net636),
    .A1(\cpu.icache.r_tag[2][18] ));
 sg13g2_a22oi_1 _15462_ (.Y(_08730_),
    .B1(net556),
    .B2(\cpu.icache.r_tag[6][18] ),
    .A2(_08597_),
    .A1(\cpu.icache.r_tag[3][18] ));
 sg13g2_mux2_1 _15463_ (.A0(\cpu.icache.r_tag[5][18] ),
    .A1(\cpu.icache.r_tag[7][18] ),
    .S(net946),
    .X(_08731_));
 sg13g2_buf_2 _15464_ (.A(net943),
    .X(_08732_));
 sg13g2_a22oi_1 _15465_ (.Y(_08733_),
    .B1(_08731_),
    .B2(_08732_),
    .A2(_08673_),
    .A1(\cpu.icache.r_tag[4][18] ));
 sg13g2_or2_1 _15466_ (.X(_08734_),
    .B(_08733_),
    .A(net823));
 sg13g2_nand4_1 _15467_ (.B(_08729_),
    .C(_08730_),
    .A(net452),
    .Y(_08735_),
    .D(_08734_));
 sg13g2_o21ai_1 _15468_ (.B1(_08735_),
    .Y(_08736_),
    .A1(\cpu.icache.r_tag[0][18] ),
    .A2(net416));
 sg13g2_xnor2_1 _15469_ (.Y(_08737_),
    .A(net414),
    .B(_08736_));
 sg13g2_buf_2 _15470_ (.A(\cpu.ex.pc[9] ),
    .X(_08738_));
 sg13g2_mux2_1 _15471_ (.A0(\cpu.icache.r_tag[7][9] ),
    .A1(\cpu.icache.r_tag[3][9] ),
    .S(net1064),
    .X(_08739_));
 sg13g2_a22oi_1 _15472_ (.Y(_08740_),
    .B1(_08603_),
    .B2(_08739_),
    .A2(net717),
    .A1(\cpu.icache.r_tag[2][9] ));
 sg13g2_a22oi_1 _15473_ (.Y(_08741_),
    .B1(_08665_),
    .B2(\cpu.icache.r_tag[6][9] ),
    .A2(_08584_),
    .A1(\cpu.icache.r_tag[5][9] ));
 sg13g2_a22oi_1 _15474_ (.Y(_08742_),
    .B1(_08705_),
    .B2(\cpu.icache.r_tag[4][9] ),
    .A2(net639),
    .A1(\cpu.icache.r_tag[1][9] ));
 sg13g2_nand4_1 _15475_ (.B(_08740_),
    .C(_08741_),
    .A(net504),
    .Y(_08743_),
    .D(_08742_));
 sg13g2_o21ai_1 _15476_ (.B1(_08743_),
    .Y(_08744_),
    .A1(\cpu.icache.r_tag[0][9] ),
    .A2(net503));
 sg13g2_xnor2_1 _15477_ (.Y(_08745_),
    .A(_08738_),
    .B(_08744_));
 sg13g2_buf_2 _15478_ (.A(\cpu.ex.pc[11] ),
    .X(_08746_));
 sg13g2_buf_1 _15479_ (.A(net639),
    .X(_08747_));
 sg13g2_a22oi_1 _15480_ (.Y(_08748_),
    .B1(net553),
    .B2(\cpu.icache.r_tag[1][11] ),
    .A2(_08584_),
    .A1(\cpu.icache.r_tag[5][11] ));
 sg13g2_a22oi_1 _15481_ (.Y(_08749_),
    .B1(net638),
    .B2(\cpu.icache.r_tag[3][11] ),
    .A2(_08578_),
    .A1(\cpu.icache.r_tag[2][11] ));
 sg13g2_mux2_1 _15482_ (.A0(\cpu.icache.r_tag[4][11] ),
    .A1(\cpu.icache.r_tag[6][11] ),
    .S(net1063),
    .X(_08750_));
 sg13g2_a22oi_1 _15483_ (.Y(_08751_),
    .B1(_08750_),
    .B2(_08566_),
    .A2(_08603_),
    .A1(\cpu.icache.r_tag[7][11] ));
 sg13g2_or2_1 _15484_ (.X(_08752_),
    .B(_08751_),
    .A(net947));
 sg13g2_nand4_1 _15485_ (.B(_08748_),
    .C(_08749_),
    .A(net504),
    .Y(_08753_),
    .D(_08752_));
 sg13g2_o21ai_1 _15486_ (.B1(_08753_),
    .Y(_08754_),
    .A1(\cpu.icache.r_tag[0][11] ),
    .A2(net503));
 sg13g2_xnor2_1 _15487_ (.Y(_08755_),
    .A(_08746_),
    .B(_08754_));
 sg13g2_nor2_1 _15488_ (.A(_08745_),
    .B(_08755_),
    .Y(_08756_));
 sg13g2_buf_1 _15489_ (.A(\cpu.ex.pc[8] ),
    .X(_08757_));
 sg13g2_inv_1 _15490_ (.Y(_08758_),
    .A(_08757_));
 sg13g2_buf_1 _15491_ (.A(_08758_),
    .X(_08759_));
 sg13g2_mux2_1 _15492_ (.A0(\cpu.icache.r_tag[7][8] ),
    .A1(\cpu.icache.r_tag[3][8] ),
    .S(net1064),
    .X(_08760_));
 sg13g2_a22oi_1 _15493_ (.Y(_08761_),
    .B1(net637),
    .B2(_08760_),
    .A2(net641),
    .A1(\cpu.icache.r_tag[2][8] ));
 sg13g2_buf_1 _15494_ (.A(_08705_),
    .X(_08762_));
 sg13g2_a22oi_1 _15495_ (.Y(_08763_),
    .B1(net811),
    .B2(\cpu.icache.r_tag[4][8] ),
    .A2(net635),
    .A1(\cpu.icache.r_tag[6][8] ));
 sg13g2_a22oi_1 _15496_ (.Y(_08764_),
    .B1(net555),
    .B2(\cpu.icache.r_tag[1][8] ),
    .A2(net640),
    .A1(\cpu.icache.r_tag[5][8] ));
 sg13g2_nand4_1 _15497_ (.B(_08761_),
    .C(_08763_),
    .A(net503),
    .Y(_08765_),
    .D(_08764_));
 sg13g2_o21ai_1 _15498_ (.B1(_08765_),
    .Y(_08766_),
    .A1(\cpu.icache.r_tag[0][8] ),
    .A2(net453));
 sg13g2_xnor2_1 _15499_ (.Y(_08767_),
    .A(net940),
    .B(_08766_));
 sg13g2_inv_1 _15500_ (.Y(_08768_),
    .A(\cpu.ex.pc[6] ));
 sg13g2_a22oi_1 _15501_ (.Y(_08769_),
    .B1(net811),
    .B2(\cpu.icache.r_tag[4][6] ),
    .A2(net555),
    .A1(\cpu.icache.r_tag[1][6] ));
 sg13g2_a22oi_1 _15502_ (.Y(_08770_),
    .B1(net635),
    .B2(\cpu.icache.r_tag[6][6] ),
    .A2(net640),
    .A1(\cpu.icache.r_tag[5][6] ));
 sg13g2_mux2_1 _15503_ (.A0(\cpu.icache.r_tag[7][6] ),
    .A1(\cpu.icache.r_tag[3][6] ),
    .S(net1064),
    .X(_08771_));
 sg13g2_a22oi_1 _15504_ (.Y(_08772_),
    .B1(net637),
    .B2(_08771_),
    .A2(net641),
    .A1(\cpu.icache.r_tag[2][6] ));
 sg13g2_nand4_1 _15505_ (.B(_08769_),
    .C(_08770_),
    .A(net503),
    .Y(_08773_),
    .D(_08772_));
 sg13g2_o21ai_1 _15506_ (.B1(_08773_),
    .Y(_08774_),
    .A1(\cpu.icache.r_tag[0][6] ),
    .A2(net453));
 sg13g2_xnor2_1 _15507_ (.Y(_08775_),
    .A(_08768_),
    .B(_08774_));
 sg13g2_and3_1 _15508_ (.X(_08776_),
    .A(_08756_),
    .B(_08767_),
    .C(_08775_));
 sg13g2_buf_1 _15509_ (.A(\cpu.ex.pc[7] ),
    .X(_08777_));
 sg13g2_inv_1 _15510_ (.Y(_08778_),
    .A(_08777_));
 sg13g2_buf_1 _15511_ (.A(_08778_),
    .X(_08779_));
 sg13g2_buf_1 _15512_ (.A(net717),
    .X(_08780_));
 sg13g2_a22oi_1 _15513_ (.Y(_08781_),
    .B1(_08703_),
    .B2(\cpu.icache.r_tag[1][7] ),
    .A2(net634),
    .A1(\cpu.icache.r_tag[2][7] ));
 sg13g2_a22oi_1 _15514_ (.Y(_08782_),
    .B1(net811),
    .B2(\cpu.icache.r_tag[4][7] ),
    .A2(_08708_),
    .A1(\cpu.icache.r_tag[3][7] ));
 sg13g2_nor2_1 _15515_ (.A(net1126),
    .B(net948),
    .Y(_08783_));
 sg13g2_buf_2 _15516_ (.A(_08783_),
    .X(_08784_));
 sg13g2_mux2_1 _15517_ (.A0(\cpu.icache.r_tag[5][7] ),
    .A1(\cpu.icache.r_tag[7][7] ),
    .S(net1063),
    .X(_08785_));
 sg13g2_a22oi_1 _15518_ (.Y(_08786_),
    .B1(_08785_),
    .B2(net943),
    .A2(_08784_),
    .A1(\cpu.icache.r_tag[6][7] ));
 sg13g2_or2_1 _15519_ (.X(_08787_),
    .B(_08786_),
    .A(net947));
 sg13g2_nand4_1 _15520_ (.B(_08781_),
    .C(_08782_),
    .A(_08574_),
    .Y(_08788_),
    .D(_08787_));
 sg13g2_o21ai_1 _15521_ (.B1(_08788_),
    .Y(_08789_),
    .A1(\cpu.icache.r_tag[0][7] ),
    .A2(net453));
 sg13g2_xnor2_1 _15522_ (.Y(_08790_),
    .A(net939),
    .B(_08789_));
 sg13g2_buf_1 _15523_ (.A(\cpu.ex.pc[10] ),
    .X(_08791_));
 sg13g2_a22oi_1 _15524_ (.Y(_08792_),
    .B1(net553),
    .B2(\cpu.icache.r_tag[1][10] ),
    .A2(net634),
    .A1(\cpu.icache.r_tag[2][10] ));
 sg13g2_a22oi_1 _15525_ (.Y(_08793_),
    .B1(net811),
    .B2(\cpu.icache.r_tag[4][10] ),
    .A2(_08596_),
    .A1(\cpu.icache.r_tag[3][10] ));
 sg13g2_mux2_1 _15526_ (.A0(\cpu.icache.r_tag[5][10] ),
    .A1(\cpu.icache.r_tag[7][10] ),
    .S(_08605_),
    .X(_08794_));
 sg13g2_a22oi_1 _15527_ (.Y(_08795_),
    .B1(_08794_),
    .B2(net943),
    .A2(_08784_),
    .A1(\cpu.icache.r_tag[6][10] ));
 sg13g2_or2_1 _15528_ (.X(_08796_),
    .B(_08795_),
    .A(_08600_));
 sg13g2_nand4_1 _15529_ (.B(_08792_),
    .C(_08793_),
    .A(net504),
    .Y(_08797_),
    .D(_08796_));
 sg13g2_o21ai_1 _15530_ (.B1(_08797_),
    .Y(_08798_),
    .A1(\cpu.icache.r_tag[0][10] ),
    .A2(net453));
 sg13g2_xor2_1 _15531_ (.B(_08798_),
    .A(_08791_),
    .X(_08799_));
 sg13g2_buf_1 _15532_ (.A(net812),
    .X(_08800_));
 sg13g2_buf_2 _15533_ (.A(net942),
    .X(_08801_));
 sg13g2_buf_1 _15534_ (.A(net810),
    .X(_08802_));
 sg13g2_mux4_1 _15535_ (.S0(net712),
    .A0(\cpu.icache.r_valid[4] ),
    .A1(\cpu.icache.r_valid[5] ),
    .A2(\cpu.icache.r_valid[6] ),
    .A3(\cpu.icache.r_valid[7] ),
    .S1(net711),
    .X(_08803_));
 sg13g2_mux4_1 _15536_ (.S0(net712),
    .A0(\cpu.icache.r_valid[0] ),
    .A1(\cpu.icache.r_valid[1] ),
    .A2(\cpu.icache.r_valid[2] ),
    .A3(\cpu.icache.r_valid[3] ),
    .S1(net711),
    .X(_08804_));
 sg13g2_mux2_1 _15537_ (.A0(_08803_),
    .A1(_08804_),
    .S(_08562_),
    .X(_08805_));
 sg13g2_buf_1 _15538_ (.A(\cpu.ex.pc[5] ),
    .X(_08806_));
 sg13g2_inv_1 _15539_ (.Y(_08807_),
    .A(_08806_));
 sg13g2_buf_1 _15540_ (.A(_08807_),
    .X(_08808_));
 sg13g2_a22oi_1 _15541_ (.Y(_08809_),
    .B1(net553),
    .B2(\cpu.icache.r_tag[1][5] ),
    .A2(net640),
    .A1(\cpu.icache.r_tag[5][5] ));
 sg13g2_a22oi_1 _15542_ (.Y(_08810_),
    .B1(net811),
    .B2(\cpu.icache.r_tag[4][5] ),
    .A2(_08780_),
    .A1(\cpu.icache.r_tag[2][5] ));
 sg13g2_mux2_1 _15543_ (.A0(\cpu.icache.r_tag[7][5] ),
    .A1(\cpu.icache.r_tag[3][5] ),
    .S(_08599_),
    .X(_08811_));
 sg13g2_nor2_1 _15544_ (.A(net1126),
    .B(net1064),
    .Y(_08812_));
 sg13g2_a22oi_1 _15545_ (.Y(_08813_),
    .B1(_08812_),
    .B2(\cpu.icache.r_tag[6][5] ),
    .A2(_08811_),
    .A1(net943));
 sg13g2_nand2b_1 _15546_ (.Y(_08814_),
    .B(net810),
    .A_N(_08813_));
 sg13g2_nand4_1 _15547_ (.B(_08809_),
    .C(_08810_),
    .A(_08571_),
    .Y(_08815_),
    .D(_08814_));
 sg13g2_o21ai_1 _15548_ (.B1(_08815_),
    .Y(_08816_),
    .A1(\cpu.icache.r_tag[0][5] ),
    .A2(net501));
 sg13g2_xnor2_1 _15549_ (.Y(_08817_),
    .A(net938),
    .B(_08816_));
 sg13g2_and4_1 _15550_ (.A(_08790_),
    .B(_08799_),
    .C(_08805_),
    .D(_08817_),
    .X(_08818_));
 sg13g2_nand4_1 _15551_ (.B(_08737_),
    .C(_08776_),
    .A(_08713_),
    .Y(_08819_),
    .D(_08818_));
 sg13g2_mux4_1 _15552_ (.S0(_08529_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][2] ),
    .S1(_08551_),
    .X(_08820_));
 sg13g2_mux4_1 _15553_ (.S0(_08529_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][2] ),
    .S1(net951),
    .X(_08821_));
 sg13g2_mux4_1 _15554_ (.S0(net827),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][2] ),
    .S1(net951),
    .X(_08822_));
 sg13g2_mux4_1 _15555_ (.S0(net827),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][2] ),
    .S1(net951),
    .X(_08823_));
 sg13g2_mux4_1 _15556_ (.S0(net1065),
    .A0(_08820_),
    .A1(_08821_),
    .A2(_08822_),
    .A3(_08823_),
    .S1(net1067),
    .X(_08824_));
 sg13g2_nand2b_1 _15557_ (.Y(_08825_),
    .B(net1068),
    .A_N(_08824_));
 sg13g2_mux4_1 _15558_ (.S0(net719),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][2] ),
    .S1(net816),
    .X(_08826_));
 sg13g2_mux4_1 _15559_ (.S0(net719),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][2] ),
    .S1(net816),
    .X(_08827_));
 sg13g2_mux4_1 _15560_ (.S0(net714),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][2] ),
    .S1(net816),
    .X(_08828_));
 sg13g2_mux4_1 _15561_ (.S0(net719),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][2] ),
    .S1(net816),
    .X(_08829_));
 sg13g2_mux4_1 _15562_ (.S0(net952),
    .A0(_08826_),
    .A1(_08827_),
    .A2(_08828_),
    .A3(_08829_),
    .S1(net1067),
    .X(_08830_));
 sg13g2_nor2_1 _15563_ (.A(net815),
    .B(_08695_),
    .Y(_08831_));
 sg13g2_a22oi_1 _15564_ (.Y(_08832_),
    .B1(_08830_),
    .B2(_08831_),
    .A2(_08825_),
    .A1(net815));
 sg13g2_buf_1 _15565_ (.A(_08832_),
    .X(_08833_));
 sg13g2_a22oi_1 _15566_ (.Y(_08834_),
    .B1(net635),
    .B2(\cpu.icache.r_tag[6][14] ),
    .A2(_08579_),
    .A1(\cpu.icache.r_tag[2][14] ));
 sg13g2_a22oi_1 _15567_ (.Y(_08835_),
    .B1(_08708_),
    .B2(\cpu.icache.r_tag[3][14] ),
    .A2(_08747_),
    .A1(\cpu.icache.r_tag[1][14] ));
 sg13g2_mux2_1 _15568_ (.A0(\cpu.icache.r_tag[5][14] ),
    .A1(\cpu.icache.r_tag[7][14] ),
    .S(_08605_),
    .X(_08836_));
 sg13g2_a22oi_1 _15569_ (.Y(_08837_),
    .B1(_08836_),
    .B2(net943),
    .A2(_08673_),
    .A1(\cpu.icache.r_tag[4][14] ));
 sg13g2_or2_1 _15570_ (.X(_08838_),
    .B(_08837_),
    .A(_08600_));
 sg13g2_nand3_1 _15571_ (.B(_08835_),
    .C(_08838_),
    .A(_08834_),
    .Y(_08839_));
 sg13g2_mux2_1 _15572_ (.A0(\cpu.icache.r_tag[0][14] ),
    .A1(_08839_),
    .S(net453),
    .X(_08840_));
 sg13g2_xnor2_1 _15573_ (.Y(_08841_),
    .A(_08833_),
    .B(_08840_));
 sg13g2_mux4_1 _15574_ (.S0(net821),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][10] ),
    .S1(net945),
    .X(_08842_));
 sg13g2_mux4_1 _15575_ (.S0(net821),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][10] ),
    .S1(net945),
    .X(_08843_));
 sg13g2_mux4_1 _15576_ (.S0(net826),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][10] ),
    .S1(_08616_),
    .X(_08844_));
 sg13g2_mux4_1 _15577_ (.S0(_08614_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][10] ),
    .S1(_08616_),
    .X(_08845_));
 sg13g2_mux4_1 _15578_ (.S0(net953),
    .A0(_08842_),
    .A1(_08843_),
    .A2(_08844_),
    .A3(_08845_),
    .S1(net1065),
    .X(_08846_));
 sg13g2_mux4_1 _15579_ (.S0(net821),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][10] ),
    .S1(net945),
    .X(_08847_));
 sg13g2_mux4_1 _15580_ (.S0(net821),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][10] ),
    .S1(net945),
    .X(_08848_));
 sg13g2_mux4_1 _15581_ (.S0(net826),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][10] ),
    .S1(net954),
    .X(_08849_));
 sg13g2_mux4_1 _15582_ (.S0(net826),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][10] ),
    .S1(net945),
    .X(_08850_));
 sg13g2_mux4_1 _15583_ (.S0(net953),
    .A0(_08847_),
    .A1(_08848_),
    .A2(_08849_),
    .A3(_08850_),
    .S1(net1065),
    .X(_08851_));
 sg13g2_mux2_1 _15584_ (.A0(_08846_),
    .A1(_08851_),
    .S(net1067),
    .X(_08852_));
 sg13g2_nand2b_1 _15585_ (.Y(_08853_),
    .B(_08852_),
    .A_N(net1062));
 sg13g2_buf_1 _15586_ (.A(_08853_),
    .X(_08854_));
 sg13g2_a22oi_1 _15587_ (.Y(_08855_),
    .B1(_08762_),
    .B2(\cpu.icache.r_tag[4][22] ),
    .A2(_08703_),
    .A1(\cpu.icache.r_tag[1][22] ));
 sg13g2_a22oi_1 _15588_ (.Y(_08856_),
    .B1(net635),
    .B2(\cpu.icache.r_tag[6][22] ),
    .A2(_08585_),
    .A1(\cpu.icache.r_tag[5][22] ));
 sg13g2_mux2_1 _15589_ (.A0(\cpu.icache.r_tag[7][22] ),
    .A1(\cpu.icache.r_tag[3][22] ),
    .S(net1064),
    .X(_08857_));
 sg13g2_a22oi_1 _15590_ (.Y(_08858_),
    .B1(_08604_),
    .B2(_08857_),
    .A2(_08579_),
    .A1(\cpu.icache.r_tag[2][22] ));
 sg13g2_nand4_1 _15591_ (.B(_08855_),
    .C(_08856_),
    .A(_08574_),
    .Y(_08859_),
    .D(_08858_));
 sg13g2_o21ai_1 _15592_ (.B1(_08859_),
    .Y(_08860_),
    .A1(\cpu.icache.r_tag[0][22] ),
    .A2(_08572_));
 sg13g2_xor2_1 _15593_ (.B(_08860_),
    .A(net449),
    .X(_08861_));
 sg13g2_mux4_1 _15594_ (.S0(net1070),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][11] ),
    .S1(net1066),
    .X(_08862_));
 sg13g2_mux4_1 _15595_ (.S0(_08528_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][11] ),
    .S1(_08536_),
    .X(_08863_));
 sg13g2_mux4_1 _15596_ (.S0(net1070),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][11] ),
    .S1(net1130),
    .X(_08864_));
 sg13g2_mux4_1 _15597_ (.S0(net1070),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][11] ),
    .S1(net1066),
    .X(_08865_));
 sg13g2_mux4_1 _15598_ (.S0(net1071),
    .A0(_08862_),
    .A1(_08863_),
    .A2(_08864_),
    .A3(_08865_),
    .S1(_08545_),
    .X(_08866_));
 sg13g2_mux4_1 _15599_ (.S0(net1070),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][11] ),
    .S1(net1066),
    .X(_08867_));
 sg13g2_mux4_1 _15600_ (.S0(net1070),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][11] ),
    .S1(net1066),
    .X(_08868_));
 sg13g2_mux4_1 _15601_ (.S0(net1070),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][11] ),
    .S1(net1130),
    .X(_08869_));
 sg13g2_mux4_1 _15602_ (.S0(net1070),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][11] ),
    .S1(net1130),
    .X(_08870_));
 sg13g2_mux4_1 _15603_ (.S0(net1071),
    .A0(_08867_),
    .A1(_08868_),
    .A2(_08869_),
    .A3(_08870_),
    .S1(_08453_),
    .X(_08871_));
 sg13g2_mux2_1 _15604_ (.A0(_08866_),
    .A1(_08871_),
    .S(net1129),
    .X(_08872_));
 sg13g2_nand2b_1 _15605_ (.Y(_08873_),
    .B(_08872_),
    .A_N(net1062));
 sg13g2_buf_2 _15606_ (.A(_08873_),
    .X(_08874_));
 sg13g2_nand2_1 _15607_ (.Y(_08875_),
    .A(\cpu.icache.r_tag[2][23] ),
    .B(net636));
 sg13g2_a22oi_1 _15608_ (.Y(_08876_),
    .B1(_08762_),
    .B2(\cpu.icache.r_tag[4][23] ),
    .A2(_08666_),
    .A1(\cpu.icache.r_tag[6][23] ));
 sg13g2_nor2_2 _15609_ (.A(net948),
    .B(_08593_),
    .Y(_08877_));
 sg13g2_a22oi_1 _15610_ (.Y(_08878_),
    .B1(_08877_),
    .B2(\cpu.icache.r_tag[3][23] ),
    .A2(net949),
    .A1(\cpu.icache.r_tag[5][23] ));
 sg13g2_nor2_1 _15611_ (.A(net822),
    .B(_08878_),
    .Y(_08879_));
 sg13g2_a221oi_1 _15612_ (.B2(\cpu.icache.r_tag[7][23] ),
    .C1(_08879_),
    .B1(_08700_),
    .A1(\cpu.icache.r_tag[1][23] ),
    .Y(_08880_),
    .A2(_08747_));
 sg13g2_nand4_1 _15613_ (.B(_08875_),
    .C(_08876_),
    .A(_08661_),
    .Y(_08881_),
    .D(_08880_));
 sg13g2_o21ai_1 _15614_ (.B1(_08881_),
    .Y(_08882_),
    .A1(\cpu.icache.r_tag[0][23] ),
    .A2(net453));
 sg13g2_xor2_1 _15615_ (.B(_08882_),
    .A(_08874_),
    .X(_08883_));
 sg13g2_mux4_1 _15616_ (.S0(net826),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][7] ),
    .S1(_08537_),
    .X(_08884_));
 sg13g2_mux4_1 _15617_ (.S0(net826),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][7] ),
    .S1(net954),
    .X(_08885_));
 sg13g2_mux4_1 _15618_ (.S0(_08528_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][7] ),
    .S1(_08537_),
    .X(_08886_));
 sg13g2_mux4_1 _15619_ (.S0(_08534_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][7] ),
    .S1(net954),
    .X(_08887_));
 sg13g2_mux4_1 _15620_ (.S0(net953),
    .A0(_08884_),
    .A1(_08885_),
    .A2(_08886_),
    .A3(_08887_),
    .S1(net1065),
    .X(_08888_));
 sg13g2_mux4_1 _15621_ (.S0(net826),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][7] ),
    .S1(net954),
    .X(_08889_));
 sg13g2_mux4_1 _15622_ (.S0(net826),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][7] ),
    .S1(net954),
    .X(_08890_));
 sg13g2_mux4_1 _15623_ (.S0(_08528_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][7] ),
    .S1(net954),
    .X(_08891_));
 sg13g2_mux4_1 _15624_ (.S0(_08528_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][7] ),
    .S1(net954),
    .X(_08892_));
 sg13g2_mux4_1 _15625_ (.S0(net953),
    .A0(_08889_),
    .A1(_08890_),
    .A2(_08891_),
    .A3(_08892_),
    .S1(net1065),
    .X(_08893_));
 sg13g2_mux2_1 _15626_ (.A0(_08888_),
    .A1(_08893_),
    .S(net1067),
    .X(_08894_));
 sg13g2_nand2b_1 _15627_ (.Y(_08895_),
    .B(_08894_),
    .A_N(net1062));
 sg13g2_buf_1 _15628_ (.A(_08895_),
    .X(_08896_));
 sg13g2_and2_1 _15629_ (.A(\cpu.icache.r_tag[3][19] ),
    .B(_08596_),
    .X(_08897_));
 sg13g2_a221oi_1 _15630_ (.B2(\cpu.icache.r_tag[6][19] ),
    .C1(_08897_),
    .B1(_08666_),
    .A1(\cpu.icache.r_tag[1][19] ),
    .Y(_08898_),
    .A2(net639));
 sg13g2_a22oi_1 _15631_ (.Y(_08899_),
    .B1(net811),
    .B2(\cpu.icache.r_tag[4][19] ),
    .A2(_08780_),
    .A1(\cpu.icache.r_tag[2][19] ));
 sg13g2_a22oi_1 _15632_ (.Y(_08900_),
    .B1(_08700_),
    .B2(\cpu.icache.r_tag[7][19] ),
    .A2(_08584_),
    .A1(\cpu.icache.r_tag[5][19] ));
 sg13g2_nand4_1 _15633_ (.B(_08898_),
    .C(_08899_),
    .A(_08571_),
    .Y(_08901_),
    .D(_08900_));
 sg13g2_o21ai_1 _15634_ (.B1(_08901_),
    .Y(_08902_),
    .A1(\cpu.icache.r_tag[0][19] ),
    .A2(_08661_));
 sg13g2_xnor2_1 _15635_ (.Y(_08903_),
    .A(net448),
    .B(_08902_));
 sg13g2_inv_1 _15636_ (.Y(_08904_),
    .A(_08903_));
 sg13g2_nor4_1 _15637_ (.A(_08841_),
    .B(_08861_),
    .C(_08883_),
    .D(_08904_),
    .Y(_08905_));
 sg13g2_mux4_1 _15638_ (.S0(net714),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][5] ),
    .S1(net817),
    .X(_08906_));
 sg13g2_mux4_1 _15639_ (.S0(net714),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][5] ),
    .S1(net817),
    .X(_08907_));
 sg13g2_mux4_1 _15640_ (.S0(net713),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][5] ),
    .S1(net813),
    .X(_08908_));
 sg13g2_mux4_1 _15641_ (.S0(net713),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][5] ),
    .S1(net813),
    .X(_08909_));
 sg13g2_mux4_1 _15642_ (.S0(_08693_),
    .A0(_08906_),
    .A1(_08907_),
    .A2(_08908_),
    .A3(_08909_),
    .S1(net941),
    .X(_08910_));
 sg13g2_mux4_1 _15643_ (.S0(_08686_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][5] ),
    .S1(net817),
    .X(_08911_));
 sg13g2_mux4_1 _15644_ (.S0(net714),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][5] ),
    .S1(net817),
    .X(_08912_));
 sg13g2_mux4_1 _15645_ (.S0(net715),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][5] ),
    .S1(net820),
    .X(_08913_));
 sg13g2_mux4_1 _15646_ (.S0(net715),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][5] ),
    .S1(net813),
    .X(_08914_));
 sg13g2_mux4_1 _15647_ (.S0(_08693_),
    .A0(_08911_),
    .A1(_08912_),
    .A2(_08913_),
    .A3(_08914_),
    .S1(net941),
    .X(_08915_));
 sg13g2_mux2_1 _15648_ (.A0(_08910_),
    .A1(_08915_),
    .S(net955),
    .X(_08916_));
 sg13g2_nand2b_1 _15649_ (.Y(_08917_),
    .B(_08916_),
    .A_N(net1062));
 sg13g2_buf_2 _15650_ (.A(_08917_),
    .X(_08918_));
 sg13g2_a22oi_1 _15651_ (.Y(_08919_),
    .B1(net556),
    .B2(\cpu.icache.r_tag[6][17] ),
    .A2(_08580_),
    .A1(\cpu.icache.r_tag[2][17] ));
 sg13g2_a22oi_1 _15652_ (.Y(_08920_),
    .B1(net814),
    .B2(\cpu.icache.r_tag[4][17] ),
    .A2(net558),
    .A1(\cpu.icache.r_tag[1][17] ));
 sg13g2_mux2_1 _15653_ (.A0(\cpu.icache.r_tag[7][17] ),
    .A1(\cpu.icache.r_tag[3][17] ),
    .S(net947),
    .X(_08921_));
 sg13g2_a22oi_1 _15654_ (.Y(_08922_),
    .B1(_08921_),
    .B2(net810),
    .A2(net949),
    .A1(\cpu.icache.r_tag[5][17] ));
 sg13g2_nand2b_1 _15655_ (.Y(_08923_),
    .B(net712),
    .A_N(_08922_));
 sg13g2_nand4_1 _15656_ (.B(_08919_),
    .C(_08920_),
    .A(net452),
    .Y(_08924_),
    .D(_08923_));
 sg13g2_o21ai_1 _15657_ (.B1(_08924_),
    .Y(_08925_),
    .A1(\cpu.icache.r_tag[0][17] ),
    .A2(_08573_));
 sg13g2_xnor2_1 _15658_ (.Y(_08926_),
    .A(net413),
    .B(_08925_));
 sg13g2_mux4_1 _15659_ (.S0(_08714_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][8] ),
    .S1(net817),
    .X(_08927_));
 sg13g2_mux4_1 _15660_ (.S0(_08686_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][8] ),
    .S1(_08687_),
    .X(_08928_));
 sg13g2_mux4_1 _15661_ (.S0(net715),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][8] ),
    .S1(net820),
    .X(_08929_));
 sg13g2_mux4_1 _15662_ (.S0(net715),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][8] ),
    .S1(_08715_),
    .X(_08930_));
 sg13g2_mux4_1 _15663_ (.S0(net815),
    .A0(_08927_),
    .A1(_08928_),
    .A2(_08929_),
    .A3(_08930_),
    .S1(net941),
    .X(_08931_));
 sg13g2_mux4_1 _15664_ (.S0(net713),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][8] ),
    .S1(net813),
    .X(_08932_));
 sg13g2_mux4_1 _15665_ (.S0(net713),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][8] ),
    .S1(_08687_),
    .X(_08933_));
 sg13g2_mux4_1 _15666_ (.S0(net715),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][8] ),
    .S1(net820),
    .X(_08934_));
 sg13g2_mux4_1 _15667_ (.S0(net715),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][8] ),
    .S1(net820),
    .X(_08935_));
 sg13g2_mux4_1 _15668_ (.S0(net824),
    .A0(_08932_),
    .A1(_08933_),
    .A2(_08934_),
    .A3(_08935_),
    .S1(net952),
    .X(_08936_));
 sg13g2_mux2_1 _15669_ (.A0(_08931_),
    .A1(_08936_),
    .S(net955),
    .X(_08937_));
 sg13g2_nand2b_1 _15670_ (.Y(_08938_),
    .B(_08937_),
    .A_N(net1062));
 sg13g2_buf_1 _15671_ (.A(_08938_),
    .X(_08939_));
 sg13g2_a22oi_1 _15672_ (.Y(_08940_),
    .B1(_08667_),
    .B2(\cpu.icache.r_tag[6][20] ),
    .A2(_08662_),
    .A1(\cpu.icache.r_tag[2][20] ));
 sg13g2_a22oi_1 _15673_ (.Y(_08941_),
    .B1(_08706_),
    .B2(\cpu.icache.r_tag[4][20] ),
    .A2(_08590_),
    .A1(\cpu.icache.r_tag[1][20] ));
 sg13g2_mux2_1 _15674_ (.A0(\cpu.icache.r_tag[7][20] ),
    .A1(\cpu.icache.r_tag[3][20] ),
    .S(net947),
    .X(_08942_));
 sg13g2_a22oi_1 _15675_ (.Y(_08943_),
    .B1(_08942_),
    .B2(net810),
    .A2(net949),
    .A1(\cpu.icache.r_tag[5][20] ));
 sg13g2_nand2b_1 _15676_ (.Y(_08944_),
    .B(net712),
    .A_N(_08943_));
 sg13g2_nand4_1 _15677_ (.B(_08940_),
    .C(_08941_),
    .A(_08575_),
    .Y(_08945_),
    .D(_08944_));
 sg13g2_o21ai_1 _15678_ (.B1(_08945_),
    .Y(_08946_),
    .A1(\cpu.icache.r_tag[0][20] ),
    .A2(_08573_));
 sg13g2_xnor2_1 _15679_ (.Y(_08947_),
    .A(net412),
    .B(_08946_));
 sg13g2_mux4_1 _15680_ (.S0(net713),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][9] ),
    .S1(net813),
    .X(_08948_));
 sg13g2_mux4_1 _15681_ (.S0(_08714_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][9] ),
    .S1(_08715_),
    .X(_08949_));
 sg13g2_mux4_1 _15682_ (.S0(_08615_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][9] ),
    .S1(net819),
    .X(_08950_));
 sg13g2_mux4_1 _15683_ (.S0(net716),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][9] ),
    .S1(_08622_),
    .X(_08951_));
 sg13g2_mux4_1 _15684_ (.S0(net824),
    .A0(_08948_),
    .A1(_08949_),
    .A2(_08950_),
    .A3(_08951_),
    .S1(_08546_),
    .X(_08952_));
 sg13g2_mux4_1 _15685_ (.S0(_08619_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][9] ),
    .S1(_08617_),
    .X(_08953_));
 sg13g2_mux4_1 _15686_ (.S0(_08619_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][9] ),
    .S1(_08617_),
    .X(_08954_));
 sg13g2_mux4_1 _15687_ (.S0(net718),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][9] ),
    .S1(net819),
    .X(_08955_));
 sg13g2_mux4_1 _15688_ (.S0(net716),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][9] ),
    .S1(net819),
    .X(_08956_));
 sg13g2_mux4_1 _15689_ (.S0(net824),
    .A0(_08953_),
    .A1(_08954_),
    .A2(_08955_),
    .A3(_08956_),
    .S1(net952),
    .X(_08957_));
 sg13g2_mux2_1 _15690_ (.A0(_08952_),
    .A1(_08957_),
    .S(_08532_),
    .X(_08958_));
 sg13g2_nand2b_1 _15691_ (.Y(_08959_),
    .B(_08958_),
    .A_N(net1062));
 sg13g2_buf_1 _15692_ (.A(_08959_),
    .X(_08960_));
 sg13g2_a22oi_1 _15693_ (.Y(_08961_),
    .B1(_08590_),
    .B2(\cpu.icache.r_tag[1][21] ),
    .A2(_08662_),
    .A1(\cpu.icache.r_tag[2][21] ));
 sg13g2_a22oi_1 _15694_ (.Y(_08962_),
    .B1(_08597_),
    .B2(\cpu.icache.r_tag[3][21] ),
    .A2(_08585_),
    .A1(\cpu.icache.r_tag[5][21] ));
 sg13g2_mux2_1 _15695_ (.A0(\cpu.icache.r_tag[4][21] ),
    .A1(\cpu.icache.r_tag[6][21] ),
    .S(_08606_),
    .X(_08963_));
 sg13g2_a22oi_1 _15696_ (.Y(_08964_),
    .B1(_08963_),
    .B2(net822),
    .A2(_08604_),
    .A1(\cpu.icache.r_tag[7][21] ));
 sg13g2_or2_1 _15697_ (.X(_08965_),
    .B(_08964_),
    .A(_08601_));
 sg13g2_nand3_1 _15698_ (.B(_08962_),
    .C(_08965_),
    .A(_08961_),
    .Y(_08966_));
 sg13g2_mux2_1 _15699_ (.A0(\cpu.icache.r_tag[0][21] ),
    .A1(_08966_),
    .S(_08575_),
    .X(_08967_));
 sg13g2_xor2_1 _15700_ (.B(_08967_),
    .A(net411),
    .X(_08968_));
 sg13g2_nand4_1 _15701_ (.B(_08926_),
    .C(_08947_),
    .A(_08905_),
    .Y(_08969_),
    .D(_08968_));
 sg13g2_nor3_2 _15702_ (.A(_08643_),
    .B(_08819_),
    .C(_08969_),
    .Y(_08970_));
 sg13g2_and3_1 _15703_ (.X(_08971_),
    .A(_08374_),
    .B(_08527_),
    .C(_08970_));
 sg13g2_buf_2 _15704_ (.A(_08971_),
    .X(_08972_));
 sg13g2_buf_1 _15705_ (.A(_08972_),
    .X(_08973_));
 sg13g2_buf_1 _15706_ (.A(_08972_),
    .X(_08974_));
 sg13g2_buf_1 _15707_ (.A(\cpu.ex.pc[1] ),
    .X(_08975_));
 sg13g2_buf_1 _15708_ (.A(_08975_),
    .X(_08976_));
 sg13g2_buf_1 _15709_ (.A(net1060),
    .X(_08977_));
 sg13g2_buf_1 _15710_ (.A(net937),
    .X(_08978_));
 sg13g2_and2_1 _15711_ (.A(net1128),
    .B(_08568_),
    .X(_08979_));
 sg13g2_buf_2 _15712_ (.A(_08979_),
    .X(_08980_));
 sg13g2_buf_1 _15713_ (.A(_08980_),
    .X(_08981_));
 sg13g2_mux2_1 _15714_ (.A0(\cpu.icache.r_data[7][16] ),
    .A1(\cpu.icache.r_data[3][16] ),
    .S(net823),
    .X(_08982_));
 sg13g2_a22oi_1 _15715_ (.Y(_08983_),
    .B1(_08982_),
    .B2(net711),
    .A2(net949),
    .A1(\cpu.icache.r_data[5][16] ));
 sg13g2_nand2b_1 _15716_ (.Y(_08984_),
    .B(net712),
    .A_N(_08983_));
 sg13g2_a22oi_1 _15717_ (.Y(_08985_),
    .B1(net814),
    .B2(\cpu.icache.r_data[4][16] ),
    .A2(net502),
    .A1(\cpu.icache.r_data[1][16] ));
 sg13g2_a22oi_1 _15718_ (.Y(_08986_),
    .B1(net556),
    .B2(\cpu.icache.r_data[6][16] ),
    .A2(net559),
    .A1(\cpu.icache.r_data[2][16] ));
 sg13g2_nand3_1 _15719_ (.B(_08985_),
    .C(_08986_),
    .A(_08984_),
    .Y(_08987_));
 sg13g2_a21oi_1 _15720_ (.A1(\cpu.icache.r_data[0][16] ),
    .A2(net499),
    .Y(_08988_),
    .B1(_08987_));
 sg13g2_nand2b_1 _15721_ (.Y(_08989_),
    .B(net499),
    .A_N(\cpu.icache.r_data[0][0] ));
 sg13g2_mux2_1 _15722_ (.A0(\cpu.icache.r_data[7][0] ),
    .A1(\cpu.icache.r_data[3][0] ),
    .S(net823),
    .X(_08990_));
 sg13g2_a22oi_1 _15723_ (.Y(_08991_),
    .B1(net637),
    .B2(_08990_),
    .A2(net559),
    .A1(\cpu.icache.r_data[2][0] ));
 sg13g2_buf_1 _15724_ (.A(net640),
    .X(_08992_));
 sg13g2_a22oi_1 _15725_ (.Y(_08993_),
    .B1(net556),
    .B2(\cpu.icache.r_data[6][0] ),
    .A2(net552),
    .A1(\cpu.icache.r_data[5][0] ));
 sg13g2_a22oi_1 _15726_ (.Y(_08994_),
    .B1(net814),
    .B2(\cpu.icache.r_data[4][0] ),
    .A2(net502),
    .A1(\cpu.icache.r_data[1][0] ));
 sg13g2_nand4_1 _15727_ (.B(_08991_),
    .C(_08993_),
    .A(net416),
    .Y(_08995_),
    .D(_08994_));
 sg13g2_a21oi_1 _15728_ (.A1(_08989_),
    .A2(_08995_),
    .Y(_08996_),
    .B1(net809));
 sg13g2_a21oi_1 _15729_ (.A1(net809),
    .A2(_08988_),
    .Y(_08997_),
    .B1(_08996_));
 sg13g2_buf_1 _15730_ (.A(_08997_),
    .X(_08998_));
 sg13g2_a22oi_1 _15731_ (.Y(_08999_),
    .B1(net814),
    .B2(\cpu.icache.r_data[4][1] ),
    .A2(net559),
    .A1(\cpu.icache.r_data[2][1] ));
 sg13g2_buf_1 _15732_ (.A(net557),
    .X(_09000_));
 sg13g2_a22oi_1 _15733_ (.Y(_09001_),
    .B1(net498),
    .B2(\cpu.icache.r_data[3][1] ),
    .A2(net502),
    .A1(\cpu.icache.r_data[1][1] ));
 sg13g2_mux2_1 _15734_ (.A0(\cpu.icache.r_data[5][1] ),
    .A1(\cpu.icache.r_data[7][1] ),
    .S(net946),
    .X(_09002_));
 sg13g2_a22oi_1 _15735_ (.Y(_09003_),
    .B1(_09002_),
    .B2(net812),
    .A2(_08784_),
    .A1(\cpu.icache.r_data[6][1] ));
 sg13g2_or2_1 _15736_ (.X(_09004_),
    .B(_09003_),
    .A(net823));
 sg13g2_nand3_1 _15737_ (.B(_09001_),
    .C(_09004_),
    .A(_08999_),
    .Y(_09005_));
 sg13g2_mux2_1 _15738_ (.A0(\cpu.icache.r_data[0][1] ),
    .A1(_09005_),
    .S(net416),
    .X(_09006_));
 sg13g2_buf_1 _15739_ (.A(net814),
    .X(_09007_));
 sg13g2_a22oi_1 _15740_ (.Y(_09008_),
    .B1(net710),
    .B2(\cpu.icache.r_data[4][17] ),
    .A2(net502),
    .A1(\cpu.icache.r_data[1][17] ));
 sg13g2_a22oi_1 _15741_ (.Y(_09009_),
    .B1(_08700_),
    .B2(\cpu.icache.r_data[7][17] ),
    .A2(net559),
    .A1(\cpu.icache.r_data[2][17] ));
 sg13g2_a22oi_1 _15742_ (.Y(_09010_),
    .B1(_08877_),
    .B2(\cpu.icache.r_data[3][17] ),
    .A2(net949),
    .A1(\cpu.icache.r_data[5][17] ));
 sg13g2_inv_1 _15743_ (.Y(_09011_),
    .A(_09010_));
 sg13g2_inv_1 _15744_ (.Y(_09012_),
    .A(_08975_));
 sg13g2_buf_1 _15745_ (.A(_09012_),
    .X(_09013_));
 sg13g2_a221oi_1 _15746_ (.B2(_08800_),
    .C1(net936),
    .B1(_09011_),
    .A1(\cpu.icache.r_data[6][17] ),
    .Y(_09014_),
    .A2(net556));
 sg13g2_nand2_1 _15747_ (.Y(_09015_),
    .A(\cpu.icache.r_data[0][17] ),
    .B(net499));
 sg13g2_nand4_1 _15748_ (.B(_09009_),
    .C(_09014_),
    .A(_09008_),
    .Y(_09016_),
    .D(_09015_));
 sg13g2_o21ai_1 _15749_ (.B1(_09016_),
    .Y(_09017_),
    .A1(net937),
    .A2(_09006_));
 sg13g2_buf_1 _15750_ (.A(_09017_),
    .X(_09018_));
 sg13g2_nand2_1 _15751_ (.Y(_09019_),
    .A(net212),
    .B(net240));
 sg13g2_buf_2 _15752_ (.A(_09019_),
    .X(_09020_));
 sg13g2_nor2_1 _15753_ (.A(_00204_),
    .B(_08569_),
    .Y(_09021_));
 sg13g2_mux2_1 _15754_ (.A0(\cpu.icache.r_data[5][31] ),
    .A1(\cpu.icache.r_data[7][31] ),
    .S(net1063),
    .X(_09022_));
 sg13g2_a22oi_1 _15755_ (.Y(_09023_),
    .B1(_09022_),
    .B2(net1061),
    .A2(_08784_),
    .A1(\cpu.icache.r_data[6][31] ));
 sg13g2_nor2_1 _15756_ (.A(net1064),
    .B(_09023_),
    .Y(_09024_));
 sg13g2_a22oi_1 _15757_ (.Y(_09025_),
    .B1(_08595_),
    .B2(\cpu.icache.r_data[3][31] ),
    .A2(_08588_),
    .A1(\cpu.icache.r_data[1][31] ));
 sg13g2_a22oi_1 _15758_ (.Y(_09026_),
    .B1(_08705_),
    .B2(\cpu.icache.r_data[4][31] ),
    .A2(_08577_),
    .A1(\cpu.icache.r_data[2][31] ));
 sg13g2_nand2_1 _15759_ (.Y(_09027_),
    .A(_09025_),
    .B(_09026_));
 sg13g2_nor3_1 _15760_ (.A(_09021_),
    .B(_09024_),
    .C(_09027_),
    .Y(_09028_));
 sg13g2_nand2_1 _15761_ (.Y(_09029_),
    .A(\cpu.icache.r_data[6][15] ),
    .B(_08665_));
 sg13g2_a22oi_1 _15762_ (.Y(_09030_),
    .B1(_08700_),
    .B2(\cpu.icache.r_data[7][15] ),
    .A2(_08588_),
    .A1(\cpu.icache.r_data[1][15] ));
 sg13g2_a22oi_1 _15763_ (.Y(_09031_),
    .B1(_08877_),
    .B2(\cpu.icache.r_data[3][15] ),
    .A2(_08581_),
    .A1(\cpu.icache.r_data[5][15] ));
 sg13g2_nand2b_1 _15764_ (.Y(_09032_),
    .B(_08669_),
    .A_N(_09031_));
 sg13g2_a22oi_1 _15765_ (.Y(_09033_),
    .B1(_08705_),
    .B2(\cpu.icache.r_data[4][15] ),
    .A2(_08577_),
    .A1(\cpu.icache.r_data[2][15] ));
 sg13g2_nand4_1 _15766_ (.B(_09030_),
    .C(_09032_),
    .A(_09029_),
    .Y(_09034_),
    .D(_09033_));
 sg13g2_nand2_1 _15767_ (.Y(_09035_),
    .A(_00203_),
    .B(_08980_));
 sg13g2_o21ai_1 _15768_ (.B1(_09035_),
    .Y(_09036_),
    .A1(_08980_),
    .A2(_09034_));
 sg13g2_mux2_1 _15769_ (.A0(_09028_),
    .A1(_09036_),
    .S(_09012_),
    .X(_09037_));
 sg13g2_buf_1 _15770_ (.A(_09037_),
    .X(_09038_));
 sg13g2_inv_1 _15771_ (.Y(_09039_),
    .A(_09038_));
 sg13g2_buf_1 _15772_ (.A(_09039_),
    .X(_09040_));
 sg13g2_nor2_1 _15773_ (.A(_00202_),
    .B(net560),
    .Y(_09041_));
 sg13g2_mux2_1 _15774_ (.A0(\cpu.icache.r_data[4][30] ),
    .A1(\cpu.icache.r_data[6][30] ),
    .S(net942),
    .X(_09042_));
 sg13g2_a22oi_1 _15775_ (.Y(_09043_),
    .B1(_09042_),
    .B2(net950),
    .A2(_08603_),
    .A1(\cpu.icache.r_data[7][30] ));
 sg13g2_nor2_1 _15776_ (.A(net947),
    .B(_09043_),
    .Y(_09044_));
 sg13g2_a22oi_1 _15777_ (.Y(_09045_),
    .B1(net638),
    .B2(\cpu.icache.r_data[3][30] ),
    .A2(net639),
    .A1(\cpu.icache.r_data[1][30] ));
 sg13g2_a22oi_1 _15778_ (.Y(_09046_),
    .B1(_08584_),
    .B2(\cpu.icache.r_data[5][30] ),
    .A2(net717),
    .A1(\cpu.icache.r_data[2][30] ));
 sg13g2_nand2_1 _15779_ (.Y(_09047_),
    .A(_09045_),
    .B(_09046_));
 sg13g2_nor3_1 _15780_ (.A(_09041_),
    .B(_09044_),
    .C(_09047_),
    .Y(_09048_));
 sg13g2_nand2_1 _15781_ (.Y(_09049_),
    .A(_00201_),
    .B(_08980_));
 sg13g2_a22oi_1 _15782_ (.Y(_09050_),
    .B1(net639),
    .B2(\cpu.icache.r_data[1][14] ),
    .A2(_08584_),
    .A1(\cpu.icache.r_data[5][14] ));
 sg13g2_a22oi_1 _15783_ (.Y(_09051_),
    .B1(_08705_),
    .B2(\cpu.icache.r_data[4][14] ),
    .A2(net717),
    .A1(\cpu.icache.r_data[2][14] ));
 sg13g2_mux2_1 _15784_ (.A0(\cpu.icache.r_data[7][14] ),
    .A1(\cpu.icache.r_data[3][14] ),
    .S(net1128),
    .X(_09052_));
 sg13g2_a22oi_1 _15785_ (.Y(_09053_),
    .B1(_09052_),
    .B2(net1061),
    .A2(_08812_),
    .A1(\cpu.icache.r_data[6][14] ));
 sg13g2_nand2b_1 _15786_ (.Y(_09054_),
    .B(net946),
    .A_N(_09053_));
 sg13g2_nand4_1 _15787_ (.B(_09050_),
    .C(_09051_),
    .A(net560),
    .Y(_09055_),
    .D(_09054_));
 sg13g2_a21oi_1 _15788_ (.A1(_09049_),
    .A2(_09055_),
    .Y(_09056_),
    .B1(net1060));
 sg13g2_a21oi_1 _15789_ (.A1(net937),
    .A2(_09048_),
    .Y(_09057_),
    .B1(_09056_));
 sg13g2_buf_1 _15790_ (.A(_09057_),
    .X(_09058_));
 sg13g2_and2_1 _15791_ (.A(_08671_),
    .B(\cpu.icache.r_data[6][13] ),
    .X(_09059_));
 sg13g2_a21oi_1 _15792_ (.A1(_08592_),
    .A2(\cpu.icache.r_data[4][13] ),
    .Y(_09060_),
    .B1(_09059_));
 sg13g2_nor2_1 _15793_ (.A(_08566_),
    .B(net942),
    .Y(_09061_));
 sg13g2_a22oi_1 _15794_ (.Y(_09062_),
    .B1(_08603_),
    .B2(\cpu.icache.r_data[7][13] ),
    .A2(_09061_),
    .A1(\cpu.icache.r_data[5][13] ));
 sg13g2_o21ai_1 _15795_ (.B1(_09062_),
    .Y(_09063_),
    .A1(net812),
    .A2(_09060_));
 sg13g2_buf_1 _15796_ (.A(_08593_),
    .X(_09064_));
 sg13g2_buf_1 _15797_ (.A(net935),
    .X(_09065_));
 sg13g2_a22oi_1 _15798_ (.Y(_09066_),
    .B1(net638),
    .B2(\cpu.icache.r_data[3][13] ),
    .A2(net634),
    .A1(\cpu.icache.r_data[2][13] ));
 sg13g2_inv_1 _15799_ (.Y(_09067_),
    .A(_09066_));
 sg13g2_a221oi_1 _15800_ (.B2(_09065_),
    .C1(_09067_),
    .B1(_09063_),
    .A1(\cpu.icache.r_data[1][13] ),
    .Y(_09068_),
    .A2(net558));
 sg13g2_nor2_1 _15801_ (.A(\cpu.icache.r_data[0][13] ),
    .B(net501),
    .Y(_09069_));
 sg13g2_a21oi_1 _15802_ (.A1(_08572_),
    .A2(_09068_),
    .Y(_09070_),
    .B1(_09069_));
 sg13g2_nand2_1 _15803_ (.Y(_09071_),
    .A(\cpu.icache.r_data[0][29] ),
    .B(_08980_));
 sg13g2_mux4_1 _15804_ (.S0(net943),
    .A0(\cpu.icache.r_data[4][29] ),
    .A1(\cpu.icache.r_data[5][29] ),
    .A2(\cpu.icache.r_data[6][29] ),
    .A3(\cpu.icache.r_data[7][29] ),
    .S1(net810),
    .X(_09072_));
 sg13g2_nand2_1 _15805_ (.Y(_09073_),
    .A(net935),
    .B(_09072_));
 sg13g2_nand2_1 _15806_ (.Y(_09074_),
    .A(\cpu.icache.r_data[2][29] ),
    .B(net636));
 sg13g2_a22oi_1 _15807_ (.Y(_09075_),
    .B1(net557),
    .B2(\cpu.icache.r_data[3][29] ),
    .A2(net555),
    .A1(\cpu.icache.r_data[1][29] ));
 sg13g2_nand4_1 _15808_ (.B(_09073_),
    .C(_09074_),
    .A(_09071_),
    .Y(_09076_),
    .D(_09075_));
 sg13g2_and2_1 _15809_ (.A(net1060),
    .B(_09076_),
    .X(_09077_));
 sg13g2_a21o_1 _15810_ (.A2(_09070_),
    .A1(net936),
    .B1(_09077_),
    .X(_09078_));
 sg13g2_buf_1 _15811_ (.A(_09078_),
    .X(_09079_));
 sg13g2_nor2_1 _15812_ (.A(_09058_),
    .B(_09079_),
    .Y(_09080_));
 sg13g2_buf_1 _15813_ (.A(_09080_),
    .X(_09081_));
 sg13g2_nand2_1 _15814_ (.Y(_09082_),
    .A(net239),
    .B(_09081_));
 sg13g2_buf_1 _15815_ (.A(_09082_),
    .X(_09083_));
 sg13g2_nor2_2 _15816_ (.A(_09020_),
    .B(net152),
    .Y(_09084_));
 sg13g2_nor2_1 _15817_ (.A(_00206_),
    .B(net503),
    .Y(_09085_));
 sg13g2_mux2_1 _15818_ (.A0(\cpu.icache.r_data[7][26] ),
    .A1(\cpu.icache.r_data[3][26] ),
    .S(net1064),
    .X(_09086_));
 sg13g2_a22oi_1 _15819_ (.Y(_09087_),
    .B1(_09086_),
    .B2(_08801_),
    .A2(_08582_),
    .A1(\cpu.icache.r_data[5][26] ));
 sg13g2_nor2_1 _15820_ (.A(net822),
    .B(_09087_),
    .Y(_09088_));
 sg13g2_a22oi_1 _15821_ (.Y(_09089_),
    .B1(net811),
    .B2(\cpu.icache.r_data[4][26] ),
    .A2(net641),
    .A1(\cpu.icache.r_data[2][26] ));
 sg13g2_a22oi_1 _15822_ (.Y(_09090_),
    .B1(net635),
    .B2(\cpu.icache.r_data[6][26] ),
    .A2(net555),
    .A1(\cpu.icache.r_data[1][26] ));
 sg13g2_nand2_1 _15823_ (.Y(_09091_),
    .A(_09089_),
    .B(_09090_));
 sg13g2_nor3_1 _15824_ (.A(_09085_),
    .B(_09088_),
    .C(_09091_),
    .Y(_09092_));
 sg13g2_nand2_1 _15825_ (.Y(_09093_),
    .A(_00205_),
    .B(net499));
 sg13g2_mux4_1 _15826_ (.S0(_08670_),
    .A0(\cpu.icache.r_data[4][10] ),
    .A1(\cpu.icache.r_data[5][10] ),
    .A2(\cpu.icache.r_data[6][10] ),
    .A3(\cpu.icache.r_data[7][10] ),
    .S1(net946),
    .X(_09094_));
 sg13g2_nand2_1 _15827_ (.Y(_09095_),
    .A(net935),
    .B(_09094_));
 sg13g2_a22oi_1 _15828_ (.Y(_09096_),
    .B1(net554),
    .B2(\cpu.icache.r_data[3][10] ),
    .A2(net634),
    .A1(\cpu.icache.r_data[2][10] ));
 sg13g2_nand2_1 _15829_ (.Y(_09097_),
    .A(\cpu.icache.r_data[1][10] ),
    .B(net555));
 sg13g2_nand4_1 _15830_ (.B(_09095_),
    .C(_09096_),
    .A(net503),
    .Y(_09098_),
    .D(_09097_));
 sg13g2_a21oi_1 _15831_ (.A1(_09093_),
    .A2(_09098_),
    .Y(_09099_),
    .B1(net1060));
 sg13g2_a21oi_1 _15832_ (.A1(net937),
    .A2(_09092_),
    .Y(_09100_),
    .B1(_09099_));
 sg13g2_buf_2 _15833_ (.A(_09100_),
    .X(_09101_));
 sg13g2_buf_1 _15834_ (.A(_09101_),
    .X(_09102_));
 sg13g2_mux4_1 _15835_ (.S0(_08732_),
    .A0(\cpu.icache.r_data[4][27] ),
    .A1(\cpu.icache.r_data[5][27] ),
    .A2(\cpu.icache.r_data[6][27] ),
    .A3(\cpu.icache.r_data[7][27] ),
    .S1(net711),
    .X(_09103_));
 sg13g2_and2_1 _15836_ (.A(\cpu.icache.r_data[1][27] ),
    .B(net553),
    .X(_09104_));
 sg13g2_a221oi_1 _15837_ (.B2(\cpu.icache.r_data[3][27] ),
    .C1(_09104_),
    .B1(net554),
    .A1(\cpu.icache.r_data[2][27] ),
    .Y(_09105_),
    .A2(net641));
 sg13g2_o21ai_1 _15838_ (.B1(_09105_),
    .Y(_09106_),
    .A1(_00208_),
    .A2(net501));
 sg13g2_a21oi_1 _15839_ (.A1(_09065_),
    .A2(_09103_),
    .Y(_09107_),
    .B1(_09106_));
 sg13g2_nand2_1 _15840_ (.Y(_09108_),
    .A(_00207_),
    .B(net499));
 sg13g2_and2_1 _15841_ (.A(\cpu.icache.r_data[3][11] ),
    .B(net638),
    .X(_09109_));
 sg13g2_a221oi_1 _15842_ (.B2(\cpu.icache.r_data[6][11] ),
    .C1(_09109_),
    .B1(net635),
    .A1(\cpu.icache.r_data[1][11] ),
    .Y(_09110_),
    .A2(net555));
 sg13g2_a22oi_1 _15843_ (.Y(_09111_),
    .B1(_08706_),
    .B2(\cpu.icache.r_data[4][11] ),
    .A2(net641),
    .A1(\cpu.icache.r_data[2][11] ));
 sg13g2_a22oi_1 _15844_ (.Y(_09112_),
    .B1(_08700_),
    .B2(\cpu.icache.r_data[7][11] ),
    .A2(net640),
    .A1(\cpu.icache.r_data[5][11] ));
 sg13g2_nand4_1 _15845_ (.B(_09110_),
    .C(_09111_),
    .A(net501),
    .Y(_09113_),
    .D(_09112_));
 sg13g2_a21oi_1 _15846_ (.A1(_09108_),
    .A2(_09113_),
    .Y(_09114_),
    .B1(net937));
 sg13g2_a21oi_1 _15847_ (.A1(net937),
    .A2(_09107_),
    .Y(_09115_),
    .B1(_09114_));
 sg13g2_buf_1 _15848_ (.A(_09115_),
    .X(_09116_));
 sg13g2_inv_2 _15849_ (.Y(_09117_),
    .A(_09116_));
 sg13g2_nand4_1 _15850_ (.B(_09084_),
    .C(net238),
    .A(net119),
    .Y(_09118_),
    .D(_09117_));
 sg13g2_o21ai_1 _15851_ (.B1(_09118_),
    .Y(_00016_),
    .A1(_08373_),
    .A2(_08973_));
 sg13g2_buf_1 _15852_ (.A(\cpu.dec.r_op[6] ),
    .X(_09119_));
 sg13g2_buf_1 _15853_ (.A(_09119_),
    .X(_09120_));
 sg13g2_inv_2 _15854_ (.Y(_09121_),
    .A(net1059));
 sg13g2_mux4_1 _15855_ (.S0(net812),
    .A0(\cpu.icache.r_data[4][22] ),
    .A1(\cpu.icache.r_data[5][22] ),
    .A2(\cpu.icache.r_data[6][22] ),
    .A3(\cpu.icache.r_data[7][22] ),
    .S1(net810),
    .X(_09122_));
 sg13g2_and2_1 _15856_ (.A(\cpu.icache.r_data[1][22] ),
    .B(net639),
    .X(_09123_));
 sg13g2_a221oi_1 _15857_ (.B2(\cpu.icache.r_data[3][22] ),
    .C1(_09123_),
    .B1(net554),
    .A1(\cpu.icache.r_data[2][22] ),
    .Y(_09124_),
    .A2(net634));
 sg13g2_o21ai_1 _15858_ (.B1(_09124_),
    .Y(_09125_),
    .A1(_00212_),
    .A2(net504));
 sg13g2_a21oi_1 _15859_ (.A1(net808),
    .A2(_09122_),
    .Y(_09126_),
    .B1(_09125_));
 sg13g2_nand2_1 _15860_ (.Y(_09127_),
    .A(_00211_),
    .B(_08980_));
 sg13g2_a22oi_1 _15861_ (.Y(_09128_),
    .B1(net640),
    .B2(\cpu.icache.r_data[5][6] ),
    .A2(net634),
    .A1(\cpu.icache.r_data[2][6] ));
 sg13g2_a22oi_1 _15862_ (.Y(_09129_),
    .B1(net554),
    .B2(\cpu.icache.r_data[3][6] ),
    .A2(net553),
    .A1(\cpu.icache.r_data[1][6] ));
 sg13g2_mux2_1 _15863_ (.A0(\cpu.icache.r_data[4][6] ),
    .A1(\cpu.icache.r_data[6][6] ),
    .S(net1063),
    .X(_09130_));
 sg13g2_a22oi_1 _15864_ (.Y(_09131_),
    .B1(_09130_),
    .B2(net950),
    .A2(_08603_),
    .A1(\cpu.icache.r_data[7][6] ));
 sg13g2_or2_1 _15865_ (.X(_09132_),
    .B(_09131_),
    .A(net947));
 sg13g2_nand4_1 _15866_ (.B(_09128_),
    .C(_09129_),
    .A(net504),
    .Y(_09133_),
    .D(_09132_));
 sg13g2_a21oi_1 _15867_ (.A1(_09127_),
    .A2(_09133_),
    .Y(_09134_),
    .B1(net1060));
 sg13g2_a21oi_1 _15868_ (.A1(net809),
    .A2(_09126_),
    .Y(_09135_),
    .B1(_09134_));
 sg13g2_buf_2 _15869_ (.A(_09135_),
    .X(_09136_));
 sg13g2_mux4_1 _15870_ (.S0(net812),
    .A0(\cpu.icache.r_data[4][21] ),
    .A1(\cpu.icache.r_data[5][21] ),
    .A2(\cpu.icache.r_data[6][21] ),
    .A3(\cpu.icache.r_data[7][21] ),
    .S1(net711),
    .X(_09137_));
 sg13g2_and2_1 _15871_ (.A(\cpu.icache.r_data[1][21] ),
    .B(net553),
    .X(_09138_));
 sg13g2_a221oi_1 _15872_ (.B2(\cpu.icache.r_data[3][21] ),
    .C1(_09138_),
    .B1(net554),
    .A1(\cpu.icache.r_data[2][21] ),
    .Y(_09139_),
    .A2(net641));
 sg13g2_o21ai_1 _15873_ (.B1(_09139_),
    .Y(_09140_),
    .A1(_00210_),
    .A2(net501));
 sg13g2_a21oi_1 _15874_ (.A1(net808),
    .A2(_09137_),
    .Y(_09141_),
    .B1(_09140_));
 sg13g2_nand2_1 _15875_ (.Y(_09142_),
    .A(_00209_),
    .B(net499));
 sg13g2_mux4_1 _15876_ (.S0(_08670_),
    .A0(\cpu.icache.r_data[4][5] ),
    .A1(\cpu.icache.r_data[5][5] ),
    .A2(\cpu.icache.r_data[6][5] ),
    .A3(\cpu.icache.r_data[7][5] ),
    .S1(net810),
    .X(_09143_));
 sg13g2_nand2_1 _15877_ (.Y(_09144_),
    .A(net808),
    .B(_09143_));
 sg13g2_a22oi_1 _15878_ (.Y(_09145_),
    .B1(net557),
    .B2(\cpu.icache.r_data[3][5] ),
    .A2(net636),
    .A1(\cpu.icache.r_data[2][5] ));
 sg13g2_nand2_1 _15879_ (.Y(_09146_),
    .A(\cpu.icache.r_data[1][5] ),
    .B(net558));
 sg13g2_nand4_1 _15880_ (.B(_09144_),
    .C(_09145_),
    .A(net501),
    .Y(_09147_),
    .D(_09146_));
 sg13g2_nand3_1 _15881_ (.B(_09142_),
    .C(_09147_),
    .A(net936),
    .Y(_09148_));
 sg13g2_o21ai_1 _15882_ (.B1(_09148_),
    .Y(_09149_),
    .A1(net936),
    .A2(_09141_));
 sg13g2_buf_1 _15883_ (.A(_09149_),
    .X(_09150_));
 sg13g2_buf_1 _15884_ (.A(_09150_),
    .X(_09151_));
 sg13g2_nor2_1 _15885_ (.A(_09136_),
    .B(net211),
    .Y(_09152_));
 sg13g2_inv_1 _15886_ (.Y(_09153_),
    .A(_09101_));
 sg13g2_nor2_1 _15887_ (.A(_09153_),
    .B(_09117_),
    .Y(_09154_));
 sg13g2_nand4_1 _15888_ (.B(_09084_),
    .C(_09152_),
    .A(net119),
    .Y(_09155_),
    .D(_09154_));
 sg13g2_o21ai_1 _15889_ (.B1(_09155_),
    .Y(_00017_),
    .A1(_09121_),
    .A2(_08973_));
 sg13g2_buf_2 _15890_ (.A(\cpu.dec.r_op[4] ),
    .X(_09156_));
 sg13g2_buf_1 _15891_ (.A(_09156_),
    .X(_09157_));
 sg13g2_buf_2 _15892_ (.A(_08833_),
    .X(_09158_));
 sg13g2_xor2_1 _15893_ (.B(_08840_),
    .A(net410),
    .X(_09159_));
 sg13g2_nand4_1 _15894_ (.B(_09159_),
    .C(_08926_),
    .A(_08737_),
    .Y(_09160_),
    .D(_08947_));
 sg13g2_or2_1 _15895_ (.X(_09161_),
    .B(_09160_),
    .A(_08643_));
 sg13g2_nand2b_1 _15896_ (.Y(_09162_),
    .B(_08968_),
    .A_N(_08883_));
 sg13g2_nand3_1 _15897_ (.B(_08790_),
    .C(_08805_),
    .A(_08756_),
    .Y(_09163_));
 sg13g2_nand4_1 _15898_ (.B(_08775_),
    .C(_08799_),
    .A(_08767_),
    .Y(_09164_),
    .D(_08817_));
 sg13g2_nor3_1 _15899_ (.A(_08904_),
    .B(_09163_),
    .C(_09164_),
    .Y(_09165_));
 sg13g2_nand2_1 _15900_ (.Y(_09166_),
    .A(_08713_),
    .B(_09165_));
 sg13g2_nor4_2 _15901_ (.A(_08861_),
    .B(_09161_),
    .C(_09162_),
    .Y(_09167_),
    .D(_09166_));
 sg13g2_nand3_1 _15902_ (.B(_08527_),
    .C(_09167_),
    .A(_08374_),
    .Y(_09168_));
 sg13g2_buf_1 _15903_ (.A(_09168_),
    .X(_09169_));
 sg13g2_buf_1 _15904_ (.A(_09169_),
    .X(_09170_));
 sg13g2_buf_1 _15905_ (.A(net108),
    .X(_09171_));
 sg13g2_a21o_1 _15906_ (.A2(_09126_),
    .A1(_08977_),
    .B1(_09134_),
    .X(_09172_));
 sg13g2_buf_1 _15907_ (.A(_09172_),
    .X(_09173_));
 sg13g2_inv_2 _15908_ (.Y(_09174_),
    .A(_09150_));
 sg13g2_nand2_2 _15909_ (.Y(_09175_),
    .A(net281),
    .B(_09174_));
 sg13g2_inv_1 _15910_ (.Y(_09176_),
    .A(_00213_));
 sg13g2_and2_1 _15911_ (.A(_08606_),
    .B(\cpu.icache.r_data[6][12] ),
    .X(_09177_));
 sg13g2_a21oi_1 _15912_ (.A1(_08592_),
    .A2(\cpu.icache.r_data[4][12] ),
    .Y(_09178_),
    .B1(_09177_));
 sg13g2_a22oi_1 _15913_ (.Y(_09179_),
    .B1(net637),
    .B2(\cpu.icache.r_data[7][12] ),
    .A2(_09061_),
    .A1(\cpu.icache.r_data[5][12] ));
 sg13g2_o21ai_1 _15914_ (.B1(_09179_),
    .Y(_09180_),
    .A1(net812),
    .A2(_09178_));
 sg13g2_nand2_1 _15915_ (.Y(_09181_),
    .A(net808),
    .B(_09180_));
 sg13g2_nand2_1 _15916_ (.Y(_09182_),
    .A(\cpu.icache.r_data[1][12] ),
    .B(net502));
 sg13g2_a22oi_1 _15917_ (.Y(_09183_),
    .B1(net557),
    .B2(\cpu.icache.r_data[3][12] ),
    .A2(net636),
    .A1(\cpu.icache.r_data[2][12] ));
 sg13g2_nand4_1 _15918_ (.B(_09181_),
    .C(_09182_),
    .A(net452),
    .Y(_09184_),
    .D(_09183_));
 sg13g2_o21ai_1 _15919_ (.B1(_09184_),
    .Y(_09185_),
    .A1(_09176_),
    .A2(net416));
 sg13g2_mux4_1 _15920_ (.S0(_08800_),
    .A0(\cpu.icache.r_data[4][28] ),
    .A1(\cpu.icache.r_data[5][28] ),
    .A2(\cpu.icache.r_data[6][28] ),
    .A3(\cpu.icache.r_data[7][28] ),
    .S1(_08802_),
    .X(_09186_));
 sg13g2_and2_1 _15921_ (.A(\cpu.icache.r_data[1][28] ),
    .B(net558),
    .X(_09187_));
 sg13g2_a221oi_1 _15922_ (.B2(\cpu.icache.r_data[3][28] ),
    .C1(_09187_),
    .B1(net557),
    .A1(\cpu.icache.r_data[2][28] ),
    .Y(_09188_),
    .A2(net636));
 sg13g2_o21ai_1 _15923_ (.B1(_09188_),
    .Y(_09189_),
    .A1(_00214_),
    .A2(net452));
 sg13g2_a21oi_1 _15924_ (.A1(net808),
    .A2(_09186_),
    .Y(_09190_),
    .B1(_09189_));
 sg13g2_mux2_1 _15925_ (.A0(_09185_),
    .A1(_09190_),
    .S(net937),
    .X(_09191_));
 sg13g2_buf_1 _15926_ (.A(_09191_),
    .X(_09192_));
 sg13g2_buf_1 _15927_ (.A(_09192_),
    .X(_09193_));
 sg13g2_buf_1 _15928_ (.A(_09193_),
    .X(_09194_));
 sg13g2_buf_1 _15929_ (.A(_09038_),
    .X(_09195_));
 sg13g2_nor3_1 _15930_ (.A(net280),
    .B(_09058_),
    .C(_09079_),
    .Y(_09196_));
 sg13g2_buf_2 _15931_ (.A(_09196_),
    .X(_09197_));
 sg13g2_buf_1 _15932_ (.A(_09197_),
    .X(_09198_));
 sg13g2_inv_1 _15933_ (.Y(_09199_),
    .A(net240));
 sg13g2_nand2_1 _15934_ (.Y(_09200_),
    .A(net212),
    .B(_09199_));
 sg13g2_buf_1 _15935_ (.A(_09200_),
    .X(_09201_));
 sg13g2_nor3_2 _15936_ (.A(_09153_),
    .B(_09117_),
    .C(net151),
    .Y(_09202_));
 sg13g2_nand2_1 _15937_ (.Y(_09203_),
    .A(net179),
    .B(_09202_));
 sg13g2_nor4_1 _15938_ (.A(net108),
    .B(_09175_),
    .C(net180),
    .D(_09203_),
    .Y(_09204_));
 sg13g2_a21o_1 _15939_ (.A2(net92),
    .A1(net1058),
    .B1(_09204_),
    .X(_00015_));
 sg13g2_nand2_1 _15940_ (.Y(_09205_),
    .A(_09151_),
    .B(net180));
 sg13g2_nand3_1 _15941_ (.B(net281),
    .C(_09154_),
    .A(_09084_),
    .Y(_09206_));
 sg13g2_mux4_1 _15942_ (.S0(net1061),
    .A0(\cpu.icache.r_data[4][3] ),
    .A1(\cpu.icache.r_data[5][3] ),
    .A2(\cpu.icache.r_data[6][3] ),
    .A3(\cpu.icache.r_data[7][3] ),
    .S1(net942),
    .X(_09207_));
 sg13g2_nand2_1 _15943_ (.Y(_09208_),
    .A(net935),
    .B(_09207_));
 sg13g2_a22oi_1 _15944_ (.Y(_09209_),
    .B1(net638),
    .B2(\cpu.icache.r_data[3][3] ),
    .A2(net717),
    .A1(\cpu.icache.r_data[2][3] ));
 sg13g2_nand2_1 _15945_ (.Y(_09210_),
    .A(\cpu.icache.r_data[1][3] ),
    .B(net553));
 sg13g2_and4_1 _15946_ (.A(net504),
    .B(_09208_),
    .C(_09209_),
    .D(_09210_),
    .X(_09211_));
 sg13g2_a21oi_1 _15947_ (.A1(_00217_),
    .A2(net499),
    .Y(_09212_),
    .B1(_09211_));
 sg13g2_nor2_1 _15948_ (.A(_00218_),
    .B(net504),
    .Y(_09213_));
 sg13g2_mux2_1 _15949_ (.A0(\cpu.icache.r_data[4][19] ),
    .A1(\cpu.icache.r_data[6][19] ),
    .S(net942),
    .X(_09214_));
 sg13g2_a22oi_1 _15950_ (.Y(_09215_),
    .B1(_09214_),
    .B2(net822),
    .A2(net637),
    .A1(\cpu.icache.r_data[7][19] ));
 sg13g2_nor2_1 _15951_ (.A(net823),
    .B(_09215_),
    .Y(_09216_));
 sg13g2_a22oi_1 _15952_ (.Y(_09217_),
    .B1(net554),
    .B2(\cpu.icache.r_data[3][19] ),
    .A2(net553),
    .A1(\cpu.icache.r_data[1][19] ));
 sg13g2_a22oi_1 _15953_ (.Y(_09218_),
    .B1(_08584_),
    .B2(\cpu.icache.r_data[5][19] ),
    .A2(net634),
    .A1(\cpu.icache.r_data[2][19] ));
 sg13g2_nand2_1 _15954_ (.Y(_09219_),
    .A(_09217_),
    .B(_09218_));
 sg13g2_or4_1 _15955_ (.A(net936),
    .B(_09213_),
    .C(_09216_),
    .D(_09219_),
    .X(_09220_));
 sg13g2_o21ai_1 _15956_ (.B1(_09220_),
    .Y(_09221_),
    .A1(net1060),
    .A2(_09212_));
 sg13g2_buf_2 _15957_ (.A(_09221_),
    .X(_09222_));
 sg13g2_nor2_1 _15958_ (.A(_00216_),
    .B(net416),
    .Y(_09223_));
 sg13g2_mux2_1 _15959_ (.A0(\cpu.icache.r_data[7][18] ),
    .A1(\cpu.icache.r_data[3][18] ),
    .S(net823),
    .X(_09224_));
 sg13g2_a22oi_1 _15960_ (.Y(_09225_),
    .B1(_09224_),
    .B2(_08802_),
    .A2(net949),
    .A1(\cpu.icache.r_data[5][18] ));
 sg13g2_nor2_1 _15961_ (.A(_08608_),
    .B(_09225_),
    .Y(_09226_));
 sg13g2_a22oi_1 _15962_ (.Y(_09227_),
    .B1(net814),
    .B2(\cpu.icache.r_data[4][18] ),
    .A2(net559),
    .A1(\cpu.icache.r_data[2][18] ));
 sg13g2_a22oi_1 _15963_ (.Y(_09228_),
    .B1(net556),
    .B2(\cpu.icache.r_data[6][18] ),
    .A2(net502),
    .A1(\cpu.icache.r_data[1][18] ));
 sg13g2_nand2_1 _15964_ (.Y(_09229_),
    .A(_09227_),
    .B(_09228_));
 sg13g2_nor3_1 _15965_ (.A(_09223_),
    .B(_09226_),
    .C(_09229_),
    .Y(_09230_));
 sg13g2_nand2_1 _15966_ (.Y(_09231_),
    .A(_00215_),
    .B(net499));
 sg13g2_mux4_1 _15967_ (.S0(net812),
    .A0(\cpu.icache.r_data[4][2] ),
    .A1(\cpu.icache.r_data[5][2] ),
    .A2(\cpu.icache.r_data[6][2] ),
    .A3(\cpu.icache.r_data[7][2] ),
    .S1(net810),
    .X(_09232_));
 sg13g2_nand2_1 _15968_ (.Y(_09233_),
    .A(net808),
    .B(_09232_));
 sg13g2_a22oi_1 _15969_ (.Y(_09234_),
    .B1(net498),
    .B2(\cpu.icache.r_data[3][2] ),
    .A2(net559),
    .A1(\cpu.icache.r_data[2][2] ));
 sg13g2_nand2_1 _15970_ (.Y(_09235_),
    .A(\cpu.icache.r_data[1][2] ),
    .B(net502));
 sg13g2_nand4_1 _15971_ (.B(_09233_),
    .C(_09234_),
    .A(net416),
    .Y(_09236_),
    .D(_09235_));
 sg13g2_a21oi_1 _15972_ (.A1(_09231_),
    .A2(_09236_),
    .Y(_09237_),
    .B1(net937));
 sg13g2_a21oi_1 _15973_ (.A1(_08978_),
    .A2(_09230_),
    .Y(_09238_),
    .B1(_09237_));
 sg13g2_buf_1 _15974_ (.A(_09238_),
    .X(_09239_));
 sg13g2_inv_1 _15975_ (.Y(_09240_),
    .A(net209));
 sg13g2_nor2_1 _15976_ (.A(_09222_),
    .B(_09240_),
    .Y(_09241_));
 sg13g2_mux4_1 _15977_ (.S0(net1061),
    .A0(\cpu.icache.r_data[4][4] ),
    .A1(\cpu.icache.r_data[5][4] ),
    .A2(\cpu.icache.r_data[6][4] ),
    .A3(\cpu.icache.r_data[7][4] ),
    .S1(net946),
    .X(_09242_));
 sg13g2_nand2_1 _15978_ (.Y(_09243_),
    .A(_09064_),
    .B(_09242_));
 sg13g2_a22oi_1 _15979_ (.Y(_09244_),
    .B1(net554),
    .B2(\cpu.icache.r_data[3][4] ),
    .A2(net634),
    .A1(\cpu.icache.r_data[2][4] ));
 sg13g2_nand2_1 _15980_ (.Y(_09245_),
    .A(\cpu.icache.r_data[1][4] ),
    .B(net555));
 sg13g2_and4_1 _15981_ (.A(net503),
    .B(_09243_),
    .C(_09244_),
    .D(_09245_),
    .X(_09246_));
 sg13g2_a21oi_1 _15982_ (.A1(_00219_),
    .A2(_08981_),
    .Y(_09247_),
    .B1(_09246_));
 sg13g2_a22oi_1 _15983_ (.Y(_09248_),
    .B1(net558),
    .B2(\cpu.icache.r_data[1][20] ),
    .A2(net636),
    .A1(\cpu.icache.r_data[2][20] ));
 sg13g2_a22oi_1 _15984_ (.Y(_09249_),
    .B1(net814),
    .B2(\cpu.icache.r_data[4][20] ),
    .A2(_08700_),
    .A1(\cpu.icache.r_data[7][20] ));
 sg13g2_a22oi_1 _15985_ (.Y(_09250_),
    .B1(_08877_),
    .B2(\cpu.icache.r_data[3][20] ),
    .A2(net949),
    .A1(\cpu.icache.r_data[5][20] ));
 sg13g2_nand2b_1 _15986_ (.Y(_09251_),
    .B(net812),
    .A_N(_09250_));
 sg13g2_a21oi_1 _15987_ (.A1(\cpu.icache.r_data[6][20] ),
    .A2(net635),
    .Y(_09252_),
    .B1(net936));
 sg13g2_and4_1 _15988_ (.A(_09248_),
    .B(_09249_),
    .C(_09251_),
    .D(_09252_),
    .X(_09253_));
 sg13g2_o21ai_1 _15989_ (.B1(_09253_),
    .Y(_09254_),
    .A1(_00220_),
    .A2(net452));
 sg13g2_o21ai_1 _15990_ (.B1(_09254_),
    .Y(_09255_),
    .A1(_08977_),
    .A2(_09247_));
 sg13g2_buf_1 _15991_ (.A(_09255_),
    .X(_09256_));
 sg13g2_nand3_1 _15992_ (.B(_09150_),
    .C(_09256_),
    .A(net281),
    .Y(_09257_));
 sg13g2_buf_1 _15993_ (.A(_09257_),
    .X(_09258_));
 sg13g2_nor2_1 _15994_ (.A(net210),
    .B(_09258_),
    .Y(_09259_));
 sg13g2_nand4_1 _15995_ (.B(_09202_),
    .C(_09241_),
    .A(_09198_),
    .Y(_09260_),
    .D(_09259_));
 sg13g2_o21ai_1 _15996_ (.B1(_09260_),
    .Y(_09261_),
    .A1(_09205_),
    .A2(_09206_));
 sg13g2_buf_1 _15997_ (.A(\cpu.dec.r_op[3] ),
    .X(_09262_));
 sg13g2_buf_1 _15998_ (.A(net1125),
    .X(_09263_));
 sg13g2_buf_2 _15999_ (.A(net108),
    .X(_09264_));
 sg13g2_mux2_1 _16000_ (.A0(_09261_),
    .A1(net1057),
    .S(net91),
    .X(_00014_));
 sg13g2_buf_1 _16001_ (.A(\cpu.spi.r_count[7] ),
    .X(_09265_));
 sg13g2_buf_1 _16002_ (.A(\cpu.spi.r_count[3] ),
    .X(_09266_));
 sg13g2_buf_1 _16003_ (.A(\cpu.spi.r_count[0] ),
    .X(_09267_));
 sg13g2_buf_1 _16004_ (.A(\cpu.spi.r_count[1] ),
    .X(_09268_));
 sg13g2_nor2_1 _16005_ (.A(_09267_),
    .B(_09268_),
    .Y(_09269_));
 sg13g2_nand2b_1 _16006_ (.Y(_09270_),
    .B(_09269_),
    .A_N(\cpu.spi.r_count[2] ));
 sg13g2_nor3_1 _16007_ (.A(_09266_),
    .B(\cpu.spi.r_count[4] ),
    .C(_09270_),
    .Y(_09271_));
 sg13g2_nor2b_1 _16008_ (.A(\cpu.spi.r_count[5] ),
    .B_N(_09271_),
    .Y(_09272_));
 sg13g2_nor2b_1 _16009_ (.A(\cpu.spi.r_count[6] ),
    .B_N(_09272_),
    .Y(_09273_));
 sg13g2_nand2b_1 _16010_ (.Y(_09274_),
    .B(_09273_),
    .A_N(_09265_));
 sg13g2_buf_1 _16011_ (.A(_09274_),
    .X(_09275_));
 sg13g2_buf_1 _16012_ (.A(net497),
    .X(_09276_));
 sg13g2_buf_2 _16013_ (.A(\cpu.addr[6] ),
    .X(_09277_));
 sg13g2_buf_1 _16014_ (.A(\cpu.addr[8] ),
    .X(_09278_));
 sg13g2_buf_1 _16015_ (.A(_09278_),
    .X(_09279_));
 sg13g2_buf_2 _16016_ (.A(\cpu.addr[7] ),
    .X(_09280_));
 sg13g2_nor2b_1 _16017_ (.A(net1056),
    .B_N(_09280_),
    .Y(_09281_));
 sg13g2_nand2_1 _16018_ (.Y(_09282_),
    .A(_09277_),
    .B(_09281_));
 sg13g2_buf_1 _16019_ (.A(_09282_),
    .X(_09283_));
 sg13g2_buf_2 _16020_ (.A(\cpu.dec.r_trap ),
    .X(_09284_));
 sg13g2_buf_1 _16021_ (.A(\cpu.ex.r_ie ),
    .X(_09285_));
 sg13g2_inv_1 _16022_ (.Y(_09286_),
    .A(_09285_));
 sg13g2_buf_2 _16023_ (.A(\cpu.gpio.r_enable_in[0] ),
    .X(_09287_));
 sg13g2_buf_2 _16024_ (.A(ui_in[0]),
    .X(_09288_));
 sg13g2_buf_2 _16025_ (.A(\cpu.gpio.r_enable_in[7] ),
    .X(_09289_));
 sg13g2_buf_2 _16026_ (.A(ui_in[7]),
    .X(_09290_));
 sg13g2_a22oi_1 _16027_ (.Y(_09291_),
    .B1(_09289_),
    .B2(_09290_),
    .A2(_09288_),
    .A1(_09287_));
 sg13g2_buf_1 _16028_ (.A(uio_in[4]),
    .X(_09292_));
 sg13g2_buf_2 _16029_ (.A(\cpu.gpio.r_enable_io[7] ),
    .X(_09293_));
 sg13g2_buf_2 _16030_ (.A(uio_in[7]),
    .X(_09294_));
 sg13g2_a22oi_1 _16031_ (.Y(_09295_),
    .B1(_09293_),
    .B2(_09294_),
    .A2(_09292_),
    .A1(\cpu.gpio.r_enable_io[4] ));
 sg13g2_buf_1 _16032_ (.A(\cpu.gpio.r_enable_in[3] ),
    .X(_09296_));
 sg13g2_buf_8 _16033_ (.A(ui_in[3]),
    .X(_09297_));
 sg13g2_buf_1 _16034_ (.A(\cpu.gpio.r_enable_in[6] ),
    .X(_09298_));
 sg13g2_buf_2 _16035_ (.A(ui_in[6]),
    .X(_09299_));
 sg13g2_a22oi_1 _16036_ (.Y(_09300_),
    .B1(_09298_),
    .B2(_09299_),
    .A2(_09297_),
    .A1(_09296_));
 sg13g2_buf_1 _16037_ (.A(\cpu.gpio.r_enable_in[1] ),
    .X(_09301_));
 sg13g2_buf_8 _16038_ (.A(ui_in[1]),
    .X(_09302_));
 sg13g2_buf_1 _16039_ (.A(\cpu.gpio.r_enable_in[4] ),
    .X(_09303_));
 sg13g2_buf_2 _16040_ (.A(ui_in[4]),
    .X(_09304_));
 sg13g2_a22oi_1 _16041_ (.Y(_09305_),
    .B1(_09303_),
    .B2(_09304_),
    .A2(_09302_),
    .A1(_09301_));
 sg13g2_and4_1 _16042_ (.A(_09291_),
    .B(_09295_),
    .C(_09300_),
    .D(_09305_),
    .X(_09306_));
 sg13g2_buf_1 _16043_ (.A(\cpu.gpio.r_enable_in[2] ),
    .X(_09307_));
 sg13g2_buf_2 _16044_ (.A(ui_in[2]),
    .X(_09308_));
 sg13g2_buf_1 _16045_ (.A(\cpu.gpio.r_enable_in[5] ),
    .X(_09309_));
 sg13g2_buf_2 _16046_ (.A(ui_in[5]),
    .X(_09310_));
 sg13g2_a22oi_1 _16047_ (.Y(_09311_),
    .B1(_09309_),
    .B2(_09310_),
    .A2(_09308_),
    .A1(_09307_));
 sg13g2_buf_1 _16048_ (.A(\cpu.gpio.r_enable_io[5] ),
    .X(_09312_));
 sg13g2_buf_2 _16049_ (.A(uio_in[5]),
    .X(_09313_));
 sg13g2_buf_1 _16050_ (.A(\cpu.gpio.r_enable_io[6] ),
    .X(_09314_));
 sg13g2_buf_1 _16051_ (.A(uio_in[6]),
    .X(_09315_));
 sg13g2_a22oi_1 _16052_ (.Y(_09316_),
    .B1(_09314_),
    .B2(_09315_),
    .A2(_09313_),
    .A1(_09312_));
 sg13g2_and2_1 _16053_ (.A(_09311_),
    .B(_09316_),
    .X(_09317_));
 sg13g2_buf_2 _16054_ (.A(\cpu.intr.r_enable[4] ),
    .X(_09318_));
 sg13g2_inv_1 _16055_ (.Y(_09319_),
    .A(_09318_));
 sg13g2_a21oi_2 _16056_ (.B1(_09319_),
    .Y(_09320_),
    .A2(_09317_),
    .A1(_09306_));
 sg13g2_buf_1 _16057_ (.A(\cpu.intr.r_timer ),
    .X(_09321_));
 sg13g2_buf_1 _16058_ (.A(\cpu.intr.spi_intr ),
    .X(_09322_));
 sg13g2_buf_1 _16059_ (.A(\cpu.intr.r_enable[5] ),
    .X(_09323_));
 sg13g2_a22oi_1 _16060_ (.Y(_09324_),
    .B1(_09322_),
    .B2(_09323_),
    .A2(\cpu.intr.r_enable[2] ),
    .A1(_09321_));
 sg13g2_buf_1 _16061_ (.A(\cpu.intr.r_enable[1] ),
    .X(_09325_));
 sg13g2_buf_1 _16062_ (.A(\cpu.intr.r_swi ),
    .X(_09326_));
 sg13g2_a22oi_1 _16063_ (.Y(_09327_),
    .B1(\cpu.intr.r_enable[3] ),
    .B2(_09326_),
    .A2(_09325_),
    .A1(\cpu.intr.r_clock ));
 sg13g2_buf_2 _16064_ (.A(\cpu.uart.r_x_int ),
    .X(_09328_));
 sg13g2_buf_2 _16065_ (.A(\cpu.uart.r_r_int ),
    .X(_09329_));
 sg13g2_o21ai_1 _16066_ (.B1(\cpu.intr.r_enable[0] ),
    .Y(_09330_),
    .A1(_09328_),
    .A2(_09329_));
 sg13g2_nand3_1 _16067_ (.B(_09327_),
    .C(_09330_),
    .A(_09324_),
    .Y(_09331_));
 sg13g2_buf_2 _16068_ (.A(_09331_),
    .X(_09332_));
 sg13g2_nor2_1 _16069_ (.A(_09320_),
    .B(_09332_),
    .Y(_09333_));
 sg13g2_nor2_1 _16070_ (.A(_09286_),
    .B(_09333_),
    .Y(_09334_));
 sg13g2_and2_1 _16071_ (.A(_08452_),
    .B(_09334_),
    .X(_09335_));
 sg13g2_nor4_1 _16072_ (.A(_09284_),
    .B(_08431_),
    .C(_08525_),
    .D(_09335_),
    .Y(_09336_));
 sg13g2_buf_2 _16073_ (.A(_09336_),
    .X(_09337_));
 sg13g2_buf_2 _16074_ (.A(\cpu.addr[3] ),
    .X(_09338_));
 sg13g2_buf_1 _16075_ (.A(_09338_),
    .X(_09339_));
 sg13g2_buf_1 _16076_ (.A(net1055),
    .X(_09340_));
 sg13g2_buf_1 _16077_ (.A(_09340_),
    .X(_09341_));
 sg13g2_buf_1 _16078_ (.A(net807),
    .X(_09342_));
 sg13g2_buf_1 _16079_ (.A(net708),
    .X(_09343_));
 sg13g2_buf_2 _16080_ (.A(net633),
    .X(_09344_));
 sg13g2_buf_2 _16081_ (.A(net551),
    .X(_09345_));
 sg13g2_buf_2 _16082_ (.A(\cpu.addr[2] ),
    .X(_09346_));
 sg13g2_buf_8 _16083_ (.A(_09346_),
    .X(_09347_));
 sg13g2_inv_2 _16084_ (.Y(_09348_),
    .A(net1054));
 sg13g2_buf_1 _16085_ (.A(_09348_),
    .X(_09349_));
 sg13g2_buf_1 _16086_ (.A(\cpu.addr[1] ),
    .X(_09350_));
 sg13g2_inv_2 _16087_ (.Y(_09351_),
    .A(_09350_));
 sg13g2_buf_1 _16088_ (.A(_09351_),
    .X(_09352_));
 sg13g2_nand2_1 _16089_ (.Y(_09353_),
    .A(net806),
    .B(net933));
 sg13g2_nor3_1 _16090_ (.A(_00197_),
    .B(net496),
    .C(_09353_),
    .Y(_09354_));
 sg13g2_nand2_1 _16091_ (.Y(_09355_),
    .A(_09337_),
    .B(_09354_));
 sg13g2_inv_1 _16092_ (.Y(_09356_),
    .A(_08500_));
 sg13g2_buf_1 _16093_ (.A(_08432_),
    .X(_09357_));
 sg13g2_buf_1 _16094_ (.A(_08498_),
    .X(_09358_));
 sg13g2_nor2_1 _16095_ (.A(_09358_),
    .B(_08500_),
    .Y(_09359_));
 sg13g2_a21oi_1 _16096_ (.A1(net1052),
    .A2(net1053),
    .Y(_09360_),
    .B1(_09359_));
 sg13g2_nand2_1 _16097_ (.Y(_09361_),
    .A(_08499_),
    .B(_09360_));
 sg13g2_o21ai_1 _16098_ (.B1(_09361_),
    .Y(_09362_),
    .A1(_09356_),
    .A2(net1053));
 sg13g2_buf_2 _16099_ (.A(_09362_),
    .X(_09363_));
 sg13g2_nor3_2 _16100_ (.A(_09283_),
    .B(_09355_),
    .C(_09363_),
    .Y(_09364_));
 sg13g2_buf_1 _16101_ (.A(\cpu.spi.r_state[1] ),
    .X(_09365_));
 sg13g2_inv_1 _16102_ (.Y(_09366_),
    .A(net1124));
 sg13g2_nand3b_1 _16103_ (.B(_09337_),
    .C(_08393_),
    .Y(_09367_),
    .A_N(net957));
 sg13g2_buf_2 _16104_ (.A(_09367_),
    .X(_09368_));
 sg13g2_or2_1 _16105_ (.X(_09369_),
    .B(_09368_),
    .A(net709));
 sg13g2_buf_1 _16106_ (.A(_09369_),
    .X(_09370_));
 sg13g2_nor2_1 _16107_ (.A(net496),
    .B(_09370_),
    .Y(_09371_));
 sg13g2_buf_1 _16108_ (.A(_09371_),
    .X(_09372_));
 sg13g2_nor2_1 _16109_ (.A(_09366_),
    .B(_09372_),
    .Y(_09373_));
 sg13g2_buf_1 _16110_ (.A(_09373_),
    .X(_09374_));
 sg13g2_buf_1 _16111_ (.A(\cpu.spi.r_state[3] ),
    .X(_09375_));
 sg13g2_a21oi_1 _16112_ (.A1(_09364_),
    .A2(_09374_),
    .Y(_09376_),
    .B1(_09375_));
 sg13g2_buf_2 _16113_ (.A(\cpu.spi.r_state[0] ),
    .X(_09377_));
 sg13g2_buf_1 _16114_ (.A(net1054),
    .X(_09378_));
 sg13g2_buf_1 _16115_ (.A(net932),
    .X(_09379_));
 sg13g2_buf_1 _16116_ (.A(_09350_),
    .X(_09380_));
 sg13g2_nor2_1 _16117_ (.A(net805),
    .B(net1051),
    .Y(_09381_));
 sg13g2_buf_1 _16118_ (.A(_09381_),
    .X(_09382_));
 sg13g2_nand2_1 _16119_ (.Y(_09383_),
    .A(net632),
    .B(_09372_));
 sg13g2_nand2b_1 _16120_ (.Y(_09384_),
    .B(net1),
    .A_N(r_reset));
 sg13g2_buf_2 _16121_ (.A(_09384_),
    .X(_09385_));
 sg13g2_buf_1 _16122_ (.A(_09385_),
    .X(_09386_));
 sg13g2_a21oi_1 _16123_ (.A1(_09377_),
    .A2(_09383_),
    .Y(_09387_),
    .B1(net931));
 sg13g2_o21ai_1 _16124_ (.B1(_09387_),
    .Y(_00029_),
    .A1(net447),
    .A2(_09376_));
 sg13g2_buf_2 _16125_ (.A(_09386_),
    .X(_09388_));
 sg13g2_buf_1 _16126_ (.A(net804),
    .X(_09389_));
 sg13g2_buf_1 _16127_ (.A(net707),
    .X(_09390_));
 sg13g2_inv_1 _16128_ (.Y(_09391_),
    .A(_09364_));
 sg13g2_nor2b_1 _16129_ (.A(_09265_),
    .B_N(_09273_),
    .Y(_09392_));
 sg13g2_buf_1 _16130_ (.A(_09392_),
    .X(_09393_));
 sg13g2_buf_1 _16131_ (.A(_09393_),
    .X(_09394_));
 sg13g2_buf_1 _16132_ (.A(\cpu.spi.r_bits[0] ),
    .X(_09395_));
 sg13g2_buf_1 _16133_ (.A(\cpu.spi.r_bits[1] ),
    .X(_09396_));
 sg13g2_nor3_1 _16134_ (.A(_09395_),
    .B(_09396_),
    .C(\cpu.spi.r_bits[2] ),
    .Y(_09397_));
 sg13g2_buf_1 _16135_ (.A(\cpu.spi.r_timeout_count[7] ),
    .X(_09398_));
 sg13g2_buf_1 _16136_ (.A(\cpu.spi.r_timeout_count[0] ),
    .X(_09399_));
 sg13g2_buf_1 _16137_ (.A(\cpu.spi.r_timeout_count[1] ),
    .X(_09400_));
 sg13g2_or3_1 _16138_ (.A(_09399_),
    .B(_09400_),
    .C(\cpu.spi.r_timeout_count[2] ),
    .X(_09401_));
 sg13g2_buf_1 _16139_ (.A(_09401_),
    .X(_09402_));
 sg13g2_or2_1 _16140_ (.X(_09403_),
    .B(_09402_),
    .A(\cpu.spi.r_timeout_count[3] ));
 sg13g2_buf_1 _16141_ (.A(_09403_),
    .X(_09404_));
 sg13g2_or2_1 _16142_ (.X(_09405_),
    .B(_09404_),
    .A(\cpu.spi.r_timeout_count[4] ));
 sg13g2_buf_1 _16143_ (.A(_09405_),
    .X(_09406_));
 sg13g2_or2_1 _16144_ (.X(_09407_),
    .B(_09406_),
    .A(\cpu.spi.r_timeout_count[5] ));
 sg13g2_buf_1 _16145_ (.A(_09407_),
    .X(_09408_));
 sg13g2_or2_1 _16146_ (.X(_09409_),
    .B(_09408_),
    .A(\cpu.spi.r_timeout_count[6] ));
 sg13g2_buf_1 _16147_ (.A(_09409_),
    .X(_09410_));
 sg13g2_buf_1 _16148_ (.A(\cpu.spi.r_searching ),
    .X(_09411_));
 sg13g2_o21ai_1 _16149_ (.B1(_09411_),
    .Y(_09412_),
    .A1(_09398_),
    .A2(_09410_));
 sg13g2_nand2_1 _16150_ (.Y(_09413_),
    .A(_09397_),
    .B(_09412_));
 sg13g2_buf_1 _16151_ (.A(\cpu.spi.r_in[3] ),
    .X(_09414_));
 sg13g2_buf_1 _16152_ (.A(\cpu.spi.r_in[6] ),
    .X(_09415_));
 sg13g2_buf_1 _16153_ (.A(\cpu.spi.r_in[1] ),
    .X(_09416_));
 sg13g2_buf_1 _16154_ (.A(\cpu.spi.r_in[0] ),
    .X(_09417_));
 sg13g2_nand2_1 _16155_ (.Y(_09418_),
    .A(_09416_),
    .B(_09417_));
 sg13g2_nand3_1 _16156_ (.B(_09415_),
    .C(_09418_),
    .A(_09414_),
    .Y(_09419_));
 sg13g2_buf_1 _16157_ (.A(\cpu.spi.r_in[2] ),
    .X(_09420_));
 sg13g2_buf_1 _16158_ (.A(\cpu.spi.r_in[5] ),
    .X(_09421_));
 sg13g2_buf_1 _16159_ (.A(\cpu.spi.r_in[4] ),
    .X(_09422_));
 sg13g2_nand4_1 _16160_ (.B(_09421_),
    .C(_09422_),
    .A(_09420_),
    .Y(_09423_),
    .D(\cpu.spi.r_in[7] ));
 sg13g2_nor2_1 _16161_ (.A(_09419_),
    .B(_09423_),
    .Y(_09424_));
 sg13g2_o21ai_1 _16162_ (.B1(_09411_),
    .Y(_09425_),
    .A1(_00222_),
    .A2(_09424_));
 sg13g2_nand2_1 _16163_ (.Y(_09426_),
    .A(_09413_),
    .B(_09425_));
 sg13g2_nand2_1 _16164_ (.Y(_09427_),
    .A(net446),
    .B(_09426_));
 sg13g2_inv_1 _16165_ (.Y(_09428_),
    .A(_09427_));
 sg13g2_buf_1 _16166_ (.A(\cpu.spi.r_state[6] ),
    .X(_09429_));
 sg13g2_buf_1 _16167_ (.A(_09429_),
    .X(_09430_));
 sg13g2_a22oi_1 _16168_ (.Y(_09431_),
    .B1(_09428_),
    .B2(net1050),
    .A2(_09374_),
    .A1(_09391_));
 sg13g2_nor2_1 _16169_ (.A(net631),
    .B(_09431_),
    .Y(_00030_));
 sg13g2_buf_1 _16170_ (.A(net1124),
    .X(_09432_));
 sg13g2_buf_1 _16171_ (.A(_09372_),
    .X(_09433_));
 sg13g2_buf_1 _16172_ (.A(net107),
    .X(_09434_));
 sg13g2_a21oi_1 _16173_ (.A1(net1049),
    .A2(_09434_),
    .Y(_09435_),
    .B1(\cpu.spi.r_state[5] ));
 sg13g2_buf_2 _16174_ (.A(\cpu.spi.r_state[4] ),
    .X(_09436_));
 sg13g2_inv_1 _16175_ (.Y(_09437_),
    .A(_09429_));
 sg13g2_nor2_1 _16176_ (.A(_09437_),
    .B(_09426_),
    .Y(_09438_));
 sg13g2_nor3_1 _16177_ (.A(_09436_),
    .B(net447),
    .C(_09438_),
    .Y(_09439_));
 sg13g2_buf_1 _16178_ (.A(\cpu.spi.r_state[2] ),
    .X(_09440_));
 sg13g2_nor2b_1 _16179_ (.A(r_reset),
    .B_N(net1),
    .Y(_09441_));
 sg13g2_buf_1 _16180_ (.A(_09441_),
    .X(_09442_));
 sg13g2_buf_2 _16181_ (.A(_09442_),
    .X(_09443_));
 sg13g2_buf_2 _16182_ (.A(net930),
    .X(_09444_));
 sg13g2_buf_2 _16183_ (.A(net803),
    .X(_09445_));
 sg13g2_o21ai_1 _16184_ (.B1(net706),
    .Y(_09446_),
    .A1(net1123),
    .A2(net446));
 sg13g2_a21oi_1 _16185_ (.A1(_09435_),
    .A2(_09439_),
    .Y(_00031_),
    .B1(_09446_));
 sg13g2_buf_1 _16186_ (.A(net804),
    .X(_09447_));
 sg13g2_nor3_1 _16187_ (.A(net705),
    .B(_09394_),
    .C(_09376_),
    .Y(_00032_));
 sg13g2_inv_1 _16188_ (.Y(_09448_),
    .A(_09383_));
 sg13g2_a22oi_1 _16189_ (.Y(_09449_),
    .B1(_09276_),
    .B2(_09436_),
    .A2(_09448_),
    .A1(_09377_));
 sg13g2_nor2_1 _16190_ (.A(net631),
    .B(_09449_),
    .Y(_00033_));
 sg13g2_nor3_1 _16191_ (.A(net705),
    .B(net446),
    .C(_09435_),
    .Y(_00034_));
 sg13g2_nand2_1 _16192_ (.Y(_09450_),
    .A(net1050),
    .B(net447));
 sg13g2_nand2_1 _16193_ (.Y(_09451_),
    .A(net1123),
    .B(net446));
 sg13g2_buf_1 _16194_ (.A(net804),
    .X(_09452_));
 sg13g2_buf_1 _16195_ (.A(_09452_),
    .X(_09453_));
 sg13g2_a21oi_1 _16196_ (.A1(_09450_),
    .A2(_09451_),
    .Y(_00035_),
    .B1(_09453_));
 sg13g2_buf_2 _16197_ (.A(\cpu.ex.r_mult_off[0] ),
    .X(_09454_));
 sg13g2_buf_1 _16198_ (.A(\cpu.dec.mult ),
    .X(_09455_));
 sg13g2_nand3b_1 _16199_ (.B(\cpu.dec.iready ),
    .C(_00199_),
    .Y(_09456_),
    .A_N(\cpu.ex.r_branch_stall ));
 sg13g2_buf_2 _16200_ (.A(_09456_),
    .X(_09457_));
 sg13g2_nor2_1 _16201_ (.A(_09385_),
    .B(_09457_),
    .Y(_09458_));
 sg13g2_buf_2 _16202_ (.A(_09458_),
    .X(_09459_));
 sg13g2_and2_1 _16203_ (.A(_09455_),
    .B(_09459_),
    .X(_09460_));
 sg13g2_buf_1 _16204_ (.A(_09460_),
    .X(_09461_));
 sg13g2_and2_1 _16205_ (.A(\cpu.dec.div ),
    .B(_09459_),
    .X(_09462_));
 sg13g2_buf_2 _16206_ (.A(_09462_),
    .X(_09463_));
 sg13g2_nor2_1 _16207_ (.A(net629),
    .B(_09463_),
    .Y(_09464_));
 sg13g2_buf_1 _16208_ (.A(_09464_),
    .X(_09465_));
 sg13g2_nand2_2 _16209_ (.Y(\cpu.ex.c_mult_off[0] ),
    .A(_09454_),
    .B(net495));
 sg13g2_buf_1 _16210_ (.A(\cpu.ex.r_div_running ),
    .X(_09466_));
 sg13g2_buf_2 _16211_ (.A(\cpu.ex.r_mult_off[1] ),
    .X(_09467_));
 sg13g2_buf_1 _16212_ (.A(\cpu.ex.r_mult_off[2] ),
    .X(_09468_));
 sg13g2_nor2_2 _16213_ (.A(_09454_),
    .B(_09467_),
    .Y(_09469_));
 sg13g2_nand2b_1 _16214_ (.Y(_09470_),
    .B(_09469_),
    .A_N(_09468_));
 sg13g2_xor2_1 _16215_ (.B(_09470_),
    .A(\cpu.ex.r_mult_off[3] ),
    .X(_09471_));
 sg13g2_nand2_1 _16216_ (.Y(_09472_),
    .A(net495),
    .B(_09471_));
 sg13g2_buf_1 _16217_ (.A(_09472_),
    .X(\cpu.ex.c_mult_off[3] ));
 sg13g2_nor4_2 _16218_ (.A(_09467_),
    .B(_09468_),
    .C(\cpu.ex.c_mult_off[0] ),
    .Y(_09473_),
    .D(\cpu.ex.c_mult_off[3] ));
 sg13g2_buf_1 _16219_ (.A(_09463_),
    .X(_09474_));
 sg13g2_o21ai_1 _16220_ (.B1(_09442_),
    .Y(_09475_),
    .A1(_09466_),
    .A2(_09474_));
 sg13g2_a21oi_1 _16221_ (.A1(_09466_),
    .A2(_09473_),
    .Y(\cpu.ex.c_div_running ),
    .B1(_09475_));
 sg13g2_buf_1 _16222_ (.A(\cpu.ex.r_mult_running ),
    .X(_09476_));
 sg13g2_inv_1 _16223_ (.Y(_09477_),
    .A(net1122));
 sg13g2_nand2_1 _16224_ (.Y(_09478_),
    .A(_09455_),
    .B(_09459_));
 sg13g2_buf_1 _16225_ (.A(_09478_),
    .X(_09479_));
 sg13g2_nand2_1 _16226_ (.Y(_09480_),
    .A(_09477_),
    .B(net628));
 sg13g2_buf_1 _16227_ (.A(_09480_),
    .X(_09481_));
 sg13g2_nand2_1 _16228_ (.Y(_09482_),
    .A(_09442_),
    .B(_09481_));
 sg13g2_a21oi_1 _16229_ (.A1(net1122),
    .A2(_09473_),
    .Y(\cpu.ex.c_mult_running ),
    .B1(_09482_));
 sg13g2_inv_1 _16230_ (.Y(_09483_),
    .A(\cpu.qspi.r_state[17] ));
 sg13g2_inv_1 _16231_ (.Y(_09484_),
    .A(net1069));
 sg13g2_buf_1 _16232_ (.A(_09484_),
    .X(_09485_));
 sg13g2_buf_1 _16233_ (.A(\cpu.dcache.flush_write ),
    .X(_09486_));
 sg13g2_inv_1 _16234_ (.Y(_09487_),
    .A(_09486_));
 sg13g2_mux4_1 _16235_ (.S0(net805),
    .A0(\cpu.dcache.r_valid[4] ),
    .A1(\cpu.dcache.r_valid[5] ),
    .A2(\cpu.dcache.r_valid[6] ),
    .A3(\cpu.dcache.r_valid[7] ),
    .S1(net708),
    .X(_09488_));
 sg13g2_mux4_1 _16236_ (.S0(net805),
    .A0(\cpu.dcache.r_valid[0] ),
    .A1(\cpu.dcache.r_valid[1] ),
    .A2(\cpu.dcache.r_valid[2] ),
    .A3(\cpu.dcache.r_valid[3] ),
    .S1(net807),
    .X(_09489_));
 sg13g2_buf_2 _16237_ (.A(\cpu.addr[4] ),
    .X(_09490_));
 sg13g2_inv_4 _16238_ (.A(net1121),
    .Y(_09491_));
 sg13g2_mux2_1 _16239_ (.A0(_09488_),
    .A1(_09489_),
    .S(_09491_),
    .X(_09492_));
 sg13g2_mux4_1 _16240_ (.S0(net805),
    .A0(\cpu.dcache.r_dirty[4] ),
    .A1(\cpu.dcache.r_dirty[5] ),
    .A2(\cpu.dcache.r_dirty[6] ),
    .A3(\cpu.dcache.r_dirty[7] ),
    .S1(_09342_),
    .X(_09493_));
 sg13g2_mux4_1 _16241_ (.S0(net805),
    .A0(\cpu.dcache.r_dirty[0] ),
    .A1(\cpu.dcache.r_dirty[1] ),
    .A2(\cpu.dcache.r_dirty[2] ),
    .A3(\cpu.dcache.r_dirty[3] ),
    .S1(_09342_),
    .X(_09494_));
 sg13g2_buf_1 _16242_ (.A(_09491_),
    .X(_09495_));
 sg13g2_mux2_1 _16243_ (.A0(_09493_),
    .A1(_09494_),
    .S(net929),
    .X(_09496_));
 sg13g2_nand3_1 _16244_ (.B(_09492_),
    .C(_09496_),
    .A(_09337_),
    .Y(_09497_));
 sg13g2_buf_1 _16245_ (.A(_09497_),
    .X(_09498_));
 sg13g2_and2_1 _16246_ (.A(_09487_),
    .B(_09498_),
    .X(_09499_));
 sg13g2_buf_2 _16247_ (.A(_00227_),
    .X(_09500_));
 sg13g2_and3_1 _16248_ (.X(_09501_),
    .A(net1054),
    .B(_09339_),
    .C(_09500_));
 sg13g2_buf_2 _16249_ (.A(_09501_),
    .X(_09502_));
 sg13g2_buf_1 _16250_ (.A(_09502_),
    .X(_09503_));
 sg13g2_buf_1 _16251_ (.A(net704),
    .X(_09504_));
 sg13g2_nand2b_1 _16252_ (.Y(_09505_),
    .B(net1121),
    .A_N(net1054));
 sg13g2_nor2_1 _16253_ (.A(net934),
    .B(_09505_),
    .Y(_09506_));
 sg13g2_buf_1 _16254_ (.A(_09506_),
    .X(_09507_));
 sg13g2_buf_1 _16255_ (.A(net703),
    .X(_09508_));
 sg13g2_a22oi_1 _16256_ (.Y(_09509_),
    .B1(net626),
    .B2(\cpu.dcache.r_tag[4][14] ),
    .A2(_09504_),
    .A1(\cpu.dcache.r_tag[3][14] ));
 sg13g2_nor3_2 _16257_ (.A(_09348_),
    .B(_09491_),
    .C(net934),
    .Y(_09510_));
 sg13g2_buf_1 _16258_ (.A(_09510_),
    .X(_09511_));
 sg13g2_nand2_1 _16259_ (.Y(_09512_),
    .A(\cpu.dcache.r_tag[5][14] ),
    .B(net702));
 sg13g2_nor2b_1 _16260_ (.A(_09346_),
    .B_N(_09338_),
    .Y(_09513_));
 sg13g2_buf_1 _16261_ (.A(_09513_),
    .X(_09514_));
 sg13g2_and2_1 _16262_ (.A(_09500_),
    .B(net928),
    .X(_09515_));
 sg13g2_buf_2 _16263_ (.A(_09515_),
    .X(_09516_));
 sg13g2_buf_1 _16264_ (.A(_09516_),
    .X(_09517_));
 sg13g2_buf_1 _16265_ (.A(net625),
    .X(_09518_));
 sg13g2_inv_1 _16266_ (.Y(_09519_),
    .A(net1055));
 sg13g2_nor2_1 _16267_ (.A(_09519_),
    .B(_09505_),
    .Y(_09520_));
 sg13g2_buf_1 _16268_ (.A(_09520_),
    .X(_09521_));
 sg13g2_a22oi_1 _16269_ (.Y(_09522_),
    .B1(net701),
    .B2(\cpu.dcache.r_tag[6][14] ),
    .A2(_09518_),
    .A1(\cpu.dcache.r_tag[2][14] ));
 sg13g2_nor2b_1 _16270_ (.A(net1055),
    .B_N(_09500_),
    .Y(_09523_));
 sg13g2_and2_1 _16271_ (.A(net932),
    .B(_09523_),
    .X(_09524_));
 sg13g2_buf_1 _16272_ (.A(_09524_),
    .X(_09525_));
 sg13g2_buf_1 _16273_ (.A(net700),
    .X(_09526_));
 sg13g2_nand2_1 _16274_ (.Y(_09527_),
    .A(_09347_),
    .B(net1055));
 sg13g2_nor2_1 _16275_ (.A(_09491_),
    .B(_09527_),
    .Y(_09528_));
 sg13g2_buf_1 _16276_ (.A(_09528_),
    .X(_09529_));
 sg13g2_nand3b_1 _16277_ (.B(_09500_),
    .C(net1054),
    .Y(_09530_),
    .A_N(net1055));
 sg13g2_buf_1 _16278_ (.A(_09530_),
    .X(_09531_));
 sg13g2_nor2_1 _16279_ (.A(net1121),
    .B(net1055),
    .Y(_09532_));
 sg13g2_buf_2 _16280_ (.A(_09532_),
    .X(_09533_));
 sg13g2_nand2_1 _16281_ (.Y(_09534_),
    .A(_09531_),
    .B(_09533_));
 sg13g2_buf_1 _16282_ (.A(_09534_),
    .X(_09535_));
 sg13g2_nor2_1 _16283_ (.A(_00245_),
    .B(net623),
    .Y(_09536_));
 sg13g2_a221oi_1 _16284_ (.B2(\cpu.dcache.r_tag[7][14] ),
    .C1(_09536_),
    .B1(net699),
    .A1(\cpu.dcache.r_tag[1][14] ),
    .Y(_09537_),
    .A2(_09526_));
 sg13g2_nand4_1 _16285_ (.B(_09512_),
    .C(_09522_),
    .A(_09509_),
    .Y(_09538_),
    .D(_09537_));
 sg13g2_buf_1 _16286_ (.A(net956),
    .X(_09539_));
 sg13g2_buf_2 _16287_ (.A(net801),
    .X(_09540_));
 sg13g2_buf_1 _16288_ (.A(net698),
    .X(_09541_));
 sg13g2_buf_8 _16289_ (.A(net1073),
    .X(_09542_));
 sg13g2_buf_8 _16290_ (.A(net927),
    .X(_09543_));
 sg13g2_buf_8 _16291_ (.A(_09543_),
    .X(_09544_));
 sg13g2_buf_2 _16292_ (.A(net1072),
    .X(_09545_));
 sg13g2_buf_2 _16293_ (.A(_09545_),
    .X(_09546_));
 sg13g2_mux4_1 _16294_ (.S0(net697),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][2] ),
    .S1(net800),
    .X(_09547_));
 sg13g2_mux4_1 _16295_ (.S0(_09544_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][2] ),
    .S1(net800),
    .X(_09548_));
 sg13g2_buf_8 _16296_ (.A(_09543_),
    .X(_09549_));
 sg13g2_buf_2 _16297_ (.A(_09545_),
    .X(_09550_));
 sg13g2_mux4_1 _16298_ (.S0(net696),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][2] ),
    .S1(net799),
    .X(_09551_));
 sg13g2_buf_2 _16299_ (.A(_09545_),
    .X(_09552_));
 sg13g2_mux4_1 _16300_ (.S0(_09549_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][2] ),
    .S1(net798),
    .X(_09553_));
 sg13g2_mux4_1 _16301_ (.S0(_08497_),
    .A0(_09547_),
    .A1(_09548_),
    .A2(_09551_),
    .A3(_09553_),
    .S1(_08377_),
    .X(_09554_));
 sg13g2_nand2_1 _16302_ (.Y(_09555_),
    .A(net1068),
    .B(_09554_));
 sg13g2_buf_8 _16303_ (.A(_09543_),
    .X(_09556_));
 sg13g2_buf_2 _16304_ (.A(_09545_),
    .X(_09557_));
 sg13g2_mux4_1 _16305_ (.S0(net695),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][2] ),
    .S1(net797),
    .X(_09558_));
 sg13g2_mux4_1 _16306_ (.S0(net695),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][2] ),
    .S1(_09557_),
    .X(_09559_));
 sg13g2_mux4_1 _16307_ (.S0(net697),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][2] ),
    .S1(net800),
    .X(_09560_));
 sg13g2_mux4_1 _16308_ (.S0(net697),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][2] ),
    .S1(_09546_),
    .X(_09561_));
 sg13g2_mux4_1 _16309_ (.S0(_08497_),
    .A0(_09558_),
    .A1(_09559_),
    .A2(_09560_),
    .A3(_09561_),
    .S1(net1075),
    .X(_09562_));
 sg13g2_o21ai_1 _16310_ (.B1(net622),
    .Y(_09563_),
    .A1(_08695_),
    .A2(_09562_));
 sg13g2_o21ai_1 _16311_ (.B1(_09563_),
    .Y(_09564_),
    .A1(net622),
    .A2(_09555_));
 sg13g2_buf_1 _16312_ (.A(_09564_),
    .X(_09565_));
 sg13g2_xnor2_1 _16313_ (.Y(_09566_),
    .A(_09538_),
    .B(net409));
 sg13g2_nor2_1 _16314_ (.A(_08388_),
    .B(_08398_),
    .Y(_09567_));
 sg13g2_buf_1 _16315_ (.A(_09567_),
    .X(_09568_));
 sg13g2_buf_8 _16316_ (.A(_09543_),
    .X(_09569_));
 sg13g2_buf_2 _16317_ (.A(_09545_),
    .X(_09570_));
 sg13g2_mux4_1 _16318_ (.S0(net694),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][5] ),
    .S1(net795),
    .X(_09571_));
 sg13g2_mux4_1 _16319_ (.S0(net694),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][5] ),
    .S1(net797),
    .X(_09572_));
 sg13g2_buf_8 _16320_ (.A(_09543_),
    .X(_09573_));
 sg13g2_mux4_1 _16321_ (.S0(_09573_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][5] ),
    .S1(_09552_),
    .X(_09574_));
 sg13g2_mux4_1 _16322_ (.S0(_09573_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][5] ),
    .S1(net800),
    .X(_09575_));
 sg13g2_buf_1 _16323_ (.A(_08428_),
    .X(_09576_));
 sg13g2_buf_2 _16324_ (.A(net794),
    .X(_09577_));
 sg13g2_mux4_1 _16325_ (.S0(net692),
    .A0(_09571_),
    .A1(_09572_),
    .A2(_09574_),
    .A3(_09575_),
    .S1(net698),
    .X(_09578_));
 sg13g2_nand2_1 _16326_ (.Y(_09579_),
    .A(net796),
    .B(_09578_));
 sg13g2_buf_1 _16327_ (.A(_08497_),
    .X(_09580_));
 sg13g2_mux4_1 _16328_ (.S0(net697),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][5] ),
    .S1(_09546_),
    .X(_09581_));
 sg13g2_mux4_1 _16329_ (.S0(net694),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][5] ),
    .S1(net795),
    .X(_09582_));
 sg13g2_mux4_1 _16330_ (.S0(net693),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][5] ),
    .S1(net798),
    .X(_09583_));
 sg13g2_mux4_1 _16331_ (.S0(net693),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][5] ),
    .S1(_09552_),
    .X(_09584_));
 sg13g2_mux4_1 _16332_ (.S0(_09577_),
    .A0(_09581_),
    .A1(_09582_),
    .A2(_09583_),
    .A3(_09584_),
    .S1(net801),
    .X(_09585_));
 sg13g2_nand2_1 _16333_ (.Y(_09586_),
    .A(net691),
    .B(_09585_));
 sg13g2_a21oi_2 _16334_ (.B1(_08644_),
    .Y(_09587_),
    .A2(_09586_),
    .A1(_09579_));
 sg13g2_buf_1 _16335_ (.A(_09587_),
    .X(_09588_));
 sg13g2_a22oi_1 _16336_ (.Y(_09589_),
    .B1(net701),
    .B2(\cpu.dcache.r_tag[6][17] ),
    .A2(_09511_),
    .A1(\cpu.dcache.r_tag[5][17] ));
 sg13g2_nand2_1 _16337_ (.Y(_09590_),
    .A(\cpu.dcache.r_tag[7][17] ),
    .B(net699));
 sg13g2_a22oi_1 _16338_ (.Y(_09591_),
    .B1(_09518_),
    .B2(\cpu.dcache.r_tag[2][17] ),
    .A2(net626),
    .A1(\cpu.dcache.r_tag[4][17] ));
 sg13g2_nor2_1 _16339_ (.A(_00248_),
    .B(net623),
    .Y(_09592_));
 sg13g2_a221oi_1 _16340_ (.B2(\cpu.dcache.r_tag[3][17] ),
    .C1(_09592_),
    .B1(net704),
    .A1(\cpu.dcache.r_tag[1][17] ),
    .Y(_09593_),
    .A2(net624));
 sg13g2_nand4_1 _16341_ (.B(_09590_),
    .C(_09591_),
    .A(_09589_),
    .Y(_09594_),
    .D(_09593_));
 sg13g2_xnor2_1 _16342_ (.Y(_09595_),
    .A(net408),
    .B(_09594_));
 sg13g2_mux4_1 _16343_ (.S0(_09556_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][11] ),
    .S1(net797),
    .X(_09596_));
 sg13g2_mux4_1 _16344_ (.S0(net695),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][11] ),
    .S1(net797),
    .X(_09597_));
 sg13g2_mux4_1 _16345_ (.S0(net697),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][11] ),
    .S1(net800),
    .X(_09598_));
 sg13g2_mux4_1 _16346_ (.S0(net697),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][11] ),
    .S1(net800),
    .X(_09599_));
 sg13g2_mux4_1 _16347_ (.S0(net692),
    .A0(_09596_),
    .A1(_09597_),
    .A2(_09598_),
    .A3(_09599_),
    .S1(net698),
    .X(_09600_));
 sg13g2_nand2_1 _16348_ (.Y(_09601_),
    .A(net796),
    .B(_09600_));
 sg13g2_mux4_1 _16349_ (.S0(_09569_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][11] ),
    .S1(_09570_),
    .X(_09602_));
 sg13g2_mux4_1 _16350_ (.S0(_09569_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][11] ),
    .S1(_09570_),
    .X(_09603_));
 sg13g2_mux4_1 _16351_ (.S0(net693),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][11] ),
    .S1(net798),
    .X(_09604_));
 sg13g2_mux4_1 _16352_ (.S0(net693),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][11] ),
    .S1(net798),
    .X(_09605_));
 sg13g2_mux4_1 _16353_ (.S0(net692),
    .A0(_09602_),
    .A1(_09603_),
    .A2(_09604_),
    .A3(_09605_),
    .S1(net698),
    .X(_09606_));
 sg13g2_nand2_1 _16354_ (.Y(_09607_),
    .A(net691),
    .B(_09606_));
 sg13g2_a21oi_2 _16355_ (.B1(_08644_),
    .Y(_09608_),
    .A2(_09607_),
    .A1(_09601_));
 sg13g2_buf_2 _16356_ (.A(_09608_),
    .X(_09609_));
 sg13g2_and2_1 _16357_ (.A(_09531_),
    .B(_09533_),
    .X(_09610_));
 sg13g2_buf_2 _16358_ (.A(_09610_),
    .X(_09611_));
 sg13g2_nand2b_1 _16359_ (.Y(_09612_),
    .B(_09611_),
    .A_N(_00251_));
 sg13g2_buf_1 _16360_ (.A(net1121),
    .X(_09613_));
 sg13g2_and2_1 _16361_ (.A(net807),
    .B(\cpu.dcache.r_tag[6][23] ),
    .X(_09614_));
 sg13g2_a21oi_1 _16362_ (.A1(_09519_),
    .A2(\cpu.dcache.r_tag[4][23] ),
    .Y(_09615_),
    .B1(_09614_));
 sg13g2_nand3_1 _16363_ (.B(net807),
    .C(\cpu.dcache.r_tag[7][23] ),
    .A(net805),
    .Y(_09616_));
 sg13g2_o21ai_1 _16364_ (.B1(_09616_),
    .Y(_09617_),
    .A1(net805),
    .A2(_09615_));
 sg13g2_nand2_1 _16365_ (.Y(_09618_),
    .A(net1048),
    .B(_09617_));
 sg13g2_a22oi_1 _16366_ (.Y(_09619_),
    .B1(_09504_),
    .B2(\cpu.dcache.r_tag[3][23] ),
    .A2(net624),
    .A1(\cpu.dcache.r_tag[1][23] ));
 sg13g2_a22oi_1 _16367_ (.Y(_09620_),
    .B1(net702),
    .B2(\cpu.dcache.r_tag[5][23] ),
    .A2(_09517_),
    .A1(\cpu.dcache.r_tag[2][23] ));
 sg13g2_nand4_1 _16368_ (.B(_09618_),
    .C(_09619_),
    .A(_09612_),
    .Y(_09621_),
    .D(_09620_));
 sg13g2_xnor2_1 _16369_ (.Y(_09622_),
    .A(_09609_),
    .B(_09621_));
 sg13g2_buf_1 _16370_ (.A(net623),
    .X(_09623_));
 sg13g2_mux2_1 _16371_ (.A0(\cpu.dcache.r_tag[4][15] ),
    .A1(\cpu.dcache.r_tag[6][15] ),
    .S(net807),
    .X(_09624_));
 sg13g2_nor2_2 _16372_ (.A(_09348_),
    .B(net807),
    .Y(_09625_));
 sg13g2_a22oi_1 _16373_ (.Y(_09626_),
    .B1(_09625_),
    .B2(\cpu.dcache.r_tag[5][15] ),
    .A2(_09624_),
    .A1(_09348_));
 sg13g2_nand2b_1 _16374_ (.Y(_09627_),
    .B(net1048),
    .A_N(_09626_));
 sg13g2_a22oi_1 _16375_ (.Y(_09628_),
    .B1(net699),
    .B2(\cpu.dcache.r_tag[7][15] ),
    .A2(net625),
    .A1(\cpu.dcache.r_tag[2][15] ));
 sg13g2_a22oi_1 _16376_ (.Y(_09629_),
    .B1(net704),
    .B2(\cpu.dcache.r_tag[3][15] ),
    .A2(net624),
    .A1(\cpu.dcache.r_tag[1][15] ));
 sg13g2_and3_1 _16377_ (.X(_09630_),
    .A(_09627_),
    .B(_09628_),
    .C(_09629_));
 sg13g2_o21ai_1 _16378_ (.B1(_09630_),
    .Y(_09631_),
    .A1(_00246_),
    .A2(net548));
 sg13g2_buf_1 _16379_ (.A(_08377_),
    .X(_09632_));
 sg13g2_buf_8 _16380_ (.A(_09543_),
    .X(_09633_));
 sg13g2_buf_2 _16381_ (.A(_09545_),
    .X(_09634_));
 sg13g2_mux4_1 _16382_ (.S0(net690),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][3] ),
    .S1(net793),
    .X(_09635_));
 sg13g2_mux4_1 _16383_ (.S0(_09633_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][3] ),
    .S1(net793),
    .X(_09636_));
 sg13g2_buf_8 _16384_ (.A(net927),
    .X(_09637_));
 sg13g2_mux4_1 _16385_ (.S0(net792),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][3] ),
    .S1(net793),
    .X(_09638_));
 sg13g2_mux4_1 _16386_ (.S0(net690),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][3] ),
    .S1(_09634_),
    .X(_09639_));
 sg13g2_mux4_1 _16387_ (.S0(_08497_),
    .A0(_09635_),
    .A1(_09636_),
    .A2(_09638_),
    .A3(_09639_),
    .S1(net801),
    .X(_09640_));
 sg13g2_nand2_1 _16388_ (.Y(_09641_),
    .A(net1132),
    .B(_09640_));
 sg13g2_mux4_1 _16389_ (.S0(net696),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][3] ),
    .S1(net799),
    .X(_09642_));
 sg13g2_mux4_1 _16390_ (.S0(net693),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][3] ),
    .S1(net798),
    .X(_09643_));
 sg13g2_mux4_1 _16391_ (.S0(net690),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][3] ),
    .S1(net793),
    .X(_09644_));
 sg13g2_mux4_1 _16392_ (.S0(net690),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][3] ),
    .S1(_09634_),
    .X(_09645_));
 sg13g2_mux4_1 _16393_ (.S0(_08497_),
    .A0(_09642_),
    .A1(_09643_),
    .A2(_09644_),
    .A3(_09645_),
    .S1(net801),
    .X(_09646_));
 sg13g2_o21ai_1 _16394_ (.B1(net1075),
    .Y(_09647_),
    .A1(_08695_),
    .A2(_09646_));
 sg13g2_o21ai_1 _16395_ (.B1(_09647_),
    .Y(_09648_),
    .A1(net926),
    .A2(_09641_));
 sg13g2_buf_1 _16396_ (.A(_09648_),
    .X(_09649_));
 sg13g2_xnor2_1 _16397_ (.Y(_09650_),
    .A(_09631_),
    .B(_09649_));
 sg13g2_nand4_1 _16398_ (.B(_09595_),
    .C(_09622_),
    .A(_09566_),
    .Y(_09651_),
    .D(_09650_));
 sg13g2_buf_2 _16399_ (.A(net1072),
    .X(_09652_));
 sg13g2_mux4_1 _16400_ (.S0(net792),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][7] ),
    .S1(net925),
    .X(_09653_));
 sg13g2_mux4_1 _16401_ (.S0(net792),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][7] ),
    .S1(net925),
    .X(_09654_));
 sg13g2_mux4_1 _16402_ (.S0(net792),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][7] ),
    .S1(net925),
    .X(_09655_));
 sg13g2_mux4_1 _16403_ (.S0(net792),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][7] ),
    .S1(net925),
    .X(_09656_));
 sg13g2_mux4_1 _16404_ (.S0(net794),
    .A0(_09653_),
    .A1(_09654_),
    .A2(_09655_),
    .A3(_09656_),
    .S1(_09539_),
    .X(_09657_));
 sg13g2_nand2_1 _16405_ (.Y(_09658_),
    .A(net796),
    .B(_09657_));
 sg13g2_mux4_1 _16406_ (.S0(net792),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][7] ),
    .S1(_09652_),
    .X(_09659_));
 sg13g2_mux4_1 _16407_ (.S0(net792),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][7] ),
    .S1(net925),
    .X(_09660_));
 sg13g2_mux4_1 _16408_ (.S0(_09637_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][7] ),
    .S1(_09652_),
    .X(_09661_));
 sg13g2_mux4_1 _16409_ (.S0(_09637_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][7] ),
    .S1(net925),
    .X(_09662_));
 sg13g2_mux4_1 _16410_ (.S0(net794),
    .A0(_09659_),
    .A1(_09660_),
    .A2(_09661_),
    .A3(_09662_),
    .S1(net801),
    .X(_09663_));
 sg13g2_nand2_1 _16411_ (.Y(_09664_),
    .A(net691),
    .B(_09663_));
 sg13g2_a21oi_2 _16412_ (.B1(_08644_),
    .Y(_09665_),
    .A2(_09664_),
    .A1(_09658_));
 sg13g2_buf_2 _16413_ (.A(_09665_),
    .X(_09666_));
 sg13g2_inv_1 _16414_ (.Y(_09667_),
    .A(_09666_));
 sg13g2_nor2_1 _16415_ (.A(_00250_),
    .B(net548),
    .Y(_09668_));
 sg13g2_mux2_1 _16416_ (.A0(\cpu.dcache.r_tag[5][19] ),
    .A1(\cpu.dcache.r_tag[7][19] ),
    .S(net807),
    .X(_09669_));
 sg13g2_nor2_1 _16417_ (.A(net1054),
    .B(net934),
    .Y(_09670_));
 sg13g2_buf_1 _16418_ (.A(_09670_),
    .X(_09671_));
 sg13g2_a22oi_1 _16419_ (.Y(_09672_),
    .B1(_09671_),
    .B2(\cpu.dcache.r_tag[4][19] ),
    .A2(_09669_),
    .A1(_09379_));
 sg13g2_nor2_1 _16420_ (.A(_09491_),
    .B(_09672_),
    .Y(_09673_));
 sg13g2_a22oi_1 _16421_ (.Y(_09674_),
    .B1(net701),
    .B2(\cpu.dcache.r_tag[6][19] ),
    .A2(net704),
    .A1(\cpu.dcache.r_tag[3][19] ));
 sg13g2_a22oi_1 _16422_ (.Y(_09675_),
    .B1(net625),
    .B2(\cpu.dcache.r_tag[2][19] ),
    .A2(net624),
    .A1(\cpu.dcache.r_tag[1][19] ));
 sg13g2_nand2_1 _16423_ (.Y(_09676_),
    .A(_09674_),
    .B(_09675_));
 sg13g2_nor3_1 _16424_ (.A(_09668_),
    .B(_09673_),
    .C(_09676_),
    .Y(_09677_));
 sg13g2_xnor2_1 _16425_ (.Y(_09678_),
    .A(_09667_),
    .B(_09677_));
 sg13g2_buf_8 _16426_ (.A(_09543_),
    .X(_09679_));
 sg13g2_buf_1 _16427_ (.A(net925),
    .X(_09680_));
 sg13g2_mux4_1 _16428_ (.S0(_09679_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][4] ),
    .S1(_09680_),
    .X(_09681_));
 sg13g2_buf_8 _16429_ (.A(net792),
    .X(_09682_));
 sg13g2_mux4_1 _16430_ (.S0(net687),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][4] ),
    .S1(net791),
    .X(_09683_));
 sg13g2_buf_2 _16431_ (.A(net925),
    .X(_09684_));
 sg13g2_mux4_1 _16432_ (.S0(net688),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][4] ),
    .S1(net790),
    .X(_09685_));
 sg13g2_mux4_1 _16433_ (.S0(net688),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][4] ),
    .S1(net790),
    .X(_09686_));
 sg13g2_mux4_1 _16434_ (.S0(net692),
    .A0(_09681_),
    .A1(_09683_),
    .A2(_09685_),
    .A3(_09686_),
    .S1(net698),
    .X(_09687_));
 sg13g2_nand2_1 _16435_ (.Y(_09688_),
    .A(net796),
    .B(_09687_));
 sg13g2_mux4_1 _16436_ (.S0(net688),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][4] ),
    .S1(net790),
    .X(_09689_));
 sg13g2_mux4_1 _16437_ (.S0(_09679_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][4] ),
    .S1(_09684_),
    .X(_09690_));
 sg13g2_mux4_1 _16438_ (.S0(_09556_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][4] ),
    .S1(net797),
    .X(_09691_));
 sg13g2_mux4_1 _16439_ (.S0(net695),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][4] ),
    .S1(net797),
    .X(_09692_));
 sg13g2_mux4_1 _16440_ (.S0(net692),
    .A0(_09689_),
    .A1(_09690_),
    .A2(_09691_),
    .A3(_09692_),
    .S1(net698),
    .X(_09693_));
 sg13g2_nand2_1 _16441_ (.Y(_09694_),
    .A(net691),
    .B(_09693_));
 sg13g2_a21oi_1 _16442_ (.A1(_09688_),
    .A2(_09694_),
    .Y(_09695_),
    .B1(_08645_));
 sg13g2_buf_1 _16443_ (.A(_09695_),
    .X(_09696_));
 sg13g2_buf_1 _16444_ (.A(net624),
    .X(_09697_));
 sg13g2_buf_1 _16445_ (.A(_09533_),
    .X(_09698_));
 sg13g2_a22oi_1 _16446_ (.Y(_09699_),
    .B1(_09528_),
    .B2(\cpu.dcache.r_tag[7][16] ),
    .A2(_09502_),
    .A1(\cpu.dcache.r_tag[3][16] ));
 sg13g2_a22oi_1 _16447_ (.Y(_09700_),
    .B1(_09510_),
    .B2(\cpu.dcache.r_tag[5][16] ),
    .A2(_09516_),
    .A1(\cpu.dcache.r_tag[2][16] ));
 sg13g2_a22oi_1 _16448_ (.Y(_09701_),
    .B1(_09520_),
    .B2(\cpu.dcache.r_tag[6][16] ),
    .A2(net703),
    .A1(\cpu.dcache.r_tag[4][16] ));
 sg13g2_nand3_1 _16449_ (.B(_09700_),
    .C(_09701_),
    .A(_09699_),
    .Y(_09702_));
 sg13g2_nand2_1 _16450_ (.Y(_09703_),
    .A(_00247_),
    .B(_09533_));
 sg13g2_o21ai_1 _16451_ (.B1(_09703_),
    .Y(_09704_),
    .A1(_09698_),
    .A2(_09702_));
 sg13g2_o21ai_1 _16452_ (.B1(net547),
    .Y(_09705_),
    .A1(\cpu.dcache.r_tag[1][16] ),
    .A2(_09702_));
 sg13g2_o21ai_1 _16453_ (.B1(_09705_),
    .Y(_09706_),
    .A1(net547),
    .A2(_09704_));
 sg13g2_xnor2_1 _16454_ (.Y(_09707_),
    .A(net406),
    .B(_09706_));
 sg13g2_nand2_1 _16455_ (.Y(_09708_),
    .A(_09678_),
    .B(_09707_));
 sg13g2_mux4_1 _16456_ (.S0(net693),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][6] ),
    .S1(net798),
    .X(_09709_));
 sg13g2_mux4_1 _16457_ (.S0(net697),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][6] ),
    .S1(net800),
    .X(_09710_));
 sg13g2_mux4_1 _16458_ (.S0(net696),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][6] ),
    .S1(net799),
    .X(_09711_));
 sg13g2_mux4_1 _16459_ (.S0(net696),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][6] ),
    .S1(net799),
    .X(_09712_));
 sg13g2_mux4_1 _16460_ (.S0(net794),
    .A0(_09709_),
    .A1(_09710_),
    .A2(_09711_),
    .A3(_09712_),
    .S1(net801),
    .X(_09713_));
 sg13g2_nand2_1 _16461_ (.Y(_09714_),
    .A(net796),
    .B(_09713_));
 sg13g2_mux4_1 _16462_ (.S0(net693),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][6] ),
    .S1(net798),
    .X(_09715_));
 sg13g2_mux4_1 _16463_ (.S0(net693),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][6] ),
    .S1(net798),
    .X(_09716_));
 sg13g2_mux4_1 _16464_ (.S0(_09633_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][6] ),
    .S1(_09550_),
    .X(_09717_));
 sg13g2_mux4_1 _16465_ (.S0(_09549_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][6] ),
    .S1(_09550_),
    .X(_09718_));
 sg13g2_mux4_1 _16466_ (.S0(net794),
    .A0(_09715_),
    .A1(_09716_),
    .A2(_09717_),
    .A3(_09718_),
    .S1(_09539_),
    .X(_09719_));
 sg13g2_nand2_1 _16467_ (.Y(_09720_),
    .A(net691),
    .B(_09719_));
 sg13g2_a21oi_2 _16468_ (.B1(_08644_),
    .Y(_09721_),
    .A2(_09720_),
    .A1(_09714_));
 sg13g2_buf_1 _16469_ (.A(_09721_),
    .X(_09722_));
 sg13g2_a22oi_1 _16470_ (.Y(_09723_),
    .B1(_09508_),
    .B2(\cpu.dcache.r_tag[4][18] ),
    .A2(_09503_),
    .A1(\cpu.dcache.r_tag[3][18] ));
 sg13g2_nand2_1 _16471_ (.Y(_09724_),
    .A(\cpu.dcache.r_tag[7][18] ),
    .B(net699));
 sg13g2_a22oi_1 _16472_ (.Y(_09725_),
    .B1(_09521_),
    .B2(\cpu.dcache.r_tag[6][18] ),
    .A2(net625),
    .A1(\cpu.dcache.r_tag[2][18] ));
 sg13g2_nor2_1 _16473_ (.A(_00249_),
    .B(net623),
    .Y(_09726_));
 sg13g2_a221oi_1 _16474_ (.B2(\cpu.dcache.r_tag[5][18] ),
    .C1(_09726_),
    .B1(net702),
    .A1(\cpu.dcache.r_tag[1][18] ),
    .Y(_09727_),
    .A2(net624));
 sg13g2_nand4_1 _16475_ (.B(_09724_),
    .C(_09725_),
    .A(_09723_),
    .Y(_09728_),
    .D(_09727_));
 sg13g2_xnor2_1 _16476_ (.Y(_09729_),
    .A(net405),
    .B(_09728_));
 sg13g2_mux4_1 _16477_ (.S0(net688),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][8] ),
    .S1(net790),
    .X(_09730_));
 sg13g2_mux4_1 _16478_ (.S0(net688),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][8] ),
    .S1(net790),
    .X(_09731_));
 sg13g2_mux4_1 _16479_ (.S0(net694),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][8] ),
    .S1(net795),
    .X(_09732_));
 sg13g2_mux4_1 _16480_ (.S0(net695),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][8] ),
    .S1(net797),
    .X(_09733_));
 sg13g2_mux4_1 _16481_ (.S0(net692),
    .A0(_09730_),
    .A1(_09731_),
    .A2(_09732_),
    .A3(_09733_),
    .S1(net698),
    .X(_09734_));
 sg13g2_nand2_1 _16482_ (.Y(_09735_),
    .A(_09568_),
    .B(_09734_));
 sg13g2_mux4_1 _16483_ (.S0(net695),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][8] ),
    .S1(net790),
    .X(_09736_));
 sg13g2_mux4_1 _16484_ (.S0(net688),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][8] ),
    .S1(net790),
    .X(_09737_));
 sg13g2_mux4_1 _16485_ (.S0(net694),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][8] ),
    .S1(net795),
    .X(_09738_));
 sg13g2_mux4_1 _16486_ (.S0(net694),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][8] ),
    .S1(net795),
    .X(_09739_));
 sg13g2_mux4_1 _16487_ (.S0(net692),
    .A0(_09736_),
    .A1(_09737_),
    .A2(_09738_),
    .A3(_09739_),
    .S1(net698),
    .X(_09740_));
 sg13g2_nand2_1 _16488_ (.Y(_09741_),
    .A(net691),
    .B(_09740_));
 sg13g2_a21oi_2 _16489_ (.B1(_08645_),
    .Y(_09742_),
    .A2(_09741_),
    .A1(_09735_));
 sg13g2_buf_1 _16490_ (.A(_09742_),
    .X(_09743_));
 sg13g2_and2_1 _16491_ (.A(\cpu.dcache.r_tag[3][20] ),
    .B(net704),
    .X(_09744_));
 sg13g2_a221oi_1 _16492_ (.B2(\cpu.dcache.r_tag[6][20] ),
    .C1(_09744_),
    .B1(net701),
    .A1(\cpu.dcache.r_tag[4][20] ),
    .Y(_09745_),
    .A2(_09508_));
 sg13g2_a22oi_1 _16493_ (.Y(_09746_),
    .B1(net702),
    .B2(\cpu.dcache.r_tag[5][20] ),
    .A2(net624),
    .A1(\cpu.dcache.r_tag[1][20] ));
 sg13g2_a22oi_1 _16494_ (.Y(_09747_),
    .B1(net699),
    .B2(\cpu.dcache.r_tag[7][20] ),
    .A2(net625),
    .A1(\cpu.dcache.r_tag[2][20] ));
 sg13g2_nand4_1 _16495_ (.B(_09745_),
    .C(_09746_),
    .A(_09623_),
    .Y(_09748_),
    .D(_09747_));
 sg13g2_o21ai_1 _16496_ (.B1(_09748_),
    .Y(_09749_),
    .A1(\cpu.dcache.r_tag[0][20] ),
    .A2(net548));
 sg13g2_xor2_1 _16497_ (.B(_09749_),
    .A(net404),
    .X(_09750_));
 sg13g2_nand2_1 _16498_ (.Y(_09751_),
    .A(_09729_),
    .B(_09750_));
 sg13g2_nor3_1 _16499_ (.A(_09651_),
    .B(_09708_),
    .C(_09751_),
    .Y(_09752_));
 sg13g2_buf_2 _16500_ (.A(net927),
    .X(_09753_));
 sg13g2_buf_2 _16501_ (.A(net1072),
    .X(_09754_));
 sg13g2_mux4_1 _16502_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][0] ),
    .S1(net924),
    .X(_09755_));
 sg13g2_mux4_1 _16503_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][0] ),
    .S1(net924),
    .X(_09756_));
 sg13g2_mux4_1 _16504_ (.S0(net927),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][0] ),
    .S1(net1072),
    .X(_09757_));
 sg13g2_mux4_1 _16505_ (.S0(net927),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][0] ),
    .S1(_08422_),
    .X(_09758_));
 sg13g2_mux4_1 _16506_ (.S0(_08428_),
    .A0(_09755_),
    .A1(_09756_),
    .A2(_09757_),
    .A3(_09758_),
    .S1(net956),
    .X(_09759_));
 sg13g2_mux4_1 _16507_ (.S0(net927),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][0] ),
    .S1(net1072),
    .X(_09760_));
 sg13g2_mux4_1 _16508_ (.S0(net927),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][0] ),
    .S1(net924),
    .X(_09761_));
 sg13g2_mux4_1 _16509_ (.S0(net927),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][0] ),
    .S1(_08422_),
    .X(_09762_));
 sg13g2_mux4_1 _16510_ (.S0(_09542_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][0] ),
    .S1(net1072),
    .X(_09763_));
 sg13g2_mux4_1 _16511_ (.S0(_08428_),
    .A0(_09760_),
    .A1(_09761_),
    .A2(_09762_),
    .A3(_09763_),
    .S1(net956),
    .X(_09764_));
 sg13g2_mux2_1 _16512_ (.A0(_09759_),
    .A1(_09764_),
    .S(net691),
    .X(_09765_));
 sg13g2_nand2_1 _16513_ (.Y(_09766_),
    .A(net1132),
    .B(_09765_));
 sg13g2_o21ai_1 _16514_ (.B1(_09766_),
    .Y(_09767_),
    .A1(_08531_),
    .A2(_08400_));
 sg13g2_buf_1 _16515_ (.A(_09767_),
    .X(_09768_));
 sg13g2_buf_1 _16516_ (.A(_09611_),
    .X(_09769_));
 sg13g2_a22oi_1 _16517_ (.Y(_09770_),
    .B1(net625),
    .B2(\cpu.dcache.r_tag[2][12] ),
    .A2(net700),
    .A1(\cpu.dcache.r_tag[1][12] ));
 sg13g2_a22oi_1 _16518_ (.Y(_09771_),
    .B1(net703),
    .B2(\cpu.dcache.r_tag[4][12] ),
    .A2(_09503_),
    .A1(\cpu.dcache.r_tag[3][12] ));
 sg13g2_mux2_1 _16519_ (.A0(\cpu.dcache.r_tag[5][12] ),
    .A1(\cpu.dcache.r_tag[7][12] ),
    .S(net934),
    .X(_09772_));
 sg13g2_a22oi_1 _16520_ (.Y(_09773_),
    .B1(_09772_),
    .B2(net932),
    .A2(net928),
    .A1(\cpu.dcache.r_tag[6][12] ));
 sg13g2_nand2b_1 _16521_ (.Y(_09774_),
    .B(net1048),
    .A_N(_09773_));
 sg13g2_and4_1 _16522_ (.A(_09535_),
    .B(_09770_),
    .C(_09771_),
    .D(_09774_),
    .X(_09775_));
 sg13g2_a21oi_1 _16523_ (.A1(_00243_),
    .A2(net546),
    .Y(_09776_),
    .B1(_09775_));
 sg13g2_xor2_1 _16524_ (.B(_09776_),
    .A(net403),
    .X(_09777_));
 sg13g2_nand2b_1 _16525_ (.Y(_09778_),
    .B(_09611_),
    .A_N(_00244_));
 sg13g2_a22oi_1 _16526_ (.Y(_09779_),
    .B1(net701),
    .B2(\cpu.dcache.r_tag[6][13] ),
    .A2(net704),
    .A1(\cpu.dcache.r_tag[3][13] ));
 sg13g2_a22oi_1 _16527_ (.Y(_09780_),
    .B1(_09529_),
    .B2(\cpu.dcache.r_tag[7][13] ),
    .A2(net703),
    .A1(\cpu.dcache.r_tag[4][13] ));
 sg13g2_a22oi_1 _16528_ (.Y(_09781_),
    .B1(net702),
    .B2(\cpu.dcache.r_tag[5][13] ),
    .A2(net625),
    .A1(\cpu.dcache.r_tag[2][13] ));
 sg13g2_nand4_1 _16529_ (.B(_09779_),
    .C(_09780_),
    .A(_09778_),
    .Y(_09782_),
    .D(_09781_));
 sg13g2_a21oi_1 _16530_ (.A1(\cpu.dcache.r_tag[1][13] ),
    .A2(net547),
    .Y(_09783_),
    .B1(_09782_));
 sg13g2_mux4_1 _16531_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][1] ),
    .S1(net924),
    .X(_09784_));
 sg13g2_mux4_1 _16532_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][1] ),
    .S1(_09545_),
    .X(_09785_));
 sg13g2_mux4_1 _16533_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][1] ),
    .S1(net924),
    .X(_09786_));
 sg13g2_mux4_1 _16534_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][1] ),
    .S1(net924),
    .X(_09787_));
 sg13g2_mux4_1 _16535_ (.S0(_09576_),
    .A0(_09784_),
    .A1(_09785_),
    .A2(_09786_),
    .A3(_09787_),
    .S1(_08405_),
    .X(_09788_));
 sg13g2_mux4_1 _16536_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][1] ),
    .S1(net924),
    .X(_09789_));
 sg13g2_mux4_1 _16537_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][1] ),
    .S1(net924),
    .X(_09790_));
 sg13g2_mux4_1 _16538_ (.S0(_09753_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][1] ),
    .S1(_09754_),
    .X(_09791_));
 sg13g2_mux4_1 _16539_ (.S0(_09753_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][1] ),
    .S1(_09754_),
    .X(_09792_));
 sg13g2_mux4_1 _16540_ (.S0(_08428_),
    .A0(_09789_),
    .A1(_09790_),
    .A2(_09791_),
    .A3(_09792_),
    .S1(_08405_),
    .X(_09793_));
 sg13g2_mux2_1 _16541_ (.A0(_09788_),
    .A1(_09793_),
    .S(_09580_),
    .X(_09794_));
 sg13g2_nand2_1 _16542_ (.Y(_09795_),
    .A(net1132),
    .B(_09794_));
 sg13g2_o21ai_1 _16543_ (.B1(_09795_),
    .Y(_09796_),
    .A1(net1068),
    .A2(_08404_));
 sg13g2_buf_1 _16544_ (.A(_09796_),
    .X(_09797_));
 sg13g2_xnor2_1 _16545_ (.Y(_09798_),
    .A(_09783_),
    .B(net402));
 sg13g2_nor2_1 _16546_ (.A(_09777_),
    .B(_09798_),
    .Y(_09799_));
 sg13g2_inv_1 _16547_ (.Y(_09800_),
    .A(_00242_));
 sg13g2_mux2_1 _16548_ (.A0(\cpu.dcache.r_tag[5][11] ),
    .A1(\cpu.dcache.r_tag[7][11] ),
    .S(_09340_),
    .X(_09801_));
 sg13g2_a22oi_1 _16549_ (.Y(_09802_),
    .B1(_09801_),
    .B2(net932),
    .A2(net689),
    .A1(\cpu.dcache.r_tag[4][11] ));
 sg13g2_nand2b_1 _16550_ (.Y(_09803_),
    .B(net1048),
    .A_N(_09802_));
 sg13g2_a22oi_1 _16551_ (.Y(_09804_),
    .B1(_09516_),
    .B2(\cpu.dcache.r_tag[2][11] ),
    .A2(_09502_),
    .A1(\cpu.dcache.r_tag[3][11] ));
 sg13g2_a22oi_1 _16552_ (.Y(_09805_),
    .B1(net701),
    .B2(\cpu.dcache.r_tag[6][11] ),
    .A2(net700),
    .A1(\cpu.dcache.r_tag[1][11] ));
 sg13g2_nand3_1 _16553_ (.B(_09804_),
    .C(_09805_),
    .A(_09803_),
    .Y(_09806_));
 sg13g2_a21oi_1 _16554_ (.A1(_09800_),
    .A2(_09611_),
    .Y(_09807_),
    .B1(_09806_));
 sg13g2_xor2_1 _16555_ (.B(_09807_),
    .A(_00241_),
    .X(_09808_));
 sg13g2_nand2b_1 _16556_ (.Y(_09809_),
    .B(_09611_),
    .A_N(_00232_));
 sg13g2_and2_1 _16557_ (.A(net934),
    .B(\cpu.dcache.r_tag[6][6] ),
    .X(_09810_));
 sg13g2_a21oi_1 _16558_ (.A1(_09519_),
    .A2(\cpu.dcache.r_tag[4][6] ),
    .Y(_09811_),
    .B1(_09810_));
 sg13g2_nand3_1 _16559_ (.B(_09341_),
    .C(\cpu.dcache.r_tag[7][6] ),
    .A(_09378_),
    .Y(_09812_));
 sg13g2_o21ai_1 _16560_ (.B1(_09812_),
    .Y(_09813_),
    .A1(net932),
    .A2(_09811_));
 sg13g2_nand2_1 _16561_ (.Y(_09814_),
    .A(net1048),
    .B(_09813_));
 sg13g2_a22oi_1 _16562_ (.Y(_09815_),
    .B1(net704),
    .B2(\cpu.dcache.r_tag[3][6] ),
    .A2(net700),
    .A1(\cpu.dcache.r_tag[1][6] ));
 sg13g2_a22oi_1 _16563_ (.Y(_09816_),
    .B1(net702),
    .B2(\cpu.dcache.r_tag[5][6] ),
    .A2(_09517_),
    .A1(\cpu.dcache.r_tag[2][6] ));
 sg13g2_nand4_1 _16564_ (.B(_09814_),
    .C(_09815_),
    .A(_09809_),
    .Y(_09817_),
    .D(_09816_));
 sg13g2_xnor2_1 _16565_ (.Y(_09818_),
    .A(_00231_),
    .B(_09817_));
 sg13g2_nand2_1 _16566_ (.Y(_09819_),
    .A(\cpu.dcache.r_tag[7][10] ),
    .B(_09529_));
 sg13g2_a22oi_1 _16567_ (.Y(_09820_),
    .B1(_09510_),
    .B2(\cpu.dcache.r_tag[5][10] ),
    .A2(_09502_),
    .A1(\cpu.dcache.r_tag[3][10] ));
 sg13g2_a22oi_1 _16568_ (.Y(_09821_),
    .B1(_09520_),
    .B2(\cpu.dcache.r_tag[6][10] ),
    .A2(net703),
    .A1(\cpu.dcache.r_tag[4][10] ));
 sg13g2_a22oi_1 _16569_ (.Y(_09822_),
    .B1(_09516_),
    .B2(\cpu.dcache.r_tag[2][10] ),
    .A2(net700),
    .A1(\cpu.dcache.r_tag[1][10] ));
 sg13g2_nand4_1 _16570_ (.B(_09820_),
    .C(_09821_),
    .A(_09819_),
    .Y(_09823_),
    .D(_09822_));
 sg13g2_nand2_1 _16571_ (.Y(_09824_),
    .A(_00240_),
    .B(_09611_));
 sg13g2_o21ai_1 _16572_ (.B1(_09824_),
    .Y(_09825_),
    .A1(_09611_),
    .A2(_09823_));
 sg13g2_xor2_1 _16573_ (.B(_09825_),
    .A(_00239_),
    .X(_09826_));
 sg13g2_nor3_1 _16574_ (.A(_09808_),
    .B(_09818_),
    .C(_09826_),
    .Y(_09827_));
 sg13g2_buf_1 _16575_ (.A(_00229_),
    .X(_09828_));
 sg13g2_inv_1 _16576_ (.Y(_09829_),
    .A(\cpu.dcache.r_tag[6][5] ));
 sg13g2_nand3b_1 _16577_ (.B(net1121),
    .C(net1055),
    .Y(_09830_),
    .A_N(_09346_));
 sg13g2_buf_2 _16578_ (.A(_09830_),
    .X(_09831_));
 sg13g2_nand4_1 _16579_ (.B(_09339_),
    .C(_09500_),
    .A(net1054),
    .Y(_09832_),
    .D(\cpu.dcache.r_tag[3][5] ));
 sg13g2_o21ai_1 _16580_ (.B1(_09832_),
    .Y(_09833_),
    .A1(_09829_),
    .A2(_09831_));
 sg13g2_inv_1 _16581_ (.Y(_09834_),
    .A(\cpu.dcache.r_tag[5][5] ));
 sg13g2_nand3b_1 _16582_ (.B(\cpu.addr[4] ),
    .C(_09346_),
    .Y(_09835_),
    .A_N(_09338_));
 sg13g2_buf_2 _16583_ (.A(_09835_),
    .X(_09836_));
 sg13g2_nand4_1 _16584_ (.B(net1121),
    .C(net1055),
    .A(net1054),
    .Y(_09837_),
    .D(\cpu.dcache.r_tag[7][5] ));
 sg13g2_o21ai_1 _16585_ (.B1(_09837_),
    .Y(_09838_),
    .A1(_09834_),
    .A2(_09836_));
 sg13g2_nor2b_1 _16586_ (.A(_09347_),
    .B_N(net1121),
    .Y(_09839_));
 sg13g2_and3_1 _16587_ (.X(_09840_),
    .A(_09519_),
    .B(\cpu.dcache.r_tag[4][5] ),
    .C(_09839_));
 sg13g2_and3_1 _16588_ (.X(_09841_),
    .A(_09500_),
    .B(\cpu.dcache.r_tag[2][5] ),
    .C(net928));
 sg13g2_or4_1 _16589_ (.A(_09833_),
    .B(_09838_),
    .C(_09840_),
    .D(_09841_),
    .X(_09842_));
 sg13g2_nand2_1 _16590_ (.Y(_09843_),
    .A(_00230_),
    .B(_09533_));
 sg13g2_o21ai_1 _16591_ (.B1(_09843_),
    .Y(_09844_),
    .A1(_09533_),
    .A2(_09842_));
 sg13g2_o21ai_1 _16592_ (.B1(net700),
    .Y(_09845_),
    .A1(\cpu.dcache.r_tag[1][5] ),
    .A2(_09842_));
 sg13g2_o21ai_1 _16593_ (.B1(_09845_),
    .Y(_09846_),
    .A1(_09526_),
    .A2(_09844_));
 sg13g2_xnor2_1 _16594_ (.Y(_09847_),
    .A(net1120),
    .B(_09846_));
 sg13g2_inv_1 _16595_ (.Y(_09848_),
    .A(_00234_));
 sg13g2_a22oi_1 _16596_ (.Y(_09849_),
    .B1(_09516_),
    .B2(\cpu.dcache.r_tag[2][7] ),
    .A2(net700),
    .A1(\cpu.dcache.r_tag[1][7] ));
 sg13g2_a22oi_1 _16597_ (.Y(_09850_),
    .B1(net703),
    .B2(\cpu.dcache.r_tag[4][7] ),
    .A2(_09502_),
    .A1(\cpu.dcache.r_tag[3][7] ));
 sg13g2_mux2_1 _16598_ (.A0(\cpu.dcache.r_tag[5][7] ),
    .A1(\cpu.dcache.r_tag[7][7] ),
    .S(net934),
    .X(_09851_));
 sg13g2_a22oi_1 _16599_ (.Y(_09852_),
    .B1(_09851_),
    .B2(net932),
    .A2(net928),
    .A1(\cpu.dcache.r_tag[6][7] ));
 sg13g2_nand2b_1 _16600_ (.Y(_09853_),
    .B(net1121),
    .A_N(_09852_));
 sg13g2_nand4_1 _16601_ (.B(_09849_),
    .C(_09850_),
    .A(_09534_),
    .Y(_09854_),
    .D(_09853_));
 sg13g2_o21ai_1 _16602_ (.B1(_09854_),
    .Y(_09855_),
    .A1(_09848_),
    .A2(net623));
 sg13g2_xor2_1 _16603_ (.B(_09855_),
    .A(_00233_),
    .X(_09856_));
 sg13g2_inv_1 _16604_ (.Y(_09857_),
    .A(_00238_));
 sg13g2_a22oi_1 _16605_ (.Y(_09858_),
    .B1(_09516_),
    .B2(\cpu.dcache.r_tag[2][9] ),
    .A2(_09525_),
    .A1(\cpu.dcache.r_tag[1][9] ));
 sg13g2_a22oi_1 _16606_ (.Y(_09859_),
    .B1(net703),
    .B2(\cpu.dcache.r_tag[4][9] ),
    .A2(_09502_),
    .A1(\cpu.dcache.r_tag[3][9] ));
 sg13g2_mux2_1 _16607_ (.A0(\cpu.dcache.r_tag[5][9] ),
    .A1(\cpu.dcache.r_tag[7][9] ),
    .S(net934),
    .X(_09860_));
 sg13g2_a22oi_1 _16608_ (.Y(_09861_),
    .B1(_09860_),
    .B2(net932),
    .A2(net928),
    .A1(\cpu.dcache.r_tag[6][9] ));
 sg13g2_nand2b_1 _16609_ (.Y(_09862_),
    .B(_09490_),
    .A_N(_09861_));
 sg13g2_nand4_1 _16610_ (.B(_09858_),
    .C(_09859_),
    .A(net623),
    .Y(_09863_),
    .D(_09862_));
 sg13g2_o21ai_1 _16611_ (.B1(_09863_),
    .Y(_09864_),
    .A1(_09857_),
    .A2(net623));
 sg13g2_xor2_1 _16612_ (.B(_09864_),
    .A(_00237_),
    .X(_09865_));
 sg13g2_buf_2 _16613_ (.A(_00235_),
    .X(_09866_));
 sg13g2_inv_1 _16614_ (.Y(_09867_),
    .A(_00236_));
 sg13g2_a22oi_1 _16615_ (.Y(_09868_),
    .B1(_09516_),
    .B2(\cpu.dcache.r_tag[2][8] ),
    .A2(net700),
    .A1(\cpu.dcache.r_tag[1][8] ));
 sg13g2_a22oi_1 _16616_ (.Y(_09869_),
    .B1(_09507_),
    .B2(\cpu.dcache.r_tag[4][8] ),
    .A2(_09502_),
    .A1(\cpu.dcache.r_tag[3][8] ));
 sg13g2_mux2_1 _16617_ (.A0(\cpu.dcache.r_tag[5][8] ),
    .A1(\cpu.dcache.r_tag[7][8] ),
    .S(net934),
    .X(_09870_));
 sg13g2_a22oi_1 _16618_ (.Y(_09871_),
    .B1(_09870_),
    .B2(net932),
    .A2(_09514_),
    .A1(\cpu.dcache.r_tag[6][8] ));
 sg13g2_nand2b_1 _16619_ (.Y(_09872_),
    .B(_09613_),
    .A_N(_09871_));
 sg13g2_nand4_1 _16620_ (.B(_09868_),
    .C(_09869_),
    .A(_09535_),
    .Y(_09873_),
    .D(_09872_));
 sg13g2_o21ai_1 _16621_ (.B1(_09873_),
    .Y(_09874_),
    .A1(_09867_),
    .A2(net623));
 sg13g2_xor2_1 _16622_ (.B(_09874_),
    .A(_09866_),
    .X(_09875_));
 sg13g2_nor4_1 _16623_ (.A(_09847_),
    .B(_09856_),
    .C(_09865_),
    .D(_09875_),
    .Y(_09876_));
 sg13g2_mux4_1 _16624_ (.S0(net696),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][9] ),
    .S1(net799),
    .X(_09877_));
 sg13g2_mux4_1 _16625_ (.S0(net696),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][9] ),
    .S1(net799),
    .X(_09878_));
 sg13g2_mux4_1 _16626_ (.S0(net690),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][9] ),
    .S1(net793),
    .X(_09879_));
 sg13g2_mux4_1 _16627_ (.S0(net690),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][9] ),
    .S1(net793),
    .X(_09880_));
 sg13g2_mux4_1 _16628_ (.S0(net794),
    .A0(_09877_),
    .A1(_09878_),
    .A2(_09879_),
    .A3(_09880_),
    .S1(net801),
    .X(_09881_));
 sg13g2_nand2_1 _16629_ (.Y(_09882_),
    .A(net796),
    .B(_09881_));
 sg13g2_mux4_1 _16630_ (.S0(net696),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][9] ),
    .S1(net799),
    .X(_09883_));
 sg13g2_mux4_1 _16631_ (.S0(net696),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][9] ),
    .S1(net799),
    .X(_09884_));
 sg13g2_mux4_1 _16632_ (.S0(net690),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][9] ),
    .S1(net793),
    .X(_09885_));
 sg13g2_mux4_1 _16633_ (.S0(net690),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][9] ),
    .S1(net793),
    .X(_09886_));
 sg13g2_mux4_1 _16634_ (.S0(net794),
    .A0(_09883_),
    .A1(_09884_),
    .A2(_09885_),
    .A3(_09886_),
    .S1(net801),
    .X(_09887_));
 sg13g2_nand2_1 _16635_ (.Y(_09888_),
    .A(net691),
    .B(_09887_));
 sg13g2_a21oi_1 _16636_ (.A1(_09882_),
    .A2(_09888_),
    .Y(_09889_),
    .B1(_08644_));
 sg13g2_buf_1 _16637_ (.A(_09889_),
    .X(_09890_));
 sg13g2_a22oi_1 _16638_ (.Y(_09891_),
    .B1(_09521_),
    .B2(\cpu.dcache.r_tag[6][21] ),
    .A2(_09511_),
    .A1(\cpu.dcache.r_tag[5][21] ));
 sg13g2_a22oi_1 _16639_ (.Y(_09892_),
    .B1(_09516_),
    .B2(\cpu.dcache.r_tag[2][21] ),
    .A2(_09502_),
    .A1(\cpu.dcache.r_tag[3][21] ));
 sg13g2_a22oi_1 _16640_ (.Y(_09893_),
    .B1(_09528_),
    .B2(\cpu.dcache.r_tag[7][21] ),
    .A2(net703),
    .A1(\cpu.dcache.r_tag[4][21] ));
 sg13g2_nand3_1 _16641_ (.B(_09892_),
    .C(_09893_),
    .A(_09891_),
    .Y(_09894_));
 sg13g2_nand2b_1 _16642_ (.Y(_09895_),
    .B(net686),
    .A_N(\cpu.dcache.r_tag[0][21] ));
 sg13g2_o21ai_1 _16643_ (.B1(_09895_),
    .Y(_09896_),
    .A1(_09698_),
    .A2(_09894_));
 sg13g2_o21ai_1 _16644_ (.B1(_09697_),
    .Y(_09897_),
    .A1(\cpu.dcache.r_tag[1][21] ),
    .A2(_09894_));
 sg13g2_o21ai_1 _16645_ (.B1(_09897_),
    .Y(_09898_),
    .A1(net547),
    .A2(_09896_));
 sg13g2_xnor2_1 _16646_ (.Y(_09899_),
    .A(net401),
    .B(_09898_));
 sg13g2_mux4_1 _16647_ (.S0(net688),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][10] ),
    .S1(_09684_),
    .X(_09900_));
 sg13g2_mux4_1 _16648_ (.S0(net688),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][10] ),
    .S1(net790),
    .X(_09901_));
 sg13g2_mux4_1 _16649_ (.S0(net694),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][10] ),
    .S1(net795),
    .X(_09902_));
 sg13g2_mux4_1 _16650_ (.S0(net694),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][10] ),
    .S1(net795),
    .X(_09903_));
 sg13g2_mux4_1 _16651_ (.S0(_09577_),
    .A0(_09900_),
    .A1(_09901_),
    .A2(_09902_),
    .A3(_09903_),
    .S1(_09540_),
    .X(_09904_));
 sg13g2_nand2_1 _16652_ (.Y(_09905_),
    .A(net796),
    .B(_09904_));
 sg13g2_mux4_1 _16653_ (.S0(net695),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][10] ),
    .S1(_09557_),
    .X(_09906_));
 sg13g2_mux4_1 _16654_ (.S0(net695),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][10] ),
    .S1(net797),
    .X(_09907_));
 sg13g2_mux4_1 _16655_ (.S0(_09544_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][10] ),
    .S1(net800),
    .X(_09908_));
 sg13g2_mux4_1 _16656_ (.S0(net697),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][10] ),
    .S1(net795),
    .X(_09909_));
 sg13g2_mux4_1 _16657_ (.S0(net692),
    .A0(_09906_),
    .A1(_09907_),
    .A2(_09908_),
    .A3(_09909_),
    .S1(_09540_),
    .X(_09910_));
 sg13g2_nand2_1 _16658_ (.Y(_09911_),
    .A(_09580_),
    .B(_09910_));
 sg13g2_a21oi_2 _16659_ (.B1(_08644_),
    .Y(_09912_),
    .A2(_09911_),
    .A1(_09905_));
 sg13g2_buf_1 _16660_ (.A(_09912_),
    .X(_09913_));
 sg13g2_mux2_1 _16661_ (.A0(\cpu.dcache.r_tag[5][22] ),
    .A1(\cpu.dcache.r_tag[7][22] ),
    .S(net807),
    .X(_09914_));
 sg13g2_a22oi_1 _16662_ (.Y(_09915_),
    .B1(_09914_),
    .B2(_09379_),
    .A2(_09671_),
    .A1(\cpu.dcache.r_tag[4][22] ));
 sg13g2_nand2b_1 _16663_ (.Y(_09916_),
    .B(_09613_),
    .A_N(_09915_));
 sg13g2_a22oi_1 _16664_ (.Y(_09917_),
    .B1(net625),
    .B2(\cpu.dcache.r_tag[2][22] ),
    .A2(net704),
    .A1(\cpu.dcache.r_tag[3][22] ));
 sg13g2_a22oi_1 _16665_ (.Y(_09918_),
    .B1(net701),
    .B2(\cpu.dcache.r_tag[6][22] ),
    .A2(net624),
    .A1(\cpu.dcache.r_tag[1][22] ));
 sg13g2_nand3_1 _16666_ (.B(_09917_),
    .C(_09918_),
    .A(_09916_),
    .Y(_09919_));
 sg13g2_a21oi_1 _16667_ (.A1(\cpu.dcache.r_tag[0][22] ),
    .A2(net546),
    .Y(_09920_),
    .B1(_09919_));
 sg13g2_xor2_1 _16668_ (.B(_09920_),
    .A(net400),
    .X(_09921_));
 sg13g2_and4_1 _16669_ (.A(_09827_),
    .B(_09876_),
    .C(_09899_),
    .D(_09921_),
    .X(_09922_));
 sg13g2_nand4_1 _16670_ (.B(_09752_),
    .C(_09799_),
    .A(_09492_),
    .Y(_09923_),
    .D(_09922_));
 sg13g2_buf_1 _16671_ (.A(_09923_),
    .X(_09924_));
 sg13g2_inv_1 _16672_ (.Y(_09925_),
    .A(_09799_));
 sg13g2_nand4_1 _16673_ (.B(_09827_),
    .C(_09876_),
    .A(_09622_),
    .Y(_09926_),
    .D(_09899_));
 sg13g2_nand4_1 _16674_ (.B(_09595_),
    .C(_09650_),
    .A(_09566_),
    .Y(_09927_),
    .D(_09729_));
 sg13g2_nand4_1 _16675_ (.B(_09707_),
    .C(_09750_),
    .A(_09678_),
    .Y(_09928_),
    .D(_09921_));
 sg13g2_nor4_1 _16676_ (.A(_09925_),
    .B(_09926_),
    .C(_09927_),
    .D(_09928_),
    .Y(_09929_));
 sg13g2_a21oi_1 _16677_ (.A1(_09487_),
    .A2(_09929_),
    .Y(_09930_),
    .B1(_09498_));
 sg13g2_a21oi_1 _16678_ (.A1(_09499_),
    .A2(_09924_),
    .Y(_09931_),
    .B1(_09930_));
 sg13g2_nand2b_1 _16679_ (.Y(_09932_),
    .B(_09337_),
    .A_N(_08393_));
 sg13g2_a21oi_1 _16680_ (.A1(net957),
    .A2(_09363_),
    .Y(_09933_),
    .B1(_09932_));
 sg13g2_nand2b_1 _16681_ (.Y(_09934_),
    .B(_09933_),
    .A_N(_09931_));
 sg13g2_o21ai_1 _16682_ (.B1(_09934_),
    .Y(_09935_),
    .A1(net802),
    .A2(_08970_));
 sg13g2_nor2_1 _16683_ (.A(_09483_),
    .B(_09935_),
    .Y(_09936_));
 sg13g2_inv_1 _16684_ (.Y(_09937_),
    .A(_09936_));
 sg13g2_buf_1 _16685_ (.A(\cpu.qspi.r_state[7] ),
    .X(_09938_));
 sg13g2_buf_1 _16686_ (.A(\cpu.qspi.r_ind ),
    .X(_09939_));
 sg13g2_buf_1 _16687_ (.A(_00252_),
    .X(_09940_));
 sg13g2_buf_1 _16688_ (.A(\cpu.qspi.r_count[0] ),
    .X(_09941_));
 sg13g2_buf_2 _16689_ (.A(\cpu.qspi.r_count[1] ),
    .X(_09942_));
 sg13g2_buf_1 _16690_ (.A(\cpu.qspi.r_count[2] ),
    .X(_09943_));
 sg13g2_nor4_2 _16691_ (.A(_09941_),
    .B(_09942_),
    .C(_09943_),
    .Y(_09944_),
    .D(\cpu.qspi.r_count[3] ));
 sg13g2_and2_1 _16692_ (.A(_09940_),
    .B(_09944_),
    .X(_09945_));
 sg13g2_buf_1 _16693_ (.A(_09945_),
    .X(_09946_));
 sg13g2_buf_2 _16694_ (.A(\cpu.qspi.r_state[2] ),
    .X(_09947_));
 sg13g2_buf_1 _16695_ (.A(\cpu.qspi.r_state[1] ),
    .X(_09948_));
 sg13g2_a221oi_1 _16696_ (.B2(_09947_),
    .C1(_09948_),
    .B1(_09946_),
    .A1(_09938_),
    .Y(_09949_),
    .A2(_09939_));
 sg13g2_a21oi_1 _16697_ (.A1(_09937_),
    .A2(_09949_),
    .Y(_00026_),
    .B1(net630));
 sg13g2_buf_1 _16698_ (.A(\cpu.qspi.r_state[16] ),
    .X(_09950_));
 sg13g2_nand2_1 _16699_ (.Y(_09951_),
    .A(_09940_),
    .B(_09944_));
 sg13g2_buf_1 _16700_ (.A(_09951_),
    .X(_09952_));
 sg13g2_nand2_1 _16701_ (.Y(_09953_),
    .A(_09950_),
    .B(net788));
 sg13g2_buf_2 _16702_ (.A(\cpu.qspi.r_state[8] ),
    .X(_09954_));
 sg13g2_nand2_1 _16703_ (.Y(_09955_),
    .A(net802),
    .B(_09930_));
 sg13g2_buf_2 _16704_ (.A(_09955_),
    .X(_09956_));
 sg13g2_inv_1 _16705_ (.Y(_09957_),
    .A(_09956_));
 sg13g2_nand2_1 _16706_ (.Y(_09958_),
    .A(_09954_),
    .B(_09957_));
 sg13g2_a21oi_1 _16707_ (.A1(_09953_),
    .A2(_09958_),
    .Y(_00025_),
    .B1(net630));
 sg13g2_buf_1 _16708_ (.A(\cpu.qspi.r_state[4] ),
    .X(_09959_));
 sg13g2_buf_1 _16709_ (.A(\cpu.qspi.r_state[9] ),
    .X(_09960_));
 sg13g2_a21oi_1 _16710_ (.A1(_09959_),
    .A2(_09946_),
    .Y(_09961_),
    .B1(_09960_));
 sg13g2_nor2_1 _16711_ (.A(net631),
    .B(_09961_),
    .Y(_00022_));
 sg13g2_buf_1 _16712_ (.A(\cpu.qspi.r_state[12] ),
    .X(_09962_));
 sg13g2_buf_1 _16713_ (.A(_09962_),
    .X(_09963_));
 sg13g2_inv_1 _16714_ (.Y(_09964_),
    .A(_00277_));
 sg13g2_a21oi_1 _16715_ (.A1(net1047),
    .A2(net788),
    .Y(_09965_),
    .B1(_09964_));
 sg13g2_nor2_1 _16716_ (.A(net631),
    .B(_09965_),
    .Y(_00023_));
 sg13g2_inv_1 _16717_ (.Y(_09966_),
    .A(\cpu.qspi.r_rom_mode[1] ));
 sg13g2_buf_1 _16718_ (.A(\cpu.qspi.r_rom_mode[0] ),
    .X(_09967_));
 sg13g2_inv_1 _16719_ (.Y(_09968_),
    .A(_09609_));
 sg13g2_or2_1 _16720_ (.X(_09969_),
    .B(_08874_),
    .A(net802));
 sg13g2_o21ai_1 _16721_ (.B1(_09969_),
    .Y(_09970_),
    .A1(net1069),
    .A2(_09968_));
 sg13g2_inv_1 _16722_ (.Y(_09971_),
    .A(_09970_));
 sg13g2_nor2_1 _16723_ (.A(_09967_),
    .B(_09971_),
    .Y(_09972_));
 sg13g2_a21oi_1 _16724_ (.A1(_09967_),
    .A2(_09956_),
    .Y(_09973_),
    .B1(_09972_));
 sg13g2_nor2_1 _16725_ (.A(_09966_),
    .B(_09973_),
    .Y(_09974_));
 sg13g2_buf_2 _16726_ (.A(_09974_),
    .X(_09975_));
 sg13g2_nor3_1 _16727_ (.A(_09967_),
    .B(\cpu.qspi.r_rom_mode[1] ),
    .C(_09971_),
    .Y(_09976_));
 sg13g2_buf_2 _16728_ (.A(_09976_),
    .X(_09977_));
 sg13g2_nor2_1 _16729_ (.A(_09977_),
    .B(_09975_),
    .Y(_09978_));
 sg13g2_buf_2 _16730_ (.A(_09978_),
    .X(_09979_));
 sg13g2_and2_1 _16731_ (.A(\cpu.qspi.r_quad[2] ),
    .B(_09977_),
    .X(_09980_));
 sg13g2_a221oi_1 _16732_ (.B2(\cpu.qspi.r_quad[0] ),
    .C1(_09980_),
    .B1(_09979_),
    .A1(\cpu.qspi.r_quad[1] ),
    .Y(_09981_),
    .A2(_09975_));
 sg13g2_buf_2 _16733_ (.A(_09981_),
    .X(_09982_));
 sg13g2_nand2_1 _16734_ (.Y(_09983_),
    .A(\cpu.qspi.r_state[17] ),
    .B(_09935_));
 sg13g2_inv_1 _16735_ (.Y(_09984_),
    .A(_09983_));
 sg13g2_a22oi_1 _16736_ (.Y(_09985_),
    .B1(_09982_),
    .B2(_09984_),
    .A2(net788),
    .A1(_09959_));
 sg13g2_nor2_1 _16737_ (.A(net631),
    .B(_09985_),
    .Y(_00028_));
 sg13g2_nand2_1 _16738_ (.Y(_09986_),
    .A(_09947_),
    .B(_09952_));
 sg13g2_buf_1 _16739_ (.A(\cpu.qspi.r_state[14] ),
    .X(_09987_));
 sg13g2_nand2_1 _16740_ (.Y(_09988_),
    .A(net1119),
    .B(_09946_));
 sg13g2_a21oi_1 _16741_ (.A1(_09986_),
    .A2(_09988_),
    .Y(_00027_),
    .B1(net630));
 sg13g2_inv_1 _16742_ (.Y(_09989_),
    .A(_09938_));
 sg13g2_buf_1 _16743_ (.A(net803),
    .X(_09990_));
 sg13g2_o21ai_1 _16744_ (.B1(net685),
    .Y(_00021_),
    .A1(_09989_),
    .A2(_09939_));
 sg13g2_buf_1 _16745_ (.A(\cpu.dec.r_op[10] ),
    .X(_09991_));
 sg13g2_buf_1 _16746_ (.A(_09991_),
    .X(_09992_));
 sg13g2_inv_1 _16747_ (.Y(_09993_),
    .A(net1046));
 sg13g2_buf_1 _16748_ (.A(_08972_),
    .X(_09994_));
 sg13g2_nor2_1 _16749_ (.A(_09101_),
    .B(_09116_),
    .Y(_09995_));
 sg13g2_nand3_1 _16750_ (.B(_09084_),
    .C(_09995_),
    .A(_08974_),
    .Y(_09996_));
 sg13g2_o21ai_1 _16751_ (.B1(_09996_),
    .Y(_00011_),
    .A1(_09993_),
    .A2(net118));
 sg13g2_buf_2 _16752_ (.A(\cpu.dec.r_op[1] ),
    .X(_09997_));
 sg13g2_buf_1 _16753_ (.A(_09169_),
    .X(_09998_));
 sg13g2_nand2_1 _16754_ (.Y(_09999_),
    .A(_09154_),
    .B(_09259_));
 sg13g2_inv_1 _16755_ (.Y(_10000_),
    .A(_09999_));
 sg13g2_inv_1 _16756_ (.Y(_10001_),
    .A(_09222_));
 sg13g2_a21o_1 _16757_ (.A2(_08988_),
    .A1(_08978_),
    .B1(_08996_),
    .X(_10002_));
 sg13g2_buf_2 _16758_ (.A(_10002_),
    .X(_10003_));
 sg13g2_nor2_1 _16759_ (.A(_10003_),
    .B(_09018_),
    .Y(_10004_));
 sg13g2_buf_1 _16760_ (.A(_10004_),
    .X(_10005_));
 sg13g2_nand2_1 _16761_ (.Y(_10006_),
    .A(net150),
    .B(net209));
 sg13g2_nor2_1 _16762_ (.A(_10001_),
    .B(_10006_),
    .Y(_10007_));
 sg13g2_inv_2 _16763_ (.Y(_10008_),
    .A(net210));
 sg13g2_nor3_1 _16764_ (.A(net281),
    .B(_09151_),
    .C(_10008_),
    .Y(_10009_));
 sg13g2_a22oi_1 _16765_ (.Y(_10010_),
    .B1(_10009_),
    .B2(_09202_),
    .A2(_10007_),
    .A1(_10000_));
 sg13g2_nor3_1 _16766_ (.A(net106),
    .B(net152),
    .C(_10010_),
    .Y(_10011_));
 sg13g2_a21o_1 _16767_ (.A2(net92),
    .A1(_09997_),
    .B1(_10011_),
    .X(_00012_));
 sg13g2_buf_1 _16768_ (.A(_08998_),
    .X(_10012_));
 sg13g2_buf_1 _16769_ (.A(_09116_),
    .X(_10013_));
 sg13g2_buf_1 _16770_ (.A(net240),
    .X(_10014_));
 sg13g2_buf_1 _16771_ (.A(_10014_),
    .X(_10015_));
 sg13g2_nand3_1 _16772_ (.B(net238),
    .C(_10009_),
    .A(net177),
    .Y(_10016_));
 sg13g2_o21ai_1 _16773_ (.B1(_10016_),
    .Y(_10017_),
    .A1(net177),
    .A2(net238));
 sg13g2_nand4_1 _16774_ (.B(net179),
    .C(_10013_),
    .A(_10012_),
    .Y(_10018_),
    .D(_10017_));
 sg13g2_buf_1 _16775_ (.A(\cpu.dec.r_op[9] ),
    .X(_10019_));
 sg13g2_buf_1 _16776_ (.A(_10019_),
    .X(_10020_));
 sg13g2_buf_1 _16777_ (.A(net108),
    .X(_10021_));
 sg13g2_nand2_1 _16778_ (.Y(_10022_),
    .A(net1045),
    .B(net89));
 sg13g2_o21ai_1 _16779_ (.B1(_10022_),
    .Y(_00020_),
    .A1(net92),
    .A2(_10018_));
 sg13g2_buf_1 _16780_ (.A(\cpu.dec.r_op[8] ),
    .X(_10023_));
 sg13g2_inv_1 _16781_ (.Y(_10024_),
    .A(net1118));
 sg13g2_buf_1 _16782_ (.A(_09058_),
    .X(_10025_));
 sg13g2_a21oi_1 _16783_ (.A1(net936),
    .A2(_09070_),
    .Y(_10026_),
    .B1(_09077_));
 sg13g2_nand2_1 _16784_ (.Y(_10027_),
    .A(net280),
    .B(_10026_));
 sg13g2_buf_1 _16785_ (.A(_10027_),
    .X(_10028_));
 sg13g2_nor2_1 _16786_ (.A(net279),
    .B(_10028_),
    .Y(_10029_));
 sg13g2_buf_1 _16787_ (.A(_10029_),
    .X(_10030_));
 sg13g2_nor2_1 _16788_ (.A(_08998_),
    .B(_09018_),
    .Y(_10031_));
 sg13g2_buf_2 _16789_ (.A(_10031_),
    .X(_10032_));
 sg13g2_nand3_1 _16790_ (.B(_10030_),
    .C(_10032_),
    .A(net119),
    .Y(_10033_));
 sg13g2_o21ai_1 _16791_ (.B1(_10033_),
    .Y(_00019_),
    .A1(net1044),
    .A2(net118));
 sg13g2_buf_1 _16792_ (.A(\cpu.qspi.r_state[5] ),
    .X(_10034_));
 sg13g2_a21oi_1 _16793_ (.A1(net1119),
    .A2(net788),
    .Y(_10035_),
    .B1(_10034_));
 sg13g2_nor2_1 _16794_ (.A(net631),
    .B(_10035_),
    .Y(_00024_));
 sg13g2_buf_1 _16795_ (.A(\cpu.dec.r_op[2] ),
    .X(_10036_));
 sg13g2_buf_1 _16796_ (.A(net1117),
    .X(_10037_));
 sg13g2_inv_1 _16797_ (.Y(_10038_),
    .A(net1043));
 sg13g2_o21ai_1 _16798_ (.B1(_09102_),
    .Y(_10039_),
    .A1(net281),
    .A2(_09205_));
 sg13g2_nand4_1 _16799_ (.B(_09084_),
    .C(net208),
    .A(_08974_),
    .Y(_10040_),
    .D(_10039_));
 sg13g2_o21ai_1 _16800_ (.B1(_10040_),
    .Y(_00013_),
    .A1(_10038_),
    .A2(_09994_));
 sg13g2_nor3_1 _16801_ (.A(net152),
    .B(net151),
    .C(_09999_),
    .Y(_10041_));
 sg13g2_nor2_1 _16802_ (.A(_09222_),
    .B(net209),
    .Y(_10042_));
 sg13g2_nor3_1 _16803_ (.A(net281),
    .B(_09203_),
    .C(_09205_),
    .Y(_10043_));
 sg13g2_a21oi_1 _16804_ (.A1(_10041_),
    .A2(_10042_),
    .Y(_10044_),
    .B1(_10043_));
 sg13g2_buf_1 _16805_ (.A(\cpu.dec.r_op[7] ),
    .X(_10045_));
 sg13g2_nand2_1 _16806_ (.Y(_10046_),
    .A(_10045_),
    .B(_10021_));
 sg13g2_o21ai_1 _16807_ (.B1(_10046_),
    .Y(_00018_),
    .A1(_09171_),
    .A2(_10044_));
 sg13g2_buf_1 _16808_ (.A(\cpu.uart.r_div[11] ),
    .X(_10047_));
 sg13g2_nor3_1 _16809_ (.A(\cpu.uart.r_div[0] ),
    .B(\cpu.uart.r_div[1] ),
    .C(\cpu.uart.r_div[2] ),
    .Y(_10048_));
 sg13g2_nor2b_1 _16810_ (.A(\cpu.uart.r_div[3] ),
    .B_N(_10048_),
    .Y(_10049_));
 sg13g2_nor2b_1 _16811_ (.A(\cpu.uart.r_div[4] ),
    .B_N(_10049_),
    .Y(_10050_));
 sg13g2_nor2b_1 _16812_ (.A(\cpu.uart.r_div[5] ),
    .B_N(_10050_),
    .Y(_10051_));
 sg13g2_nor2b_1 _16813_ (.A(\cpu.uart.r_div[6] ),
    .B_N(_10051_),
    .Y(_10052_));
 sg13g2_nand2b_1 _16814_ (.Y(_10053_),
    .B(_10052_),
    .A_N(\cpu.uart.r_div[7] ));
 sg13g2_nor2_1 _16815_ (.A(\cpu.uart.r_div[8] ),
    .B(_10053_),
    .Y(_10054_));
 sg13g2_nand2b_1 _16816_ (.Y(_10055_),
    .B(_10054_),
    .A_N(\cpu.uart.r_div[9] ));
 sg13g2_buf_1 _16817_ (.A(_10055_),
    .X(_10056_));
 sg13g2_nor3_1 _16818_ (.A(_10047_),
    .B(\cpu.uart.r_div[10] ),
    .C(_10056_),
    .Y(_10057_));
 sg13g2_buf_1 _16819_ (.A(_10057_),
    .X(_10058_));
 sg13g2_nor2_1 _16820_ (.A(net931),
    .B(net348),
    .Y(_10059_));
 sg13g2_buf_1 _16821_ (.A(_10059_),
    .X(_10060_));
 sg13g2_buf_1 _16822_ (.A(_10060_),
    .X(_10061_));
 sg13g2_mux2_1 _16823_ (.A0(\cpu.uart.r_div_value[0] ),
    .A1(_00279_),
    .S(net205),
    .X(_00079_));
 sg13g2_xnor2_1 _16824_ (.Y(_10062_),
    .A(\cpu.uart.r_div[0] ),
    .B(\cpu.uart.r_div[1] ));
 sg13g2_mux2_1 _16825_ (.A0(\cpu.uart.r_div_value[1] ),
    .A1(_10062_),
    .S(net205),
    .X(_00082_));
 sg13g2_o21ai_1 _16826_ (.B1(\cpu.uart.r_div[2] ),
    .Y(_10063_),
    .A1(\cpu.uart.r_div[0] ),
    .A2(\cpu.uart.r_div[1] ));
 sg13g2_nor2b_1 _16827_ (.A(_10048_),
    .B_N(_10063_),
    .Y(_10064_));
 sg13g2_nor2_1 _16828_ (.A(\cpu.uart.r_div_value[2] ),
    .B(net237),
    .Y(_10065_));
 sg13g2_a21oi_1 _16829_ (.A1(_10061_),
    .A2(_10064_),
    .Y(_00083_),
    .B1(_10065_));
 sg13g2_xnor2_1 _16830_ (.Y(_10066_),
    .A(\cpu.uart.r_div[3] ),
    .B(_10048_));
 sg13g2_nor2_1 _16831_ (.A(\cpu.uart.r_div_value[3] ),
    .B(net237),
    .Y(_10067_));
 sg13g2_a21oi_1 _16832_ (.A1(_10061_),
    .A2(_10066_),
    .Y(_00084_),
    .B1(_10067_));
 sg13g2_xnor2_1 _16833_ (.Y(_10068_),
    .A(\cpu.uart.r_div[4] ),
    .B(_10049_));
 sg13g2_nor2_1 _16834_ (.A(\cpu.uart.r_div_value[4] ),
    .B(net237),
    .Y(_10069_));
 sg13g2_a21oi_1 _16835_ (.A1(net205),
    .A2(_10068_),
    .Y(_00085_),
    .B1(_10069_));
 sg13g2_xnor2_1 _16836_ (.Y(_10070_),
    .A(\cpu.uart.r_div[5] ),
    .B(_10050_));
 sg13g2_nor2_1 _16837_ (.A(\cpu.uart.r_div_value[5] ),
    .B(net237),
    .Y(_10071_));
 sg13g2_a21oi_1 _16838_ (.A1(net205),
    .A2(_10070_),
    .Y(_00086_),
    .B1(_10071_));
 sg13g2_xnor2_1 _16839_ (.Y(_10072_),
    .A(\cpu.uart.r_div[6] ),
    .B(_10051_));
 sg13g2_nor2_1 _16840_ (.A(\cpu.uart.r_div_value[6] ),
    .B(net237),
    .Y(_10073_));
 sg13g2_a21oi_1 _16841_ (.A1(net205),
    .A2(_10072_),
    .Y(_00087_),
    .B1(_10073_));
 sg13g2_xnor2_1 _16842_ (.Y(_10074_),
    .A(\cpu.uart.r_div[7] ),
    .B(_10052_));
 sg13g2_nor2_1 _16843_ (.A(\cpu.uart.r_div_value[7] ),
    .B(net237),
    .Y(_10075_));
 sg13g2_a21oi_1 _16844_ (.A1(net205),
    .A2(_10074_),
    .Y(_00088_),
    .B1(_10075_));
 sg13g2_xor2_1 _16845_ (.B(_10053_),
    .A(\cpu.uart.r_div[8] ),
    .X(_10076_));
 sg13g2_nor2_1 _16846_ (.A(\cpu.uart.r_div_value[8] ),
    .B(net237),
    .Y(_10077_));
 sg13g2_a21oi_1 _16847_ (.A1(net205),
    .A2(_10076_),
    .Y(_00089_),
    .B1(_10077_));
 sg13g2_xnor2_1 _16848_ (.Y(_10078_),
    .A(\cpu.uart.r_div[9] ),
    .B(_10054_));
 sg13g2_nor2_1 _16849_ (.A(\cpu.uart.r_div_value[9] ),
    .B(net237),
    .Y(_10079_));
 sg13g2_a21oi_1 _16850_ (.A1(net205),
    .A2(_10078_),
    .Y(_00090_),
    .B1(_10079_));
 sg13g2_buf_1 _16851_ (.A(\cpu.uart.r_div_value[10] ),
    .X(_10080_));
 sg13g2_inv_1 _16852_ (.Y(_10081_),
    .A(_10080_));
 sg13g2_nand2_1 _16853_ (.Y(_10082_),
    .A(net803),
    .B(_10056_));
 sg13g2_o21ai_1 _16854_ (.B1(_10082_),
    .Y(_10083_),
    .A1(_10047_),
    .A2(_10080_));
 sg13g2_inv_1 _16855_ (.Y(_10084_),
    .A(\cpu.uart.r_div[10] ));
 sg13g2_nor3_1 _16856_ (.A(_10084_),
    .B(net804),
    .C(_10056_),
    .Y(_10085_));
 sg13g2_a221oi_1 _16857_ (.B2(_10084_),
    .C1(_10085_),
    .B1(_10083_),
    .A1(_10081_),
    .Y(_00080_),
    .A2(net707));
 sg13g2_nor2_1 _16858_ (.A(\cpu.uart.r_div[10] ),
    .B(_10056_),
    .Y(_10086_));
 sg13g2_nand2_1 _16859_ (.Y(_10087_),
    .A(_10047_),
    .B(net706));
 sg13g2_o21ai_1 _16860_ (.B1(\cpu.uart.r_div_value[11] ),
    .Y(_10088_),
    .A1(net804),
    .A2(net348));
 sg13g2_o21ai_1 _16861_ (.B1(_10088_),
    .Y(_00081_),
    .A1(_10086_),
    .A2(_10087_));
 sg13g2_buf_1 _16862_ (.A(\cpu.intr.r_timer_count[14] ),
    .X(_10089_));
 sg13g2_buf_1 _16863_ (.A(\cpu.intr.r_timer_count[11] ),
    .X(_10090_));
 sg13g2_buf_1 _16864_ (.A(\cpu.intr.r_timer_count[8] ),
    .X(_10091_));
 sg13g2_buf_2 _16865_ (.A(\cpu.intr.r_timer_count[1] ),
    .X(_10092_));
 sg13g2_nor3_1 _16866_ (.A(_10092_),
    .B(\cpu.intr.r_timer_count[0] ),
    .C(\cpu.intr.r_timer_count[2] ),
    .Y(_10093_));
 sg13g2_nor2b_1 _16867_ (.A(\cpu.intr.r_timer_count[3] ),
    .B_N(_10093_),
    .Y(_10094_));
 sg13g2_nor2b_1 _16868_ (.A(\cpu.intr.r_timer_count[4] ),
    .B_N(_10094_),
    .Y(_10095_));
 sg13g2_nor2b_1 _16869_ (.A(\cpu.intr.r_timer_count[5] ),
    .B_N(_10095_),
    .Y(_10096_));
 sg13g2_nor2b_1 _16870_ (.A(\cpu.intr.r_timer_count[6] ),
    .B_N(_10096_),
    .Y(_10097_));
 sg13g2_nand2b_1 _16871_ (.Y(_10098_),
    .B(_10097_),
    .A_N(\cpu.intr.r_timer_count[7] ));
 sg13g2_nor3_2 _16872_ (.A(\cpu.intr.r_timer_count[9] ),
    .B(_10091_),
    .C(_10098_),
    .Y(_10099_));
 sg13g2_nand2b_1 _16873_ (.Y(_10100_),
    .B(_10099_),
    .A_N(\cpu.intr.r_timer_count[10] ));
 sg13g2_nor3_2 _16874_ (.A(_10090_),
    .B(\cpu.intr.r_timer_count[12] ),
    .C(_10100_),
    .Y(_10101_));
 sg13g2_nand2b_1 _16875_ (.Y(_10102_),
    .B(_10101_),
    .A_N(\cpu.intr.r_timer_count[13] ));
 sg13g2_nor3_2 _16876_ (.A(\cpu.intr.r_timer_count[15] ),
    .B(_10089_),
    .C(_10102_),
    .Y(_10103_));
 sg13g2_buf_1 _16877_ (.A(\cpu.intr.r_timer_count[17] ),
    .X(_10104_));
 sg13g2_buf_1 _16878_ (.A(\cpu.intr.r_timer_count[16] ),
    .X(_10105_));
 sg13g2_buf_1 _16879_ (.A(\cpu.intr.r_timer_count[23] ),
    .X(_10106_));
 sg13g2_buf_1 _16880_ (.A(\cpu.intr.r_timer_count[18] ),
    .X(_10107_));
 sg13g2_buf_1 _16881_ (.A(\cpu.intr.r_timer_count[19] ),
    .X(_10108_));
 sg13g2_buf_1 _16882_ (.A(\cpu.intr.r_timer_count[20] ),
    .X(_10109_));
 sg13g2_nor4_1 _16883_ (.A(_10107_),
    .B(_10108_),
    .C(_10109_),
    .D(\cpu.intr.r_timer_count[21] ),
    .Y(_10110_));
 sg13g2_nand2b_1 _16884_ (.Y(_10111_),
    .B(_10110_),
    .A_N(\cpu.intr.r_timer_count[22] ));
 sg13g2_nor4_2 _16885_ (.A(_10104_),
    .B(_10105_),
    .C(_10106_),
    .Y(_10112_),
    .D(_10111_));
 sg13g2_nand2_1 _16886_ (.Y(_10113_),
    .A(_10103_),
    .B(_10112_));
 sg13g2_buf_2 _16887_ (.A(_10113_),
    .X(_10114_));
 sg13g2_buf_1 _16888_ (.A(net1051),
    .X(_10115_));
 sg13g2_buf_1 _16889_ (.A(_10115_),
    .X(_10116_));
 sg13g2_buf_1 _16890_ (.A(net787),
    .X(_10117_));
 sg13g2_buf_1 _16891_ (.A(net699),
    .X(_10118_));
 sg13g2_buf_1 _16892_ (.A(net621),
    .X(_10119_));
 sg13g2_buf_1 _16893_ (.A(net545),
    .X(_10120_));
 sg13g2_buf_1 _16894_ (.A(net494),
    .X(_10121_));
 sg13g2_buf_1 _16895_ (.A(\cpu.addr[5] ),
    .X(_10122_));
 sg13g2_buf_1 _16896_ (.A(_10122_),
    .X(_10123_));
 sg13g2_nor3_2 _16897_ (.A(net1042),
    .B(net1056),
    .C(_09280_),
    .Y(_10124_));
 sg13g2_nand2_1 _16898_ (.Y(_10125_),
    .A(_09277_),
    .B(_10124_));
 sg13g2_buf_1 _16899_ (.A(_10125_),
    .X(_10126_));
 sg13g2_nor2_1 _16900_ (.A(_09368_),
    .B(net683),
    .Y(_10127_));
 sg13g2_buf_1 _16901_ (.A(_10127_),
    .X(_10128_));
 sg13g2_nand3_1 _16902_ (.B(net445),
    .C(_10128_),
    .A(net684),
    .Y(_10129_));
 sg13g2_buf_2 _16903_ (.A(_10129_),
    .X(_10130_));
 sg13g2_nand2_1 _16904_ (.Y(_10131_),
    .A(_10114_),
    .B(_10130_));
 sg13g2_buf_1 _16905_ (.A(_10131_),
    .X(_10132_));
 sg13g2_buf_1 _16906_ (.A(_10132_),
    .X(_10133_));
 sg13g2_mux2_1 _16907_ (.A0(_00285_),
    .A1(\cpu.intr.r_timer_reload[0] ),
    .S(_10133_),
    .X(_00055_));
 sg13g2_buf_1 _16908_ (.A(_10132_),
    .X(_10134_));
 sg13g2_xor2_1 _16909_ (.B(\cpu.intr.r_timer_count[0] ),
    .A(_10092_),
    .X(_10135_));
 sg13g2_nand2_1 _16910_ (.Y(_10136_),
    .A(\cpu.intr.r_timer_reload[1] ),
    .B(_10133_));
 sg13g2_o21ai_1 _16911_ (.B1(_10136_),
    .Y(_00066_),
    .A1(net75),
    .A2(_10135_));
 sg13g2_o21ai_1 _16912_ (.B1(\cpu.intr.r_timer_count[2] ),
    .Y(_10137_),
    .A1(_10092_),
    .A2(\cpu.intr.r_timer_count[0] ));
 sg13g2_nor2b_1 _16913_ (.A(_10093_),
    .B_N(_10137_),
    .Y(_10138_));
 sg13g2_nand2_1 _16914_ (.Y(_10139_),
    .A(\cpu.intr.r_timer_reload[2] ),
    .B(net76));
 sg13g2_o21ai_1 _16915_ (.B1(_10139_),
    .Y(_00071_),
    .A1(_10134_),
    .A2(_10138_));
 sg13g2_xnor2_1 _16916_ (.Y(_10140_),
    .A(\cpu.intr.r_timer_count[3] ),
    .B(_10093_));
 sg13g2_nand2_1 _16917_ (.Y(_10141_),
    .A(\cpu.intr.r_timer_reload[3] ),
    .B(net76));
 sg13g2_o21ai_1 _16918_ (.B1(_10141_),
    .Y(_00072_),
    .A1(net75),
    .A2(_10140_));
 sg13g2_xnor2_1 _16919_ (.Y(_10142_),
    .A(\cpu.intr.r_timer_count[4] ),
    .B(_10094_));
 sg13g2_nand2_1 _16920_ (.Y(_10143_),
    .A(\cpu.intr.r_timer_reload[4] ),
    .B(net76));
 sg13g2_o21ai_1 _16921_ (.B1(_10143_),
    .Y(_00073_),
    .A1(net75),
    .A2(_10142_));
 sg13g2_xnor2_1 _16922_ (.Y(_10144_),
    .A(\cpu.intr.r_timer_count[5] ),
    .B(_10095_));
 sg13g2_buf_1 _16923_ (.A(_10132_),
    .X(_10145_));
 sg13g2_nand2_1 _16924_ (.Y(_10146_),
    .A(\cpu.intr.r_timer_reload[5] ),
    .B(net74));
 sg13g2_o21ai_1 _16925_ (.B1(_10146_),
    .Y(_00074_),
    .A1(net75),
    .A2(_10144_));
 sg13g2_xnor2_1 _16926_ (.Y(_10147_),
    .A(\cpu.intr.r_timer_count[6] ),
    .B(_10096_));
 sg13g2_nand2_1 _16927_ (.Y(_10148_),
    .A(\cpu.intr.r_timer_reload[6] ),
    .B(net74));
 sg13g2_o21ai_1 _16928_ (.B1(_10148_),
    .Y(_00075_),
    .A1(_10134_),
    .A2(_10147_));
 sg13g2_xnor2_1 _16929_ (.Y(_10149_),
    .A(\cpu.intr.r_timer_count[7] ),
    .B(_10097_));
 sg13g2_nand2_1 _16930_ (.Y(_10150_),
    .A(\cpu.intr.r_timer_reload[7] ),
    .B(_10145_));
 sg13g2_o21ai_1 _16931_ (.B1(_10150_),
    .Y(_00076_),
    .A1(net75),
    .A2(_10149_));
 sg13g2_xor2_1 _16932_ (.B(_10098_),
    .A(_10091_),
    .X(_10151_));
 sg13g2_nand2_1 _16933_ (.Y(_10152_),
    .A(\cpu.intr.r_timer_reload[8] ),
    .B(net74));
 sg13g2_o21ai_1 _16934_ (.B1(_10152_),
    .Y(_00077_),
    .A1(net75),
    .A2(_10151_));
 sg13g2_o21ai_1 _16935_ (.B1(\cpu.intr.r_timer_count[9] ),
    .Y(_10153_),
    .A1(_10091_),
    .A2(_10098_));
 sg13g2_nor2b_1 _16936_ (.A(_10099_),
    .B_N(_10153_),
    .Y(_10154_));
 sg13g2_nand2_1 _16937_ (.Y(_10155_),
    .A(\cpu.intr.r_timer_reload[9] ),
    .B(_10145_));
 sg13g2_o21ai_1 _16938_ (.B1(_10155_),
    .Y(_00078_),
    .A1(net75),
    .A2(_10154_));
 sg13g2_xnor2_1 _16939_ (.Y(_10156_),
    .A(\cpu.intr.r_timer_count[10] ),
    .B(_10099_));
 sg13g2_nand2_1 _16940_ (.Y(_10157_),
    .A(\cpu.intr.r_timer_reload[10] ),
    .B(net74));
 sg13g2_o21ai_1 _16941_ (.B1(_10157_),
    .Y(_00056_),
    .A1(net75),
    .A2(_10156_));
 sg13g2_xor2_1 _16942_ (.B(_10100_),
    .A(_10090_),
    .X(_10158_));
 sg13g2_nand2_1 _16943_ (.Y(_10159_),
    .A(\cpu.intr.r_timer_reload[11] ),
    .B(net74));
 sg13g2_o21ai_1 _16944_ (.B1(_10159_),
    .Y(_00057_),
    .A1(net76),
    .A2(_10158_));
 sg13g2_o21ai_1 _16945_ (.B1(\cpu.intr.r_timer_count[12] ),
    .Y(_10160_),
    .A1(_10090_),
    .A2(_10100_));
 sg13g2_nor2b_1 _16946_ (.A(_10101_),
    .B_N(_10160_),
    .Y(_10161_));
 sg13g2_nand2_1 _16947_ (.Y(_10162_),
    .A(\cpu.intr.r_timer_reload[12] ),
    .B(net74));
 sg13g2_o21ai_1 _16948_ (.B1(_10162_),
    .Y(_00058_),
    .A1(net76),
    .A2(_10161_));
 sg13g2_xnor2_1 _16949_ (.Y(_10163_),
    .A(\cpu.intr.r_timer_count[13] ),
    .B(_10101_));
 sg13g2_nand2_1 _16950_ (.Y(_10164_),
    .A(\cpu.intr.r_timer_reload[13] ),
    .B(net74));
 sg13g2_o21ai_1 _16951_ (.B1(_10164_),
    .Y(_00059_),
    .A1(net76),
    .A2(_10163_));
 sg13g2_xor2_1 _16952_ (.B(_10102_),
    .A(_10089_),
    .X(_10165_));
 sg13g2_nand2_1 _16953_ (.Y(_10166_),
    .A(\cpu.intr.r_timer_reload[14] ),
    .B(net74));
 sg13g2_o21ai_1 _16954_ (.B1(_10166_),
    .Y(_00060_),
    .A1(net76),
    .A2(_10165_));
 sg13g2_o21ai_1 _16955_ (.B1(\cpu.intr.r_timer_count[15] ),
    .Y(_10167_),
    .A1(_10089_),
    .A2(_10102_));
 sg13g2_nor2b_1 _16956_ (.A(_10103_),
    .B_N(_10167_),
    .Y(_10168_));
 sg13g2_nand2_1 _16957_ (.Y(_10169_),
    .A(\cpu.intr.r_timer_reload[15] ),
    .B(_10132_));
 sg13g2_o21ai_1 _16958_ (.B1(_10169_),
    .Y(_00061_),
    .A1(net76),
    .A2(_10168_));
 sg13g2_buf_1 _16959_ (.A(net933),
    .X(_10170_));
 sg13g2_buf_1 _16960_ (.A(net786),
    .X(_10171_));
 sg13g2_buf_1 _16961_ (.A(net682),
    .X(_10172_));
 sg13g2_buf_1 _16962_ (.A(net805),
    .X(_10173_));
 sg13g2_buf_1 _16963_ (.A(net681),
    .X(_10174_));
 sg13g2_buf_1 _16964_ (.A(net1048),
    .X(_10175_));
 sg13g2_buf_1 _16965_ (.A(net922),
    .X(_10176_));
 sg13g2_nand3_1 _16966_ (.B(net785),
    .C(net496),
    .A(net619),
    .Y(_10177_));
 sg13g2_buf_1 _16967_ (.A(_10177_),
    .X(_10178_));
 sg13g2_nor4_1 _16968_ (.A(net620),
    .B(_09368_),
    .C(_10178_),
    .D(_10126_),
    .Y(_10179_));
 sg13g2_buf_1 _16969_ (.A(_10179_),
    .X(_10180_));
 sg13g2_buf_1 _16970_ (.A(_10180_),
    .X(_10181_));
 sg13g2_inv_1 _16971_ (.Y(_10182_),
    .A(\cpu.intr.r_timer_reload[16] ));
 sg13g2_a21oi_1 _16972_ (.A1(_10182_),
    .A2(_10112_),
    .Y(_10183_),
    .B1(_10105_));
 sg13g2_nor2b_1 _16973_ (.A(_10103_),
    .B_N(_10105_),
    .Y(_10184_));
 sg13g2_a21oi_1 _16974_ (.A1(_10103_),
    .A2(_10183_),
    .Y(_10185_),
    .B1(_10184_));
 sg13g2_buf_1 _16975_ (.A(\cpu.dcache.wdata[0] ),
    .X(_10186_));
 sg13g2_buf_1 _16976_ (.A(_10186_),
    .X(_10187_));
 sg13g2_nand2_1 _16977_ (.Y(_10188_),
    .A(_10187_),
    .B(net148));
 sg13g2_o21ai_1 _16978_ (.B1(_10188_),
    .Y(_00062_),
    .A1(net133),
    .A2(_10185_));
 sg13g2_nand2b_1 _16979_ (.Y(_10189_),
    .B(_10112_),
    .A_N(\cpu.intr.r_timer_reload[17] ));
 sg13g2_nor2b_1 _16980_ (.A(_10105_),
    .B_N(_10103_),
    .Y(_10190_));
 sg13g2_nor2b_1 _16981_ (.A(_10104_),
    .B_N(_10190_),
    .Y(_10191_));
 sg13g2_nor2b_1 _16982_ (.A(_10190_),
    .B_N(_10104_),
    .Y(_10192_));
 sg13g2_a21oi_1 _16983_ (.A1(_10189_),
    .A2(_10191_),
    .Y(_10193_),
    .B1(_10192_));
 sg13g2_buf_2 _16984_ (.A(\cpu.dcache.wdata[1] ),
    .X(_10194_));
 sg13g2_buf_1 _16985_ (.A(_10194_),
    .X(_10195_));
 sg13g2_buf_1 _16986_ (.A(_10195_),
    .X(_10196_));
 sg13g2_nand2_1 _16987_ (.Y(_10197_),
    .A(net921),
    .B(net148));
 sg13g2_o21ai_1 _16988_ (.B1(_10197_),
    .Y(_00063_),
    .A1(net133),
    .A2(_10193_));
 sg13g2_xnor2_1 _16989_ (.Y(_10198_),
    .A(_10107_),
    .B(_10191_));
 sg13g2_o21ai_1 _16990_ (.B1(_10130_),
    .Y(_10199_),
    .A1(\cpu.intr.r_timer_reload[18] ),
    .A2(_10114_));
 sg13g2_buf_1 _16991_ (.A(\cpu.dcache.wdata[2] ),
    .X(_10200_));
 sg13g2_buf_1 _16992_ (.A(_10200_),
    .X(_10201_));
 sg13g2_buf_1 _16993_ (.A(net1039),
    .X(_10202_));
 sg13g2_nand2_1 _16994_ (.Y(_10203_),
    .A(net920),
    .B(net148));
 sg13g2_o21ai_1 _16995_ (.B1(_10203_),
    .Y(_00064_),
    .A1(_10198_),
    .A2(_10199_));
 sg13g2_nand2b_1 _16996_ (.Y(_10204_),
    .B(_10190_),
    .A_N(_10104_));
 sg13g2_nor2_1 _16997_ (.A(_10107_),
    .B(_10204_),
    .Y(_10205_));
 sg13g2_xnor2_1 _16998_ (.Y(_10206_),
    .A(_10108_),
    .B(_10205_));
 sg13g2_o21ai_1 _16999_ (.B1(_10130_),
    .Y(_10207_),
    .A1(\cpu.intr.r_timer_reload[19] ),
    .A2(_10114_));
 sg13g2_buf_1 _17000_ (.A(\cpu.dcache.wdata[3] ),
    .X(_10208_));
 sg13g2_buf_1 _17001_ (.A(net1116),
    .X(_10209_));
 sg13g2_nand2_1 _17002_ (.Y(_10210_),
    .A(_10209_),
    .B(net148));
 sg13g2_o21ai_1 _17003_ (.B1(_10210_),
    .Y(_00065_),
    .A1(_10206_),
    .A2(_10207_));
 sg13g2_nor3_1 _17004_ (.A(_10107_),
    .B(_10108_),
    .C(_10204_),
    .Y(_10211_));
 sg13g2_xor2_1 _17005_ (.B(_10211_),
    .A(_10109_),
    .X(_10212_));
 sg13g2_o21ai_1 _17006_ (.B1(_10212_),
    .Y(_10213_),
    .A1(\cpu.intr.r_timer_reload[20] ),
    .A2(_10114_));
 sg13g2_buf_2 _17007_ (.A(\cpu.dcache.wdata[4] ),
    .X(_10214_));
 sg13g2_buf_1 _17008_ (.A(_10214_),
    .X(_10215_));
 sg13g2_nand2_1 _17009_ (.Y(_10216_),
    .A(net1037),
    .B(net148));
 sg13g2_o21ai_1 _17010_ (.B1(_10216_),
    .Y(_00067_),
    .A1(net133),
    .A2(_10213_));
 sg13g2_nor2b_1 _17011_ (.A(_10109_),
    .B_N(_10211_),
    .Y(_10217_));
 sg13g2_xnor2_1 _17012_ (.Y(_10218_),
    .A(\cpu.intr.r_timer_count[21] ),
    .B(_10217_));
 sg13g2_o21ai_1 _17013_ (.B1(_10130_),
    .Y(_10219_),
    .A1(\cpu.intr.r_timer_reload[21] ),
    .A2(_10114_));
 sg13g2_buf_2 _17014_ (.A(\cpu.dcache.wdata[5] ),
    .X(_10220_));
 sg13g2_buf_1 _17015_ (.A(_10220_),
    .X(_10221_));
 sg13g2_nand2_1 _17016_ (.Y(_10222_),
    .A(net1036),
    .B(net148));
 sg13g2_o21ai_1 _17017_ (.B1(_10222_),
    .Y(_00068_),
    .A1(_10218_),
    .A2(_10219_));
 sg13g2_nand2_1 _17018_ (.Y(_10223_),
    .A(_10110_),
    .B(_10191_));
 sg13g2_xor2_1 _17019_ (.B(_10223_),
    .A(\cpu.intr.r_timer_count[22] ),
    .X(_10224_));
 sg13g2_o21ai_1 _17020_ (.B1(_10130_),
    .Y(_10225_),
    .A1(\cpu.intr.r_timer_reload[22] ),
    .A2(_10114_));
 sg13g2_buf_2 _17021_ (.A(\cpu.dcache.wdata[6] ),
    .X(_10226_));
 sg13g2_buf_1 _17022_ (.A(_10226_),
    .X(_10227_));
 sg13g2_nand2_1 _17023_ (.Y(_10228_),
    .A(net1035),
    .B(net148));
 sg13g2_o21ai_1 _17024_ (.B1(_10228_),
    .Y(_00069_),
    .A1(_10224_),
    .A2(_10225_));
 sg13g2_buf_2 _17025_ (.A(\cpu.dcache.wdata[7] ),
    .X(_10229_));
 sg13g2_buf_1 _17026_ (.A(_10229_),
    .X(_10230_));
 sg13g2_nor2b_1 _17027_ (.A(_10106_),
    .B_N(\cpu.intr.r_timer_reload[23] ),
    .Y(_10231_));
 sg13g2_nor2_1 _17028_ (.A(_10111_),
    .B(_10204_),
    .Y(_10232_));
 sg13g2_mux2_1 _17029_ (.A0(_10106_),
    .A1(_10231_),
    .S(_10232_),
    .X(_10233_));
 sg13g2_mux2_1 _17030_ (.A0(net1034),
    .A1(_10233_),
    .S(_10130_),
    .X(_00070_));
 sg13g2_buf_1 _17031_ (.A(net626),
    .X(_10234_));
 sg13g2_buf_1 _17032_ (.A(net544),
    .X(_10235_));
 sg13g2_buf_1 _17033_ (.A(net493),
    .X(_10236_));
 sg13g2_nand2_1 _17034_ (.Y(_10237_),
    .A(net444),
    .B(_10128_));
 sg13g2_buf_1 _17035_ (.A(_10237_),
    .X(_10238_));
 sg13g2_buf_1 _17036_ (.A(net117),
    .X(_10239_));
 sg13g2_buf_1 _17037_ (.A(net620),
    .X(_10240_));
 sg13g2_buf_1 _17038_ (.A(net1041),
    .X(_10241_));
 sg13g2_nand2_1 _17039_ (.Y(_10242_),
    .A(net543),
    .B(net919));
 sg13g2_nand2_1 _17040_ (.Y(_10243_),
    .A(_00286_),
    .B(_10239_));
 sg13g2_o21ai_1 _17041_ (.B1(_10243_),
    .Y(_00036_),
    .A1(_10239_),
    .A2(_10242_));
 sg13g2_buf_1 _17042_ (.A(net1040),
    .X(_10244_));
 sg13g2_buf_1 _17043_ (.A(net684),
    .X(_10245_));
 sg13g2_buf_2 _17044_ (.A(net618),
    .X(_10246_));
 sg13g2_nor2_1 _17045_ (.A(net542),
    .B(net117),
    .Y(_10247_));
 sg13g2_buf_1 _17046_ (.A(_10247_),
    .X(_10248_));
 sg13g2_buf_1 _17047_ (.A(_10248_),
    .X(_10249_));
 sg13g2_buf_1 _17048_ (.A(_10248_),
    .X(_10250_));
 sg13g2_nand2_1 _17049_ (.Y(_10251_),
    .A(_09348_),
    .B(net1051));
 sg13g2_buf_1 _17050_ (.A(_10251_),
    .X(_10252_));
 sg13g2_nor3_1 _17051_ (.A(net929),
    .B(net633),
    .C(_10252_),
    .Y(_10253_));
 sg13g2_buf_1 _17052_ (.A(_10253_),
    .X(_10254_));
 sg13g2_buf_1 _17053_ (.A(_10254_),
    .X(_10255_));
 sg13g2_buf_1 _17054_ (.A(net443),
    .X(_10256_));
 sg13g2_and2_1 _17055_ (.A(_10128_),
    .B(net399),
    .X(_10257_));
 sg13g2_buf_1 _17056_ (.A(_10257_),
    .X(_10258_));
 sg13g2_buf_1 _17057_ (.A(_10258_),
    .X(_10259_));
 sg13g2_buf_1 _17058_ (.A(\cpu.intr.r_clock_count[0] ),
    .X(_10260_));
 sg13g2_buf_2 _17059_ (.A(\cpu.intr.r_clock_count[1] ),
    .X(_10261_));
 sg13g2_xnor2_1 _17060_ (.Y(_10262_),
    .A(_10260_),
    .B(_10261_));
 sg13g2_nor3_1 _17061_ (.A(net72),
    .B(net104),
    .C(_10262_),
    .Y(_10263_));
 sg13g2_a21o_1 _17062_ (.A2(net73),
    .A1(net918),
    .B1(_10263_),
    .X(_00043_));
 sg13g2_buf_1 _17063_ (.A(net1039),
    .X(_10264_));
 sg13g2_buf_1 _17064_ (.A(\cpu.intr.r_clock_count[2] ),
    .X(_10265_));
 sg13g2_nand2_1 _17065_ (.Y(_10266_),
    .A(_10260_),
    .B(_10261_));
 sg13g2_xor2_1 _17066_ (.B(_10266_),
    .A(_10265_),
    .X(_10267_));
 sg13g2_nor3_1 _17067_ (.A(net72),
    .B(_10259_),
    .C(_10267_),
    .Y(_10268_));
 sg13g2_a21o_1 _17068_ (.A2(net73),
    .A1(net917),
    .B1(_10268_),
    .X(_00044_));
 sg13g2_buf_1 _17069_ (.A(net1116),
    .X(_10269_));
 sg13g2_buf_2 _17070_ (.A(\cpu.intr.r_clock_count[3] ),
    .X(_10270_));
 sg13g2_nand2_1 _17071_ (.Y(_10271_),
    .A(_10261_),
    .B(_10265_));
 sg13g2_nor2_1 _17072_ (.A(_00286_),
    .B(_10271_),
    .Y(_10272_));
 sg13g2_xnor2_1 _17073_ (.Y(_10273_),
    .A(_10270_),
    .B(_10272_));
 sg13g2_nor3_1 _17074_ (.A(net72),
    .B(_10259_),
    .C(_10273_),
    .Y(_10274_));
 sg13g2_a21o_1 _17075_ (.A2(net73),
    .A1(net1033),
    .B1(_10274_),
    .X(_00045_));
 sg13g2_buf_1 _17076_ (.A(_10214_),
    .X(_10275_));
 sg13g2_buf_1 _17077_ (.A(_10258_),
    .X(_10276_));
 sg13g2_buf_2 _17078_ (.A(\cpu.intr.r_clock_count[4] ),
    .X(_10277_));
 sg13g2_and4_1 _17079_ (.A(_10260_),
    .B(_10261_),
    .C(_10265_),
    .D(_10270_),
    .X(_10278_));
 sg13g2_buf_1 _17080_ (.A(_10278_),
    .X(_10279_));
 sg13g2_xnor2_1 _17081_ (.Y(_10280_),
    .A(_10277_),
    .B(_10279_));
 sg13g2_nor3_1 _17082_ (.A(net72),
    .B(net103),
    .C(_10280_),
    .Y(_10281_));
 sg13g2_a21o_1 _17083_ (.A2(net73),
    .A1(net1032),
    .B1(_10281_),
    .X(_00046_));
 sg13g2_buf_1 _17084_ (.A(net1036),
    .X(_10282_));
 sg13g2_buf_2 _17085_ (.A(\cpu.intr.r_clock_count[5] ),
    .X(_10283_));
 sg13g2_and3_1 _17086_ (.X(_10284_),
    .A(_10270_),
    .B(_10277_),
    .C(_10272_));
 sg13g2_buf_1 _17087_ (.A(_10284_),
    .X(_10285_));
 sg13g2_xnor2_1 _17088_ (.Y(_10286_),
    .A(_10283_),
    .B(_10285_));
 sg13g2_nor3_1 _17089_ (.A(_10250_),
    .B(net103),
    .C(_10286_),
    .Y(_10287_));
 sg13g2_a21o_1 _17090_ (.A2(_10249_),
    .A1(net916),
    .B1(_10287_),
    .X(_00047_));
 sg13g2_buf_1 _17091_ (.A(_10226_),
    .X(_10288_));
 sg13g2_buf_2 _17092_ (.A(\cpu.intr.r_clock_count[6] ),
    .X(_10289_));
 sg13g2_nand3_1 _17093_ (.B(_10283_),
    .C(_10279_),
    .A(_10277_),
    .Y(_10290_));
 sg13g2_xor2_1 _17094_ (.B(_10290_),
    .A(_10289_),
    .X(_10291_));
 sg13g2_nor3_1 _17095_ (.A(_10250_),
    .B(_10276_),
    .C(_10291_),
    .Y(_10292_));
 sg13g2_a21o_1 _17096_ (.A2(_10249_),
    .A1(net1031),
    .B1(_10292_),
    .X(_00048_));
 sg13g2_buf_1 _17097_ (.A(\cpu.intr.r_clock_count[7] ),
    .X(_10293_));
 sg13g2_nand3_1 _17098_ (.B(_10289_),
    .C(_10285_),
    .A(_10283_),
    .Y(_10294_));
 sg13g2_xor2_1 _17099_ (.B(_10294_),
    .A(_10293_),
    .X(_10295_));
 sg13g2_nor3_1 _17100_ (.A(_10248_),
    .B(net103),
    .C(_10295_),
    .Y(_10296_));
 sg13g2_a21o_1 _17101_ (.A2(net73),
    .A1(net1034),
    .B1(_10296_),
    .X(_00049_));
 sg13g2_buf_2 _17102_ (.A(\cpu.intr.r_clock_count[8] ),
    .X(_10297_));
 sg13g2_nand2_1 _17103_ (.Y(_10298_),
    .A(_10277_),
    .B(_10279_));
 sg13g2_nand3_1 _17104_ (.B(_10289_),
    .C(_10293_),
    .A(_10283_),
    .Y(_10299_));
 sg13g2_nor2_1 _17105_ (.A(_10298_),
    .B(_10299_),
    .Y(_10300_));
 sg13g2_xnor2_1 _17106_ (.Y(_10301_),
    .A(_10297_),
    .B(_10300_));
 sg13g2_buf_2 _17107_ (.A(\cpu.dcache.wdata[8] ),
    .X(_10302_));
 sg13g2_a21oi_1 _17108_ (.A1(net543),
    .A2(_10302_),
    .Y(_10303_),
    .B1(net105));
 sg13g2_a21oi_1 _17109_ (.A1(net105),
    .A2(_10301_),
    .Y(_00050_),
    .B1(_10303_));
 sg13g2_buf_2 _17110_ (.A(\cpu.intr.r_clock_count[9] ),
    .X(_10304_));
 sg13g2_nand2_1 _17111_ (.Y(_10305_),
    .A(_10297_),
    .B(_10300_));
 sg13g2_xor2_1 _17112_ (.B(_10305_),
    .A(_10304_),
    .X(_10306_));
 sg13g2_buf_2 _17113_ (.A(\cpu.dcache.wdata[9] ),
    .X(_10307_));
 sg13g2_a21oi_1 _17114_ (.A1(net543),
    .A2(_10307_),
    .Y(_10308_),
    .B1(net117));
 sg13g2_a21oi_1 _17115_ (.A1(net105),
    .A2(_10306_),
    .Y(_00051_),
    .B1(_10308_));
 sg13g2_buf_1 _17116_ (.A(\cpu.intr.r_clock_count[10] ),
    .X(_10309_));
 sg13g2_nand3_1 _17117_ (.B(_10304_),
    .C(_10300_),
    .A(_10297_),
    .Y(_10310_));
 sg13g2_xor2_1 _17118_ (.B(_10310_),
    .A(_10309_),
    .X(_10311_));
 sg13g2_buf_2 _17119_ (.A(\cpu.dcache.wdata[10] ),
    .X(_10312_));
 sg13g2_a21oi_1 _17120_ (.A1(net543),
    .A2(_10312_),
    .Y(_10313_),
    .B1(net117));
 sg13g2_a21oi_1 _17121_ (.A1(net105),
    .A2(_10311_),
    .Y(_00037_),
    .B1(_10313_));
 sg13g2_buf_1 _17122_ (.A(\cpu.intr.r_clock_count[11] ),
    .X(_10314_));
 sg13g2_nand3_1 _17123_ (.B(_10304_),
    .C(_10309_),
    .A(_10297_),
    .Y(_10315_));
 sg13g2_nor2_1 _17124_ (.A(_10299_),
    .B(_10315_),
    .Y(_10316_));
 sg13g2_nand2_1 _17125_ (.Y(_10317_),
    .A(_10285_),
    .B(_10316_));
 sg13g2_xor2_1 _17126_ (.B(_10317_),
    .A(_10314_),
    .X(_10318_));
 sg13g2_buf_2 _17127_ (.A(\cpu.dcache.wdata[11] ),
    .X(_10319_));
 sg13g2_a21oi_1 _17128_ (.A1(net543),
    .A2(_10319_),
    .Y(_10320_),
    .B1(net117));
 sg13g2_a21oi_1 _17129_ (.A1(net105),
    .A2(_10318_),
    .Y(_00038_),
    .B1(_10320_));
 sg13g2_buf_1 _17130_ (.A(\cpu.intr.r_clock_count[12] ),
    .X(_10321_));
 sg13g2_nand4_1 _17131_ (.B(_10314_),
    .C(_10279_),
    .A(_10277_),
    .Y(_10322_),
    .D(_10316_));
 sg13g2_xor2_1 _17132_ (.B(_10322_),
    .A(_10321_),
    .X(_10323_));
 sg13g2_buf_2 _17133_ (.A(\cpu.dcache.wdata[12] ),
    .X(_10324_));
 sg13g2_a21oi_1 _17134_ (.A1(net543),
    .A2(_10324_),
    .Y(_10325_),
    .B1(net117));
 sg13g2_a21oi_1 _17135_ (.A1(net105),
    .A2(_10323_),
    .Y(_00039_),
    .B1(_10325_));
 sg13g2_buf_2 _17136_ (.A(\cpu.dcache.wdata[13] ),
    .X(_10326_));
 sg13g2_buf_2 _17137_ (.A(\cpu.intr.r_clock_count[13] ),
    .X(_10327_));
 sg13g2_nand3_1 _17138_ (.B(_10277_),
    .C(_10272_),
    .A(_10270_),
    .Y(_10328_));
 sg13g2_nand3_1 _17139_ (.B(_10321_),
    .C(_10316_),
    .A(_10314_),
    .Y(_10329_));
 sg13g2_nor2_1 _17140_ (.A(_10328_),
    .B(_10329_),
    .Y(_10330_));
 sg13g2_xnor2_1 _17141_ (.Y(_10331_),
    .A(_10327_),
    .B(_10330_));
 sg13g2_nor3_1 _17142_ (.A(_10248_),
    .B(net103),
    .C(_10331_),
    .Y(_10332_));
 sg13g2_a21o_1 _17143_ (.A2(net72),
    .A1(_10326_),
    .B1(_10332_),
    .X(_00040_));
 sg13g2_buf_2 _17144_ (.A(\cpu.intr.r_clock_count[14] ),
    .X(_10333_));
 sg13g2_inv_1 _17145_ (.Y(_10334_),
    .A(_10327_));
 sg13g2_or2_1 _17146_ (.X(_10335_),
    .B(_10329_),
    .A(_10298_));
 sg13g2_buf_1 _17147_ (.A(_10335_),
    .X(_10336_));
 sg13g2_nor2_1 _17148_ (.A(_10334_),
    .B(_10336_),
    .Y(_10337_));
 sg13g2_xnor2_1 _17149_ (.Y(_10338_),
    .A(_10333_),
    .B(_10337_));
 sg13g2_buf_2 _17150_ (.A(\cpu.dcache.wdata[14] ),
    .X(_10339_));
 sg13g2_a21oi_1 _17151_ (.A1(net543),
    .A2(_10339_),
    .Y(_10340_),
    .B1(net117));
 sg13g2_a21oi_1 _17152_ (.A1(net105),
    .A2(_10338_),
    .Y(_00041_),
    .B1(_10340_));
 sg13g2_buf_2 _17153_ (.A(\cpu.intr.r_clock_count[15] ),
    .X(_10341_));
 sg13g2_nand3_1 _17154_ (.B(_10333_),
    .C(_10330_),
    .A(_10327_),
    .Y(_10342_));
 sg13g2_xor2_1 _17155_ (.B(_10342_),
    .A(_10341_),
    .X(_10343_));
 sg13g2_buf_2 _17156_ (.A(\cpu.dcache.wdata[15] ),
    .X(_10344_));
 sg13g2_a21oi_1 _17157_ (.A1(net543),
    .A2(_10344_),
    .Y(_10345_),
    .B1(net117));
 sg13g2_a21oi_1 _17158_ (.A1(net105),
    .A2(_10343_),
    .Y(_00042_),
    .B1(_10345_));
 sg13g2_buf_1 _17159_ (.A(\cpu.ex.r_mult[0] ),
    .X(_10346_));
 sg13g2_buf_1 _17160_ (.A(\cpu.ex.r_wb_valid ),
    .X(_10347_));
 sg13g2_inv_1 _17161_ (.Y(_10348_),
    .A(net1115));
 sg13g2_buf_8 _17162_ (.A(\cpu.ex.r_wb_addr[1] ),
    .X(_10349_));
 sg13g2_buf_8 _17163_ (.A(\cpu.ex.r_wb_addr[0] ),
    .X(_10350_));
 sg13g2_nand2_1 _17164_ (.Y(_10351_),
    .A(net1114),
    .B(net1113));
 sg13g2_buf_2 _17165_ (.A(\cpu.ex.r_wb_addr[3] ),
    .X(_10352_));
 sg13g2_buf_1 _17166_ (.A(\cpu.ex.r_wb_addr[2] ),
    .X(_10353_));
 sg13g2_inv_1 _17167_ (.Y(_10354_),
    .A(net1111));
 sg13g2_nor2_1 _17168_ (.A(net1112),
    .B(_10354_),
    .Y(_10355_));
 sg13g2_inv_1 _17169_ (.Y(_10356_),
    .A(_10355_));
 sg13g2_nor3_1 _17170_ (.A(_10348_),
    .B(_10351_),
    .C(_10356_),
    .Y(_10357_));
 sg13g2_buf_1 _17171_ (.A(_10357_),
    .X(_10358_));
 sg13g2_buf_1 _17172_ (.A(\cpu.ex.r_set_cc ),
    .X(_10359_));
 sg13g2_nand2_2 _17173_ (.Y(_10360_),
    .A(net1115),
    .B(_10359_));
 sg13g2_nor2b_1 _17174_ (.A(_10358_),
    .B_N(_10360_),
    .Y(_10361_));
 sg13g2_buf_1 _17175_ (.A(_10361_),
    .X(_10362_));
 sg13g2_nor2_2 _17176_ (.A(_09466_),
    .B(net1122),
    .Y(_10363_));
 sg13g2_nand2_2 _17177_ (.Y(_10364_),
    .A(net495),
    .B(_10363_));
 sg13g2_nand2_1 _17178_ (.Y(_10365_),
    .A(_10362_),
    .B(_10364_));
 sg13g2_buf_1 _17179_ (.A(_10365_),
    .X(_10366_));
 sg13g2_buf_1 _17180_ (.A(_10366_),
    .X(_10367_));
 sg13g2_nand2_1 _17181_ (.Y(_10368_),
    .A(_10346_),
    .B(net278));
 sg13g2_buf_2 _17182_ (.A(\cpu.dec.r_rs2_pc ),
    .X(_10369_));
 sg13g2_buf_1 _17183_ (.A(_10369_),
    .X(_10370_));
 sg13g2_buf_1 _17184_ (.A(\cpu.dec.r_rs2_inv ),
    .X(_10371_));
 sg13g2_buf_1 _17185_ (.A(\cpu.dec.needs_rs2 ),
    .X(_10372_));
 sg13g2_buf_1 _17186_ (.A(_10372_),
    .X(_10373_));
 sg13g2_buf_1 _17187_ (.A(net1029),
    .X(_10374_));
 sg13g2_or4_1 _17188_ (.A(net1114),
    .B(net1113),
    .C(\cpu.ex.r_wb_addr[3] ),
    .D(net1111),
    .X(_10375_));
 sg13g2_buf_1 _17189_ (.A(_10375_),
    .X(_10376_));
 sg13g2_buf_8 _17190_ (.A(\cpu.dec.r_rs2[2] ),
    .X(_10377_));
 sg13g2_xnor2_1 _17191_ (.Y(_10378_),
    .A(net1111),
    .B(_10377_));
 sg13g2_buf_8 _17192_ (.A(\cpu.dec.r_rs2[1] ),
    .X(_10379_));
 sg13g2_xnor2_1 _17193_ (.Y(_10380_),
    .A(net1114),
    .B(net1110));
 sg13g2_nand4_1 _17194_ (.B(_10376_),
    .C(_10378_),
    .A(net1115),
    .Y(_10381_),
    .D(_10380_));
 sg13g2_buf_8 _17195_ (.A(\cpu.dec.r_rs2[3] ),
    .X(_10382_));
 sg13g2_xor2_1 _17196_ (.B(_10382_),
    .A(net1112),
    .X(_10383_));
 sg13g2_buf_8 _17197_ (.A(\cpu.dec.r_rs2[0] ),
    .X(_10384_));
 sg13g2_xor2_1 _17198_ (.B(_10384_),
    .A(net1113),
    .X(_10385_));
 sg13g2_or2_1 _17199_ (.X(_10386_),
    .B(_10385_),
    .A(_10383_));
 sg13g2_nor2_1 _17200_ (.A(_10381_),
    .B(_10386_),
    .Y(_10387_));
 sg13g2_buf_2 _17201_ (.A(_10387_),
    .X(_10388_));
 sg13g2_buf_8 _17202_ (.A(_10388_),
    .X(_10389_));
 sg13g2_and4_1 _17203_ (.A(net1115),
    .B(_10376_),
    .C(_10378_),
    .D(_10380_),
    .X(_10390_));
 sg13g2_buf_8 _17204_ (.A(_10390_),
    .X(_10391_));
 sg13g2_nor2_1 _17205_ (.A(_10383_),
    .B(_10385_),
    .Y(_10392_));
 sg13g2_nor2_1 _17206_ (.A(_10384_),
    .B(net1110),
    .Y(_10393_));
 sg13g2_buf_2 _17207_ (.A(_10393_),
    .X(_10394_));
 sg13g2_buf_8 _17208_ (.A(_10382_),
    .X(_10395_));
 sg13g2_nor2_1 _17209_ (.A(net1028),
    .B(_10377_),
    .Y(_10396_));
 sg13g2_buf_2 _17210_ (.A(_10396_),
    .X(_10397_));
 sg13g2_a22oi_1 _17211_ (.Y(_10398_),
    .B1(_10394_),
    .B2(_10397_),
    .A2(_10392_),
    .A1(_10391_));
 sg13g2_buf_8 _17212_ (.A(_10398_),
    .X(_10399_));
 sg13g2_buf_8 _17213_ (.A(_10384_),
    .X(_10400_));
 sg13g2_buf_8 _17214_ (.A(_10377_),
    .X(_10401_));
 sg13g2_nor2b_2 _17215_ (.A(net1027),
    .B_N(net1026),
    .Y(_10402_));
 sg13g2_inv_1 _17216_ (.Y(_10403_),
    .A(\cpu.ex.r_12[15] ));
 sg13g2_nand2b_1 _17217_ (.Y(_10404_),
    .B(net1028),
    .A_N(net1110));
 sg13g2_buf_2 _17218_ (.A(_10404_),
    .X(_10405_));
 sg13g2_buf_8 _17219_ (.A(net1028),
    .X(_10406_));
 sg13g2_buf_1 _17220_ (.A(net914),
    .X(_10407_));
 sg13g2_buf_1 _17221_ (.A(net784),
    .X(_10408_));
 sg13g2_buf_8 _17222_ (.A(net1110),
    .X(_10409_));
 sg13g2_buf_8 _17223_ (.A(_10409_),
    .X(_10410_));
 sg13g2_buf_8 _17224_ (.A(net913),
    .X(_10411_));
 sg13g2_buf_8 _17225_ (.A(net783),
    .X(_10412_));
 sg13g2_nand3b_1 _17226_ (.B(net679),
    .C(\cpu.ex.r_stmp[15] ),
    .Y(_10413_),
    .A_N(net680));
 sg13g2_o21ai_1 _17227_ (.B1(_10413_),
    .Y(_10414_),
    .A1(_10403_),
    .A2(_10405_));
 sg13g2_buf_1 _17228_ (.A(\cpu.ex.mmu_read[15] ),
    .X(_10415_));
 sg13g2_buf_8 _17229_ (.A(_10401_),
    .X(_10416_));
 sg13g2_buf_8 _17230_ (.A(net912),
    .X(_10417_));
 sg13g2_buf_8 _17231_ (.A(net782),
    .X(_10418_));
 sg13g2_buf_8 _17232_ (.A(net678),
    .X(_10419_));
 sg13g2_buf_1 _17233_ (.A(net617),
    .X(_10420_));
 sg13g2_mux2_1 _17234_ (.A0(\cpu.ex.r_lr[15] ),
    .A1(_10415_),
    .S(net539),
    .X(_10421_));
 sg13g2_buf_8 _17235_ (.A(net1027),
    .X(_10422_));
 sg13g2_nor2_1 _17236_ (.A(net1110),
    .B(_10382_),
    .Y(_10423_));
 sg13g2_buf_1 _17237_ (.A(_10423_),
    .X(_10424_));
 sg13g2_and2_1 _17238_ (.A(net911),
    .B(net910),
    .X(_10425_));
 sg13g2_buf_8 _17239_ (.A(net1027),
    .X(_10426_));
 sg13g2_nor2b_1 _17240_ (.A(net913),
    .B_N(net909),
    .Y(_10427_));
 sg13g2_buf_2 _17241_ (.A(_10427_),
    .X(_10428_));
 sg13g2_and2_1 _17242_ (.A(_10395_),
    .B(net1026),
    .X(_10429_));
 sg13g2_buf_1 _17243_ (.A(_10429_),
    .X(_10430_));
 sg13g2_and3_1 _17244_ (.X(_10431_),
    .A(\cpu.ex.r_13[15] ),
    .B(_10428_),
    .C(net781));
 sg13g2_a221oi_1 _17245_ (.B2(_10425_),
    .C1(_10431_),
    .B1(_10421_),
    .A1(_10402_),
    .Y(_10432_),
    .A2(_10414_));
 sg13g2_nand2b_1 _17246_ (.Y(_10433_),
    .B(net1025),
    .A_N(net1027));
 sg13g2_buf_1 _17247_ (.A(_10433_),
    .X(_10434_));
 sg13g2_nand2_1 _17248_ (.Y(_10435_),
    .A(net914),
    .B(_10418_));
 sg13g2_nor2_1 _17249_ (.A(_10434_),
    .B(_10435_),
    .Y(_10436_));
 sg13g2_nand2_1 _17250_ (.Y(_10437_),
    .A(\cpu.ex.r_14[15] ),
    .B(_10436_));
 sg13g2_buf_8 _17251_ (.A(net1028),
    .X(_10438_));
 sg13g2_nand2b_1 _17252_ (.Y(_10439_),
    .B(net908),
    .A_N(net1026));
 sg13g2_buf_2 _17253_ (.A(_10439_),
    .X(_10440_));
 sg13g2_nor2_1 _17254_ (.A(_10434_),
    .B(_10440_),
    .Y(_10441_));
 sg13g2_buf_8 _17255_ (.A(net909),
    .X(_10442_));
 sg13g2_buf_8 _17256_ (.A(net780),
    .X(_10443_));
 sg13g2_buf_8 _17257_ (.A(net677),
    .X(_10444_));
 sg13g2_buf_8 _17258_ (.A(net616),
    .X(_10445_));
 sg13g2_mux2_1 _17259_ (.A0(\cpu.ex.r_8[15] ),
    .A1(\cpu.ex.r_9[15] ),
    .S(net538),
    .X(_10446_));
 sg13g2_nor2_2 _17260_ (.A(net678),
    .B(_10405_),
    .Y(_10447_));
 sg13g2_a22oi_1 _17261_ (.Y(_10448_),
    .B1(_10446_),
    .B2(_10447_),
    .A2(_10441_),
    .A1(\cpu.ex.r_10[15] ));
 sg13g2_buf_1 _17262_ (.A(\cpu.ex.r_sp[15] ),
    .X(_10449_));
 sg13g2_nor3_1 _17263_ (.A(net677),
    .B(net784),
    .C(net678),
    .Y(_10450_));
 sg13g2_mux4_1 _17264_ (.S0(net539),
    .A0(\cpu.ex.r_epc[15] ),
    .A1(\cpu.ex.r_mult[31] ),
    .A2(\cpu.ex.r_11[15] ),
    .A3(\cpu.ex.r_15[15] ),
    .S1(net680),
    .X(_10451_));
 sg13g2_a22oi_1 _17265_ (.Y(_10452_),
    .B1(_10451_),
    .B2(net538),
    .A2(_10450_),
    .A1(_10449_));
 sg13g2_nand2b_1 _17266_ (.Y(_10453_),
    .B(net679),
    .A_N(_10452_));
 sg13g2_nand4_1 _17267_ (.B(_10437_),
    .C(_10448_),
    .A(_10432_),
    .Y(_10454_),
    .D(_10453_));
 sg13g2_a22oi_1 _17268_ (.Y(_10455_),
    .B1(net540),
    .B2(_10454_),
    .A2(net541),
    .A1(net926));
 sg13g2_nor2_1 _17269_ (.A(net915),
    .B(\cpu.dec.imm[15] ),
    .Y(_10456_));
 sg13g2_a21oi_1 _17270_ (.A1(net915),
    .A2(_10455_),
    .Y(_10457_),
    .B1(_10456_));
 sg13g2_nor2_1 _17271_ (.A(_10371_),
    .B(_10457_),
    .Y(_10458_));
 sg13g2_nand2_1 _17272_ (.Y(_10459_),
    .A(net941),
    .B(net1030));
 sg13g2_o21ai_1 _17273_ (.B1(_10459_),
    .Y(_10460_),
    .A1(net1030),
    .A2(_10458_));
 sg13g2_buf_2 _17274_ (.A(_10460_),
    .X(_10461_));
 sg13g2_buf_1 _17275_ (.A(_00299_),
    .X(_10462_));
 sg13g2_buf_1 _17276_ (.A(net550),
    .X(_10463_));
 sg13g2_nor2_1 _17277_ (.A(_10462_),
    .B(net491),
    .Y(_10464_));
 sg13g2_buf_1 _17278_ (.A(_10464_),
    .X(_10465_));
 sg13g2_nor2b_1 _17279_ (.A(_10461_),
    .B_N(_10465_),
    .Y(_10466_));
 sg13g2_buf_1 _17280_ (.A(_10466_),
    .X(_10467_));
 sg13g2_nand2_1 _17281_ (.Y(_10468_),
    .A(\cpu.dec.div ),
    .B(_09459_));
 sg13g2_buf_1 _17282_ (.A(_10468_),
    .X(_10469_));
 sg13g2_buf_1 _17283_ (.A(net615),
    .X(_10470_));
 sg13g2_buf_1 _17284_ (.A(_00300_),
    .X(_10471_));
 sg13g2_inv_2 _17285_ (.Y(_10472_),
    .A(_10471_));
 sg13g2_nor2_1 _17286_ (.A(_10369_),
    .B(_10371_),
    .Y(_10473_));
 sg13g2_buf_1 _17287_ (.A(_10473_),
    .X(_10474_));
 sg13g2_buf_1 _17288_ (.A(_10474_),
    .X(_10475_));
 sg13g2_inv_1 _17289_ (.Y(_10476_),
    .A(_10400_));
 sg13g2_buf_1 _17290_ (.A(_10476_),
    .X(_10477_));
 sg13g2_buf_8 _17291_ (.A(net778),
    .X(_10478_));
 sg13g2_buf_1 _17292_ (.A(net676),
    .X(_10479_));
 sg13g2_buf_1 _17293_ (.A(\cpu.ex.r_mult[28] ),
    .X(_10480_));
 sg13g2_and2_1 _17294_ (.A(net913),
    .B(net782),
    .X(_10481_));
 sg13g2_buf_1 _17295_ (.A(_10481_),
    .X(_10482_));
 sg13g2_buf_2 _17296_ (.A(\cpu.ex.mmu_read[12] ),
    .X(_10483_));
 sg13g2_mux2_1 _17297_ (.A0(\cpu.ex.r_lr[12] ),
    .A1(_10483_),
    .S(net678),
    .X(_10484_));
 sg13g2_inv_2 _17298_ (.Y(_10485_),
    .A(net913));
 sg13g2_buf_1 _17299_ (.A(_10485_),
    .X(_10486_));
 sg13g2_a22oi_1 _17300_ (.Y(_10487_),
    .B1(_10484_),
    .B2(net675),
    .A2(net613),
    .A1(_10480_));
 sg13g2_nand3_1 _17301_ (.B(net676),
    .C(net613),
    .A(\cpu.ex.r_stmp[12] ),
    .Y(_10488_));
 sg13g2_o21ai_1 _17302_ (.B1(_10488_),
    .Y(_10489_),
    .A1(net614),
    .A2(_10487_));
 sg13g2_nand3_1 _17303_ (.B(net675),
    .C(_10402_),
    .A(\cpu.ex.r_12[12] ),
    .Y(_10490_));
 sg13g2_inv_2 _17304_ (.Y(_10491_),
    .A(net1026));
 sg13g2_buf_1 _17305_ (.A(_10491_),
    .X(_10492_));
 sg13g2_and2_1 _17306_ (.A(net909),
    .B(net913),
    .X(_10493_));
 sg13g2_buf_2 _17307_ (.A(_10493_),
    .X(_10494_));
 sg13g2_nand3_1 _17308_ (.B(net777),
    .C(_10494_),
    .A(\cpu.ex.r_11[12] ),
    .Y(_10495_));
 sg13g2_nand3_1 _17309_ (.B(_10490_),
    .C(_10495_),
    .A(net680),
    .Y(_10496_));
 sg13g2_o21ai_1 _17310_ (.B1(_10496_),
    .Y(_10497_),
    .A1(net680),
    .A2(_10489_));
 sg13g2_nand3_1 _17311_ (.B(net1028),
    .C(_10377_),
    .A(_10384_),
    .Y(_10498_));
 sg13g2_buf_1 _17312_ (.A(_10498_),
    .X(_10499_));
 sg13g2_buf_1 _17313_ (.A(\cpu.ex.r_sp[12] ),
    .X(_10500_));
 sg13g2_nand2_1 _17314_ (.Y(_10501_),
    .A(_10500_),
    .B(_10450_));
 sg13g2_o21ai_1 _17315_ (.B1(_10501_),
    .Y(_10502_),
    .A1(_00270_),
    .A2(_10499_));
 sg13g2_nor2b_1 _17316_ (.A(_10382_),
    .B_N(_10379_),
    .Y(_10503_));
 sg13g2_buf_1 _17317_ (.A(_10503_),
    .X(_10504_));
 sg13g2_and2_1 _17318_ (.A(net1027),
    .B(_10504_),
    .X(_10505_));
 sg13g2_buf_1 _17319_ (.A(_10505_),
    .X(_10506_));
 sg13g2_nor2b_1 _17320_ (.A(net1110),
    .B_N(net1028),
    .Y(_10507_));
 sg13g2_buf_1 _17321_ (.A(_10507_),
    .X(_10508_));
 sg13g2_buf_8 _17322_ (.A(net776),
    .X(_10509_));
 sg13g2_and3_1 _17323_ (.X(_10510_),
    .A(\cpu.ex.r_8[12] ),
    .B(net676),
    .C(net674));
 sg13g2_a21o_1 _17324_ (.A2(_10506_),
    .A1(\cpu.ex.r_epc[12] ),
    .B1(_10510_),
    .X(_10511_));
 sg13g2_nor2b_1 _17325_ (.A(_10384_),
    .B_N(net1110),
    .Y(_10512_));
 sg13g2_buf_2 _17326_ (.A(_10512_),
    .X(_10513_));
 sg13g2_a22oi_1 _17327_ (.Y(_10514_),
    .B1(_10513_),
    .B2(\cpu.ex.r_10[12] ),
    .A2(_10428_),
    .A1(\cpu.ex.r_9[12] ));
 sg13g2_nand3b_1 _17328_ (.B(net783),
    .C(\cpu.ex.r_14[12] ),
    .Y(_10515_),
    .A_N(net677));
 sg13g2_nand3b_1 _17329_ (.B(net677),
    .C(\cpu.ex.r_13[12] ),
    .Y(_10516_),
    .A_N(net783));
 sg13g2_a21o_1 _17330_ (.A2(_10516_),
    .A1(_10515_),
    .B1(_10435_),
    .X(_10517_));
 sg13g2_o21ai_1 _17331_ (.B1(_10517_),
    .Y(_10518_),
    .A1(_10440_),
    .A2(_10514_));
 sg13g2_a221oi_1 _17332_ (.B2(net777),
    .C1(_10518_),
    .B1(_10511_),
    .A1(net679),
    .Y(_10519_),
    .A2(_10502_));
 sg13g2_nand2_1 _17333_ (.Y(_10520_),
    .A(_10394_),
    .B(_10397_));
 sg13g2_o21ai_1 _17334_ (.B1(_10520_),
    .Y(_10521_),
    .A1(_10381_),
    .A2(_10386_));
 sg13g2_buf_1 _17335_ (.A(_10521_),
    .X(_10522_));
 sg13g2_a21o_1 _17336_ (.A2(_10519_),
    .A1(_10497_),
    .B1(net536),
    .X(_10523_));
 sg13g2_nand2_1 _17337_ (.Y(_10524_),
    .A(net687),
    .B(net541));
 sg13g2_nand3_1 _17338_ (.B(_10523_),
    .C(_10524_),
    .A(net915),
    .Y(_10525_));
 sg13g2_o21ai_1 _17339_ (.B1(_10525_),
    .Y(_10526_),
    .A1(net915),
    .A2(\cpu.dec.imm[12] ));
 sg13g2_inv_1 _17340_ (.Y(_10527_),
    .A(_10369_));
 sg13g2_buf_1 _17341_ (.A(_10527_),
    .X(_10528_));
 sg13g2_nor2_1 _17342_ (.A(_08534_),
    .B(net906),
    .Y(_10529_));
 sg13g2_a21o_1 _17343_ (.A2(_10526_),
    .A1(_10475_),
    .B1(_10529_),
    .X(_10530_));
 sg13g2_buf_1 _17344_ (.A(_10530_),
    .X(_10531_));
 sg13g2_buf_1 _17345_ (.A(_10531_),
    .X(_10532_));
 sg13g2_xnor2_1 _17346_ (.Y(_10533_),
    .A(_10472_),
    .B(net176));
 sg13g2_or2_1 _17347_ (.X(_10534_),
    .B(_10371_),
    .A(_10369_));
 sg13g2_buf_2 _17348_ (.A(_10534_),
    .X(_10535_));
 sg13g2_nand2b_1 _17349_ (.Y(_10536_),
    .B(net613),
    .A_N(_00271_));
 sg13g2_nor2_1 _17350_ (.A(net1025),
    .B(net1026),
    .Y(_10537_));
 sg13g2_buf_2 _17351_ (.A(_10537_),
    .X(_10538_));
 sg13g2_nand2_1 _17352_ (.Y(_10539_),
    .A(\cpu.ex.r_8[13] ),
    .B(_10538_));
 sg13g2_buf_1 _17353_ (.A(\cpu.ex.r_mult[29] ),
    .X(_10540_));
 sg13g2_buf_1 _17354_ (.A(\cpu.ex.mmu_read[13] ),
    .X(_10541_));
 sg13g2_buf_1 _17355_ (.A(_10541_),
    .X(_10542_));
 sg13g2_mux2_1 _17356_ (.A0(\cpu.ex.r_lr[13] ),
    .A1(_10542_),
    .S(net617),
    .X(_10543_));
 sg13g2_a22oi_1 _17357_ (.Y(_10544_),
    .B1(_10543_),
    .B2(net675),
    .A2(net613),
    .A1(_10540_));
 sg13g2_buf_1 _17358_ (.A(\cpu.ex.r_sp[13] ),
    .X(_10545_));
 sg13g2_nor2b_1 _17359_ (.A(net617),
    .B_N(net679),
    .Y(_10546_));
 sg13g2_nand2_1 _17360_ (.Y(_10547_),
    .A(_10545_),
    .B(_10546_));
 sg13g2_inv_2 _17361_ (.Y(_10548_),
    .A(net784));
 sg13g2_mux4_1 _17362_ (.S0(net614),
    .A0(_10536_),
    .A1(_10539_),
    .A2(_10544_),
    .A3(_10547_),
    .S1(_10548_),
    .X(_10549_));
 sg13g2_mux2_1 _17363_ (.A0(\cpu.ex.r_9[13] ),
    .A1(\cpu.ex.r_13[13] ),
    .S(net617),
    .X(_10550_));
 sg13g2_a22oi_1 _17364_ (.Y(_10551_),
    .B1(_10550_),
    .B2(net675),
    .A2(_10546_),
    .A1(\cpu.ex.r_11[13] ));
 sg13g2_nand3b_1 _17365_ (.B(_10408_),
    .C(net538),
    .Y(_10552_),
    .A_N(_10551_));
 sg13g2_nand3b_1 _17366_ (.B(net617),
    .C(\cpu.ex.r_stmp[13] ),
    .Y(_10553_),
    .A_N(_10408_));
 sg13g2_nand3b_1 _17367_ (.B(net680),
    .C(\cpu.ex.r_10[13] ),
    .Y(_10554_),
    .A_N(net617));
 sg13g2_a21oi_1 _17368_ (.A1(_10553_),
    .A2(_10554_),
    .Y(_10555_),
    .B1(net675));
 sg13g2_and3_1 _17369_ (.X(_10556_),
    .A(\cpu.ex.r_12[13] ),
    .B(net539),
    .C(net674));
 sg13g2_o21ai_1 _17370_ (.B1(net614),
    .Y(_10557_),
    .A1(_10555_),
    .A2(_10556_));
 sg13g2_nand3_1 _17371_ (.B(net538),
    .C(_10397_),
    .A(\cpu.ex.r_epc[13] ),
    .Y(_10558_));
 sg13g2_nand3_1 _17372_ (.B(net614),
    .C(net781),
    .A(\cpu.ex.r_14[13] ),
    .Y(_10559_));
 sg13g2_a21o_1 _17373_ (.A2(_10559_),
    .A1(_10558_),
    .B1(_10486_),
    .X(_10560_));
 sg13g2_nand4_1 _17374_ (.B(_10552_),
    .C(_10557_),
    .A(_10549_),
    .Y(_10561_),
    .D(_10560_));
 sg13g2_a22oi_1 _17375_ (.Y(_10562_),
    .B1(net540),
    .B2(_10561_),
    .A2(net541),
    .A1(net791));
 sg13g2_nor2_1 _17376_ (.A(net915),
    .B(\cpu.dec.imm[13] ),
    .Y(_10563_));
 sg13g2_a21oi_1 _17377_ (.A1(_10374_),
    .A2(_10562_),
    .Y(_10564_),
    .B1(_10563_));
 sg13g2_nor2_1 _17378_ (.A(_10535_),
    .B(_10564_),
    .Y(_10565_));
 sg13g2_a21oi_1 _17379_ (.A1(_08631_),
    .A2(net1030),
    .Y(_10566_),
    .B1(_10565_));
 sg13g2_buf_8 _17380_ (.A(_10566_),
    .X(_10567_));
 sg13g2_nand2_1 _17381_ (.Y(_10568_),
    .A(_10480_),
    .B(net175));
 sg13g2_buf_1 _17382_ (.A(_10471_),
    .X(_10569_));
 sg13g2_or4_1 _17383_ (.A(_10480_),
    .B(net1023),
    .C(_10531_),
    .D(_10566_),
    .X(_10570_));
 sg13g2_o21ai_1 _17384_ (.B1(_10570_),
    .Y(_10571_),
    .A1(_10533_),
    .A2(_10568_));
 sg13g2_buf_1 _17385_ (.A(_10480_),
    .X(_10572_));
 sg13g2_o21ai_1 _17386_ (.B1(net615),
    .Y(_10573_),
    .A1(net1022),
    .A2(_10472_));
 sg13g2_a21oi_1 _17387_ (.A1(_10475_),
    .A2(_10526_),
    .Y(_10574_),
    .B1(_10529_));
 sg13g2_buf_1 _17388_ (.A(_10574_),
    .X(_10575_));
 sg13g2_nor2_1 _17389_ (.A(_10575_),
    .B(net175),
    .Y(_10576_));
 sg13g2_a22oi_1 _17390_ (.Y(_10577_),
    .B1(_10573_),
    .B2(_10576_),
    .A2(_10571_),
    .A1(net537));
 sg13g2_buf_1 _17391_ (.A(_10577_),
    .X(_10578_));
 sg13g2_o21ai_1 _17392_ (.B1(net175),
    .Y(_10579_),
    .A1(_10569_),
    .A2(_10575_));
 sg13g2_nor3_1 _17393_ (.A(_10569_),
    .B(_10575_),
    .C(net175),
    .Y(_10580_));
 sg13g2_a21o_1 _17394_ (.A2(_10579_),
    .A1(net1022),
    .B1(_10580_),
    .X(_10581_));
 sg13g2_inv_1 _17395_ (.Y(_10582_),
    .A(_10581_));
 sg13g2_inv_1 _17396_ (.Y(_10583_),
    .A(_08544_));
 sg13g2_buf_1 _17397_ (.A(\cpu.ex.mmu_read[14] ),
    .X(_10584_));
 sg13g2_mux2_1 _17398_ (.A0(\cpu.ex.r_lr[14] ),
    .A1(net1109),
    .S(net539),
    .X(_10585_));
 sg13g2_a22oi_1 _17399_ (.Y(_10586_),
    .B1(_10585_),
    .B2(net675),
    .A2(_10546_),
    .A1(\cpu.ex.r_epc[14] ));
 sg13g2_nor2b_1 _17400_ (.A(net1026),
    .B_N(_10395_),
    .Y(_10587_));
 sg13g2_buf_2 _17401_ (.A(_10587_),
    .X(_10588_));
 sg13g2_nand3_1 _17402_ (.B(net679),
    .C(_10588_),
    .A(\cpu.ex.r_11[14] ),
    .Y(_10589_));
 sg13g2_o21ai_1 _17403_ (.B1(_10589_),
    .Y(_10590_),
    .A1(net680),
    .A2(_10586_));
 sg13g2_nand2_1 _17404_ (.Y(_10591_),
    .A(net538),
    .B(_10590_));
 sg13g2_and2_1 _17405_ (.A(\cpu.ex.r_9[14] ),
    .B(net538),
    .X(_10592_));
 sg13g2_nor2b_1 _17406_ (.A(net538),
    .B_N(\cpu.ex.r_stmp[14] ),
    .Y(_10593_));
 sg13g2_buf_8 _17407_ (.A(net912),
    .X(_10594_));
 sg13g2_and2_1 _17408_ (.A(net775),
    .B(net907),
    .X(_10595_));
 sg13g2_buf_1 _17409_ (.A(_10595_),
    .X(_10596_));
 sg13g2_a22oi_1 _17410_ (.Y(_10597_),
    .B1(_10593_),
    .B2(_10596_),
    .A2(_10592_),
    .A1(_10447_));
 sg13g2_buf_1 _17411_ (.A(net907),
    .X(_10598_));
 sg13g2_buf_1 _17412_ (.A(\cpu.ex.r_sp[14] ),
    .X(_10599_));
 sg13g2_a22oi_1 _17413_ (.Y(_10600_),
    .B1(net774),
    .B2(_10599_),
    .A2(net674),
    .A1(\cpu.ex.r_8[14] ));
 sg13g2_nor2_1 _17414_ (.A(net911),
    .B(net912),
    .Y(_10601_));
 sg13g2_nand2b_1 _17415_ (.Y(_10602_),
    .B(_10601_),
    .A_N(_10600_));
 sg13g2_nor2b_2 _17416_ (.A(net908),
    .B_N(net912),
    .Y(_10603_));
 sg13g2_nand3_1 _17417_ (.B(net538),
    .C(_10603_),
    .A(\cpu.ex.r_mult[30] ),
    .Y(_10604_));
 sg13g2_nand3_1 _17418_ (.B(net614),
    .C(_10588_),
    .A(\cpu.ex.r_10[14] ),
    .Y(_10605_));
 sg13g2_a21o_1 _17419_ (.A2(_10605_),
    .A1(_10604_),
    .B1(net675),
    .X(_10606_));
 sg13g2_inv_1 _17420_ (.Y(_10607_),
    .A(_00272_));
 sg13g2_mux4_1 _17421_ (.S0(net614),
    .A0(_10607_),
    .A1(\cpu.ex.r_14[14] ),
    .A2(\cpu.ex.r_13[14] ),
    .A3(\cpu.ex.r_12[14] ),
    .S1(net675),
    .X(_10608_));
 sg13g2_nand2_1 _17422_ (.Y(_10609_),
    .A(net781),
    .B(_10608_));
 sg13g2_and4_1 _17423_ (.A(_10597_),
    .B(_10602_),
    .C(_10606_),
    .D(_10609_),
    .X(_10610_));
 sg13g2_a21oi_1 _17424_ (.A1(_10591_),
    .A2(_10610_),
    .Y(_10611_),
    .B1(net536));
 sg13g2_a21o_1 _17425_ (.A2(net541),
    .A1(net622),
    .B1(_10611_),
    .X(_10612_));
 sg13g2_mux2_1 _17426_ (.A0(\cpu.dec.imm[14] ),
    .A1(_10612_),
    .S(_10374_),
    .X(_10613_));
 sg13g2_o21ai_1 _17427_ (.B1(net906),
    .Y(_10614_),
    .A1(_10371_),
    .A2(_10613_));
 sg13g2_o21ai_1 _17428_ (.B1(_10614_),
    .Y(_10615_),
    .A1(_10583_),
    .A2(net906));
 sg13g2_buf_1 _17429_ (.A(_10615_),
    .X(_10616_));
 sg13g2_a21oi_1 _17430_ (.A1(_10578_),
    .A2(_10582_),
    .Y(_10617_),
    .B1(_10616_));
 sg13g2_buf_1 _17431_ (.A(_00301_),
    .X(_10618_));
 sg13g2_nor2_1 _17432_ (.A(_08791_),
    .B(net906),
    .Y(_10619_));
 sg13g2_nand3_1 _17433_ (.B(net777),
    .C(_10494_),
    .A(\cpu.ex.r_11[10] ),
    .Y(_10620_));
 sg13g2_nand3_1 _17434_ (.B(_10486_),
    .C(_10402_),
    .A(\cpu.ex.r_12[10] ),
    .Y(_10621_));
 sg13g2_a21oi_1 _17435_ (.A1(_10620_),
    .A2(_10621_),
    .Y(_10622_),
    .B1(_10548_));
 sg13g2_nand3_1 _17436_ (.B(net616),
    .C(net910),
    .A(\cpu.ex.r_lr[10] ),
    .Y(_10623_));
 sg13g2_and2_1 _17437_ (.A(net1110),
    .B(_10382_),
    .X(_10624_));
 sg13g2_buf_1 _17438_ (.A(_10624_),
    .X(_10625_));
 sg13g2_nand3_1 _17439_ (.B(net676),
    .C(_10625_),
    .A(\cpu.ex.r_10[10] ),
    .Y(_10626_));
 sg13g2_a21oi_1 _17440_ (.A1(_10623_),
    .A2(_10626_),
    .Y(_10627_),
    .B1(net539));
 sg13g2_nand3_1 _17441_ (.B(net617),
    .C(net674),
    .A(\cpu.ex.r_13[10] ),
    .Y(_10628_));
 sg13g2_nand3_1 _17442_ (.B(net777),
    .C(net774),
    .A(\cpu.ex.r_epc[10] ),
    .Y(_10629_));
 sg13g2_a21oi_1 _17443_ (.A1(_10628_),
    .A2(_10629_),
    .Y(_10630_),
    .B1(net614));
 sg13g2_nor3_1 _17444_ (.A(_10622_),
    .B(_10627_),
    .C(_10630_),
    .Y(_10631_));
 sg13g2_nand3_1 _17445_ (.B(net616),
    .C(net674),
    .A(\cpu.ex.r_9[10] ),
    .Y(_10632_));
 sg13g2_buf_1 _17446_ (.A(\cpu.ex.r_sp[10] ),
    .X(_10633_));
 sg13g2_nand3_1 _17447_ (.B(net676),
    .C(net774),
    .A(_10633_),
    .Y(_10634_));
 sg13g2_nand3_1 _17448_ (.B(_10632_),
    .C(_10634_),
    .A(net777),
    .Y(_10635_));
 sg13g2_inv_1 _17449_ (.Y(_10636_),
    .A(_00268_));
 sg13g2_buf_1 _17450_ (.A(\cpu.ex.r_mult[26] ),
    .X(_10637_));
 sg13g2_mux2_1 _17451_ (.A0(_10636_),
    .A1(net1108),
    .S(_10548_),
    .X(_10638_));
 sg13g2_a21o_1 _17452_ (.A2(_10638_),
    .A1(_10494_),
    .B1(net777),
    .X(_10639_));
 sg13g2_a22oi_1 _17453_ (.Y(_10640_),
    .B1(_10538_),
    .B2(\cpu.ex.r_8[10] ),
    .A2(net613),
    .A1(\cpu.ex.r_14[10] ));
 sg13g2_nand3_1 _17454_ (.B(net617),
    .C(net774),
    .A(\cpu.ex.r_stmp[10] ),
    .Y(_10641_));
 sg13g2_o21ai_1 _17455_ (.B1(_10641_),
    .Y(_10642_),
    .A1(_10548_),
    .A2(_10640_));
 sg13g2_a22oi_1 _17456_ (.Y(_10643_),
    .B1(_10642_),
    .B2(net614),
    .A2(_10639_),
    .A1(_10635_));
 sg13g2_a21oi_1 _17457_ (.A1(_10631_),
    .A2(_10643_),
    .Y(_10644_),
    .B1(net536));
 sg13g2_buf_1 _17458_ (.A(\cpu.addr[10] ),
    .X(_10645_));
 sg13g2_nand2_1 _17459_ (.Y(_10646_),
    .A(net1107),
    .B(net541));
 sg13g2_nand3b_1 _17460_ (.B(_10646_),
    .C(net915),
    .Y(_10647_),
    .A_N(_10644_));
 sg13g2_inv_2 _17461_ (.Y(_10648_),
    .A(_10372_));
 sg13g2_inv_1 _17462_ (.Y(_10649_),
    .A(\cpu.dec.imm[10] ));
 sg13g2_nand2_1 _17463_ (.Y(_10650_),
    .A(_10648_),
    .B(_10649_));
 sg13g2_a21oi_1 _17464_ (.A1(_10647_),
    .A2(_10650_),
    .Y(_10651_),
    .B1(_10535_));
 sg13g2_or2_1 _17465_ (.X(_10652_),
    .B(_10651_),
    .A(_10619_));
 sg13g2_buf_1 _17466_ (.A(_10652_),
    .X(_10653_));
 sg13g2_xnor2_1 _17467_ (.Y(_10654_),
    .A(_10618_),
    .B(net204));
 sg13g2_nor2_1 _17468_ (.A(_08746_),
    .B(_10528_),
    .Y(_10655_));
 sg13g2_buf_1 _17469_ (.A(_10655_),
    .X(_10656_));
 sg13g2_nor2_1 _17470_ (.A(net777),
    .B(_10405_),
    .Y(_10657_));
 sg13g2_inv_1 _17471_ (.Y(_10658_),
    .A(\cpu.ex.r_epc[11] ));
 sg13g2_or2_1 _17472_ (.X(_10659_),
    .B(net912),
    .A(net908));
 sg13g2_nand3b_1 _17473_ (.B(_10407_),
    .C(net678),
    .Y(_10660_),
    .A_N(_00269_));
 sg13g2_o21ai_1 _17474_ (.B1(_10660_),
    .Y(_10661_),
    .A1(_10658_),
    .A2(_10659_));
 sg13g2_a221oi_1 _17475_ (.B2(_10412_),
    .C1(net676),
    .B1(_10661_),
    .A1(\cpu.ex.r_13[11] ),
    .Y(_10662_),
    .A2(_10657_));
 sg13g2_and3_1 _17476_ (.X(_10663_),
    .A(\cpu.ex.r_12[11] ),
    .B(net678),
    .C(net776));
 sg13g2_buf_1 _17477_ (.A(\cpu.ex.r_sp[11] ),
    .X(_10664_));
 sg13g2_and3_1 _17478_ (.X(_10665_),
    .A(_10664_),
    .B(_10492_),
    .C(net774));
 sg13g2_and3_1 _17479_ (.X(_10666_),
    .A(\cpu.ex.r_8[11] ),
    .B(_10485_),
    .C(_10588_));
 sg13g2_nor4_1 _17480_ (.A(net616),
    .B(_10663_),
    .C(_10665_),
    .D(_10666_),
    .Y(_10667_));
 sg13g2_nor2b_1 _17481_ (.A(_10407_),
    .B_N(net677),
    .Y(_10668_));
 sg13g2_nor2b_1 _17482_ (.A(net1027),
    .B_N(net1028),
    .Y(_10669_));
 sg13g2_a22oi_1 _17483_ (.Y(_10670_),
    .B1(_10669_),
    .B2(\cpu.ex.r_14[11] ),
    .A2(_10668_),
    .A1(\cpu.ex.r_mult[27] ));
 sg13g2_nand2b_1 _17484_ (.Y(_10671_),
    .B(net613),
    .A_N(_10670_));
 sg13g2_o21ai_1 _17485_ (.B1(_10671_),
    .Y(_10672_),
    .A1(_10662_),
    .A2(_10667_));
 sg13g2_mux2_1 _17486_ (.A0(\cpu.ex.r_9[11] ),
    .A1(\cpu.ex.r_11[11] ),
    .S(net783),
    .X(_10673_));
 sg13g2_a22oi_1 _17487_ (.Y(_10674_),
    .B1(_10673_),
    .B2(_10445_),
    .A2(_10513_),
    .A1(\cpu.ex.r_10[11] ));
 sg13g2_nand3_1 _17488_ (.B(net676),
    .C(net613),
    .A(\cpu.ex.r_stmp[11] ),
    .Y(_10675_));
 sg13g2_nand3_1 _17489_ (.B(net616),
    .C(_10538_),
    .A(\cpu.ex.r_lr[11] ),
    .Y(_10676_));
 sg13g2_a21o_1 _17490_ (.A2(_10676_),
    .A1(_10675_),
    .B1(net680),
    .X(_10677_));
 sg13g2_o21ai_1 _17491_ (.B1(_10677_),
    .Y(_10678_),
    .A1(_10440_),
    .A2(_10674_));
 sg13g2_o21ai_1 _17492_ (.B1(net540),
    .Y(_10679_),
    .A1(_10672_),
    .A2(_10678_));
 sg13g2_buf_2 _17493_ (.A(\cpu.addr[11] ),
    .X(_10680_));
 sg13g2_nand2_1 _17494_ (.Y(_10681_),
    .A(_10680_),
    .B(_10389_));
 sg13g2_nand3_1 _17495_ (.B(_10679_),
    .C(_10681_),
    .A(net915),
    .Y(_10682_));
 sg13g2_or2_1 _17496_ (.X(_10683_),
    .B(\cpu.dec.imm[11] ),
    .A(net1029));
 sg13g2_a21oi_1 _17497_ (.A1(_10682_),
    .A2(_10683_),
    .Y(_10684_),
    .B1(_10535_));
 sg13g2_buf_2 _17498_ (.A(_10684_),
    .X(_10685_));
 sg13g2_or2_1 _17499_ (.X(_10686_),
    .B(_10685_),
    .A(_10656_));
 sg13g2_buf_1 _17500_ (.A(_10686_),
    .X(_10687_));
 sg13g2_nand2_1 _17501_ (.Y(_10688_),
    .A(net1108),
    .B(net615));
 sg13g2_nor2_1 _17502_ (.A(_10687_),
    .B(_10688_),
    .Y(_10689_));
 sg13g2_inv_1 _17503_ (.Y(_10690_),
    .A(_10618_));
 sg13g2_o21ai_1 _17504_ (.B1(net615),
    .Y(_10691_),
    .A1(net1108),
    .A2(_10690_));
 sg13g2_nor2_1 _17505_ (.A(_10619_),
    .B(_10651_),
    .Y(_10692_));
 sg13g2_nor2_1 _17506_ (.A(_10656_),
    .B(_10685_),
    .Y(_10693_));
 sg13g2_nor2_1 _17507_ (.A(_10692_),
    .B(_10693_),
    .Y(_10694_));
 sg13g2_o21ai_1 _17508_ (.B1(_10690_),
    .Y(_10695_),
    .A1(_10656_),
    .A2(_10685_));
 sg13g2_nor4_1 _17509_ (.A(net1108),
    .B(net550),
    .C(net204),
    .D(_10695_),
    .Y(_10696_));
 sg13g2_a221oi_1 _17510_ (.B2(_10694_),
    .C1(_10696_),
    .B1(_10691_),
    .A1(_10654_),
    .Y(_10697_),
    .A2(_10689_));
 sg13g2_nor2b_1 _17511_ (.A(_00267_),
    .B_N(_10411_),
    .Y(_10698_));
 sg13g2_nor2b_1 _17512_ (.A(_10419_),
    .B_N(\cpu.ex.r_lr[9] ),
    .Y(_10699_));
 sg13g2_a22oi_1 _17513_ (.Y(_10700_),
    .B1(_10699_),
    .B2(net910),
    .A2(_10698_),
    .A1(net781));
 sg13g2_nand3_1 _17514_ (.B(_10419_),
    .C(net674),
    .A(\cpu.ex.r_13[9] ),
    .Y(_10701_));
 sg13g2_a21oi_1 _17515_ (.A1(_10700_),
    .A2(_10701_),
    .Y(_10702_),
    .B1(_10479_));
 sg13g2_mux2_1 _17516_ (.A0(\cpu.ex.r_epc[9] ),
    .A1(\cpu.ex.r_11[9] ),
    .S(net784),
    .X(_10703_));
 sg13g2_mux2_1 _17517_ (.A0(\cpu.ex.r_8[9] ),
    .A1(\cpu.ex.r_9[9] ),
    .S(net677),
    .X(_10704_));
 sg13g2_a22oi_1 _17518_ (.Y(_10705_),
    .B1(_10704_),
    .B2(net674),
    .A2(_10703_),
    .A1(_10494_));
 sg13g2_buf_1 _17519_ (.A(\cpu.ex.r_sp[9] ),
    .X(_10706_));
 sg13g2_nand3_1 _17520_ (.B(_10397_),
    .C(_10513_),
    .A(_10706_),
    .Y(_10707_));
 sg13g2_o21ai_1 _17521_ (.B1(_10707_),
    .Y(_10708_),
    .A1(net539),
    .A2(_10705_));
 sg13g2_nand3_1 _17522_ (.B(net616),
    .C(net774),
    .A(\cpu.ex.r_mult[25] ),
    .Y(_10709_));
 sg13g2_nand3_1 _17523_ (.B(net676),
    .C(net674),
    .A(\cpu.ex.r_12[9] ),
    .Y(_10710_));
 sg13g2_a21oi_1 _17524_ (.A1(_10709_),
    .A2(_10710_),
    .Y(_10711_),
    .B1(net777));
 sg13g2_mux2_1 _17525_ (.A0(\cpu.ex.r_10[9] ),
    .A1(\cpu.ex.r_14[9] ),
    .S(net678),
    .X(_10712_));
 sg13g2_a22oi_1 _17526_ (.Y(_10713_),
    .B1(_10712_),
    .B2(net680),
    .A2(_10603_),
    .A1(\cpu.ex.r_stmp[9] ));
 sg13g2_nor2_1 _17527_ (.A(_10434_),
    .B(_10713_),
    .Y(_10714_));
 sg13g2_nor4_1 _17528_ (.A(_10702_),
    .B(_10708_),
    .C(_10711_),
    .D(_10714_),
    .Y(_10715_));
 sg13g2_buf_1 _17529_ (.A(\cpu.addr[9] ),
    .X(_10716_));
 sg13g2_nand2_1 _17530_ (.Y(_10717_),
    .A(_10716_),
    .B(net541));
 sg13g2_o21ai_1 _17531_ (.B1(_10717_),
    .Y(_10718_),
    .A1(net536),
    .A2(_10715_));
 sg13g2_or2_1 _17532_ (.X(_10719_),
    .B(\cpu.dec.imm[9] ),
    .A(_10373_));
 sg13g2_o21ai_1 _17533_ (.B1(_10719_),
    .Y(_10720_),
    .A1(_10648_),
    .A2(_10718_));
 sg13g2_nor2_1 _17534_ (.A(_08738_),
    .B(net906),
    .Y(_10721_));
 sg13g2_a21oi_1 _17535_ (.A1(net779),
    .A2(_10720_),
    .Y(_10722_),
    .B1(_10721_));
 sg13g2_buf_1 _17536_ (.A(_10722_),
    .X(_10723_));
 sg13g2_inv_1 _17537_ (.Y(_10724_),
    .A(_00266_));
 sg13g2_mux2_1 _17538_ (.A0(\cpu.ex.r_epc[8] ),
    .A1(\cpu.ex.r_11[8] ),
    .S(net784),
    .X(_10725_));
 sg13g2_a22oi_1 _17539_ (.Y(_10726_),
    .B1(_10725_),
    .B2(_10492_),
    .A2(net781),
    .A1(_10724_));
 sg13g2_buf_1 _17540_ (.A(\cpu.ex.r_sp[8] ),
    .X(_10727_));
 sg13g2_mux2_1 _17541_ (.A0(_10727_),
    .A1(\cpu.ex.r_stmp[8] ),
    .S(net678),
    .X(_10728_));
 sg13g2_nor2_1 _17542_ (.A(net911),
    .B(net908),
    .Y(_10729_));
 sg13g2_nand2_1 _17543_ (.Y(_10730_),
    .A(_10728_),
    .B(_10729_));
 sg13g2_o21ai_1 _17544_ (.B1(_10730_),
    .Y(_10731_),
    .A1(_10479_),
    .A2(_10726_));
 sg13g2_nand2_1 _17545_ (.Y(_10732_),
    .A(net679),
    .B(_10731_));
 sg13g2_a22oi_1 _17546_ (.Y(_10733_),
    .B1(net774),
    .B2(\cpu.ex.r_mult[24] ),
    .A2(_10509_),
    .A1(\cpu.ex.r_13[8] ));
 sg13g2_and2_1 _17547_ (.A(_10400_),
    .B(net1026),
    .X(_10734_));
 sg13g2_buf_1 _17548_ (.A(_10734_),
    .X(_10735_));
 sg13g2_nor2b_1 _17549_ (.A(_10733_),
    .B_N(_10735_),
    .Y(_10736_));
 sg13g2_a22oi_1 _17550_ (.Y(_10737_),
    .B1(_10538_),
    .B2(\cpu.ex.r_8[8] ),
    .A2(_10482_),
    .A1(\cpu.ex.r_14[8] ));
 sg13g2_nor2b_1 _17551_ (.A(_10737_),
    .B_N(_10669_),
    .Y(_10738_));
 sg13g2_a22oi_1 _17552_ (.Y(_10739_),
    .B1(_10513_),
    .B2(\cpu.ex.r_10[8] ),
    .A2(_10428_),
    .A1(\cpu.ex.r_9[8] ));
 sg13g2_nor2_1 _17553_ (.A(_10440_),
    .B(_10739_),
    .Y(_10740_));
 sg13g2_nand3_1 _17554_ (.B(_10478_),
    .C(net781),
    .A(\cpu.ex.r_12[8] ),
    .Y(_10741_));
 sg13g2_nand3_1 _17555_ (.B(net616),
    .C(_10397_),
    .A(\cpu.ex.r_lr[8] ),
    .Y(_10742_));
 sg13g2_a21oi_1 _17556_ (.A1(_10741_),
    .A2(_10742_),
    .Y(_10743_),
    .B1(net679));
 sg13g2_nor4_1 _17557_ (.A(_10736_),
    .B(_10738_),
    .C(_10740_),
    .D(_10743_),
    .Y(_10744_));
 sg13g2_a21oi_1 _17558_ (.A1(_10732_),
    .A2(_10744_),
    .Y(_10745_),
    .B1(net536));
 sg13g2_nand2_1 _17559_ (.Y(_10746_),
    .A(_09278_),
    .B(_10388_));
 sg13g2_nand2_1 _17560_ (.Y(_10747_),
    .A(net1029),
    .B(_10746_));
 sg13g2_or2_1 _17561_ (.X(_10748_),
    .B(\cpu.dec.imm[8] ),
    .A(net1029));
 sg13g2_o21ai_1 _17562_ (.B1(_10748_),
    .Y(_10749_),
    .A1(_10745_),
    .A2(_10747_));
 sg13g2_nor2_1 _17563_ (.A(_08757_),
    .B(net906),
    .Y(_10750_));
 sg13g2_a21o_1 _17564_ (.A2(_10749_),
    .A1(net779),
    .B1(_10750_),
    .X(_10751_));
 sg13g2_buf_1 _17565_ (.A(_10751_),
    .X(_10752_));
 sg13g2_buf_1 _17566_ (.A(_10752_),
    .X(_10753_));
 sg13g2_buf_1 _17567_ (.A(_00303_),
    .X(_10754_));
 sg13g2_nor2_1 _17568_ (.A(net1106),
    .B(_09463_),
    .Y(_10755_));
 sg13g2_a21oi_1 _17569_ (.A1(net779),
    .A2(_10749_),
    .Y(_10756_),
    .B1(_10750_));
 sg13g2_buf_2 _17570_ (.A(_10756_),
    .X(_10757_));
 sg13g2_mux2_1 _17571_ (.A0(net1106),
    .A1(_10755_),
    .S(_10757_),
    .X(_10758_));
 sg13g2_buf_1 _17572_ (.A(_00302_),
    .X(_10759_));
 sg13g2_a22oi_1 _17573_ (.Y(_10760_),
    .B1(_10758_),
    .B2(_10759_),
    .A2(net203),
    .A1(net550));
 sg13g2_nor2_1 _17574_ (.A(_10759_),
    .B(net550),
    .Y(_10761_));
 sg13g2_buf_1 _17575_ (.A(_10761_),
    .X(_10762_));
 sg13g2_xnor2_1 _17576_ (.Y(_10763_),
    .A(net1106),
    .B(_10752_));
 sg13g2_nand3_1 _17577_ (.B(_10762_),
    .C(_10763_),
    .A(_10723_),
    .Y(_10764_));
 sg13g2_o21ai_1 _17578_ (.B1(_10764_),
    .Y(_10765_),
    .A1(_10723_),
    .A2(_10760_));
 sg13g2_nand2b_1 _17579_ (.Y(_10766_),
    .B(_10765_),
    .A_N(_10697_));
 sg13g2_buf_1 _17580_ (.A(_10766_),
    .X(_10767_));
 sg13g2_nand2_1 _17581_ (.Y(_10768_),
    .A(_10477_),
    .B(net782));
 sg13g2_a22oi_1 _17582_ (.Y(_10769_),
    .B1(net907),
    .B2(\cpu.ex.r_stmp[1] ),
    .A2(net776),
    .A1(\cpu.ex.r_12[1] ));
 sg13g2_nand3_1 _17583_ (.B(_10513_),
    .C(_10588_),
    .A(\cpu.ex.r_10[1] ),
    .Y(_10770_));
 sg13g2_o21ai_1 _17584_ (.B1(_10770_),
    .Y(_10771_),
    .A1(_10768_),
    .A2(_10769_));
 sg13g2_buf_1 _17585_ (.A(\cpu.ex.r_sp[1] ),
    .X(_10772_));
 sg13g2_and2_1 _17586_ (.A(net911),
    .B(net914),
    .X(_10773_));
 sg13g2_a22oi_1 _17587_ (.Y(_10774_),
    .B1(_10773_),
    .B2(\cpu.ex.r_11[1] ),
    .A2(_10729_),
    .A1(_10772_));
 sg13g2_inv_1 _17588_ (.Y(_10775_),
    .A(\cpu.ex.r_14[1] ));
 sg13g2_nand3b_1 _17589_ (.B(_10409_),
    .C(_10438_),
    .Y(_10776_),
    .A_N(net1027));
 sg13g2_o21ai_1 _17590_ (.B1(net782),
    .Y(_10777_),
    .A1(_10775_),
    .A2(_10776_));
 sg13g2_nand3b_1 _17591_ (.B(net783),
    .C(_10777_),
    .Y(_10778_),
    .A_N(_10774_));
 sg13g2_mux2_1 _17592_ (.A0(\cpu.ex.r_lr[1] ),
    .A1(\cpu.ex.r_9[1] ),
    .S(net908),
    .X(_10779_));
 sg13g2_and2_1 _17593_ (.A(_10538_),
    .B(_10779_),
    .X(_10780_));
 sg13g2_nand2b_1 _17594_ (.Y(_10781_),
    .B(_10406_),
    .A_N(_00259_));
 sg13g2_nand2b_1 _17595_ (.Y(_10782_),
    .B(\cpu.ex.r_mult[17] ),
    .A_N(net914));
 sg13g2_nand2_1 _17596_ (.Y(_10783_),
    .A(_10410_),
    .B(net782));
 sg13g2_a21oi_1 _17597_ (.A1(_10781_),
    .A2(_10782_),
    .Y(_10784_),
    .B1(_10783_));
 sg13g2_o21ai_1 _17598_ (.B1(_10442_),
    .Y(_10785_),
    .A1(_10780_),
    .A2(_10784_));
 sg13g2_nand3b_1 _17599_ (.B(_10778_),
    .C(_10785_),
    .Y(_10786_),
    .A_N(_10771_));
 sg13g2_nor2_1 _17600_ (.A(_10426_),
    .B(_10405_),
    .Y(_10787_));
 sg13g2_a221oi_1 _17601_ (.B2(\cpu.ex.r_8[1] ),
    .C1(net775),
    .B1(_10787_),
    .A1(\cpu.ex.r_epc[1] ),
    .Y(_10788_),
    .A2(_10506_));
 sg13g2_buf_1 _17602_ (.A(\cpu.ex.r_prev_ie ),
    .X(_10789_));
 sg13g2_and3_1 _17603_ (.X(_10790_),
    .A(\cpu.ex.r_13[1] ),
    .B(net911),
    .C(net908));
 sg13g2_a21o_1 _17604_ (.A2(_10729_),
    .A1(_10789_),
    .B1(_10790_),
    .X(_10791_));
 sg13g2_a221oi_1 _17605_ (.B2(_10485_),
    .C1(_10777_),
    .B1(_10791_),
    .A1(\cpu.ex.mmu_read[1] ),
    .Y(_10792_),
    .A2(_10425_));
 sg13g2_nor3_1 _17606_ (.A(_09351_),
    .B(_10383_),
    .C(_10385_),
    .Y(_10793_));
 sg13g2_a21oi_1 _17607_ (.A1(_10391_),
    .A2(_10793_),
    .Y(_10794_),
    .B1(_10648_));
 sg13g2_o21ai_1 _17608_ (.B1(_10794_),
    .Y(_10795_),
    .A1(_10788_),
    .A2(_10792_));
 sg13g2_buf_1 _17609_ (.A(\cpu.dec.imm[1] ),
    .X(_10796_));
 sg13g2_inv_1 _17610_ (.Y(_10797_),
    .A(_10796_));
 sg13g2_a22oi_1 _17611_ (.Y(_10798_),
    .B1(net536),
    .B2(_10794_),
    .A2(_10648_),
    .A1(_10797_));
 sg13g2_o21ai_1 _17612_ (.B1(_10798_),
    .Y(_10799_),
    .A1(_10786_),
    .A2(_10795_));
 sg13g2_buf_1 _17613_ (.A(_10799_),
    .X(_10800_));
 sg13g2_nor2_1 _17614_ (.A(_08975_),
    .B(_10527_),
    .Y(_10801_));
 sg13g2_a21o_1 _17615_ (.A2(_10800_),
    .A1(net779),
    .B1(_10801_),
    .X(_10802_));
 sg13g2_buf_2 _17616_ (.A(_10802_),
    .X(_10803_));
 sg13g2_nor2_1 _17617_ (.A(\cpu.ex.pc[2] ),
    .B(_10527_),
    .Y(_10804_));
 sg13g2_buf_1 _17618_ (.A(\cpu.dec.imm[2] ),
    .X(_10805_));
 sg13g2_nor3_1 _17619_ (.A(_10805_),
    .B(_10372_),
    .C(_10535_),
    .Y(_10806_));
 sg13g2_nor2_1 _17620_ (.A(_10804_),
    .B(_10806_),
    .Y(_10807_));
 sg13g2_nand3_1 _17621_ (.B(_10391_),
    .C(_10392_),
    .A(_09346_),
    .Y(_10808_));
 sg13g2_inv_1 _17622_ (.Y(_10809_),
    .A(_10776_));
 sg13g2_mux2_1 _17623_ (.A0(\cpu.ex.r_10[2] ),
    .A1(\cpu.ex.r_14[2] ),
    .S(net782),
    .X(_10810_));
 sg13g2_nor2b_1 _17624_ (.A(net775),
    .B_N(\cpu.ex.r_epc[2] ),
    .Y(_10811_));
 sg13g2_a22oi_1 _17625_ (.Y(_10812_),
    .B1(_10811_),
    .B2(_10506_),
    .A2(_10810_),
    .A1(_10809_));
 sg13g2_nand2b_1 _17626_ (.Y(_10813_),
    .B(net912),
    .A_N(_00260_));
 sg13g2_nand2b_1 _17627_ (.Y(_10814_),
    .B(\cpu.ex.r_11[2] ),
    .A_N(_10416_));
 sg13g2_nand3_1 _17628_ (.B(net1025),
    .C(_10438_),
    .A(_10422_),
    .Y(_10815_));
 sg13g2_a21o_1 _17629_ (.A2(_10814_),
    .A1(_10813_),
    .B1(_10815_),
    .X(_10816_));
 sg13g2_mux2_1 _17630_ (.A0(\cpu.ex.r_12[2] ),
    .A1(\cpu.ex.r_13[2] ),
    .S(_10422_),
    .X(_10817_));
 sg13g2_nand3_1 _17631_ (.B(net776),
    .C(_10817_),
    .A(_10594_),
    .Y(_10818_));
 sg13g2_buf_1 _17632_ (.A(\cpu.ex.mmu_read[2] ),
    .X(_10819_));
 sg13g2_mux2_1 _17633_ (.A0(\cpu.ex.r_lr[2] ),
    .A1(_10819_),
    .S(net912),
    .X(_10820_));
 sg13g2_nand3_1 _17634_ (.B(_10424_),
    .C(_10820_),
    .A(_10426_),
    .Y(_10821_));
 sg13g2_mux2_1 _17635_ (.A0(\cpu.ex.r_stmp[2] ),
    .A1(\cpu.ex.r_mult[18] ),
    .S(net911),
    .X(_10822_));
 sg13g2_nand3_1 _17636_ (.B(net907),
    .C(_10822_),
    .A(_10417_),
    .Y(_10823_));
 sg13g2_and4_1 _17637_ (.A(_10816_),
    .B(_10818_),
    .C(_10821_),
    .D(_10823_),
    .X(_10824_));
 sg13g2_buf_1 _17638_ (.A(\cpu.ex.r_sp[2] ),
    .X(_10825_));
 sg13g2_nor2_1 _17639_ (.A(_10659_),
    .B(_10434_),
    .Y(_10826_));
 sg13g2_nor3_1 _17640_ (.A(net778),
    .B(net913),
    .C(_10440_),
    .Y(_10827_));
 sg13g2_nand3b_1 _17641_ (.B(net782),
    .C(_08452_),
    .Y(_10828_),
    .A_N(net914));
 sg13g2_nand3b_1 _17642_ (.B(net914),
    .C(\cpu.ex.r_8[2] ),
    .Y(_10829_),
    .A_N(_10416_));
 sg13g2_or2_1 _17643_ (.X(_10830_),
    .B(net913),
    .A(net909));
 sg13g2_a21oi_1 _17644_ (.A1(_10828_),
    .A2(_10829_),
    .Y(_10831_),
    .B1(_10830_));
 sg13g2_a221oi_1 _17645_ (.B2(\cpu.ex.r_9[2] ),
    .C1(_10831_),
    .B1(_10827_),
    .A1(_10825_),
    .Y(_10832_),
    .A2(_10826_));
 sg13g2_and4_1 _17646_ (.A(_10808_),
    .B(_10812_),
    .C(_10824_),
    .D(_10832_),
    .X(_10833_));
 sg13g2_and2_1 _17647_ (.A(_10522_),
    .B(_10808_),
    .X(_10834_));
 sg13g2_nor2_2 _17648_ (.A(_10648_),
    .B(_10535_),
    .Y(_10835_));
 sg13g2_o21ai_1 _17649_ (.B1(_10835_),
    .Y(_10836_),
    .A1(_10833_),
    .A2(_10834_));
 sg13g2_nand2_1 _17650_ (.Y(_10837_),
    .A(_10807_),
    .B(_10836_));
 sg13g2_buf_2 _17651_ (.A(_10837_),
    .X(_10838_));
 sg13g2_a21oi_1 _17652_ (.A1(_10803_),
    .A2(_10838_),
    .Y(_10839_),
    .B1(net615));
 sg13g2_buf_1 _17653_ (.A(_00309_),
    .X(_10840_));
 sg13g2_inv_2 _17654_ (.Y(_10841_),
    .A(_10840_));
 sg13g2_nor3_1 _17655_ (.A(_10841_),
    .B(_10803_),
    .C(_10838_),
    .Y(_10842_));
 sg13g2_nor2_1 _17656_ (.A(_10839_),
    .B(_10842_),
    .Y(_10843_));
 sg13g2_buf_2 _17657_ (.A(_00308_),
    .X(_10844_));
 sg13g2_o21ai_1 _17658_ (.B1(_10838_),
    .Y(_10845_),
    .A1(_10841_),
    .A2(_10803_));
 sg13g2_nand2_1 _17659_ (.Y(_10846_),
    .A(_10844_),
    .B(_10845_));
 sg13g2_buf_1 _17660_ (.A(_00305_),
    .X(_10847_));
 sg13g2_inv_1 _17661_ (.Y(_10848_),
    .A(_10847_));
 sg13g2_nand2_1 _17662_ (.Y(_10849_),
    .A(_10372_),
    .B(_10474_));
 sg13g2_nand3_1 _17663_ (.B(net778),
    .C(net613),
    .A(\cpu.ex.r_stmp[5] ),
    .Y(_10850_));
 sg13g2_nand3_1 _17664_ (.B(net780),
    .C(_10538_),
    .A(\cpu.ex.r_lr[5] ),
    .Y(_10851_));
 sg13g2_a21oi_1 _17665_ (.A1(_10850_),
    .A2(_10851_),
    .Y(_10852_),
    .B1(net784));
 sg13g2_nand3_1 _17666_ (.B(_10428_),
    .C(net781),
    .A(\cpu.ex.r_13[5] ),
    .Y(_10853_));
 sg13g2_nand3_1 _17667_ (.B(_10513_),
    .C(_10588_),
    .A(\cpu.ex.r_10[5] ),
    .Y(_10854_));
 sg13g2_mux2_1 _17668_ (.A0(\cpu.ex.r_epc[5] ),
    .A1(\cpu.ex.r_mult[21] ),
    .S(net782),
    .X(_10855_));
 sg13g2_nand3_1 _17669_ (.B(net907),
    .C(_10855_),
    .A(net780),
    .Y(_10856_));
 sg13g2_nand3_1 _17670_ (.B(_10854_),
    .C(_10856_),
    .A(_10853_),
    .Y(_10857_));
 sg13g2_nand2_1 _17671_ (.Y(_10858_),
    .A(net778),
    .B(_10491_));
 sg13g2_buf_1 _17672_ (.A(\cpu.ex.r_sp[5] ),
    .X(_10859_));
 sg13g2_a22oi_1 _17673_ (.Y(_10860_),
    .B1(net907),
    .B2(_10859_),
    .A2(net776),
    .A1(\cpu.ex.r_8[5] ));
 sg13g2_nand3b_1 _17674_ (.B(net780),
    .C(\cpu.ex.r_11[5] ),
    .Y(_10861_),
    .A_N(net775));
 sg13g2_nand3b_1 _17675_ (.B(net775),
    .C(\cpu.ex.r_14[5] ),
    .Y(_10862_),
    .A_N(net909));
 sg13g2_nand2_1 _17676_ (.Y(_10863_),
    .A(net783),
    .B(net914));
 sg13g2_a21o_1 _17677_ (.A2(_10862_),
    .A1(_10861_),
    .B1(_10863_),
    .X(_10864_));
 sg13g2_o21ai_1 _17678_ (.B1(_10864_),
    .Y(_10865_),
    .A1(_10858_),
    .A2(_10860_));
 sg13g2_inv_1 _17679_ (.Y(_10866_),
    .A(_00263_));
 sg13g2_a22oi_1 _17680_ (.Y(_10867_),
    .B1(_10494_),
    .B2(_10866_),
    .A2(_10394_),
    .A1(\cpu.ex.r_12[5] ));
 sg13g2_nand4_1 _17681_ (.B(net780),
    .C(_10491_),
    .A(\cpu.ex.r_9[5] ),
    .Y(_10868_),
    .D(net776));
 sg13g2_o21ai_1 _17682_ (.B1(_10868_),
    .Y(_10869_),
    .A1(_10435_),
    .A2(_10867_));
 sg13g2_nor4_1 _17683_ (.A(_10852_),
    .B(_10857_),
    .C(_10865_),
    .D(_10869_),
    .Y(_10870_));
 sg13g2_nand2_1 _17684_ (.Y(_10871_),
    .A(_10122_),
    .B(_10388_));
 sg13g2_o21ai_1 _17685_ (.B1(_10871_),
    .Y(_10872_),
    .A1(_10522_),
    .A2(_10870_));
 sg13g2_nor2_1 _17686_ (.A(_10373_),
    .B(\cpu.dec.imm[5] ),
    .Y(_10873_));
 sg13g2_a22oi_1 _17687_ (.Y(_10874_),
    .B1(net779),
    .B2(_10873_),
    .A2(_10369_),
    .A1(_08808_));
 sg13g2_o21ai_1 _17688_ (.B1(_10874_),
    .Y(_10875_),
    .A1(_10849_),
    .A2(_10872_));
 sg13g2_buf_2 _17689_ (.A(_10875_),
    .X(_10876_));
 sg13g2_buf_8 _17690_ (.A(_10876_),
    .X(_10877_));
 sg13g2_nand3_1 _17691_ (.B(_10391_),
    .C(_10392_),
    .A(_09490_),
    .Y(_10878_));
 sg13g2_mux2_1 _17692_ (.A0(\cpu.ex.r_10[4] ),
    .A1(\cpu.ex.r_14[4] ),
    .S(net775),
    .X(_10879_));
 sg13g2_inv_1 _17693_ (.Y(_10880_),
    .A(\cpu.ex.r_9[4] ));
 sg13g2_nand2b_1 _17694_ (.Y(_10881_),
    .B(_10384_),
    .A_N(_10377_));
 sg13g2_buf_1 _17695_ (.A(_10881_),
    .X(_10882_));
 sg13g2_nand3b_1 _17696_ (.B(net775),
    .C(\cpu.ex.r_12[4] ),
    .Y(_10883_),
    .A_N(net780));
 sg13g2_o21ai_1 _17697_ (.B1(_10883_),
    .Y(_10884_),
    .A1(_10880_),
    .A2(_10882_));
 sg13g2_nand2b_1 _17698_ (.Y(_10885_),
    .B(_10418_),
    .A_N(_00262_));
 sg13g2_nand2b_1 _17699_ (.Y(_10886_),
    .B(\cpu.ex.r_11[4] ),
    .A_N(_10594_));
 sg13g2_a21oi_1 _17700_ (.A1(_10885_),
    .A2(_10886_),
    .Y(_10887_),
    .B1(_10815_));
 sg13g2_a221oi_1 _17701_ (.B2(_10508_),
    .C1(_10887_),
    .B1(_10884_),
    .A1(_10809_),
    .Y(_10888_),
    .A2(_10879_));
 sg13g2_inv_1 _17702_ (.Y(_10889_),
    .A(\cpu.ex.r_8[4] ));
 sg13g2_nand3b_1 _17703_ (.B(net775),
    .C(_08397_),
    .Y(_10890_),
    .A_N(_10406_));
 sg13g2_o21ai_1 _17704_ (.B1(_10890_),
    .Y(_10891_),
    .A1(_10889_),
    .A2(_10440_));
 sg13g2_nor2b_1 _17705_ (.A(net780),
    .B_N(\cpu.ex.r_stmp[4] ),
    .Y(_10892_));
 sg13g2_a22oi_1 _17706_ (.Y(_10893_),
    .B1(_10892_),
    .B2(_10596_),
    .A2(_10891_),
    .A1(_10394_));
 sg13g2_buf_1 _17707_ (.A(\cpu.ex.r_sp[4] ),
    .X(_10894_));
 sg13g2_inv_1 _17708_ (.Y(_10895_),
    .A(\cpu.ex.r_13[4] ));
 sg13g2_nand3b_1 _17709_ (.B(_10411_),
    .C(\cpu.ex.r_mult[20] ),
    .Y(_10896_),
    .A_N(net914));
 sg13g2_o21ai_1 _17710_ (.B1(_10896_),
    .Y(_10897_),
    .A1(_10895_),
    .A2(_10405_));
 sg13g2_mux2_1 _17711_ (.A0(\cpu.ex.r_lr[4] ),
    .A1(\cpu.ex.r_epc[4] ),
    .S(net913),
    .X(_10898_));
 sg13g2_and3_1 _17712_ (.X(_10899_),
    .A(net780),
    .B(_10397_),
    .C(_10898_));
 sg13g2_a221oi_1 _17713_ (.B2(_10897_),
    .C1(_10899_),
    .B1(_10735_),
    .A1(_10894_),
    .Y(_10900_),
    .A2(_10826_));
 sg13g2_and4_1 _17714_ (.A(_10878_),
    .B(_10888_),
    .C(_10893_),
    .D(_10900_),
    .X(_10901_));
 sg13g2_and2_1 _17715_ (.A(net536),
    .B(_10878_),
    .X(_10902_));
 sg13g2_o21ai_1 _17716_ (.B1(_10835_),
    .Y(_10903_),
    .A1(_10901_),
    .A2(_10902_));
 sg13g2_nor2_1 _17717_ (.A(net1029),
    .B(\cpu.dec.imm[4] ),
    .Y(_10904_));
 sg13g2_a22oi_1 _17718_ (.Y(_10905_),
    .B1(_10474_),
    .B2(_10904_),
    .A2(_10369_),
    .A1(_08562_));
 sg13g2_nand2_1 _17719_ (.Y(_10906_),
    .A(_10903_),
    .B(_10905_));
 sg13g2_buf_2 _17720_ (.A(_10906_),
    .X(_10907_));
 sg13g2_buf_1 _17721_ (.A(_10907_),
    .X(_10908_));
 sg13g2_buf_1 _17722_ (.A(_00306_),
    .X(_10909_));
 sg13g2_inv_2 _17723_ (.Y(_10910_),
    .A(_10909_));
 sg13g2_a22oi_1 _17724_ (.Y(_10911_),
    .B1(net235),
    .B2(_10910_),
    .A2(net236),
    .A1(_10848_));
 sg13g2_or2_1 _17725_ (.X(_10912_),
    .B(_10911_),
    .A(_09463_));
 sg13g2_buf_2 _17726_ (.A(_00307_),
    .X(_10913_));
 sg13g2_nand2_1 _17727_ (.Y(_10914_),
    .A(_09338_),
    .B(_10388_));
 sg13g2_nand3b_1 _17728_ (.B(net908),
    .C(\cpu.ex.r_9[3] ),
    .Y(_10915_),
    .A_N(net1025));
 sg13g2_nand3b_1 _17729_ (.B(net1025),
    .C(\cpu.ex.r_epc[3] ),
    .Y(_10916_),
    .A_N(net1028));
 sg13g2_a21o_1 _17730_ (.A2(_10916_),
    .A1(_10915_),
    .B1(_10882_),
    .X(_10917_));
 sg13g2_buf_1 _17731_ (.A(\cpu.ex.r_sp[3] ),
    .X(_10918_));
 sg13g2_nand3_1 _17732_ (.B(_10397_),
    .C(_10513_),
    .A(_10918_),
    .Y(_10919_));
 sg13g2_nand2b_1 _17733_ (.Y(_10920_),
    .B(net1025),
    .A_N(_00261_));
 sg13g2_nand2b_1 _17734_ (.Y(_10921_),
    .B(\cpu.ex.r_13[3] ),
    .A_N(net1025));
 sg13g2_a21o_1 _17735_ (.A2(_10921_),
    .A1(_10920_),
    .B1(_10499_),
    .X(_10922_));
 sg13g2_mux4_1 _17736_ (.S0(_10379_),
    .A0(\cpu.ex.r_8[3] ),
    .A1(\cpu.ex.r_10[3] ),
    .A2(\cpu.ex.r_12[3] ),
    .A3(\cpu.ex.r_14[3] ),
    .S1(_10401_),
    .X(_10923_));
 sg13g2_nand2_1 _17737_ (.Y(_10924_),
    .A(_10669_),
    .B(_10923_));
 sg13g2_nand4_1 _17738_ (.B(_10919_),
    .C(_10922_),
    .A(_10917_),
    .Y(_10925_),
    .D(_10924_));
 sg13g2_mux2_1 _17739_ (.A0(\cpu.ex.r_stmp[3] ),
    .A1(\cpu.ex.r_mult[19] ),
    .S(net1027),
    .X(_10926_));
 sg13g2_nand3_1 _17740_ (.B(net907),
    .C(_10926_),
    .A(net912),
    .Y(_10927_));
 sg13g2_nand4_1 _17741_ (.B(net911),
    .C(_10491_),
    .A(\cpu.ex.r_11[3] ),
    .Y(_10928_),
    .D(_10625_));
 sg13g2_nand3_1 _17742_ (.B(_10402_),
    .C(net910),
    .A(_08394_),
    .Y(_10929_));
 sg13g2_buf_1 _17743_ (.A(\cpu.ex.mmu_read[3] ),
    .X(_10930_));
 sg13g2_mux2_1 _17744_ (.A0(\cpu.ex.r_lr[3] ),
    .A1(_10930_),
    .S(net1026),
    .X(_10931_));
 sg13g2_nand3_1 _17745_ (.B(net910),
    .C(_10931_),
    .A(net911),
    .Y(_10932_));
 sg13g2_nand4_1 _17746_ (.B(_10928_),
    .C(_10929_),
    .A(_10927_),
    .Y(_10933_),
    .D(_10932_));
 sg13g2_o21ai_1 _17747_ (.B1(net540),
    .Y(_10934_),
    .A1(_10925_),
    .A2(_10933_));
 sg13g2_and3_1 _17748_ (.X(_10935_),
    .A(_10835_),
    .B(_10914_),
    .C(_10934_));
 sg13g2_buf_1 _17749_ (.A(_10935_),
    .X(_10936_));
 sg13g2_buf_1 _17750_ (.A(\cpu.dec.imm[3] ),
    .X(_10937_));
 sg13g2_nor2_1 _17751_ (.A(_10937_),
    .B(_10372_),
    .Y(_10938_));
 sg13g2_a22oi_1 _17752_ (.Y(_10939_),
    .B1(_10474_),
    .B2(_10938_),
    .A2(_10369_),
    .A1(_08563_));
 sg13g2_buf_1 _17753_ (.A(_10939_),
    .X(_10940_));
 sg13g2_inv_1 _17754_ (.Y(_10941_),
    .A(_10940_));
 sg13g2_nor2_1 _17755_ (.A(_10936_),
    .B(_10941_),
    .Y(_10942_));
 sg13g2_buf_8 _17756_ (.A(_10942_),
    .X(_10943_));
 sg13g2_o21ai_1 _17757_ (.B1(_10469_),
    .Y(_10944_),
    .A1(_10848_),
    .A2(net236));
 sg13g2_nand3_1 _17758_ (.B(_10914_),
    .C(_10934_),
    .A(_10835_),
    .Y(_10945_));
 sg13g2_buf_1 _17759_ (.A(_10945_),
    .X(_10946_));
 sg13g2_nand2_1 _17760_ (.Y(_10947_),
    .A(_10946_),
    .B(_10940_));
 sg13g2_buf_1 _17761_ (.A(_10947_),
    .X(_10948_));
 sg13g2_nand3_1 _17762_ (.B(net236),
    .C(_10907_),
    .A(net277),
    .Y(_10949_));
 sg13g2_nor2_1 _17763_ (.A(_10910_),
    .B(net235),
    .Y(_10950_));
 sg13g2_a221oi_1 _17764_ (.B2(_10949_),
    .C1(_10950_),
    .B1(_10944_),
    .A1(_10913_),
    .Y(_10951_),
    .A2(_10943_));
 sg13g2_and4_1 _17765_ (.A(_10843_),
    .B(_10846_),
    .C(_10912_),
    .D(_10951_),
    .X(_10952_));
 sg13g2_buf_1 _17766_ (.A(_10952_),
    .X(_10953_));
 sg13g2_or2_1 _17767_ (.X(_10954_),
    .B(_10806_),
    .A(_10804_));
 sg13g2_buf_1 _17768_ (.A(_10954_),
    .X(_10955_));
 sg13g2_nand3_1 _17769_ (.B(_10824_),
    .C(_10832_),
    .A(_10812_),
    .Y(_10956_));
 sg13g2_a221oi_1 _17770_ (.B2(_10956_),
    .C1(_10849_),
    .B1(net540),
    .A1(_09378_),
    .Y(_10957_),
    .A2(_10388_));
 sg13g2_buf_1 _17771_ (.A(_10957_),
    .X(_10958_));
 sg13g2_nor2_1 _17772_ (.A(_10955_),
    .B(_10958_),
    .Y(_10959_));
 sg13g2_nand2_1 _17773_ (.Y(_10960_),
    .A(_10841_),
    .B(_10803_));
 sg13g2_o21ai_1 _17774_ (.B1(_10960_),
    .Y(_10961_),
    .A1(_10844_),
    .A2(_10959_));
 sg13g2_buf_1 _17775_ (.A(\cpu.dec.imm[0] ),
    .X(_10962_));
 sg13g2_nor3_1 _17776_ (.A(_10962_),
    .B(net1029),
    .C(_10371_),
    .Y(_10963_));
 sg13g2_buf_1 _17777_ (.A(\cpu.ex.genblk3.r_prev_supmode ),
    .X(_10964_));
 sg13g2_mux2_1 _17778_ (.A0(_10964_),
    .A1(\cpu.ex.r_11[0] ),
    .S(net908),
    .X(_10965_));
 sg13g2_a221oi_1 _17779_ (.B2(_10491_),
    .C1(net778),
    .B1(_10965_),
    .A1(\cpu.ex.r_15[0] ),
    .Y(_10966_),
    .A2(_10430_));
 sg13g2_a21oi_1 _17780_ (.A1(\cpu.ex.r_stmp[0] ),
    .A2(_10603_),
    .Y(_10967_),
    .B1(net909));
 sg13g2_nor3_1 _17781_ (.A(_10485_),
    .B(_10966_),
    .C(_10967_),
    .Y(_10968_));
 sg13g2_a22oi_1 _17782_ (.Y(_10969_),
    .B1(_10601_),
    .B2(\cpu.ex.r_8[0] ),
    .A2(_10735_),
    .A1(\cpu.ex.r_13[0] ));
 sg13g2_nand4_1 _17783_ (.B(net909),
    .C(_10491_),
    .A(\cpu.ex.r_9[0] ),
    .Y(_10970_),
    .D(net776));
 sg13g2_o21ai_1 _17784_ (.B1(_10970_),
    .Y(_10971_),
    .A1(_10405_),
    .A2(_10969_));
 sg13g2_nand3_1 _17785_ (.B(_10410_),
    .C(_10588_),
    .A(\cpu.ex.r_10[0] ),
    .Y(_10972_));
 sg13g2_nand3_1 _17786_ (.B(_10485_),
    .C(_10603_),
    .A(_09285_),
    .Y(_10973_));
 sg13g2_a21oi_1 _17787_ (.A1(_10972_),
    .A2(_10973_),
    .Y(_10974_),
    .B1(_10442_));
 sg13g2_mux2_1 _17788_ (.A0(\cpu.ex.r_12[0] ),
    .A1(\cpu.ex.r_14[0] ),
    .S(net1025),
    .X(_10975_));
 sg13g2_nand3_1 _17789_ (.B(_10430_),
    .C(_10975_),
    .A(net778),
    .Y(_10976_));
 sg13g2_nand4_1 _17790_ (.B(net909),
    .C(_10417_),
    .A(\cpu.ex.r_mult[16] ),
    .Y(_10977_),
    .D(net907));
 sg13g2_nand2_1 _17791_ (.Y(_10978_),
    .A(_10976_),
    .B(_10977_));
 sg13g2_or4_1 _17792_ (.A(_10968_),
    .B(_10971_),
    .C(_10974_),
    .D(_10978_),
    .X(_10979_));
 sg13g2_nand2b_1 _17793_ (.Y(_10980_),
    .B(_10372_),
    .A_N(_10371_));
 sg13g2_a221oi_1 _17794_ (.B2(_10979_),
    .C1(_10980_),
    .B1(net540),
    .A1(_09358_),
    .Y(_10981_),
    .A2(_10388_));
 sg13g2_nor3_1 _17795_ (.A(_10369_),
    .B(_10963_),
    .C(_10981_),
    .Y(_10982_));
 sg13g2_buf_2 _17796_ (.A(_10982_),
    .X(_10983_));
 sg13g2_inv_2 _17797_ (.Y(_10984_),
    .A(_10983_));
 sg13g2_a21oi_1 _17798_ (.A1(_10469_),
    .A2(_10961_),
    .Y(_10985_),
    .B1(_10984_));
 sg13g2_a22oi_1 _17799_ (.Y(_10986_),
    .B1(_10494_),
    .B2(\cpu.ex.r_11[6] ),
    .A2(_10394_),
    .A1(\cpu.ex.r_8[6] ));
 sg13g2_nand3b_1 _17800_ (.B(net784),
    .C(\cpu.ex.r_9[6] ),
    .Y(_10987_),
    .A_N(net783));
 sg13g2_nand3b_1 _17801_ (.B(net783),
    .C(\cpu.ex.r_epc[6] ),
    .Y(_10988_),
    .A_N(net784));
 sg13g2_a21o_1 _17802_ (.A2(_10988_),
    .A1(_10987_),
    .B1(_10882_),
    .X(_10989_));
 sg13g2_o21ai_1 _17803_ (.B1(_10989_),
    .Y(_10990_),
    .A1(_10440_),
    .A2(_10986_));
 sg13g2_a21oi_1 _17804_ (.A1(\cpu.ex.r_14[6] ),
    .A2(_10436_),
    .Y(_10991_),
    .B1(_10990_));
 sg13g2_buf_1 _17805_ (.A(\cpu.ex.r_sp[6] ),
    .X(_10992_));
 sg13g2_nand2_1 _17806_ (.Y(_10993_),
    .A(_10992_),
    .B(_10450_));
 sg13g2_o21ai_1 _17807_ (.B1(_10993_),
    .Y(_10994_),
    .A1(_00264_),
    .A2(_10499_));
 sg13g2_nand3_1 _17808_ (.B(_10443_),
    .C(_10509_),
    .A(\cpu.ex.r_13[6] ),
    .Y(_10995_));
 sg13g2_nand3_1 _17809_ (.B(net778),
    .C(_10598_),
    .A(\cpu.ex.r_stmp[6] ),
    .Y(_10996_));
 sg13g2_buf_1 _17810_ (.A(\cpu.ex.r_mult[22] ),
    .X(_10997_));
 sg13g2_nand3_1 _17811_ (.B(_10443_),
    .C(net774),
    .A(_10997_),
    .Y(_10998_));
 sg13g2_nand3_1 _17812_ (.B(net778),
    .C(net776),
    .A(\cpu.ex.r_12[6] ),
    .Y(_10999_));
 sg13g2_nand4_1 _17813_ (.B(_10996_),
    .C(_10998_),
    .A(_10995_),
    .Y(_11000_),
    .D(_10999_));
 sg13g2_nand3_1 _17814_ (.B(net616),
    .C(net910),
    .A(\cpu.ex.r_lr[6] ),
    .Y(_11001_));
 sg13g2_nand3_1 _17815_ (.B(_10478_),
    .C(_10625_),
    .A(\cpu.ex.r_10[6] ),
    .Y(_11002_));
 sg13g2_a21oi_1 _17816_ (.A1(_11001_),
    .A2(_11002_),
    .Y(_11003_),
    .B1(net539));
 sg13g2_a221oi_1 _17817_ (.B2(net539),
    .C1(_11003_),
    .B1(_11000_),
    .A1(net679),
    .Y(_11004_),
    .A2(_10994_));
 sg13g2_a21oi_2 _17818_ (.B1(net536),
    .Y(_11005_),
    .A2(_11004_),
    .A1(_10991_));
 sg13g2_a21o_1 _17819_ (.A2(_10388_),
    .A1(_09277_),
    .B1(_10849_),
    .X(_11006_));
 sg13g2_nor2_1 _17820_ (.A(net1029),
    .B(\cpu.dec.imm[6] ),
    .Y(_11007_));
 sg13g2_a22oi_1 _17821_ (.Y(_11008_),
    .B1(net779),
    .B2(_11007_),
    .A2(net1030),
    .A1(_08768_));
 sg13g2_o21ai_1 _17822_ (.B1(_11008_),
    .Y(_11009_),
    .A1(_11005_),
    .A2(_11006_));
 sg13g2_buf_1 _17823_ (.A(_11009_),
    .X(_11010_));
 sg13g2_buf_1 _17824_ (.A(_11010_),
    .X(_11011_));
 sg13g2_inv_1 _17825_ (.Y(_11012_),
    .A(_10997_));
 sg13g2_buf_1 _17826_ (.A(_00304_),
    .X(_11013_));
 sg13g2_a21oi_1 _17827_ (.A1(_11012_),
    .A2(_11013_),
    .Y(_11014_),
    .B1(_09463_));
 sg13g2_nor2_1 _17828_ (.A(net234),
    .B(_11014_),
    .Y(_11015_));
 sg13g2_a22oi_1 _17829_ (.Y(_11016_),
    .B1(_10447_),
    .B2(\cpu.ex.r_9[7] ),
    .A2(_10596_),
    .A1(\cpu.ex.r_mult[23] ));
 sg13g2_a221oi_1 _17830_ (.B2(\cpu.ex.r_8[7] ),
    .C1(net677),
    .B1(_10447_),
    .A1(\cpu.ex.r_stmp[7] ),
    .Y(_11017_),
    .A2(_10596_));
 sg13g2_a21o_1 _17831_ (.A2(_11016_),
    .A1(_10444_),
    .B1(_11017_),
    .X(_11018_));
 sg13g2_a22oi_1 _17832_ (.Y(_11019_),
    .B1(_10625_),
    .B2(\cpu.ex.r_11[7] ),
    .A2(net910),
    .A1(\cpu.ex.r_lr[7] ));
 sg13g2_or2_1 _17833_ (.X(_11020_),
    .B(_11019_),
    .A(_10882_));
 sg13g2_buf_1 _17834_ (.A(\cpu.ex.r_sp[7] ),
    .X(_11021_));
 sg13g2_mux2_1 _17835_ (.A0(_11021_),
    .A1(\cpu.ex.r_epc[7] ),
    .S(net677),
    .X(_11022_));
 sg13g2_and2_1 _17836_ (.A(_10491_),
    .B(_10598_),
    .X(_11023_));
 sg13g2_and3_1 _17837_ (.X(_11024_),
    .A(\cpu.ex.r_13[7] ),
    .B(_10428_),
    .C(net781));
 sg13g2_a221oi_1 _17838_ (.B2(_11023_),
    .C1(_11024_),
    .B1(_11022_),
    .A1(\cpu.ex.r_10[7] ),
    .Y(_11025_),
    .A2(_10441_));
 sg13g2_inv_1 _17839_ (.Y(_11026_),
    .A(_00265_));
 sg13g2_a22oi_1 _17840_ (.Y(_11027_),
    .B1(_10494_),
    .B2(_11026_),
    .A2(_10394_),
    .A1(\cpu.ex.r_12[7] ));
 sg13g2_nor2_1 _17841_ (.A(_10548_),
    .B(_11027_),
    .Y(_11028_));
 sg13g2_buf_1 _17842_ (.A(\cpu.dec.user_io ),
    .X(_11029_));
 sg13g2_a22oi_1 _17843_ (.Y(_11030_),
    .B1(_10625_),
    .B2(\cpu.ex.r_14[7] ),
    .A2(net910),
    .A1(_11029_));
 sg13g2_nor2_1 _17844_ (.A(_10444_),
    .B(_11030_),
    .Y(_11031_));
 sg13g2_o21ai_1 _17845_ (.B1(_10420_),
    .Y(_11032_),
    .A1(_11028_),
    .A2(_11031_));
 sg13g2_nand4_1 _17846_ (.B(_11020_),
    .C(_11025_),
    .A(_11018_),
    .Y(_11033_),
    .D(_11032_));
 sg13g2_a221oi_1 _17847_ (.B2(_11033_),
    .C1(_10849_),
    .B1(_10399_),
    .A1(_09280_),
    .Y(_11034_),
    .A2(_10388_));
 sg13g2_or3_1 _17848_ (.A(net1029),
    .B(\cpu.dec.imm[7] ),
    .C(_10535_),
    .X(_11035_));
 sg13g2_o21ai_1 _17849_ (.B1(_11035_),
    .Y(_11036_),
    .A1(_08777_),
    .A2(net906));
 sg13g2_or2_1 _17850_ (.X(_11037_),
    .B(_11036_),
    .A(_11034_));
 sg13g2_buf_1 _17851_ (.A(_11037_),
    .X(_11038_));
 sg13g2_nand2b_1 _17852_ (.Y(_11039_),
    .B(net276),
    .A_N(_11015_));
 sg13g2_nor2_2 _17853_ (.A(_11012_),
    .B(_09463_),
    .Y(_11040_));
 sg13g2_nor2_1 _17854_ (.A(_11013_),
    .B(_09463_),
    .Y(_11041_));
 sg13g2_or2_1 _17855_ (.X(_11042_),
    .B(_11041_),
    .A(net234));
 sg13g2_nand2_1 _17856_ (.Y(_11043_),
    .A(_11040_),
    .B(_11042_));
 sg13g2_nand2_1 _17857_ (.Y(_11044_),
    .A(_11039_),
    .B(_11043_));
 sg13g2_nor2b_1 _17858_ (.A(_10985_),
    .B_N(_11044_),
    .Y(_11045_));
 sg13g2_inv_1 _17859_ (.Y(_11046_),
    .A(\cpu.ex.c_mult_off[3] ));
 sg13g2_nand2_1 _17860_ (.Y(_11047_),
    .A(_09454_),
    .B(_09467_));
 sg13g2_buf_1 _17861_ (.A(\cpu.dec.r_rs1[2] ),
    .X(_11048_));
 sg13g2_buf_8 _17862_ (.A(_11048_),
    .X(_11049_));
 sg13g2_buf_8 _17863_ (.A(_11049_),
    .X(_11050_));
 sg13g2_inv_2 _17864_ (.Y(_11051_),
    .A(net905));
 sg13g2_buf_1 _17865_ (.A(_11051_),
    .X(_11052_));
 sg13g2_buf_2 _17866_ (.A(\cpu.dec.r_rs1[0] ),
    .X(_11053_));
 sg13g2_buf_8 _17867_ (.A(_11053_),
    .X(_11054_));
 sg13g2_buf_1 _17868_ (.A(net1020),
    .X(_11055_));
 sg13g2_buf_8 _17869_ (.A(\cpu.dec.r_rs1[3] ),
    .X(_11056_));
 sg13g2_buf_8 _17870_ (.A(_11056_),
    .X(_11057_));
 sg13g2_buf_8 _17871_ (.A(net1019),
    .X(_11058_));
 sg13g2_buf_8 _17872_ (.A(net903),
    .X(_11059_));
 sg13g2_nor2b_1 _17873_ (.A(_11055_),
    .B_N(net773),
    .Y(_11060_));
 sg13g2_buf_2 _17874_ (.A(_11060_),
    .X(_11061_));
 sg13g2_nand3_1 _17875_ (.B(\cpu.ex.r_8[14] ),
    .C(_11061_),
    .A(net673),
    .Y(_11062_));
 sg13g2_buf_1 _17876_ (.A(net904),
    .X(_11063_));
 sg13g2_nor2b_1 _17877_ (.A(_11056_),
    .B_N(net1021),
    .Y(_11064_));
 sg13g2_buf_8 _17878_ (.A(_11064_),
    .X(_11065_));
 sg13g2_nand3_1 _17879_ (.B(_10584_),
    .C(_11065_),
    .A(net772),
    .Y(_11066_));
 sg13g2_buf_8 _17880_ (.A(\cpu.dec.r_rs1[1] ),
    .X(_11067_));
 sg13g2_buf_1 _17881_ (.A(_11067_),
    .X(_11068_));
 sg13g2_buf_1 _17882_ (.A(_11068_),
    .X(_11069_));
 sg13g2_a21oi_1 _17883_ (.A1(_11062_),
    .A2(_11066_),
    .Y(_11070_),
    .B1(net902));
 sg13g2_and2_1 _17884_ (.A(_11053_),
    .B(_11067_),
    .X(_11071_));
 sg13g2_buf_2 _17885_ (.A(_11071_),
    .X(_11072_));
 sg13g2_buf_1 _17886_ (.A(_11072_),
    .X(_11073_));
 sg13g2_nor2b_1 _17887_ (.A(net1021),
    .B_N(_11056_),
    .Y(_11074_));
 sg13g2_buf_2 _17888_ (.A(_11074_),
    .X(_11075_));
 sg13g2_nand3_1 _17889_ (.B(net771),
    .C(_11075_),
    .A(\cpu.ex.r_11[14] ),
    .Y(_11076_));
 sg13g2_buf_1 _17890_ (.A(net905),
    .X(_11077_));
 sg13g2_buf_1 _17891_ (.A(net770),
    .X(_11078_));
 sg13g2_nor2b_1 _17892_ (.A(_11057_),
    .B_N(_11067_),
    .Y(_11079_));
 sg13g2_buf_1 _17893_ (.A(_11079_),
    .X(_11080_));
 sg13g2_mux2_1 _17894_ (.A0(\cpu.ex.r_stmp[14] ),
    .A1(\cpu.ex.r_mult[30] ),
    .S(net904),
    .X(_11081_));
 sg13g2_nand3_1 _17895_ (.B(net769),
    .C(_11081_),
    .A(net672),
    .Y(_11082_));
 sg13g2_nor2_1 _17896_ (.A(net1019),
    .B(net1021),
    .Y(_11083_));
 sg13g2_buf_2 _17897_ (.A(_11083_),
    .X(_11084_));
 sg13g2_buf_1 _17898_ (.A(_11084_),
    .X(_11085_));
 sg13g2_nor2b_1 _17899_ (.A(_11067_),
    .B_N(_11053_),
    .Y(_11086_));
 sg13g2_buf_1 _17900_ (.A(_11086_),
    .X(_11087_));
 sg13g2_nand3_1 _17901_ (.B(net671),
    .C(net901),
    .A(\cpu.ex.r_lr[14] ),
    .Y(_11088_));
 sg13g2_nand3_1 _17902_ (.B(_11082_),
    .C(_11088_),
    .A(_11076_),
    .Y(_11089_));
 sg13g2_nor2_1 _17903_ (.A(_11053_),
    .B(_11067_),
    .Y(_11090_));
 sg13g2_buf_2 _17904_ (.A(_11090_),
    .X(_11091_));
 sg13g2_buf_1 _17905_ (.A(_11091_),
    .X(_11092_));
 sg13g2_and2_1 _17906_ (.A(net1019),
    .B(net1021),
    .X(_11093_));
 sg13g2_buf_1 _17907_ (.A(_11093_),
    .X(_11094_));
 sg13g2_nand3_1 _17908_ (.B(net768),
    .C(net767),
    .A(\cpu.ex.r_12[14] ),
    .Y(_11095_));
 sg13g2_nand3_1 _17909_ (.B(net671),
    .C(net771),
    .A(\cpu.ex.r_epc[14] ),
    .Y(_11096_));
 sg13g2_nand3_1 _17910_ (.B(net767),
    .C(net901),
    .A(\cpu.ex.r_13[14] ),
    .Y(_11097_));
 sg13g2_buf_8 _17911_ (.A(_11067_),
    .X(_11098_));
 sg13g2_nand4_1 _17912_ (.B(net1017),
    .C(net1019),
    .A(net1020),
    .Y(_11099_),
    .D(net1021));
 sg13g2_buf_1 _17913_ (.A(_11099_),
    .X(_11100_));
 sg13g2_nand2b_1 _17914_ (.Y(_11101_),
    .B(_10607_),
    .A_N(net766));
 sg13g2_nand4_1 _17915_ (.B(_11096_),
    .C(_11097_),
    .A(_11095_),
    .Y(_11102_),
    .D(_11101_));
 sg13g2_nand2b_1 _17916_ (.Y(_11103_),
    .B(net1017),
    .A_N(_11053_));
 sg13g2_buf_1 _17917_ (.A(_11103_),
    .X(_11104_));
 sg13g2_a22oi_1 _17918_ (.Y(_11105_),
    .B1(net767),
    .B2(\cpu.ex.r_14[14] ),
    .A2(net671),
    .A1(_10599_));
 sg13g2_nand3b_1 _17919_ (.B(net902),
    .C(\cpu.ex.r_10[14] ),
    .Y(_11106_),
    .A_N(net904));
 sg13g2_nand3b_1 _17920_ (.B(\cpu.ex.r_9[14] ),
    .C(net772),
    .Y(_11107_),
    .A_N(net902));
 sg13g2_nand2b_1 _17921_ (.Y(_11108_),
    .B(net1019),
    .A_N(net1021));
 sg13g2_buf_2 _17922_ (.A(_11108_),
    .X(_11109_));
 sg13g2_a21o_1 _17923_ (.A2(_11107_),
    .A1(_11106_),
    .B1(_11109_),
    .X(_11110_));
 sg13g2_o21ai_1 _17924_ (.B1(_11110_),
    .Y(_11111_),
    .A1(net765),
    .A2(_11105_));
 sg13g2_nor4_1 _17925_ (.A(_11070_),
    .B(_11089_),
    .C(_11102_),
    .D(_11111_),
    .Y(_11112_));
 sg13g2_xor2_1 _17926_ (.B(_11049_),
    .A(net1111),
    .X(_11113_));
 sg13g2_xor2_1 _17927_ (.B(_11098_),
    .A(net1114),
    .X(_11114_));
 sg13g2_xor2_1 _17928_ (.B(net1019),
    .A(net1112),
    .X(_11115_));
 sg13g2_xor2_1 _17929_ (.B(net1020),
    .A(net1113),
    .X(_11116_));
 sg13g2_nor4_1 _17930_ (.A(_11113_),
    .B(_11114_),
    .C(_11115_),
    .D(_11116_),
    .Y(_11117_));
 sg13g2_nand3_1 _17931_ (.B(_10376_),
    .C(_11117_),
    .A(net1115),
    .Y(_11118_));
 sg13g2_buf_2 _17932_ (.A(_11118_),
    .X(_11119_));
 sg13g2_buf_8 _17933_ (.A(_11119_),
    .X(_11120_));
 sg13g2_mux2_1 _17934_ (.A0(_08512_),
    .A1(_11112_),
    .S(net535),
    .X(_11121_));
 sg13g2_nand2b_1 _17935_ (.Y(_11122_),
    .B(_11121_),
    .A_N(_11047_));
 sg13g2_nand3_1 _17936_ (.B(_09467_),
    .C(_00195_),
    .A(_09454_),
    .Y(_11123_));
 sg13g2_nand4_1 _17937_ (.B(_09295_),
    .C(_09300_),
    .A(_09291_),
    .Y(_11124_),
    .D(_09305_));
 sg13g2_nand2_1 _17938_ (.Y(_11125_),
    .A(_09311_),
    .B(_09316_));
 sg13g2_buf_1 _17939_ (.A(_00273_),
    .X(_11126_));
 sg13g2_nor4_1 _17940_ (.A(_11053_),
    .B(_11067_),
    .C(_11056_),
    .D(_11048_),
    .Y(_11127_));
 sg13g2_or3_1 _17941_ (.A(_09284_),
    .B(_11126_),
    .C(_11127_),
    .X(_11128_));
 sg13g2_nor4_2 _17942_ (.A(_11124_),
    .B(_11125_),
    .C(_09332_),
    .Y(_11129_),
    .D(_11128_));
 sg13g2_nor4_1 _17943_ (.A(_09284_),
    .B(_09318_),
    .C(_11126_),
    .D(_11127_),
    .Y(_11130_));
 sg13g2_nor2b_1 _17944_ (.A(_09332_),
    .B_N(_11130_),
    .Y(_11131_));
 sg13g2_nor4_1 _17945_ (.A(_09284_),
    .B(_09285_),
    .C(_11126_),
    .D(_11127_),
    .Y(_11132_));
 sg13g2_or3_1 _17946_ (.A(_11129_),
    .B(_11131_),
    .C(_11132_),
    .X(_11133_));
 sg13g2_and3_1 _17947_ (.X(_11134_),
    .A(_08427_),
    .B(_08429_),
    .C(_11133_));
 sg13g2_buf_8 _17948_ (.A(_11134_),
    .X(_11135_));
 sg13g2_buf_1 _17949_ (.A(\cpu.br ),
    .X(_11136_));
 sg13g2_inv_2 _17950_ (.Y(_11137_),
    .A(_11136_));
 sg13g2_a21o_1 _17951_ (.A2(_11133_),
    .A1(_08434_),
    .B1(_11137_),
    .X(_11138_));
 sg13g2_buf_1 _17952_ (.A(_11138_),
    .X(_11139_));
 sg13g2_a21oi_1 _17953_ (.A1(net505),
    .A2(_11135_),
    .Y(_11140_),
    .B1(_11139_));
 sg13g2_buf_2 _17954_ (.A(_11140_),
    .X(_11141_));
 sg13g2_mux2_1 _17955_ (.A0(_11122_),
    .A1(_11123_),
    .S(_11141_),
    .X(_11142_));
 sg13g2_nand2_1 _17956_ (.Y(_11143_),
    .A(net628),
    .B(_10468_));
 sg13g2_nor2_1 _17957_ (.A(_11143_),
    .B(_09469_),
    .Y(_11144_));
 sg13g2_and2_1 _17958_ (.A(_09468_),
    .B(_11144_),
    .X(_11145_));
 sg13g2_inv_1 _17959_ (.Y(_11146_),
    .A(_00194_));
 sg13g2_buf_1 _17960_ (.A(net794),
    .X(_11147_));
 sg13g2_and3_1 _17961_ (.X(_11148_),
    .A(net1115),
    .B(_10376_),
    .C(_11117_));
 sg13g2_buf_1 _17962_ (.A(_11148_),
    .X(_11149_));
 sg13g2_buf_1 _17963_ (.A(net612),
    .X(_11150_));
 sg13g2_inv_1 _17964_ (.Y(_11151_),
    .A(net1020));
 sg13g2_buf_1 _17965_ (.A(_11151_),
    .X(_11152_));
 sg13g2_nor2_1 _17966_ (.A(net1018),
    .B(net903),
    .Y(_11153_));
 sg13g2_buf_2 _17967_ (.A(_11153_),
    .X(_11154_));
 sg13g2_and2_1 _17968_ (.A(net1017),
    .B(_11057_),
    .X(_11155_));
 sg13g2_buf_2 _17969_ (.A(_11155_),
    .X(_11156_));
 sg13g2_a22oi_1 _17970_ (.Y(_11157_),
    .B1(_11156_),
    .B2(\cpu.ex.r_15[15] ),
    .A2(_11154_),
    .A1(_10415_));
 sg13g2_nor3_1 _17971_ (.A(net764),
    .B(net673),
    .C(_11157_),
    .Y(_11158_));
 sg13g2_nand2_1 _17972_ (.Y(_11159_),
    .A(net903),
    .B(net905));
 sg13g2_nand2b_1 _17973_ (.Y(_11160_),
    .B(_11053_),
    .A_N(_11067_));
 sg13g2_buf_2 _17974_ (.A(_11160_),
    .X(_11161_));
 sg13g2_nor2_1 _17975_ (.A(_11159_),
    .B(_11161_),
    .Y(_11162_));
 sg13g2_buf_2 _17976_ (.A(_11162_),
    .X(_11163_));
 sg13g2_nor2_2 _17977_ (.A(_11109_),
    .B(_11161_),
    .Y(_11164_));
 sg13g2_a22oi_1 _17978_ (.Y(_11165_),
    .B1(_11164_),
    .B2(\cpu.ex.r_9[15] ),
    .A2(_11163_),
    .A1(\cpu.ex.r_13[15] ));
 sg13g2_and2_1 _17979_ (.A(_11091_),
    .B(net767),
    .X(_11166_));
 sg13g2_buf_1 _17980_ (.A(_11166_),
    .X(_11167_));
 sg13g2_and2_1 _17981_ (.A(_11065_),
    .B(_11072_),
    .X(_11168_));
 sg13g2_buf_8 _17982_ (.A(_11168_),
    .X(_11169_));
 sg13g2_a22oi_1 _17983_ (.Y(_11170_),
    .B1(_11169_),
    .B2(\cpu.ex.r_mult[31] ),
    .A2(_11167_),
    .A1(\cpu.ex.r_12[15] ));
 sg13g2_nand2_1 _17984_ (.Y(_11171_),
    .A(_11165_),
    .B(_11170_));
 sg13g2_nor2b_1 _17985_ (.A(net1020),
    .B_N(net1017),
    .Y(_11172_));
 sg13g2_buf_2 _17986_ (.A(_11172_),
    .X(_11173_));
 sg13g2_buf_8 _17987_ (.A(net773),
    .X(_11174_));
 sg13g2_mux4_1 _17988_ (.S0(net770),
    .A0(_10449_),
    .A1(\cpu.ex.r_stmp[15] ),
    .A2(\cpu.ex.r_10[15] ),
    .A3(\cpu.ex.r_14[15] ),
    .S1(net669),
    .X(_11175_));
 sg13g2_nand2_1 _17989_ (.Y(_11176_),
    .A(_11173_),
    .B(_11175_));
 sg13g2_nand2_1 _17990_ (.Y(_11177_),
    .A(_11054_),
    .B(net1017));
 sg13g2_nor2_1 _17991_ (.A(_11177_),
    .B(_11109_),
    .Y(_11178_));
 sg13g2_buf_2 _17992_ (.A(_11178_),
    .X(_11179_));
 sg13g2_and2_1 _17993_ (.A(_11091_),
    .B(_11075_),
    .X(_11180_));
 sg13g2_buf_2 _17994_ (.A(_11180_),
    .X(_11181_));
 sg13g2_a22oi_1 _17995_ (.Y(_11182_),
    .B1(_11181_),
    .B2(\cpu.ex.r_8[15] ),
    .A2(_11179_),
    .A1(\cpu.ex.r_11[15] ));
 sg13g2_and2_1 _17996_ (.A(_11084_),
    .B(net901),
    .X(_11183_));
 sg13g2_buf_1 _17997_ (.A(_11183_),
    .X(_11184_));
 sg13g2_nand2_1 _17998_ (.Y(_11185_),
    .A(\cpu.ex.r_lr[15] ),
    .B(_11184_));
 sg13g2_nand3_1 _17999_ (.B(net671),
    .C(net771),
    .A(\cpu.ex.r_epc[15] ),
    .Y(_11186_));
 sg13g2_nand4_1 _18000_ (.B(_11182_),
    .C(_11185_),
    .A(_11176_),
    .Y(_11187_),
    .D(_11186_));
 sg13g2_nor4_1 _18001_ (.A(net534),
    .B(_11158_),
    .C(_11171_),
    .D(_11187_),
    .Y(_11188_));
 sg13g2_a21oi_1 _18002_ (.A1(_11147_),
    .A2(net534),
    .Y(_11189_),
    .B1(_11188_));
 sg13g2_a21o_1 _18003_ (.A2(_11135_),
    .A1(net505),
    .B1(_11139_),
    .X(_11190_));
 sg13g2_buf_8 _18004_ (.A(_11190_),
    .X(_11191_));
 sg13g2_buf_8 _18005_ (.A(_11191_),
    .X(_11192_));
 sg13g2_mux2_1 _18006_ (.A0(_11146_),
    .A1(_11189_),
    .S(net347),
    .X(_11193_));
 sg13g2_buf_8 _18007_ (.A(_11193_),
    .X(_11194_));
 sg13g2_nand2_1 _18008_ (.Y(_11195_),
    .A(net495),
    .B(_09470_));
 sg13g2_a22oi_1 _18009_ (.Y(_11196_),
    .B1(_11194_),
    .B2(_11195_),
    .A2(_11145_),
    .A1(_11142_));
 sg13g2_nor2b_1 _18010_ (.A(_09454_),
    .B_N(_09467_),
    .Y(_11197_));
 sg13g2_buf_1 _18011_ (.A(_11197_),
    .X(_11198_));
 sg13g2_inv_1 _18012_ (.Y(_11199_),
    .A(net903));
 sg13g2_buf_1 _18013_ (.A(_11199_),
    .X(_11200_));
 sg13g2_nand4_1 _18014_ (.B(_11052_),
    .C(\cpu.ex.r_epc[13] ),
    .A(net668),
    .Y(_11201_),
    .D(_11073_));
 sg13g2_nor2b_1 _18015_ (.A(_00271_),
    .B_N(net770),
    .Y(_11202_));
 sg13g2_nor2b_1 _18016_ (.A(net770),
    .B_N(\cpu.ex.r_8[13] ),
    .Y(_11203_));
 sg13g2_a22oi_1 _18017_ (.Y(_11204_),
    .B1(_11203_),
    .B2(net768),
    .A2(_11202_),
    .A1(_11072_));
 sg13g2_nand3_1 _18018_ (.B(\cpu.ex.r_12[13] ),
    .C(net768),
    .A(net672),
    .Y(_11205_));
 sg13g2_a21o_1 _18019_ (.A2(_11205_),
    .A1(_11204_),
    .B1(net668),
    .X(_11206_));
 sg13g2_and2_1 _18020_ (.A(_11053_),
    .B(net1019),
    .X(_11207_));
 sg13g2_buf_1 _18021_ (.A(_11207_),
    .X(_11208_));
 sg13g2_nor2_2 _18022_ (.A(net1020),
    .B(net903),
    .Y(_11209_));
 sg13g2_a22oi_1 _18023_ (.Y(_11210_),
    .B1(_11209_),
    .B2(_10545_),
    .A2(_11208_),
    .A1(\cpu.ex.r_11[13] ));
 sg13g2_nor2b_1 _18024_ (.A(net1021),
    .B_N(net1017),
    .Y(_11211_));
 sg13g2_buf_2 _18025_ (.A(_11211_),
    .X(_11212_));
 sg13g2_nand2b_1 _18026_ (.Y(_11213_),
    .B(_11212_),
    .A_N(_11210_));
 sg13g2_nand3_1 _18027_ (.B(_11206_),
    .C(_11213_),
    .A(_11201_),
    .Y(_11214_));
 sg13g2_buf_1 _18028_ (.A(_11050_),
    .X(_11215_));
 sg13g2_and2_1 _18029_ (.A(net763),
    .B(net769),
    .X(_11216_));
 sg13g2_buf_1 _18030_ (.A(_11216_),
    .X(_11217_));
 sg13g2_nor2b_1 _18031_ (.A(_11098_),
    .B_N(net1019),
    .Y(_11218_));
 sg13g2_buf_2 _18032_ (.A(_11218_),
    .X(_11219_));
 sg13g2_and2_1 _18033_ (.A(net673),
    .B(_11219_),
    .X(_11220_));
 sg13g2_a22oi_1 _18034_ (.Y(_11221_),
    .B1(_11220_),
    .B2(\cpu.ex.r_9[13] ),
    .A2(_11217_),
    .A1(_10540_));
 sg13g2_buf_1 _18035_ (.A(net669),
    .X(_11222_));
 sg13g2_and3_1 _18036_ (.X(_11223_),
    .A(_11222_),
    .B(\cpu.ex.r_14[13] ),
    .C(_11173_));
 sg13g2_inv_1 _18037_ (.Y(_11224_),
    .A(_10541_));
 sg13g2_nor3_1 _18038_ (.A(net611),
    .B(_11224_),
    .C(_11161_),
    .Y(_11225_));
 sg13g2_o21ai_1 _18039_ (.B1(net672),
    .Y(_11226_),
    .A1(_11223_),
    .A2(_11225_));
 sg13g2_o21ai_1 _18040_ (.B1(_11226_),
    .Y(_11227_),
    .A1(_11152_),
    .A2(_11221_));
 sg13g2_nor2_1 _18041_ (.A(net905),
    .B(_11161_),
    .Y(_11228_));
 sg13g2_buf_2 _18042_ (.A(_11228_),
    .X(_11229_));
 sg13g2_nor2_2 _18043_ (.A(_11051_),
    .B(net765),
    .Y(_11230_));
 sg13g2_a22oi_1 _18044_ (.Y(_11231_),
    .B1(_11230_),
    .B2(\cpu.ex.r_stmp[13] ),
    .A2(_11229_),
    .A1(\cpu.ex.r_lr[13] ));
 sg13g2_nor2_1 _18045_ (.A(net770),
    .B(net765),
    .Y(_11232_));
 sg13g2_nor2_1 _18046_ (.A(net673),
    .B(_11161_),
    .Y(_11233_));
 sg13g2_a221oi_1 _18047_ (.B2(\cpu.ex.r_13[13] ),
    .C1(net668),
    .B1(_11233_),
    .A1(\cpu.ex.r_10[13] ),
    .Y(_11234_),
    .A2(_11232_));
 sg13g2_a21oi_1 _18048_ (.A1(net668),
    .A2(_11231_),
    .Y(_11235_),
    .B1(_11234_));
 sg13g2_nor4_1 _18049_ (.A(net534),
    .B(_11214_),
    .C(_11227_),
    .D(_11235_),
    .Y(_11236_));
 sg13g2_a21o_1 _18050_ (.A2(_11150_),
    .A1(_08404_),
    .B1(_11236_),
    .X(_11237_));
 sg13g2_nand2b_1 _18051_ (.Y(_11238_),
    .B(net902),
    .A_N(_00270_));
 sg13g2_nand2b_1 _18052_ (.Y(_11239_),
    .B(\cpu.ex.r_13[12] ),
    .A_N(net902));
 sg13g2_nand3_1 _18053_ (.B(net669),
    .C(net770),
    .A(net772),
    .Y(_11240_));
 sg13g2_a21oi_1 _18054_ (.A1(_11238_),
    .A2(_11239_),
    .Y(_11241_),
    .B1(_11240_));
 sg13g2_a21oi_1 _18055_ (.A1(_10480_),
    .A2(_11169_),
    .Y(_11242_),
    .B1(_11241_));
 sg13g2_a22oi_1 _18056_ (.Y(_11243_),
    .B1(net901),
    .B2(_10483_),
    .A2(_11173_),
    .A1(\cpu.ex.r_stmp[12] ));
 sg13g2_nand2b_1 _18057_ (.Y(_11244_),
    .B(_11065_),
    .A_N(_11243_));
 sg13g2_nor2_1 _18058_ (.A(net1017),
    .B(net905),
    .Y(_11245_));
 sg13g2_and2_1 _18059_ (.A(net1017),
    .B(net1021),
    .X(_11246_));
 sg13g2_buf_1 _18060_ (.A(_11246_),
    .X(_11247_));
 sg13g2_a22oi_1 _18061_ (.Y(_11248_),
    .B1(_11247_),
    .B2(\cpu.ex.r_14[12] ),
    .A2(_11245_),
    .A1(\cpu.ex.r_8[12] ));
 sg13g2_nand2b_1 _18062_ (.Y(_11249_),
    .B(_11061_),
    .A_N(_11248_));
 sg13g2_nand3_1 _18063_ (.B(_11244_),
    .C(_11249_),
    .A(_11242_),
    .Y(_11250_));
 sg13g2_a22oi_1 _18064_ (.Y(_11251_),
    .B1(_11219_),
    .B2(\cpu.ex.r_9[12] ),
    .A2(net769),
    .A1(\cpu.ex.r_epc[12] ));
 sg13g2_nand3_1 _18065_ (.B(_10500_),
    .C(_11173_),
    .A(net668),
    .Y(_11252_));
 sg13g2_o21ai_1 _18066_ (.B1(_11252_),
    .Y(_11253_),
    .A1(net764),
    .A2(_11251_));
 sg13g2_and2_1 _18067_ (.A(_11052_),
    .B(_11253_),
    .X(_11254_));
 sg13g2_nor2_1 _18068_ (.A(net668),
    .B(net765),
    .Y(_11255_));
 sg13g2_nor2_1 _18069_ (.A(net611),
    .B(_11161_),
    .Y(_11256_));
 sg13g2_a22oi_1 _18070_ (.Y(_11257_),
    .B1(_11256_),
    .B2(\cpu.ex.r_lr[12] ),
    .A2(_11255_),
    .A1(\cpu.ex.r_10[12] ));
 sg13g2_and3_1 _18071_ (.X(_11258_),
    .A(net672),
    .B(\cpu.ex.r_12[12] ),
    .C(net768));
 sg13g2_and3_1 _18072_ (.X(_11259_),
    .A(net673),
    .B(\cpu.ex.r_11[12] ),
    .C(net771));
 sg13g2_o21ai_1 _18073_ (.B1(net611),
    .Y(_11260_),
    .A1(_11258_),
    .A2(_11259_));
 sg13g2_o21ai_1 _18074_ (.B1(_11260_),
    .Y(_11261_),
    .A1(net672),
    .A2(_11257_));
 sg13g2_or4_1 _18075_ (.A(net534),
    .B(_11250_),
    .C(_11254_),
    .D(_11261_),
    .X(_11262_));
 sg13g2_o21ai_1 _18076_ (.B1(_11262_),
    .Y(_11263_),
    .A1(net687),
    .A2(net535));
 sg13g2_nor2b_1 _18077_ (.A(_09467_),
    .B_N(_09454_),
    .Y(_11264_));
 sg13g2_buf_1 _18078_ (.A(_11264_),
    .X(_11265_));
 sg13g2_a221oi_1 _18079_ (.B2(_11265_),
    .C1(_11141_),
    .B1(_11263_),
    .A1(_11198_),
    .Y(_11266_),
    .A2(_11237_));
 sg13g2_buf_8 _18080_ (.A(net347),
    .X(_11267_));
 sg13g2_a221oi_1 _18081_ (.B2(_00289_),
    .C1(net275),
    .B1(_11265_),
    .A1(_00196_),
    .Y(_11268_),
    .A2(_11198_));
 sg13g2_nor3_1 _18082_ (.A(_11143_),
    .B(_11266_),
    .C(_11268_),
    .Y(_11269_));
 sg13g2_or3_1 _18083_ (.A(_11046_),
    .B(_11196_),
    .C(_11269_),
    .X(_11270_));
 sg13g2_buf_1 _18084_ (.A(_11270_),
    .X(_11271_));
 sg13g2_and2_1 _18085_ (.A(_09468_),
    .B(_09469_),
    .X(_11272_));
 sg13g2_inv_1 _18086_ (.Y(_11273_),
    .A(_00290_));
 sg13g2_inv_1 _18087_ (.Y(_11274_),
    .A(_10680_));
 sg13g2_mux2_1 _18088_ (.A0(\cpu.ex.r_10[11] ),
    .A1(\cpu.ex.r_14[11] ),
    .S(_11077_),
    .X(_11275_));
 sg13g2_nor2_1 _18089_ (.A(_00269_),
    .B(net766),
    .Y(_11276_));
 sg13g2_a221oi_1 _18090_ (.B2(_11275_),
    .C1(_11276_),
    .B1(_11255_),
    .A1(\cpu.ex.r_11[11] ),
    .Y(_11277_),
    .A2(_11179_));
 sg13g2_a22oi_1 _18091_ (.Y(_11278_),
    .B1(_11169_),
    .B2(\cpu.ex.r_mult[27] ),
    .A2(_11167_),
    .A1(\cpu.ex.r_12[11] ));
 sg13g2_a22oi_1 _18092_ (.Y(_11279_),
    .B1(_11181_),
    .B2(\cpu.ex.r_8[11] ),
    .A2(_11164_),
    .A1(\cpu.ex.r_9[11] ));
 sg13g2_nand3_1 _18093_ (.B(_11278_),
    .C(_11279_),
    .A(_11277_),
    .Y(_11280_));
 sg13g2_nand2_1 _18094_ (.Y(_11281_),
    .A(net671),
    .B(net771));
 sg13g2_nand2_1 _18095_ (.Y(_11282_),
    .A(\cpu.ex.r_13[11] ),
    .B(_11163_));
 sg13g2_o21ai_1 _18096_ (.B1(_11282_),
    .Y(_11283_),
    .A1(_10658_),
    .A2(_11281_));
 sg13g2_mux2_1 _18097_ (.A0(_10664_),
    .A1(\cpu.ex.r_stmp[11] ),
    .S(net672),
    .X(_11284_));
 sg13g2_a22oi_1 _18098_ (.Y(_11285_),
    .B1(_11284_),
    .B2(_11173_),
    .A2(_11229_),
    .A1(\cpu.ex.r_lr[11] ));
 sg13g2_nor2_1 _18099_ (.A(net611),
    .B(_11285_),
    .Y(_11286_));
 sg13g2_nor4_1 _18100_ (.A(net534),
    .B(_11280_),
    .C(_11283_),
    .D(_11286_),
    .Y(_11287_));
 sg13g2_a21oi_1 _18101_ (.A1(_11274_),
    .A2(net534),
    .Y(_11288_),
    .B1(_11287_));
 sg13g2_mux2_1 _18102_ (.A0(_11273_),
    .A1(_11288_),
    .S(net347),
    .X(_11289_));
 sg13g2_buf_8 _18103_ (.A(_11289_),
    .X(_11290_));
 sg13g2_nand2_1 _18104_ (.Y(_11291_),
    .A(_11272_),
    .B(_11290_));
 sg13g2_inv_1 _18105_ (.Y(_11292_),
    .A(_00291_));
 sg13g2_nor2b_1 _18106_ (.A(net1018),
    .B_N(net763),
    .Y(_11293_));
 sg13g2_a22oi_1 _18107_ (.Y(_11294_),
    .B1(_11293_),
    .B2(\cpu.ex.r_12[10] ),
    .A2(_11212_),
    .A1(\cpu.ex.r_10[10] ));
 sg13g2_nor2b_1 _18108_ (.A(_11294_),
    .B_N(_11061_),
    .Y(_11295_));
 sg13g2_nand3_1 _18109_ (.B(net671),
    .C(net771),
    .A(\cpu.ex.r_epc[10] ),
    .Y(_11296_));
 sg13g2_nand3_1 _18110_ (.B(net671),
    .C(net901),
    .A(\cpu.ex.r_lr[10] ),
    .Y(_11297_));
 sg13g2_nand3_1 _18111_ (.B(net767),
    .C(net901),
    .A(\cpu.ex.r_13[10] ),
    .Y(_11298_));
 sg13g2_nand2b_1 _18112_ (.Y(_11299_),
    .B(_10636_),
    .A_N(net766));
 sg13g2_nand4_1 _18113_ (.B(_11297_),
    .C(_11298_),
    .A(_11296_),
    .Y(_11300_),
    .D(_11299_));
 sg13g2_a22oi_1 _18114_ (.Y(_11301_),
    .B1(_11065_),
    .B2(\cpu.ex.r_stmp[10] ),
    .A2(net671),
    .A1(_10633_));
 sg13g2_nand2_1 _18115_ (.Y(_11302_),
    .A(\cpu.ex.r_14[10] ),
    .B(net767));
 sg13g2_a21oi_1 _18116_ (.A1(_11301_),
    .A2(_11302_),
    .Y(_11303_),
    .B1(net765));
 sg13g2_nand3_1 _18117_ (.B(_11065_),
    .C(_11073_),
    .A(net1108),
    .Y(_11304_));
 sg13g2_nand3_1 _18118_ (.B(_11075_),
    .C(net901),
    .A(\cpu.ex.r_9[10] ),
    .Y(_11305_));
 sg13g2_nand3_1 _18119_ (.B(_11092_),
    .C(_11075_),
    .A(\cpu.ex.r_8[10] ),
    .Y(_11306_));
 sg13g2_nand3_1 _18120_ (.B(net771),
    .C(_11075_),
    .A(\cpu.ex.r_11[10] ),
    .Y(_11307_));
 sg13g2_nand4_1 _18121_ (.B(_11305_),
    .C(_11306_),
    .A(_11304_),
    .Y(_11308_),
    .D(_11307_));
 sg13g2_nor4_1 _18122_ (.A(_11295_),
    .B(_11300_),
    .C(_11303_),
    .D(_11308_),
    .Y(_11309_));
 sg13g2_nor2_1 _18123_ (.A(net1107),
    .B(net535),
    .Y(_11310_));
 sg13g2_a21oi_1 _18124_ (.A1(net535),
    .A2(_11309_),
    .Y(_11311_),
    .B1(_11310_));
 sg13g2_mux2_1 _18125_ (.A0(_11292_),
    .A1(_11311_),
    .S(net347),
    .X(_11312_));
 sg13g2_buf_8 _18126_ (.A(_11312_),
    .X(_11313_));
 sg13g2_nor2_1 _18127_ (.A(_09468_),
    .B(_09469_),
    .Y(_11314_));
 sg13g2_o21ai_1 _18128_ (.B1(_11314_),
    .Y(_11315_),
    .A1(_11047_),
    .A2(_11313_));
 sg13g2_buf_2 _18129_ (.A(_00292_),
    .X(_11316_));
 sg13g2_buf_1 _18130_ (.A(_00293_),
    .X(_11317_));
 sg13g2_a221oi_1 _18131_ (.B2(_11317_),
    .C1(net275),
    .B1(_11265_),
    .A1(_11316_),
    .Y(_11318_),
    .A2(_11198_));
 sg13g2_a22oi_1 _18132_ (.Y(_11319_),
    .B1(_11163_),
    .B2(\cpu.ex.r_13[8] ),
    .A2(_11179_),
    .A1(\cpu.ex.r_11[8] ));
 sg13g2_o21ai_1 _18133_ (.B1(_11319_),
    .Y(_11320_),
    .A1(_00266_),
    .A2(net766));
 sg13g2_a22oi_1 _18134_ (.Y(_11321_),
    .B1(_11230_),
    .B2(\cpu.ex.r_14[8] ),
    .A2(_11229_),
    .A1(\cpu.ex.r_9[8] ));
 sg13g2_a221oi_1 _18135_ (.B2(\cpu.ex.r_stmp[8] ),
    .C1(net611),
    .B1(_11230_),
    .A1(\cpu.ex.r_lr[8] ),
    .Y(_11322_),
    .A2(_11229_));
 sg13g2_a21oi_1 _18136_ (.A1(net611),
    .A2(_11321_),
    .Y(_11323_),
    .B1(_11322_));
 sg13g2_nand2_1 _18137_ (.Y(_11324_),
    .A(net764),
    .B(net673));
 sg13g2_a22oi_1 _18138_ (.Y(_11325_),
    .B1(_11219_),
    .B2(\cpu.ex.r_8[8] ),
    .A2(net769),
    .A1(_10727_));
 sg13g2_nand2_1 _18139_ (.Y(_11326_),
    .A(net669),
    .B(\cpu.ex.r_10[8] ));
 sg13g2_nand3b_1 _18140_ (.B(\cpu.ex.r_epc[8] ),
    .C(net904),
    .Y(_11327_),
    .A_N(net669));
 sg13g2_o21ai_1 _18141_ (.B1(_11327_),
    .Y(_11328_),
    .A1(net772),
    .A2(_11326_));
 sg13g2_and3_1 _18142_ (.X(_11329_),
    .A(\cpu.ex.r_12[8] ),
    .B(net768),
    .C(net767));
 sg13g2_a221oi_1 _18143_ (.B2(_11328_),
    .C1(_11329_),
    .B1(_11212_),
    .A1(\cpu.ex.r_mult[24] ),
    .Y(_11330_),
    .A2(_11169_));
 sg13g2_o21ai_1 _18144_ (.B1(_11330_),
    .Y(_11331_),
    .A1(_11324_),
    .A2(_11325_));
 sg13g2_or4_1 _18145_ (.A(net534),
    .B(_11320_),
    .C(_11323_),
    .D(_11331_),
    .X(_11332_));
 sg13g2_o21ai_1 _18146_ (.B1(_11332_),
    .Y(_11333_),
    .A1(_09278_),
    .A2(net535));
 sg13g2_inv_1 _18147_ (.Y(_11334_),
    .A(_00267_));
 sg13g2_a22oi_1 _18148_ (.Y(_11335_),
    .B1(net771),
    .B2(_11334_),
    .A2(net768),
    .A1(\cpu.ex.r_12[9] ));
 sg13g2_nor2_1 _18149_ (.A(_11159_),
    .B(_11335_),
    .Y(_11336_));
 sg13g2_a22oi_1 _18150_ (.Y(_11337_),
    .B1(_11075_),
    .B2(\cpu.ex.r_10[9] ),
    .A2(_11065_),
    .A1(\cpu.ex.r_stmp[9] ));
 sg13g2_nor2_1 _18151_ (.A(net765),
    .B(_11337_),
    .Y(_11338_));
 sg13g2_a22oi_1 _18152_ (.Y(_11339_),
    .B1(_11219_),
    .B2(\cpu.ex.r_8[9] ),
    .A2(_11080_),
    .A1(_10706_));
 sg13g2_nor2_1 _18153_ (.A(_11324_),
    .B(_11339_),
    .Y(_11340_));
 sg13g2_nor3_1 _18154_ (.A(_11336_),
    .B(_11338_),
    .C(_11340_),
    .Y(_11341_));
 sg13g2_a22oi_1 _18155_ (.Y(_11342_),
    .B1(_11220_),
    .B2(\cpu.ex.r_9[9] ),
    .A2(_11217_),
    .A1(\cpu.ex.r_mult[25] ));
 sg13g2_nand2b_1 _18156_ (.Y(_11343_),
    .B(net772),
    .A_N(_11342_));
 sg13g2_nand3_1 _18157_ (.B(\cpu.ex.r_14[9] ),
    .C(_11061_),
    .A(net672),
    .Y(_11344_));
 sg13g2_nand3_1 _18158_ (.B(\cpu.ex.r_epc[9] ),
    .C(_11085_),
    .A(net772),
    .Y(_11345_));
 sg13g2_nand2_1 _18159_ (.Y(_11346_),
    .A(_11344_),
    .B(_11345_));
 sg13g2_nand2b_1 _18160_ (.Y(_11347_),
    .B(net1020),
    .A_N(net905));
 sg13g2_a22oi_1 _18161_ (.Y(_11348_),
    .B1(_11156_),
    .B2(\cpu.ex.r_11[9] ),
    .A2(_11154_),
    .A1(\cpu.ex.r_lr[9] ));
 sg13g2_nor2_1 _18162_ (.A(_11347_),
    .B(_11348_),
    .Y(_11349_));
 sg13g2_a221oi_1 _18163_ (.B2(net902),
    .C1(_11349_),
    .B1(_11346_),
    .A1(\cpu.ex.r_13[9] ),
    .Y(_11350_),
    .A2(_11163_));
 sg13g2_nand4_1 _18164_ (.B(_11341_),
    .C(_11343_),
    .A(_11120_),
    .Y(_11351_),
    .D(_11350_));
 sg13g2_o21ai_1 _18165_ (.B1(_11351_),
    .Y(_11352_),
    .A1(_10716_),
    .A2(net535));
 sg13g2_a221oi_1 _18166_ (.B2(_11198_),
    .C1(_11141_),
    .B1(_11352_),
    .A1(_11265_),
    .Y(_11353_),
    .A2(_11333_));
 sg13g2_nor2_1 _18167_ (.A(_11143_),
    .B(_09471_),
    .Y(_11354_));
 sg13g2_o21ai_1 _18168_ (.B1(_11354_),
    .Y(_11355_),
    .A1(_11318_),
    .A2(_11353_));
 sg13g2_a21o_1 _18169_ (.A2(_11315_),
    .A1(_11291_),
    .B1(_11355_),
    .X(_11356_));
 sg13g2_buf_1 _18170_ (.A(_11356_),
    .X(_11357_));
 sg13g2_o21ai_1 _18171_ (.B1(net495),
    .Y(\cpu.ex.c_mult_off[2] ),
    .A1(_11272_),
    .A2(_11314_));
 sg13g2_nor2b_1 _18172_ (.A(\cpu.ex.c_mult_off[3] ),
    .B_N(\cpu.ex.c_mult_off[2] ),
    .Y(_11358_));
 sg13g2_nand2_1 _18173_ (.Y(_11359_),
    .A(_08593_),
    .B(_11136_));
 sg13g2_or3_1 _18174_ (.A(_08434_),
    .B(_08523_),
    .C(_11359_),
    .X(_11360_));
 sg13g2_or2_1 _18175_ (.X(_11361_),
    .B(_11359_),
    .A(_11135_));
 sg13g2_nand3_1 _18176_ (.B(_11084_),
    .C(_11072_),
    .A(\cpu.ex.r_epc[4] ),
    .Y(_11362_));
 sg13g2_nand2_1 _18177_ (.Y(_11363_),
    .A(\cpu.ex.r_8[4] ),
    .B(_11181_));
 sg13g2_mux2_1 _18178_ (.A0(\cpu.ex.r_lr[4] ),
    .A1(\cpu.ex.r_9[4] ),
    .S(net773),
    .X(_11364_));
 sg13g2_mux2_1 _18179_ (.A0(_08397_),
    .A1(\cpu.ex.r_12[4] ),
    .S(net903),
    .X(_11365_));
 sg13g2_and3_1 _18180_ (.X(_11366_),
    .A(_11215_),
    .B(_11091_),
    .C(_11365_));
 sg13g2_a221oi_1 _18181_ (.B2(_11364_),
    .C1(_11366_),
    .B1(_11229_),
    .A1(\cpu.ex.r_mult[20] ),
    .Y(_11367_),
    .A2(_11169_));
 sg13g2_nor2_1 _18182_ (.A(_00262_),
    .B(_11100_),
    .Y(_11368_));
 sg13g2_a21oi_1 _18183_ (.A1(\cpu.ex.r_11[4] ),
    .A2(_11179_),
    .Y(_11369_),
    .B1(_11368_));
 sg13g2_and4_1 _18184_ (.A(_11362_),
    .B(_11363_),
    .C(_11367_),
    .D(_11369_),
    .X(_11370_));
 sg13g2_mux2_1 _18185_ (.A0(_10894_),
    .A1(\cpu.ex.r_stmp[4] ),
    .S(net763),
    .X(_11371_));
 sg13g2_nand2_1 _18186_ (.Y(_11372_),
    .A(net763),
    .B(\cpu.ex.r_14[4] ));
 sg13g2_a21oi_1 _18187_ (.A1(_11174_),
    .A2(_11372_),
    .Y(_11373_),
    .B1(net765));
 sg13g2_o21ai_1 _18188_ (.B1(_11373_),
    .Y(_11374_),
    .A1(_11174_),
    .A2(_11371_));
 sg13g2_and2_1 _18189_ (.A(_11059_),
    .B(\cpu.ex.r_10[4] ),
    .X(_11375_));
 sg13g2_a22oi_1 _18190_ (.Y(_11376_),
    .B1(_11232_),
    .B2(_11375_),
    .A2(_11163_),
    .A1(\cpu.ex.r_13[4] ));
 sg13g2_and3_1 _18191_ (.X(_11377_),
    .A(_11119_),
    .B(_11374_),
    .C(_11376_));
 sg13g2_a22oi_1 _18192_ (.Y(_11378_),
    .B1(_11370_),
    .B2(_11377_),
    .A2(net612),
    .A1(_09491_));
 sg13g2_nand2_1 _18193_ (.Y(_11379_),
    .A(_11139_),
    .B(_11378_));
 sg13g2_nand3_1 _18194_ (.B(_11135_),
    .C(_11378_),
    .A(net505),
    .Y(_11380_));
 sg13g2_nand4_1 _18195_ (.B(_11361_),
    .C(_11379_),
    .A(_11360_),
    .Y(_11381_),
    .D(_11380_));
 sg13g2_buf_1 _18196_ (.A(_11381_),
    .X(_11382_));
 sg13g2_inv_2 _18197_ (.Y(_11383_),
    .A(_10122_));
 sg13g2_a22oi_1 _18198_ (.Y(_11384_),
    .B1(_11209_),
    .B2(_10859_),
    .A2(_11208_),
    .A1(\cpu.ex.r_11[5] ));
 sg13g2_nand2b_1 _18199_ (.Y(_11385_),
    .B(_11212_),
    .A_N(_11384_));
 sg13g2_mux2_1 _18200_ (.A0(\cpu.ex.r_10[5] ),
    .A1(\cpu.ex.r_14[5] ),
    .S(net763),
    .X(_11386_));
 sg13g2_a22oi_1 _18201_ (.Y(_11387_),
    .B1(_11255_),
    .B2(_11386_),
    .A2(_11167_),
    .A1(\cpu.ex.r_12[5] ));
 sg13g2_nor2_1 _18202_ (.A(_00263_),
    .B(net766),
    .Y(_11388_));
 sg13g2_nand3_1 _18203_ (.B(_11084_),
    .C(_11072_),
    .A(\cpu.ex.r_epc[5] ),
    .Y(_11389_));
 sg13g2_nor2b_1 _18204_ (.A(_11388_),
    .B_N(_11389_),
    .Y(_11390_));
 sg13g2_a22oi_1 _18205_ (.Y(_11391_),
    .B1(_11181_),
    .B2(\cpu.ex.r_8[5] ),
    .A2(_11163_),
    .A1(\cpu.ex.r_13[5] ));
 sg13g2_and4_1 _18206_ (.A(_11385_),
    .B(_11387_),
    .C(_11390_),
    .D(_11391_),
    .X(_11392_));
 sg13g2_mux2_1 _18207_ (.A0(\cpu.ex.r_stmp[5] ),
    .A1(\cpu.ex.r_mult[21] ),
    .S(net904),
    .X(_11393_));
 sg13g2_a22oi_1 _18208_ (.Y(_11394_),
    .B1(_11393_),
    .B2(_11217_),
    .A2(_11164_),
    .A1(\cpu.ex.r_9[5] ));
 sg13g2_nand2_1 _18209_ (.Y(_11395_),
    .A(\cpu.ex.r_lr[5] ),
    .B(_11184_));
 sg13g2_and3_1 _18210_ (.X(_11396_),
    .A(_11119_),
    .B(_11394_),
    .C(_11395_));
 sg13g2_a22oi_1 _18211_ (.Y(_11397_),
    .B1(_11392_),
    .B2(_11396_),
    .A2(net612),
    .A1(_11383_));
 sg13g2_buf_1 _18212_ (.A(_11397_),
    .X(_11398_));
 sg13g2_nand2_1 _18213_ (.Y(_11399_),
    .A(_11139_),
    .B(_11398_));
 sg13g2_nand3_1 _18214_ (.B(_11135_),
    .C(_11398_),
    .A(net505),
    .Y(_11400_));
 sg13g2_buf_2 _18215_ (.A(_00296_),
    .X(_11401_));
 sg13g2_nor2_1 _18216_ (.A(_11137_),
    .B(_11401_),
    .Y(_11402_));
 sg13g2_nand2b_1 _18217_ (.Y(_11403_),
    .B(_11402_),
    .A_N(_11135_));
 sg13g2_or4_1 _18218_ (.A(_11137_),
    .B(_11401_),
    .C(_08434_),
    .D(_08523_),
    .X(_11404_));
 sg13g2_nand4_1 _18219_ (.B(_11400_),
    .C(_11403_),
    .A(_11399_),
    .Y(_11405_),
    .D(_11404_));
 sg13g2_buf_2 _18220_ (.A(_11405_),
    .X(_11406_));
 sg13g2_inv_1 _18221_ (.Y(_11407_),
    .A(_00295_));
 sg13g2_nor2_1 _18222_ (.A(_09277_),
    .B(net535),
    .Y(_11408_));
 sg13g2_nand2_1 _18223_ (.Y(_11409_),
    .A(_11151_),
    .B(net763));
 sg13g2_a22oi_1 _18224_ (.Y(_11410_),
    .B1(_11219_),
    .B2(\cpu.ex.r_12[6] ),
    .A2(net769),
    .A1(\cpu.ex.r_stmp[6] ));
 sg13g2_or2_1 _18225_ (.X(_11411_),
    .B(_11410_),
    .A(_11409_));
 sg13g2_and2_1 _18226_ (.A(_11051_),
    .B(_11156_),
    .X(_11412_));
 sg13g2_mux2_1 _18227_ (.A0(\cpu.ex.r_10[6] ),
    .A1(\cpu.ex.r_11[6] ),
    .S(_11055_),
    .X(_11413_));
 sg13g2_a22oi_1 _18228_ (.Y(_11414_),
    .B1(_11412_),
    .B2(_11413_),
    .A2(_11169_),
    .A1(_10997_));
 sg13g2_a22oi_1 _18229_ (.Y(_11415_),
    .B1(_11181_),
    .B2(\cpu.ex.r_8[6] ),
    .A2(_11163_),
    .A1(\cpu.ex.r_13[6] ));
 sg13g2_nor2_1 _18230_ (.A(_00264_),
    .B(net766),
    .Y(_11416_));
 sg13g2_a21oi_1 _18231_ (.A1(\cpu.ex.r_lr[6] ),
    .A2(_11184_),
    .Y(_11417_),
    .B1(_11416_));
 sg13g2_nand4_1 _18232_ (.B(_11414_),
    .C(_11415_),
    .A(_11411_),
    .Y(_11418_),
    .D(_11417_));
 sg13g2_nand3_1 _18233_ (.B(\cpu.ex.r_9[6] ),
    .C(net901),
    .A(net611),
    .Y(_11419_));
 sg13g2_nand3_1 _18234_ (.B(_10992_),
    .C(_11173_),
    .A(net668),
    .Y(_11420_));
 sg13g2_a21oi_1 _18235_ (.A1(_11419_),
    .A2(_11420_),
    .Y(_11421_),
    .B1(_11078_));
 sg13g2_nand3_1 _18236_ (.B(\cpu.ex.r_14[6] ),
    .C(_11061_),
    .A(_11078_),
    .Y(_11422_));
 sg13g2_nand3_1 _18237_ (.B(\cpu.ex.r_epc[6] ),
    .C(_11084_),
    .A(net772),
    .Y(_11423_));
 sg13g2_inv_1 _18238_ (.Y(_11424_),
    .A(net1018));
 sg13g2_a21oi_1 _18239_ (.A1(_11422_),
    .A2(_11423_),
    .Y(_11425_),
    .B1(_11424_));
 sg13g2_or4_1 _18240_ (.A(net612),
    .B(_11418_),
    .C(_11421_),
    .D(_11425_),
    .X(_11426_));
 sg13g2_nor2b_1 _18241_ (.A(_11408_),
    .B_N(_11426_),
    .Y(_11427_));
 sg13g2_mux2_1 _18242_ (.A0(_11407_),
    .A1(_11427_),
    .S(_11191_),
    .X(_11428_));
 sg13g2_buf_8 _18243_ (.A(_11428_),
    .X(_11429_));
 sg13g2_inv_1 _18244_ (.Y(_11430_),
    .A(_00294_));
 sg13g2_nor2_1 _18245_ (.A(_09280_),
    .B(net535),
    .Y(_11431_));
 sg13g2_nor2_1 _18246_ (.A(net764),
    .B(net669),
    .Y(_11432_));
 sg13g2_a22oi_1 _18247_ (.Y(_11433_),
    .B1(_11432_),
    .B2(\cpu.ex.r_mult[23] ),
    .A2(_11061_),
    .A1(\cpu.ex.r_14[7] ));
 sg13g2_nor2b_1 _18248_ (.A(_11433_),
    .B_N(_11247_),
    .Y(_11434_));
 sg13g2_nand2_1 _18249_ (.Y(_11435_),
    .A(net764),
    .B(net611));
 sg13g2_a22oi_1 _18250_ (.Y(_11436_),
    .B1(_11293_),
    .B2(\cpu.ex.r_12[7] ),
    .A2(_11212_),
    .A1(\cpu.ex.r_10[7] ));
 sg13g2_a22oi_1 _18251_ (.Y(_11437_),
    .B1(_11087_),
    .B2(\cpu.ex.r_lr[7] ),
    .A2(_11173_),
    .A1(_11021_));
 sg13g2_nand2b_1 _18252_ (.Y(_11438_),
    .B(_11085_),
    .A_N(_11437_));
 sg13g2_o21ai_1 _18253_ (.B1(_11438_),
    .Y(_11439_),
    .A1(_11435_),
    .A2(_11436_));
 sg13g2_nand3_1 _18254_ (.B(_11029_),
    .C(net768),
    .A(net770),
    .Y(_11440_));
 sg13g2_nand3_1 _18255_ (.B(\cpu.ex.r_epc[7] ),
    .C(_11072_),
    .A(_11051_),
    .Y(_11441_));
 sg13g2_a21o_1 _18256_ (.A2(_11441_),
    .A1(_11440_),
    .B1(net669),
    .X(_11442_));
 sg13g2_and3_1 _18257_ (.X(_11443_),
    .A(net773),
    .B(\cpu.ex.r_13[7] ),
    .C(_11087_));
 sg13g2_inv_1 _18258_ (.Y(_11444_),
    .A(\cpu.ex.r_stmp[7] ));
 sg13g2_nor3_1 _18259_ (.A(net669),
    .B(_11444_),
    .C(_11104_),
    .Y(_11445_));
 sg13g2_o21ai_1 _18260_ (.B1(net672),
    .Y(_11446_),
    .A1(_11443_),
    .A2(_11445_));
 sg13g2_nor2_1 _18261_ (.A(_00265_),
    .B(net766),
    .Y(_11447_));
 sg13g2_a21oi_1 _18262_ (.A1(\cpu.ex.r_11[7] ),
    .A2(_11179_),
    .Y(_11448_),
    .B1(_11447_));
 sg13g2_a22oi_1 _18263_ (.Y(_11449_),
    .B1(_11181_),
    .B2(\cpu.ex.r_8[7] ),
    .A2(_11164_),
    .A1(\cpu.ex.r_9[7] ));
 sg13g2_nand4_1 _18264_ (.B(_11446_),
    .C(_11448_),
    .A(_11442_),
    .Y(_11450_),
    .D(_11449_));
 sg13g2_or4_1 _18265_ (.A(net612),
    .B(_11434_),
    .C(_11439_),
    .D(_11450_),
    .X(_11451_));
 sg13g2_nor2b_1 _18266_ (.A(_11431_),
    .B_N(_11451_),
    .Y(_11452_));
 sg13g2_mux2_1 _18267_ (.A0(_11430_),
    .A1(_11452_),
    .S(_11191_),
    .X(_11453_));
 sg13g2_buf_8 _18268_ (.A(_11453_),
    .X(_11454_));
 sg13g2_o21ai_1 _18269_ (.B1(net495),
    .Y(\cpu.ex.c_mult_off[1] ),
    .A1(_11198_),
    .A2(_11265_));
 sg13g2_mux4_1 _18270_ (.S0(\cpu.ex.c_mult_off[0] ),
    .A0(_11382_),
    .A1(_11406_),
    .A2(_11429_),
    .A3(_11454_),
    .S1(\cpu.ex.c_mult_off[1] ),
    .X(_11455_));
 sg13g2_nor2_1 _18271_ (.A(_11143_),
    .B(_11047_),
    .Y(_11456_));
 sg13g2_nand2_1 _18272_ (.Y(_11457_),
    .A(_09348_),
    .B(net534));
 sg13g2_nand2b_1 _18273_ (.Y(_11458_),
    .B(net905),
    .A_N(net1018));
 sg13g2_a22oi_1 _18274_ (.Y(_11459_),
    .B1(_11209_),
    .B2(net1129),
    .A2(_11208_),
    .A1(\cpu.ex.r_13[2] ));
 sg13g2_nor2_1 _18275_ (.A(_11458_),
    .B(_11459_),
    .Y(_11460_));
 sg13g2_a22oi_1 _18276_ (.Y(_11461_),
    .B1(_11247_),
    .B2(\cpu.ex.r_mult[18] ),
    .A2(_11245_),
    .A1(\cpu.ex.r_lr[2] ));
 sg13g2_nor3_1 _18277_ (.A(_11151_),
    .B(_11059_),
    .C(_11461_),
    .Y(_11462_));
 sg13g2_and3_1 _18278_ (.X(_11463_),
    .A(_10825_),
    .B(_11084_),
    .C(_11173_));
 sg13g2_inv_1 _18279_ (.Y(_11464_),
    .A(_00260_));
 sg13g2_a22oi_1 _18280_ (.Y(_11465_),
    .B1(_11094_),
    .B2(_11464_),
    .A2(_11084_),
    .A1(\cpu.ex.r_epc[2] ));
 sg13g2_nor2_1 _18281_ (.A(_11177_),
    .B(_11465_),
    .Y(_11466_));
 sg13g2_or4_1 _18282_ (.A(_11460_),
    .B(_11462_),
    .C(_11463_),
    .D(_11466_),
    .X(_11467_));
 sg13g2_a22oi_1 _18283_ (.Y(_11468_),
    .B1(_11230_),
    .B2(\cpu.ex.r_14[2] ),
    .A2(_11229_),
    .A1(\cpu.ex.r_9[2] ));
 sg13g2_inv_1 _18284_ (.Y(_11469_),
    .A(_10819_));
 sg13g2_nor4_1 _18285_ (.A(net1018),
    .B(net773),
    .C(_11051_),
    .D(_11469_),
    .Y(_11470_));
 sg13g2_and3_1 _18286_ (.X(_11471_),
    .A(_11051_),
    .B(\cpu.ex.r_11[2] ),
    .C(_11156_));
 sg13g2_o21ai_1 _18287_ (.B1(net904),
    .Y(_11472_),
    .A1(_11470_),
    .A2(_11471_));
 sg13g2_o21ai_1 _18288_ (.B1(_11472_),
    .Y(_11473_),
    .A1(_11200_),
    .A2(_11468_));
 sg13g2_mux2_1 _18289_ (.A0(\cpu.ex.r_8[2] ),
    .A1(\cpu.ex.r_12[2] ),
    .S(_11050_),
    .X(_11474_));
 sg13g2_a22oi_1 _18290_ (.Y(_11475_),
    .B1(_11474_),
    .B2(_11424_),
    .A2(_11212_),
    .A1(\cpu.ex.r_10[2] ));
 sg13g2_nand3_1 _18291_ (.B(\cpu.ex.r_stmp[2] ),
    .C(net769),
    .A(_11215_),
    .Y(_11476_));
 sg13g2_o21ai_1 _18292_ (.B1(_11476_),
    .Y(_11477_),
    .A1(_11200_),
    .A2(_11475_));
 sg13g2_and2_1 _18293_ (.A(net764),
    .B(_11477_),
    .X(_11478_));
 sg13g2_or4_1 _18294_ (.A(_11149_),
    .B(_11467_),
    .C(_11473_),
    .D(_11478_),
    .X(_11479_));
 sg13g2_buf_1 _18295_ (.A(_11479_),
    .X(_11480_));
 sg13g2_nand2_1 _18296_ (.Y(_11481_),
    .A(_11457_),
    .B(_11480_));
 sg13g2_mux2_1 _18297_ (.A0(_10918_),
    .A1(\cpu.ex.r_stmp[3] ),
    .S(net905),
    .X(_11482_));
 sg13g2_a22oi_1 _18298_ (.Y(_11483_),
    .B1(_11482_),
    .B2(net668),
    .A2(net767),
    .A1(\cpu.ex.r_14[3] ));
 sg13g2_nor2_1 _18299_ (.A(net765),
    .B(_11483_),
    .Y(_11484_));
 sg13g2_nand3b_1 _18300_ (.B(_11058_),
    .C(\cpu.ex.r_9[3] ),
    .Y(_11485_),
    .A_N(net1018));
 sg13g2_nand3b_1 _18301_ (.B(\cpu.ex.r_epc[3] ),
    .C(net1018),
    .Y(_11486_),
    .A_N(net903));
 sg13g2_a21oi_1 _18302_ (.A1(_11485_),
    .A2(_11486_),
    .Y(_11487_),
    .B1(_11347_));
 sg13g2_nand3b_1 _18303_ (.B(_11058_),
    .C(\cpu.ex.r_12[3] ),
    .Y(_11488_),
    .A_N(_11054_));
 sg13g2_nand3b_1 _18304_ (.B(_10930_),
    .C(net1020),
    .Y(_11489_),
    .A_N(net903));
 sg13g2_a21oi_1 _18305_ (.A1(_11488_),
    .A2(_11489_),
    .Y(_11490_),
    .B1(_11458_));
 sg13g2_and3_1 _18306_ (.X(_11491_),
    .A(\cpu.ex.r_8[3] ),
    .B(_11091_),
    .C(_11075_));
 sg13g2_nor2_1 _18307_ (.A(_00261_),
    .B(net766),
    .Y(_11492_));
 sg13g2_or4_1 _18308_ (.A(_11487_),
    .B(_11490_),
    .C(_11491_),
    .D(_11492_),
    .X(_11493_));
 sg13g2_a221oi_1 _18309_ (.B2(\cpu.ex.r_11[3] ),
    .C1(net770),
    .B1(_11156_),
    .A1(\cpu.ex.r_lr[3] ),
    .Y(_11494_),
    .A2(_11154_));
 sg13g2_a221oi_1 _18310_ (.B2(\cpu.ex.r_13[3] ),
    .C1(_11051_),
    .B1(_11219_),
    .A1(\cpu.ex.r_mult[19] ),
    .Y(_11495_),
    .A2(net769));
 sg13g2_nor3_1 _18311_ (.A(net764),
    .B(_11494_),
    .C(_11495_),
    .Y(_11496_));
 sg13g2_nand3_1 _18312_ (.B(_11424_),
    .C(_11065_),
    .A(_08394_),
    .Y(_11497_));
 sg13g2_nand3_1 _18313_ (.B(\cpu.ex.r_10[3] ),
    .C(_11075_),
    .A(_11069_),
    .Y(_11498_));
 sg13g2_a21oi_1 _18314_ (.A1(_11497_),
    .A2(_11498_),
    .Y(_11499_),
    .B1(_11063_));
 sg13g2_nor4_1 _18315_ (.A(_11484_),
    .B(_11493_),
    .C(_11496_),
    .D(_11499_),
    .Y(_11500_));
 sg13g2_nor2_1 _18316_ (.A(_09341_),
    .B(_11119_),
    .Y(_11501_));
 sg13g2_a21oi_2 _18317_ (.B1(_11501_),
    .Y(_11502_),
    .A2(_11500_),
    .A1(_11120_));
 sg13g2_nor2_1 _18318_ (.A(_11144_),
    .B(_11502_),
    .Y(_11503_));
 sg13g2_a21o_1 _18319_ (.A2(_11481_),
    .A1(_11456_),
    .B1(_11503_),
    .X(_11504_));
 sg13g2_a22oi_1 _18320_ (.Y(_11505_),
    .B1(_11184_),
    .B2(\cpu.ex.r_lr[1] ),
    .A2(_11179_),
    .A1(\cpu.ex.r_11[1] ));
 sg13g2_mux2_1 _18321_ (.A0(\cpu.ex.r_8[1] ),
    .A1(\cpu.ex.r_12[1] ),
    .S(net763),
    .X(_11506_));
 sg13g2_and2_1 _18322_ (.A(net773),
    .B(_11091_),
    .X(_11507_));
 sg13g2_nand3_1 _18323_ (.B(\cpu.ex.r_epc[1] ),
    .C(_11084_),
    .A(_11068_),
    .Y(_11508_));
 sg13g2_nand3_1 _18324_ (.B(\cpu.ex.r_13[1] ),
    .C(_11219_),
    .A(net763),
    .Y(_11509_));
 sg13g2_a21oi_1 _18325_ (.A1(_11508_),
    .A2(_11509_),
    .Y(_11510_),
    .B1(net764));
 sg13g2_a221oi_1 _18326_ (.B2(_11507_),
    .C1(_11510_),
    .B1(_11506_),
    .A1(\cpu.ex.r_9[1] ),
    .Y(_11511_),
    .A2(_11164_));
 sg13g2_mux2_1 _18327_ (.A0(_10772_),
    .A1(\cpu.ex.r_10[1] ),
    .S(net773),
    .X(_11512_));
 sg13g2_mux2_1 _18328_ (.A0(\cpu.ex.r_stmp[1] ),
    .A1(\cpu.ex.r_mult[17] ),
    .S(net904),
    .X(_11513_));
 sg13g2_a22oi_1 _18329_ (.Y(_11514_),
    .B1(_11513_),
    .B2(_11217_),
    .A2(_11512_),
    .A1(_11232_));
 sg13g2_and3_1 _18330_ (.X(_11515_),
    .A(_11505_),
    .B(_11511_),
    .C(_11514_));
 sg13g2_a22oi_1 _18331_ (.Y(_11516_),
    .B1(_11156_),
    .B2(\cpu.ex.r_14[1] ),
    .A2(_11154_),
    .A1(_10789_));
 sg13g2_inv_1 _18332_ (.Y(_11517_),
    .A(_00259_));
 sg13g2_a22oi_1 _18333_ (.Y(_11518_),
    .B1(_11156_),
    .B2(_11517_),
    .A2(_11154_),
    .A1(\cpu.ex.mmu_read[1] ));
 sg13g2_nand3b_1 _18334_ (.B(_11077_),
    .C(net904),
    .Y(_11519_),
    .A_N(_11518_));
 sg13g2_o21ai_1 _18335_ (.B1(_11519_),
    .Y(_11520_),
    .A1(_11409_),
    .A2(_11516_));
 sg13g2_nor2_1 _18336_ (.A(net612),
    .B(_11520_),
    .Y(_11521_));
 sg13g2_a22oi_1 _18337_ (.Y(_11522_),
    .B1(_11515_),
    .B2(_11521_),
    .A2(net612),
    .A1(_09351_));
 sg13g2_buf_1 _18338_ (.A(_11522_),
    .X(_11523_));
 sg13g2_buf_1 _18339_ (.A(_00200_),
    .X(_11524_));
 sg13g2_nor2_1 _18340_ (.A(_11137_),
    .B(_11524_),
    .Y(_11525_));
 sg13g2_o21ai_1 _18341_ (.B1(_11135_),
    .Y(_11526_),
    .A1(_08434_),
    .A2(net505));
 sg13g2_a22oi_1 _18342_ (.Y(_11527_),
    .B1(_11525_),
    .B2(_11526_),
    .A2(_11523_),
    .A1(_11191_));
 sg13g2_buf_2 _18343_ (.A(_11527_),
    .X(_11528_));
 sg13g2_and2_1 _18344_ (.A(net495),
    .B(_11198_),
    .X(_11529_));
 sg13g2_nand2b_1 _18345_ (.Y(_11530_),
    .B(net495),
    .A_N(_09469_));
 sg13g2_a22oi_1 _18346_ (.Y(_11531_),
    .B1(_11456_),
    .B2(_00297_),
    .A2(_11530_),
    .A1(_00191_));
 sg13g2_nor2_1 _18347_ (.A(net275),
    .B(_11531_),
    .Y(_11532_));
 sg13g2_a221oi_1 _18348_ (.B2(_11529_),
    .C1(_11532_),
    .B1(_11528_),
    .A1(net275),
    .Y(_11533_),
    .A2(_11504_));
 sg13g2_nor2_1 _18349_ (.A(_09467_),
    .B(\cpu.ex.c_mult_off[0] ),
    .Y(_11534_));
 sg13g2_nor2_1 _18350_ (.A(_08388_),
    .B(_11137_),
    .Y(_11535_));
 sg13g2_inv_1 _18351_ (.Y(_11536_),
    .A(_09284_));
 sg13g2_o21ai_1 _18352_ (.B1(_09285_),
    .Y(_11537_),
    .A1(_09320_),
    .A2(_09332_));
 sg13g2_and4_1 _18353_ (.A(_11536_),
    .B(_08427_),
    .C(_08429_),
    .D(_11537_),
    .X(_11538_));
 sg13g2_o21ai_1 _18354_ (.B1(_11538_),
    .Y(_11539_),
    .A1(_08434_),
    .A2(net505));
 sg13g2_buf_1 _18355_ (.A(_11539_),
    .X(_11540_));
 sg13g2_inv_1 _18356_ (.Y(_11541_),
    .A(net1052));
 sg13g2_a22oi_1 _18357_ (.Y(_11542_),
    .B1(_11072_),
    .B2(\cpu.ex.r_11[0] ),
    .A2(_11092_),
    .A1(\cpu.ex.r_8[0] ));
 sg13g2_nor2_1 _18358_ (.A(_11109_),
    .B(_11542_),
    .Y(_11543_));
 sg13g2_a22oi_1 _18359_ (.Y(_11544_),
    .B1(_11219_),
    .B2(\cpu.ex.r_9[0] ),
    .A2(net769),
    .A1(_10964_));
 sg13g2_nor2_1 _18360_ (.A(_11347_),
    .B(_11544_),
    .Y(_11545_));
 sg13g2_mux2_1 _18361_ (.A0(\cpu.ex.r_13[0] ),
    .A1(\cpu.ex.r_15[0] ),
    .S(net1018),
    .X(_11546_));
 sg13g2_a22oi_1 _18362_ (.Y(_11547_),
    .B1(_11546_),
    .B2(_11063_),
    .A2(net768),
    .A1(\cpu.ex.r_12[0] ));
 sg13g2_nor2_1 _18363_ (.A(_11159_),
    .B(_11547_),
    .Y(_11548_));
 sg13g2_nor3_1 _18364_ (.A(_11543_),
    .B(_11545_),
    .C(_11548_),
    .Y(_11549_));
 sg13g2_mux2_1 _18365_ (.A0(\cpu.ex.r_stmp[0] ),
    .A1(\cpu.ex.r_14[0] ),
    .S(net773),
    .X(_11550_));
 sg13g2_nor2_1 _18366_ (.A(_09286_),
    .B(_11409_),
    .Y(_11551_));
 sg13g2_a22oi_1 _18367_ (.Y(_11552_),
    .B1(_11551_),
    .B2(_11154_),
    .A2(_11550_),
    .A1(_11230_));
 sg13g2_nand4_1 _18368_ (.B(net902),
    .C(\cpu.ex.r_mult[16] ),
    .A(net772),
    .Y(_11553_),
    .D(_11065_));
 sg13g2_nand4_1 _18369_ (.B(net673),
    .C(\cpu.ex.r_10[0] ),
    .A(net902),
    .Y(_11554_),
    .D(_11061_));
 sg13g2_and4_1 _18370_ (.A(_11119_),
    .B(_11552_),
    .C(_11553_),
    .D(_11554_),
    .X(_11555_));
 sg13g2_a22oi_1 _18371_ (.Y(_11556_),
    .B1(_11549_),
    .B2(_11555_),
    .A2(net612),
    .A1(_11541_));
 sg13g2_buf_1 _18372_ (.A(_11556_),
    .X(_11557_));
 sg13g2_a22oi_1 _18373_ (.Y(_11558_),
    .B1(_11557_),
    .B2(_11192_),
    .A2(net398),
    .A1(_11535_));
 sg13g2_buf_1 _18374_ (.A(_11558_),
    .X(_11559_));
 sg13g2_or2_1 _18375_ (.X(_11560_),
    .B(\cpu.ex.c_mult_off[2] ),
    .A(\cpu.ex.c_mult_off[3] ));
 sg13g2_a21oi_1 _18376_ (.A1(_11534_),
    .A2(_11559_),
    .Y(_11561_),
    .B1(_11560_));
 sg13g2_a22oi_1 _18377_ (.Y(_11562_),
    .B1(_11533_),
    .B2(_11561_),
    .A2(_11455_),
    .A1(_11358_));
 sg13g2_nand3_1 _18378_ (.B(_11357_),
    .C(_11562_),
    .A(_11271_),
    .Y(_11563_));
 sg13g2_buf_8 _18379_ (.A(_11563_),
    .X(_11564_));
 sg13g2_and2_1 _18380_ (.A(_10953_),
    .B(_11044_),
    .X(_11565_));
 sg13g2_nor2_1 _18381_ (.A(_10909_),
    .B(_09463_),
    .Y(_11566_));
 sg13g2_a21oi_1 _18382_ (.A1(_10946_),
    .A2(_10940_),
    .Y(_11567_),
    .B1(_10913_));
 sg13g2_o21ai_1 _18383_ (.B1(_11567_),
    .Y(_11568_),
    .A1(_10907_),
    .A2(_11566_));
 sg13g2_a21oi_1 _18384_ (.A1(_10910_),
    .A2(_10907_),
    .Y(_11569_),
    .B1(_10848_));
 sg13g2_nand2b_1 _18385_ (.Y(_11570_),
    .B(net615),
    .A_N(_10913_));
 sg13g2_buf_1 _18386_ (.A(_11570_),
    .X(_11571_));
 sg13g2_a21oi_1 _18387_ (.A1(_10946_),
    .A2(_10940_),
    .Y(_11572_),
    .B1(_11571_));
 sg13g2_o21ai_1 _18388_ (.B1(_10910_),
    .Y(_11573_),
    .A1(_10907_),
    .A2(_11572_));
 sg13g2_a21oi_1 _18389_ (.A1(_10907_),
    .A2(_11572_),
    .Y(_11574_),
    .B1(net236));
 sg13g2_nor2_1 _18390_ (.A(_10848_),
    .B(net236),
    .Y(_11575_));
 sg13g2_a221oi_1 _18391_ (.B2(_11574_),
    .C1(_11575_),
    .B1(_11573_),
    .A1(_11568_),
    .Y(_11576_),
    .A2(_11569_));
 sg13g2_buf_2 _18392_ (.A(_11576_),
    .X(_11577_));
 sg13g2_inv_1 _18393_ (.Y(_11578_),
    .A(_11013_));
 sg13g2_a21oi_1 _18394_ (.A1(net234),
    .A2(_11577_),
    .Y(_11579_),
    .B1(_11578_));
 sg13g2_o21ai_1 _18395_ (.B1(_11040_),
    .Y(_11580_),
    .A1(net234),
    .A2(_11577_));
 sg13g2_nor2_1 _18396_ (.A(_11005_),
    .B(_11006_),
    .Y(_11581_));
 sg13g2_nor2b_1 _18397_ (.A(_11581_),
    .B_N(_11008_),
    .Y(_11582_));
 sg13g2_buf_1 _18398_ (.A(_11582_),
    .X(_11583_));
 sg13g2_buf_1 _18399_ (.A(_11583_),
    .X(_11584_));
 sg13g2_o21ai_1 _18400_ (.B1(_11012_),
    .Y(_11585_),
    .A1(_11013_),
    .A2(net202));
 sg13g2_nor2_1 _18401_ (.A(_11034_),
    .B(_11036_),
    .Y(_11586_));
 sg13g2_buf_1 _18402_ (.A(_11586_),
    .X(_11587_));
 sg13g2_nor3_1 _18403_ (.A(net550),
    .B(net273),
    .C(_11015_),
    .Y(_11588_));
 sg13g2_o21ai_1 _18404_ (.B1(_11588_),
    .Y(_11589_),
    .A1(_11577_),
    .A2(_11585_));
 sg13g2_o21ai_1 _18405_ (.B1(_11589_),
    .Y(_11590_),
    .A1(_11579_),
    .A2(_11580_));
 sg13g2_a221oi_1 _18406_ (.B2(_11565_),
    .C1(_11590_),
    .B1(_11564_),
    .A1(_10953_),
    .Y(_11591_),
    .A2(_11045_));
 sg13g2_buf_2 _18407_ (.A(_11591_),
    .X(_11592_));
 sg13g2_nand2_1 _18408_ (.Y(_11593_),
    .A(net204),
    .B(_10687_));
 sg13g2_buf_1 _18409_ (.A(_10687_),
    .X(_11594_));
 sg13g2_nor2_1 _18410_ (.A(_10618_),
    .B(net550),
    .Y(_11595_));
 sg13g2_nand2_1 _18411_ (.Y(_11596_),
    .A(net147),
    .B(_11595_));
 sg13g2_a21oi_1 _18412_ (.A1(_10759_),
    .A2(_10723_),
    .Y(_11597_),
    .B1(net1106));
 sg13g2_nor2_1 _18413_ (.A(net550),
    .B(_10757_),
    .Y(_11598_));
 sg13g2_a21o_1 _18414_ (.A2(_10720_),
    .A1(net779),
    .B1(_10721_),
    .X(_11599_));
 sg13g2_buf_1 _18415_ (.A(_11599_),
    .X(_11600_));
 sg13g2_a22oi_1 _18416_ (.Y(_11601_),
    .B1(_10762_),
    .B2(_11600_),
    .A2(_11598_),
    .A1(_11597_));
 sg13g2_a21oi_1 _18417_ (.A1(_11593_),
    .A2(_11596_),
    .Y(_11602_),
    .B1(_11601_));
 sg13g2_inv_1 _18418_ (.Y(_11603_),
    .A(net1108));
 sg13g2_nor2_1 _18419_ (.A(_11603_),
    .B(net550),
    .Y(_11604_));
 sg13g2_nand2_1 _18420_ (.Y(_11605_),
    .A(net204),
    .B(_11604_));
 sg13g2_nand3_1 _18421_ (.B(_10690_),
    .C(net615),
    .A(net1108),
    .Y(_11606_));
 sg13g2_a21oi_1 _18422_ (.A1(_11605_),
    .A2(_11606_),
    .Y(_11607_),
    .B1(_11601_));
 sg13g2_nand2_1 _18423_ (.Y(_11608_),
    .A(_10690_),
    .B(net615));
 sg13g2_inv_1 _18424_ (.Y(_11609_),
    .A(_11606_));
 sg13g2_a22oi_1 _18425_ (.Y(_11610_),
    .B1(_11609_),
    .B2(net204),
    .A2(_11604_),
    .A1(net147));
 sg13g2_o21ai_1 _18426_ (.B1(_11610_),
    .Y(_11611_),
    .A1(_11593_),
    .A2(_11608_));
 sg13g2_nor4_1 _18427_ (.A(_10581_),
    .B(_11602_),
    .C(_11607_),
    .D(_11611_),
    .Y(_11612_));
 sg13g2_o21ai_1 _18428_ (.B1(_11612_),
    .Y(_11613_),
    .A1(_10767_),
    .A2(_11592_));
 sg13g2_a21oi_1 _18429_ (.A1(_10617_),
    .A2(_11613_),
    .Y(_11614_),
    .B1(_10540_));
 sg13g2_nor2_1 _18430_ (.A(net234),
    .B(_11577_),
    .Y(_11615_));
 sg13g2_nor2_1 _18431_ (.A(_11579_),
    .B(_11615_),
    .Y(_11616_));
 sg13g2_nand4_1 _18432_ (.B(_11271_),
    .C(_11357_),
    .A(_10985_),
    .Y(_11617_),
    .D(_11562_));
 sg13g2_nand3_1 _18433_ (.B(_11042_),
    .C(_11617_),
    .A(_10953_),
    .Y(_11618_));
 sg13g2_nor3_1 _18434_ (.A(_11602_),
    .B(_11607_),
    .C(_11611_),
    .Y(_11619_));
 sg13g2_nand3b_1 _18435_ (.B(_11618_),
    .C(_11619_),
    .Y(_11620_),
    .A_N(_11616_));
 sg13g2_nand3b_1 _18436_ (.B(_10765_),
    .C(_11040_),
    .Y(_11621_),
    .A_N(_10697_));
 sg13g2_a21oi_1 _18437_ (.A1(_11619_),
    .A2(_11621_),
    .Y(_11622_),
    .B1(_10578_));
 sg13g2_nor3_1 _18438_ (.A(_10578_),
    .B(_10767_),
    .C(_11039_),
    .Y(_11623_));
 sg13g2_or2_1 _18439_ (.X(_11624_),
    .B(_11585_),
    .A(_11577_));
 sg13g2_and2_1 _18440_ (.A(_10953_),
    .B(_11617_),
    .X(_11625_));
 sg13g2_buf_1 _18441_ (.A(_11625_),
    .X(_11626_));
 sg13g2_a21o_1 _18442_ (.A2(_11624_),
    .A1(net537),
    .B1(_11626_),
    .X(_11627_));
 sg13g2_nand2_1 _18443_ (.Y(_11628_),
    .A(_10616_),
    .B(_10582_));
 sg13g2_a221oi_1 _18444_ (.B2(_11627_),
    .C1(_11628_),
    .B1(_11623_),
    .A1(_11620_),
    .Y(_11629_),
    .A2(_11622_));
 sg13g2_nor4_1 _18445_ (.A(_10616_),
    .B(_10578_),
    .C(_10767_),
    .D(_11039_),
    .Y(_11630_));
 sg13g2_a21oi_1 _18446_ (.A1(_11626_),
    .A2(_11630_),
    .Y(_11631_),
    .B1(net537));
 sg13g2_nor2_1 _18447_ (.A(net1030),
    .B(_10458_),
    .Y(_11632_));
 sg13g2_a21oi_1 _18448_ (.A1(net941),
    .A2(_10370_),
    .Y(_11633_),
    .B1(_11632_));
 sg13g2_buf_1 _18449_ (.A(_11633_),
    .X(_11634_));
 sg13g2_nor2_1 _18450_ (.A(net132),
    .B(_10465_),
    .Y(_11635_));
 sg13g2_nor4_2 _18451_ (.A(_11614_),
    .B(_11629_),
    .C(_11631_),
    .Y(_11636_),
    .D(_11635_));
 sg13g2_nor2_1 _18452_ (.A(_09466_),
    .B(_10463_),
    .Y(_11637_));
 sg13g2_buf_1 _18453_ (.A(_10653_),
    .X(_11638_));
 sg13g2_nand2b_1 _18454_ (.Y(_11639_),
    .B(_10803_),
    .A_N(_10983_));
 sg13g2_buf_2 _18455_ (.A(_11639_),
    .X(_11640_));
 sg13g2_nand2_1 _18456_ (.Y(_11641_),
    .A(_10838_),
    .B(net277));
 sg13g2_buf_2 _18457_ (.A(_11641_),
    .X(_11642_));
 sg13g2_nor2_2 _18458_ (.A(_11640_),
    .B(_11642_),
    .Y(_11643_));
 sg13g2_buf_1 _18459_ (.A(_10723_),
    .X(_11644_));
 sg13g2_inv_2 _18460_ (.Y(_11645_),
    .A(_10876_));
 sg13g2_nor4_1 _18461_ (.A(net273),
    .B(net173),
    .C(_10757_),
    .D(_11645_),
    .Y(_11646_));
 sg13g2_and4_1 _18462_ (.A(net174),
    .B(net147),
    .C(_11643_),
    .D(_11646_),
    .X(_11647_));
 sg13g2_nand2_1 _18463_ (.Y(_11648_),
    .A(_10583_),
    .B(net1030));
 sg13g2_o21ai_1 _18464_ (.B1(_11648_),
    .Y(_11649_),
    .A1(_10535_),
    .A2(_10613_));
 sg13g2_buf_1 _18465_ (.A(_11649_),
    .X(_11650_));
 sg13g2_and2_1 _18466_ (.A(_10903_),
    .B(_10905_),
    .X(_11651_));
 sg13g2_buf_2 _18467_ (.A(_11651_),
    .X(_11652_));
 sg13g2_buf_1 _18468_ (.A(_11652_),
    .X(_11653_));
 sg13g2_nor3_1 _18469_ (.A(net232),
    .B(net202),
    .C(_10461_),
    .Y(_11654_));
 sg13g2_and4_1 _18470_ (.A(_11647_),
    .B(_10576_),
    .C(net146),
    .D(_11654_),
    .X(_11655_));
 sg13g2_nor3_1 _18471_ (.A(_11637_),
    .B(_09481_),
    .C(_11655_),
    .Y(_11656_));
 sg13g2_buf_1 _18472_ (.A(_11656_),
    .X(_11657_));
 sg13g2_buf_1 _18473_ (.A(_11657_),
    .X(_11658_));
 sg13g2_o21ai_1 _18474_ (.B1(net71),
    .Y(_11659_),
    .A1(_10467_),
    .A2(_11636_));
 sg13g2_buf_1 _18475_ (.A(_10983_),
    .X(_11660_));
 sg13g2_buf_1 _18476_ (.A(_11564_),
    .X(_11661_));
 sg13g2_buf_1 _18477_ (.A(net102),
    .X(_11662_));
 sg13g2_buf_1 _18478_ (.A(net88),
    .X(_11663_));
 sg13g2_nand3_1 _18479_ (.B(net346),
    .C(net70),
    .A(_09481_),
    .Y(_11664_));
 sg13g2_nand2b_1 _18480_ (.Y(_11665_),
    .B(_10360_),
    .A_N(_10358_));
 sg13g2_buf_1 _18481_ (.A(_11665_),
    .X(_11666_));
 sg13g2_buf_1 _18482_ (.A(_11666_),
    .X(_11667_));
 sg13g2_a21o_1 _18483_ (.A2(_11664_),
    .A1(_11659_),
    .B1(_11667_),
    .X(_11668_));
 sg13g2_nand2_1 _18484_ (.Y(\cpu.ex.c_mult[0] ),
    .A(_10368_),
    .B(_11668_));
 sg13g2_buf_1 _18485_ (.A(\cpu.dec.load ),
    .X(_11669_));
 sg13g2_o21ai_1 _18486_ (.B1(_08457_),
    .Y(_11670_),
    .A1(_08431_),
    .A2(_08525_));
 sg13g2_buf_1 _18487_ (.A(_11670_),
    .X(_11671_));
 sg13g2_nor2_1 _18488_ (.A(_09385_),
    .B(_09473_),
    .Y(_11672_));
 sg13g2_or2_1 _18489_ (.X(_11673_),
    .B(_11672_),
    .A(_10363_));
 sg13g2_buf_1 _18490_ (.A(_11673_),
    .X(_11674_));
 sg13g2_nor2_1 _18491_ (.A(\cpu.ex.c_div_running ),
    .B(\cpu.ex.c_mult_running ),
    .Y(_11675_));
 sg13g2_nand2_1 _18492_ (.Y(_11676_),
    .A(_10964_),
    .B(\cpu.dec.r_swapsp ));
 sg13g2_nor3_1 _18493_ (.A(net1053),
    .B(_09385_),
    .C(_09457_),
    .Y(_11677_));
 sg13g2_buf_1 _18494_ (.A(_00258_),
    .X(_11678_));
 sg13g2_nand2_1 _18495_ (.Y(_11679_),
    .A(_11136_),
    .B(\cpu.cond[2] ));
 sg13g2_inv_2 _18496_ (.Y(_11680_),
    .A(_08499_));
 sg13g2_a21o_1 _18497_ (.A2(_11679_),
    .A1(_11678_),
    .B1(_11680_),
    .X(_11681_));
 sg13g2_buf_1 _18498_ (.A(_11681_),
    .X(_11682_));
 sg13g2_o21ai_1 _18499_ (.B1(net762),
    .Y(_11683_),
    .A1(_11136_),
    .A2(\cpu.dec.jmp ));
 sg13g2_nand4_1 _18500_ (.B(_11676_),
    .C(_11677_),
    .A(_11675_),
    .Y(_11684_),
    .D(_11683_));
 sg13g2_nand3_1 _18501_ (.B(_11674_),
    .C(_11684_),
    .A(_11671_),
    .Y(_11685_));
 sg13g2_buf_1 _18502_ (.A(_11685_),
    .X(_11686_));
 sg13g2_and2_1 _18503_ (.A(net930),
    .B(_11686_),
    .X(_11687_));
 sg13g2_buf_1 _18504_ (.A(_11687_),
    .X(_11688_));
 sg13g2_buf_1 _18505_ (.A(_11688_),
    .X(_11689_));
 sg13g2_nand2_1 _18506_ (.Y(_11690_),
    .A(_00310_),
    .B(net101));
 sg13g2_nor2_1 _18507_ (.A(_09487_),
    .B(_09498_),
    .Y(_11691_));
 sg13g2_inv_1 _18508_ (.Y(_11692_),
    .A(_09932_));
 sg13g2_o21ai_1 _18509_ (.B1(_11692_),
    .Y(_11693_),
    .A1(_09924_),
    .A2(_11691_));
 sg13g2_nor2b_2 _18510_ (.A(_09363_),
    .B_N(_11693_),
    .Y(_11694_));
 sg13g2_inv_1 _18511_ (.Y(_11695_),
    .A(_11694_));
 sg13g2_o21ai_1 _18512_ (.B1(_11690_),
    .Y(_11696_),
    .A1(net101),
    .A2(_11695_));
 sg13g2_nand2_1 _18513_ (.Y(_11697_),
    .A(net1053),
    .B(_11696_));
 sg13g2_o21ai_1 _18514_ (.B1(_11697_),
    .Y(_00054_),
    .A1(_11669_),
    .A2(_11690_));
 sg13g2_buf_1 _18515_ (.A(_09479_),
    .X(_11698_));
 sg13g2_nand2_1 _18516_ (.Y(_11699_),
    .A(_10346_),
    .B(_11698_));
 sg13g2_buf_1 _18517_ (.A(_10803_),
    .X(_11700_));
 sg13g2_and3_1 _18518_ (.X(_11701_),
    .A(_11271_),
    .B(_11357_),
    .C(_11562_));
 sg13g2_buf_1 _18519_ (.A(_11701_),
    .X(_11702_));
 sg13g2_nor2_1 _18520_ (.A(net231),
    .B(_11702_),
    .Y(_11703_));
 sg13g2_mux2_1 _18521_ (.A0(_11699_),
    .A1(_10346_),
    .S(_11703_),
    .X(_11704_));
 sg13g2_buf_1 _18522_ (.A(_09461_),
    .X(_11705_));
 sg13g2_buf_1 _18523_ (.A(net532),
    .X(_11706_));
 sg13g2_buf_1 _18524_ (.A(_11706_),
    .X(_11707_));
 sg13g2_a22oi_1 _18525_ (.Y(_11708_),
    .B1(_11703_),
    .B2(net441),
    .A2(_11657_),
    .A1(_10346_));
 sg13g2_o21ai_1 _18526_ (.B1(_11708_),
    .Y(_11709_),
    .A1(_09477_),
    .A2(_11704_));
 sg13g2_buf_1 _18527_ (.A(\cpu.ex.r_mult[1] ),
    .X(_11710_));
 sg13g2_inv_1 _18528_ (.Y(_11711_),
    .A(_11710_));
 sg13g2_a21oi_1 _18529_ (.A1(net492),
    .A2(_10364_),
    .Y(_11712_),
    .B1(_11711_));
 sg13g2_a21o_1 _18530_ (.A2(_11709_),
    .A1(net492),
    .B1(_11712_),
    .X(\cpu.ex.c_mult[1] ));
 sg13g2_nand2_1 _18531_ (.Y(_11713_),
    .A(_11710_),
    .B(net533));
 sg13g2_buf_1 _18532_ (.A(_10959_),
    .X(_11714_));
 sg13g2_o21ai_1 _18533_ (.B1(_10346_),
    .Y(_11715_),
    .A1(_08975_),
    .A2(_10528_));
 sg13g2_a21oi_1 _18534_ (.A1(net779),
    .A2(_10800_),
    .Y(_11716_),
    .B1(_11715_));
 sg13g2_nand2_1 _18535_ (.Y(_11717_),
    .A(net628),
    .B(_11716_));
 sg13g2_xnor2_1 _18536_ (.Y(_11718_),
    .A(net272),
    .B(_11717_));
 sg13g2_nand2_1 _18537_ (.Y(_11719_),
    .A(net102),
    .B(_11718_));
 sg13g2_mux2_1 _18538_ (.A0(_11710_),
    .A1(_11713_),
    .S(_11719_),
    .X(_11720_));
 sg13g2_inv_1 _18539_ (.Y(_11721_),
    .A(_11720_));
 sg13g2_nor2_1 _18540_ (.A(net533),
    .B(_11719_),
    .Y(_11722_));
 sg13g2_a221oi_1 _18541_ (.B2(net1122),
    .C1(_11722_),
    .B1(_11721_),
    .A1(_11710_),
    .Y(_11723_),
    .A2(_11657_));
 sg13g2_nand2_1 _18542_ (.Y(_11724_),
    .A(\cpu.ex.r_mult[2] ),
    .B(_10366_));
 sg13g2_o21ai_1 _18543_ (.B1(_11724_),
    .Y(\cpu.ex.c_mult[2] ),
    .A1(_11666_),
    .A2(_11723_));
 sg13g2_o21ai_1 _18544_ (.B1(_11711_),
    .Y(_11725_),
    .A1(_10955_),
    .A2(_10958_));
 sg13g2_nor3_1 _18545_ (.A(_11711_),
    .B(_10955_),
    .C(_10958_),
    .Y(_11726_));
 sg13g2_a21oi_1 _18546_ (.A1(_11716_),
    .A2(_11725_),
    .Y(_11727_),
    .B1(_11726_));
 sg13g2_buf_1 _18547_ (.A(_00120_),
    .X(_11728_));
 sg13g2_inv_1 _18548_ (.Y(_11729_),
    .A(_11728_));
 sg13g2_nor2_1 _18549_ (.A(_11729_),
    .B(_10943_),
    .Y(_11730_));
 sg13g2_buf_1 _18550_ (.A(_10948_),
    .X(_11731_));
 sg13g2_nor2_1 _18551_ (.A(_11728_),
    .B(net230),
    .Y(_11732_));
 sg13g2_a21oi_1 _18552_ (.A1(_11661_),
    .A2(_11730_),
    .Y(_11733_),
    .B1(_11732_));
 sg13g2_nor3_1 _18553_ (.A(net441),
    .B(_11727_),
    .C(_11733_),
    .Y(_11734_));
 sg13g2_buf_1 _18554_ (.A(_10943_),
    .X(_11735_));
 sg13g2_and4_1 _18555_ (.A(_11728_),
    .B(net229),
    .C(net88),
    .D(_11727_),
    .X(_11736_));
 sg13g2_nand2_1 _18556_ (.Y(_11737_),
    .A(net230),
    .B(_11727_));
 sg13g2_a221oi_1 _18557_ (.B2(_11737_),
    .C1(_11728_),
    .B1(net88),
    .A1(_09455_),
    .Y(_11738_),
    .A2(_09459_));
 sg13g2_nor3_1 _18558_ (.A(_11734_),
    .B(_11736_),
    .C(_11738_),
    .Y(_11739_));
 sg13g2_buf_1 _18559_ (.A(_11702_),
    .X(_11740_));
 sg13g2_nor2_1 _18560_ (.A(net533),
    .B(net100),
    .Y(_11741_));
 sg13g2_a22oi_1 _18561_ (.Y(_11742_),
    .B1(_11741_),
    .B2(net229),
    .A2(_11657_),
    .A1(_11729_));
 sg13g2_o21ai_1 _18562_ (.B1(_11742_),
    .Y(_11743_),
    .A1(_09477_),
    .A2(_11739_));
 sg13g2_a22oi_1 _18563_ (.Y(_11744_),
    .B1(_11743_),
    .B2(net492),
    .A2(_10367_),
    .A1(\cpu.ex.r_mult[3] ));
 sg13g2_inv_1 _18564_ (.Y(\cpu.ex.c_mult[3] ),
    .A(_11744_));
 sg13g2_inv_1 _18565_ (.Y(_11745_),
    .A(_00127_));
 sg13g2_a221oi_1 _18566_ (.B2(_11725_),
    .C1(_11726_),
    .B1(_11716_),
    .A1(_11729_),
    .Y(_11746_),
    .A2(_10943_));
 sg13g2_buf_1 _18567_ (.A(_11746_),
    .X(_11747_));
 sg13g2_nor2_1 _18568_ (.A(_11730_),
    .B(_11747_),
    .Y(_11748_));
 sg13g2_nor3_1 _18569_ (.A(_11745_),
    .B(_10908_),
    .C(_11748_),
    .Y(_11749_));
 sg13g2_or2_1 _18570_ (.X(_11750_),
    .B(_11747_),
    .A(_11730_));
 sg13g2_nor2_1 _18571_ (.A(_11745_),
    .B(_11652_),
    .Y(_11751_));
 sg13g2_nor2_1 _18572_ (.A(_00127_),
    .B(_10907_),
    .Y(_11752_));
 sg13g2_a21oi_1 _18573_ (.A1(net102),
    .A2(_11751_),
    .Y(_11753_),
    .B1(_11752_));
 sg13g2_nor2_1 _18574_ (.A(net232),
    .B(_11748_),
    .Y(_11754_));
 sg13g2_o21ai_1 _18575_ (.B1(_11745_),
    .Y(_11755_),
    .A1(net100),
    .A2(_11754_));
 sg13g2_o21ai_1 _18576_ (.B1(_11755_),
    .Y(_11756_),
    .A1(_11750_),
    .A2(_11753_));
 sg13g2_a22oi_1 _18577_ (.Y(_11757_),
    .B1(_11756_),
    .B2(net533),
    .A2(_11749_),
    .A1(net88));
 sg13g2_a22oi_1 _18578_ (.Y(_11758_),
    .B1(_11741_),
    .B2(net232),
    .A2(_11657_),
    .A1(_11745_));
 sg13g2_o21ai_1 _18579_ (.B1(_11758_),
    .Y(_11759_),
    .A1(_09477_),
    .A2(_11757_));
 sg13g2_a22oi_1 _18580_ (.Y(_11760_),
    .B1(_11759_),
    .B2(_10362_),
    .A2(_10367_),
    .A1(\cpu.ex.r_mult[4] ));
 sg13g2_inv_1 _18581_ (.Y(\cpu.ex.c_mult[4] ),
    .A(_11760_));
 sg13g2_buf_1 _18582_ (.A(_00139_),
    .X(_11761_));
 sg13g2_inv_1 _18583_ (.Y(_11762_),
    .A(_11761_));
 sg13g2_nor2_1 _18584_ (.A(_11761_),
    .B(net490),
    .Y(_11763_));
 sg13g2_a21oi_1 _18585_ (.A1(net232),
    .A2(_11748_),
    .Y(_11764_),
    .B1(_11745_));
 sg13g2_nor3_1 _18586_ (.A(_11706_),
    .B(_11754_),
    .C(_11764_),
    .Y(_11765_));
 sg13g2_xnor2_1 _18587_ (.Y(_11766_),
    .A(_10877_),
    .B(_11765_));
 sg13g2_nand2_1 _18588_ (.Y(_11767_),
    .A(_11661_),
    .B(_11766_));
 sg13g2_mux2_1 _18589_ (.A0(_11761_),
    .A1(_11763_),
    .S(_11767_),
    .X(_11768_));
 sg13g2_nor2_1 _18590_ (.A(_11698_),
    .B(_11767_),
    .Y(_11769_));
 sg13g2_a221oi_1 _18591_ (.B2(_09476_),
    .C1(_11769_),
    .B1(_11768_),
    .A1(_11762_),
    .Y(_11770_),
    .A2(_11658_));
 sg13g2_nand2_1 _18592_ (.Y(_11771_),
    .A(\cpu.ex.r_mult[5] ),
    .B(_10366_));
 sg13g2_o21ai_1 _18593_ (.B1(_11771_),
    .Y(\cpu.ex.c_mult[5] ),
    .A1(_11667_),
    .A2(_11770_));
 sg13g2_and2_1 _18594_ (.A(_11761_),
    .B(_10876_),
    .X(_11772_));
 sg13g2_or4_1 _18595_ (.A(_11730_),
    .B(_11747_),
    .C(_11751_),
    .D(_11772_),
    .X(_11773_));
 sg13g2_buf_1 _18596_ (.A(_11773_),
    .X(_11774_));
 sg13g2_nand2_1 _18597_ (.Y(_11775_),
    .A(_11761_),
    .B(_10876_));
 sg13g2_nor2_1 _18598_ (.A(_11761_),
    .B(_10877_),
    .Y(_11776_));
 sg13g2_a21oi_1 _18599_ (.A1(_11752_),
    .A2(_11775_),
    .Y(_11777_),
    .B1(_11776_));
 sg13g2_and2_1 _18600_ (.A(_11774_),
    .B(_11777_),
    .X(_11778_));
 sg13g2_buf_1 _18601_ (.A(_11778_),
    .X(_11779_));
 sg13g2_o21ai_1 _18602_ (.B1(net202),
    .Y(_11780_),
    .A1(net490),
    .A2(_11779_));
 sg13g2_or3_1 _18603_ (.A(net490),
    .B(net202),
    .C(_11779_),
    .X(_11781_));
 sg13g2_a21oi_1 _18604_ (.A1(_11780_),
    .A2(_11781_),
    .Y(_11782_),
    .B1(net100));
 sg13g2_nor2_1 _18605_ (.A(_00151_),
    .B(net629),
    .Y(_11783_));
 sg13g2_mux2_1 _18606_ (.A0(_11783_),
    .A1(_00151_),
    .S(_11782_),
    .X(_11784_));
 sg13g2_or3_1 _18607_ (.A(_11637_),
    .B(_09481_),
    .C(_11655_),
    .X(_11785_));
 sg13g2_buf_2 _18608_ (.A(_11785_),
    .X(_11786_));
 sg13g2_nor2_1 _18609_ (.A(_00151_),
    .B(_11786_),
    .Y(_11787_));
 sg13g2_a221oi_1 _18610_ (.B2(_09476_),
    .C1(_11787_),
    .B1(_11784_),
    .A1(net441),
    .Y(_11788_),
    .A2(_11782_));
 sg13g2_nor2_1 _18611_ (.A(_11666_),
    .B(_11788_),
    .Y(_11789_));
 sg13g2_a21oi_1 _18612_ (.A1(\cpu.ex.r_mult[6] ),
    .A2(net278),
    .Y(_11790_),
    .B1(_11789_));
 sg13g2_inv_1 _18613_ (.Y(\cpu.ex.c_mult[6] ),
    .A(_11790_));
 sg13g2_nand2_1 _18614_ (.Y(_11791_),
    .A(_09481_),
    .B(net492));
 sg13g2_buf_2 _18615_ (.A(_11791_),
    .X(_11792_));
 sg13g2_nor2_2 _18616_ (.A(_00163_),
    .B(net629),
    .Y(_11793_));
 sg13g2_nor2_1 _18617_ (.A(net234),
    .B(_11779_),
    .Y(_11794_));
 sg13g2_nand2_1 _18618_ (.Y(_11795_),
    .A(net234),
    .B(_11779_));
 sg13g2_a22oi_1 _18619_ (.Y(_11796_),
    .B1(_11795_),
    .B2(_11783_),
    .A2(_11794_),
    .A1(net628));
 sg13g2_xnor2_1 _18620_ (.Y(_11797_),
    .A(net273),
    .B(_11796_));
 sg13g2_nand2_1 _18621_ (.Y(_11798_),
    .A(net70),
    .B(_11797_));
 sg13g2_xor2_1 _18622_ (.B(_11798_),
    .A(_11793_),
    .X(_11799_));
 sg13g2_nor2_1 _18623_ (.A(_11666_),
    .B(_11786_),
    .Y(_11800_));
 sg13g2_buf_1 _18624_ (.A(_11800_),
    .X(_11801_));
 sg13g2_inv_1 _18625_ (.Y(_11802_),
    .A(_00163_));
 sg13g2_a22oi_1 _18626_ (.Y(_11803_),
    .B1(net62),
    .B2(_11802_),
    .A2(net278),
    .A1(\cpu.ex.r_mult[7] ));
 sg13g2_o21ai_1 _18627_ (.B1(_11803_),
    .Y(\cpu.ex.c_mult[7] ),
    .A1(_11792_),
    .A2(_11799_));
 sg13g2_buf_1 _18628_ (.A(_00164_),
    .X(_11804_));
 sg13g2_nor2_2 _18629_ (.A(_11804_),
    .B(net629),
    .Y(_11805_));
 sg13g2_buf_1 _18630_ (.A(_10757_),
    .X(_11806_));
 sg13g2_o21ai_1 _18631_ (.B1(_11783_),
    .Y(_11807_),
    .A1(_11802_),
    .A2(_11586_));
 sg13g2_nand2_1 _18632_ (.Y(_11808_),
    .A(net202),
    .B(_11793_));
 sg13g2_a22oi_1 _18633_ (.Y(_11809_),
    .B1(_11807_),
    .B2(_11808_),
    .A2(_11777_),
    .A1(_11774_));
 sg13g2_nand3_1 _18634_ (.B(net273),
    .C(_11583_),
    .A(net628),
    .Y(_11810_));
 sg13g2_a21oi_1 _18635_ (.A1(_11774_),
    .A2(_11777_),
    .Y(_11811_),
    .B1(_11810_));
 sg13g2_nor2_1 _18636_ (.A(net234),
    .B(_11807_),
    .Y(_11812_));
 sg13g2_and2_1 _18637_ (.A(net273),
    .B(_11793_),
    .X(_11813_));
 sg13g2_nor4_1 _18638_ (.A(_11809_),
    .B(_11811_),
    .C(_11812_),
    .D(_11813_),
    .Y(_11814_));
 sg13g2_buf_2 _18639_ (.A(_11814_),
    .X(_11815_));
 sg13g2_xnor2_1 _18640_ (.Y(_11816_),
    .A(net201),
    .B(_11815_));
 sg13g2_nand2_1 _18641_ (.Y(_11817_),
    .A(_11662_),
    .B(_11816_));
 sg13g2_mux2_1 _18642_ (.A0(_11804_),
    .A1(_11805_),
    .S(_11817_),
    .X(_11818_));
 sg13g2_nand3_1 _18643_ (.B(net201),
    .C(_11662_),
    .A(net441),
    .Y(_11819_));
 sg13g2_o21ai_1 _18644_ (.B1(_11819_),
    .Y(_11820_),
    .A1(_11804_),
    .A2(_11786_));
 sg13g2_a21oi_1 _18645_ (.A1(net1122),
    .A2(_11818_),
    .Y(_11821_),
    .B1(_11820_));
 sg13g2_nand2_1 _18646_ (.Y(_11822_),
    .A(\cpu.ex.r_mult[8] ),
    .B(net278));
 sg13g2_o21ai_1 _18647_ (.B1(_11822_),
    .Y(\cpu.ex.c_mult[8] ),
    .A1(net442),
    .A2(_11821_));
 sg13g2_nor2_1 _18648_ (.A(_00165_),
    .B(net629),
    .Y(_11823_));
 sg13g2_buf_1 _18649_ (.A(_11823_),
    .X(_11824_));
 sg13g2_nand2b_1 _18650_ (.Y(_11825_),
    .B(_11805_),
    .A_N(_11815_));
 sg13g2_nand2b_1 _18651_ (.Y(_11826_),
    .B(net628),
    .A_N(_11804_));
 sg13g2_buf_1 _18652_ (.A(_11826_),
    .X(_11827_));
 sg13g2_a21o_1 _18653_ (.A2(_11827_),
    .A1(_11815_),
    .B1(net203),
    .X(_11828_));
 sg13g2_buf_1 _18654_ (.A(_11600_),
    .X(_11829_));
 sg13g2_a21oi_1 _18655_ (.A1(_11825_),
    .A2(_11828_),
    .Y(_11830_),
    .B1(net172));
 sg13g2_nor2_1 _18656_ (.A(_11815_),
    .B(_11827_),
    .Y(_11831_));
 sg13g2_a21oi_2 _18657_ (.B1(net203),
    .Y(_11832_),
    .A2(_11827_),
    .A1(_11815_));
 sg13g2_nor3_1 _18658_ (.A(net173),
    .B(_11831_),
    .C(_11832_),
    .Y(_11833_));
 sg13g2_nor3_1 _18659_ (.A(net100),
    .B(_11830_),
    .C(_11833_),
    .Y(_11834_));
 sg13g2_xnor2_1 _18660_ (.Y(_11835_),
    .A(_11824_),
    .B(_11834_));
 sg13g2_inv_1 _18661_ (.Y(_11836_),
    .A(_00165_));
 sg13g2_a22oi_1 _18662_ (.Y(_11837_),
    .B1(net62),
    .B2(_11836_),
    .A2(_10366_),
    .A1(\cpu.ex.r_mult[9] ));
 sg13g2_o21ai_1 _18663_ (.B1(_11837_),
    .Y(\cpu.ex.c_mult[9] ),
    .A1(_11792_),
    .A2(_11835_));
 sg13g2_and2_1 _18664_ (.A(_09481_),
    .B(net492),
    .X(_11838_));
 sg13g2_buf_1 _18665_ (.A(_11838_),
    .X(_11839_));
 sg13g2_buf_1 _18666_ (.A(_10692_),
    .X(_11840_));
 sg13g2_and2_1 _18667_ (.A(net173),
    .B(_11824_),
    .X(_11841_));
 sg13g2_buf_1 _18668_ (.A(_11841_),
    .X(_11842_));
 sg13g2_or3_1 _18669_ (.A(_11831_),
    .B(_11832_),
    .C(_11842_),
    .X(_11843_));
 sg13g2_buf_1 _18670_ (.A(_11843_),
    .X(_11844_));
 sg13g2_or2_1 _18671_ (.X(_11845_),
    .B(_11824_),
    .A(net173));
 sg13g2_buf_1 _18672_ (.A(_11845_),
    .X(_11846_));
 sg13g2_nand2_1 _18673_ (.Y(_11847_),
    .A(_11844_),
    .B(_11846_));
 sg13g2_xnor2_1 _18674_ (.Y(_11848_),
    .A(net200),
    .B(_11847_));
 sg13g2_nand2_1 _18675_ (.Y(_11849_),
    .A(net70),
    .B(_11848_));
 sg13g2_buf_2 _18676_ (.A(_00166_),
    .X(_11850_));
 sg13g2_nor2_2 _18677_ (.A(_11850_),
    .B(net629),
    .Y(_11851_));
 sg13g2_xnor2_1 _18678_ (.Y(_11852_),
    .A(_11849_),
    .B(_11851_));
 sg13g2_nand2_1 _18679_ (.Y(_11853_),
    .A(net492),
    .B(net71));
 sg13g2_nor2_1 _18680_ (.A(_11850_),
    .B(_11853_),
    .Y(_11854_));
 sg13g2_a221oi_1 _18681_ (.B2(_11852_),
    .C1(_11854_),
    .B1(_11839_),
    .A1(\cpu.ex.r_mult[10] ),
    .Y(_11855_),
    .A2(net278));
 sg13g2_inv_1 _18682_ (.Y(\cpu.ex.c_mult[10] ),
    .A(_11855_));
 sg13g2_nand2b_1 _18683_ (.Y(_11856_),
    .B(net628),
    .A_N(_11850_));
 sg13g2_buf_1 _18684_ (.A(_11856_),
    .X(_11857_));
 sg13g2_a21oi_1 _18685_ (.A1(_11806_),
    .A2(_11805_),
    .Y(_11858_),
    .B1(_11813_));
 sg13g2_a21oi_1 _18686_ (.A1(net203),
    .A2(_11827_),
    .Y(_11859_),
    .B1(_11858_));
 sg13g2_a221oi_1 _18687_ (.B2(_11846_),
    .C1(_11842_),
    .B1(_11859_),
    .A1(net200),
    .Y(_11860_),
    .A2(_11851_));
 sg13g2_a21oi_1 _18688_ (.A1(net174),
    .A2(_11857_),
    .Y(_11861_),
    .B1(_11860_));
 sg13g2_nor2_1 _18689_ (.A(net200),
    .B(_11644_),
    .Y(_11862_));
 sg13g2_nor3_1 _18690_ (.A(_00165_),
    .B(_11850_),
    .C(_11705_),
    .Y(_11863_));
 sg13g2_o21ai_1 _18691_ (.B1(_11863_),
    .Y(_11864_),
    .A1(_11702_),
    .A2(_11862_));
 sg13g2_nor4_1 _18692_ (.A(net200),
    .B(_11600_),
    .C(_11824_),
    .D(_11857_),
    .Y(_11865_));
 sg13g2_xnor2_1 _18693_ (.Y(_11866_),
    .A(net173),
    .B(_11824_));
 sg13g2_nor3_1 _18694_ (.A(net174),
    .B(_11851_),
    .C(_11866_),
    .Y(_11867_));
 sg13g2_o21ai_1 _18695_ (.B1(_11564_),
    .Y(_11868_),
    .A1(_11865_),
    .A2(_11867_));
 sg13g2_nor2_1 _18696_ (.A(net273),
    .B(net201),
    .Y(_11869_));
 sg13g2_nor3_1 _18697_ (.A(_00163_),
    .B(_11804_),
    .C(_11705_),
    .Y(_11870_));
 sg13g2_o21ai_1 _18698_ (.B1(_11870_),
    .Y(_11871_),
    .A1(_11869_),
    .A2(_11702_));
 sg13g2_and4_1 _18699_ (.A(net276),
    .B(net201),
    .C(_11793_),
    .D(_11827_),
    .X(_11872_));
 sg13g2_xnor2_1 _18700_ (.Y(_11873_),
    .A(net201),
    .B(_11805_));
 sg13g2_nor3_1 _18701_ (.A(net276),
    .B(_11793_),
    .C(_11873_),
    .Y(_11874_));
 sg13g2_o21ai_1 _18702_ (.B1(_11564_),
    .Y(_11875_),
    .A1(_11872_),
    .A2(_11874_));
 sg13g2_a221oi_1 _18703_ (.B2(_11875_),
    .C1(_11796_),
    .B1(_11871_),
    .A1(_11864_),
    .Y(_11876_),
    .A2(_11868_));
 sg13g2_buf_1 _18704_ (.A(_11876_),
    .X(_11877_));
 sg13g2_or3_1 _18705_ (.A(_11594_),
    .B(_11861_),
    .C(_11877_),
    .X(_11878_));
 sg13g2_o21ai_1 _18706_ (.B1(_11594_),
    .Y(_11879_),
    .A1(_11861_),
    .A2(_11877_));
 sg13g2_a21oi_1 _18707_ (.A1(_11878_),
    .A2(_11879_),
    .Y(_11880_),
    .B1(net100));
 sg13g2_buf_2 _18708_ (.A(_00167_),
    .X(_11881_));
 sg13g2_nor2_1 _18709_ (.A(_11881_),
    .B(net629),
    .Y(_11882_));
 sg13g2_xnor2_1 _18710_ (.Y(_11883_),
    .A(_11880_),
    .B(_11882_));
 sg13g2_inv_1 _18711_ (.Y(_11884_),
    .A(_11881_));
 sg13g2_a22oi_1 _18712_ (.Y(_11885_),
    .B1(net62),
    .B2(_11884_),
    .A2(_10366_),
    .A1(\cpu.ex.r_mult[11] ));
 sg13g2_o21ai_1 _18713_ (.B1(_11885_),
    .Y(\cpu.ex.c_mult[11] ),
    .A1(_11792_),
    .A2(_11883_));
 sg13g2_buf_1 _18714_ (.A(_10575_),
    .X(_11886_));
 sg13g2_o21ai_1 _18715_ (.B1(_11881_),
    .Y(_11887_),
    .A1(_10656_),
    .A2(_10685_));
 sg13g2_nor3_1 _18716_ (.A(_11850_),
    .B(_10619_),
    .C(_10651_),
    .Y(_11888_));
 sg13g2_nor3_1 _18717_ (.A(_11881_),
    .B(_10656_),
    .C(_10685_),
    .Y(_11889_));
 sg13g2_a21oi_1 _18718_ (.A1(_11887_),
    .A2(_11888_),
    .Y(_11890_),
    .B1(_11889_));
 sg13g2_nor2_1 _18719_ (.A(net441),
    .B(_11890_),
    .Y(_11891_));
 sg13g2_buf_1 _18720_ (.A(_10693_),
    .X(_11892_));
 sg13g2_mux2_1 _18721_ (.A0(_11881_),
    .A1(_11882_),
    .S(_10687_),
    .X(_11893_));
 sg13g2_a22oi_1 _18722_ (.Y(_11894_),
    .B1(_11893_),
    .B2(_11850_),
    .A2(net170),
    .A1(net532));
 sg13g2_nor2b_1 _18723_ (.A(_11889_),
    .B_N(_11887_),
    .Y(_11895_));
 sg13g2_nand3_1 _18724_ (.B(_11851_),
    .C(_11895_),
    .A(net204),
    .Y(_11896_));
 sg13g2_o21ai_1 _18725_ (.B1(_11896_),
    .Y(_11897_),
    .A1(net204),
    .A2(_11894_));
 sg13g2_nand3_1 _18726_ (.B(_11846_),
    .C(_11897_),
    .A(_11844_),
    .Y(_11898_));
 sg13g2_nor2b_1 _18727_ (.A(_11891_),
    .B_N(_11898_),
    .Y(_11899_));
 sg13g2_xnor2_1 _18728_ (.Y(_11900_),
    .A(net171),
    .B(_11899_));
 sg13g2_nor2_1 _18729_ (.A(net100),
    .B(net62),
    .Y(_11901_));
 sg13g2_nand2_1 _18730_ (.Y(_11902_),
    .A(_11900_),
    .B(_11901_));
 sg13g2_buf_2 _18731_ (.A(_00168_),
    .X(_11903_));
 sg13g2_nor2_1 _18732_ (.A(net441),
    .B(_11792_),
    .Y(_11904_));
 sg13g2_nor2_1 _18733_ (.A(_11800_),
    .B(_11904_),
    .Y(_11905_));
 sg13g2_nor2_1 _18734_ (.A(_11903_),
    .B(_11905_),
    .Y(_11906_));
 sg13g2_nor2_1 _18735_ (.A(_11903_),
    .B(net532),
    .Y(_11907_));
 sg13g2_nor3_1 _18736_ (.A(net100),
    .B(_11792_),
    .C(_11907_),
    .Y(_11908_));
 sg13g2_and2_1 _18737_ (.A(\cpu.ex.r_mult[12] ),
    .B(net278),
    .X(_11909_));
 sg13g2_a21o_1 _18738_ (.A2(_11908_),
    .A1(_11900_),
    .B1(_11909_),
    .X(_11910_));
 sg13g2_a21o_1 _18739_ (.A2(_11906_),
    .A1(_11902_),
    .B1(_11910_),
    .X(\cpu.ex.c_mult[12] ));
 sg13g2_buf_1 _18740_ (.A(_00169_),
    .X(_11911_));
 sg13g2_inv_1 _18741_ (.Y(_11912_),
    .A(_11911_));
 sg13g2_a22oi_1 _18742_ (.Y(_11913_),
    .B1(_11801_),
    .B2(_11912_),
    .A2(_10366_),
    .A1(\cpu.ex.r_mult[13] ));
 sg13g2_buf_1 _18743_ (.A(_10567_),
    .X(_11914_));
 sg13g2_inv_1 _18744_ (.Y(_11915_),
    .A(_11903_));
 sg13g2_o21ai_1 _18745_ (.B1(_11889_),
    .Y(_11916_),
    .A1(_11915_),
    .A2(_11886_));
 sg13g2_nand2_1 _18746_ (.Y(_11917_),
    .A(_11915_),
    .B(_11886_));
 sg13g2_a21oi_2 _18747_ (.B1(net490),
    .Y(_11918_),
    .A2(_11917_),
    .A1(_11916_));
 sg13g2_inv_1 _18748_ (.Y(_11919_),
    .A(_11918_));
 sg13g2_nor2_1 _18749_ (.A(_11911_),
    .B(net629),
    .Y(_11920_));
 sg13g2_nor2_1 _18750_ (.A(_11792_),
    .B(_11920_),
    .Y(_11921_));
 sg13g2_nand4_1 _18751_ (.B(net88),
    .C(_11919_),
    .A(net145),
    .Y(_11922_),
    .D(_11921_));
 sg13g2_nand2_1 _18752_ (.Y(_11923_),
    .A(_08631_),
    .B(net1030));
 sg13g2_o21ai_1 _18753_ (.B1(_11923_),
    .Y(_11924_),
    .A1(_10535_),
    .A2(_10564_));
 sg13g2_buf_1 _18754_ (.A(_11924_),
    .X(_11925_));
 sg13g2_buf_1 _18755_ (.A(net199),
    .X(_11926_));
 sg13g2_nand2_1 _18756_ (.Y(_11927_),
    .A(_11912_),
    .B(net533));
 sg13g2_nor2_1 _18757_ (.A(_11792_),
    .B(_11927_),
    .Y(_11928_));
 sg13g2_nand3_1 _18758_ (.B(_11919_),
    .C(_11928_),
    .A(net169),
    .Y(_11929_));
 sg13g2_and2_1 _18759_ (.A(net102),
    .B(_11846_),
    .X(_11930_));
 sg13g2_o21ai_1 _18760_ (.B1(_11930_),
    .Y(_11931_),
    .A1(_11831_),
    .A2(_11832_));
 sg13g2_nand3b_1 _18761_ (.B(_11857_),
    .C(_11931_),
    .Y(_11932_),
    .A_N(_11842_));
 sg13g2_nor2_1 _18762_ (.A(net170),
    .B(_10575_),
    .Y(_11933_));
 sg13g2_or2_1 _18763_ (.X(_11934_),
    .B(_11933_),
    .A(_11702_));
 sg13g2_nor3_1 _18764_ (.A(_11881_),
    .B(_11903_),
    .C(net490),
    .Y(_11935_));
 sg13g2_mux2_1 _18765_ (.A0(_11903_),
    .A1(_11907_),
    .S(net176),
    .X(_11936_));
 sg13g2_a22oi_1 _18766_ (.Y(_11937_),
    .B1(_11936_),
    .B2(_11881_),
    .A2(net171),
    .A1(net490));
 sg13g2_nand4_1 _18767_ (.B(net147),
    .C(net171),
    .A(_11903_),
    .Y(_11938_),
    .D(_11882_));
 sg13g2_o21ai_1 _18768_ (.B1(_11938_),
    .Y(_11939_),
    .A1(net147),
    .A2(_11937_));
 sg13g2_a22oi_1 _18769_ (.Y(_11940_),
    .B1(_11939_),
    .B2(net102),
    .A2(_11935_),
    .A1(_11934_));
 sg13g2_nor2_1 _18770_ (.A(net174),
    .B(_11940_),
    .Y(_11941_));
 sg13g2_nor3_1 _18771_ (.A(_11831_),
    .B(_11832_),
    .C(_11842_),
    .Y(_11942_));
 sg13g2_a21oi_1 _18772_ (.A1(_11644_),
    .A2(net102),
    .Y(_11943_),
    .B1(_11824_));
 sg13g2_nor4_1 _18773_ (.A(_11942_),
    .B(_11857_),
    .C(_11940_),
    .D(_11943_),
    .Y(_11944_));
 sg13g2_a21o_1 _18774_ (.A2(_11941_),
    .A1(_11932_),
    .B1(_11944_),
    .X(_11945_));
 sg13g2_a21o_1 _18775_ (.A2(_11929_),
    .A1(_11922_),
    .B1(_11945_),
    .X(_11946_));
 sg13g2_and2_1 _18776_ (.A(_11926_),
    .B(_11921_),
    .X(_11947_));
 sg13g2_and2_1 _18777_ (.A(net88),
    .B(_11947_),
    .X(_11948_));
 sg13g2_nor2b_1 _18778_ (.A(net169),
    .B_N(_11928_),
    .Y(_11949_));
 sg13g2_o21ai_1 _18779_ (.B1(_11945_),
    .Y(_11950_),
    .A1(_11948_),
    .A2(_11949_));
 sg13g2_and3_1 _18780_ (.X(_11951_),
    .A(net88),
    .B(_11918_),
    .C(_11947_));
 sg13g2_a221oi_1 _18781_ (.B2(_11918_),
    .C1(_11951_),
    .B1(_11949_),
    .A1(net100),
    .Y(_11952_),
    .A2(_11928_));
 sg13g2_nand4_1 _18782_ (.B(_11946_),
    .C(_11950_),
    .A(_11913_),
    .Y(_11953_),
    .D(_11952_));
 sg13g2_buf_1 _18783_ (.A(_11953_),
    .X(\cpu.ex.c_mult[13] ));
 sg13g2_buf_1 _18784_ (.A(_10616_),
    .X(_11954_));
 sg13g2_nand2_1 _18785_ (.Y(_11955_),
    .A(net199),
    .B(_11920_));
 sg13g2_o21ai_1 _18786_ (.B1(_11955_),
    .Y(_11956_),
    .A1(_11912_),
    .A2(net199));
 sg13g2_a22oi_1 _18787_ (.Y(_11957_),
    .B1(_11956_),
    .B2(_11903_),
    .A2(_10567_),
    .A1(net532));
 sg13g2_xnor2_1 _18788_ (.Y(_11958_),
    .A(_11912_),
    .B(net199));
 sg13g2_nand3_1 _18789_ (.B(_11907_),
    .C(_11958_),
    .A(net176),
    .Y(_11959_));
 sg13g2_o21ai_1 _18790_ (.B1(_11959_),
    .Y(_11960_),
    .A1(net176),
    .A2(_11957_));
 sg13g2_and3_1 _18791_ (.X(_11961_),
    .A(_11846_),
    .B(_11897_),
    .C(_11960_));
 sg13g2_nor3_1 _18792_ (.A(net532),
    .B(net176),
    .C(_11890_),
    .Y(_11962_));
 sg13g2_o21ai_1 _18793_ (.B1(_11920_),
    .Y(_11963_),
    .A1(net175),
    .A2(_11962_));
 sg13g2_o21ai_1 _18794_ (.B1(net176),
    .Y(_11964_),
    .A1(net532),
    .A2(_11890_));
 sg13g2_a221oi_1 _18795_ (.B2(_11911_),
    .C1(_11903_),
    .B1(net199),
    .A1(_09455_),
    .Y(_11965_),
    .A2(_09459_));
 sg13g2_a22oi_1 _18796_ (.Y(_11966_),
    .B1(_11964_),
    .B2(_11965_),
    .A2(_11962_),
    .A1(net175));
 sg13g2_nand2_1 _18797_ (.Y(_11967_),
    .A(_11963_),
    .B(_11966_));
 sg13g2_a21oi_1 _18798_ (.A1(_11844_),
    .A2(_11961_),
    .Y(_11968_),
    .B1(_11967_));
 sg13g2_xnor2_1 _18799_ (.Y(_11969_),
    .A(net116),
    .B(_11968_));
 sg13g2_buf_2 _18800_ (.A(_00170_),
    .X(_11970_));
 sg13g2_inv_1 _18801_ (.Y(_11971_),
    .A(_11970_));
 sg13g2_nand2_1 _18802_ (.Y(_11972_),
    .A(_11971_),
    .B(net628));
 sg13g2_nand4_1 _18803_ (.B(_11839_),
    .C(_11969_),
    .A(net70),
    .Y(_11973_),
    .D(_11972_));
 sg13g2_nor2_1 _18804_ (.A(_11970_),
    .B(net532),
    .Y(_11974_));
 sg13g2_nand2_1 _18805_ (.Y(_11975_),
    .A(_11839_),
    .B(_11974_));
 sg13g2_a21o_1 _18806_ (.A2(_11969_),
    .A1(_11663_),
    .B1(_11975_),
    .X(_11976_));
 sg13g2_a22oi_1 _18807_ (.Y(_11977_),
    .B1(_11801_),
    .B2(_11971_),
    .A2(net278),
    .A1(\cpu.ex.r_mult[14] ));
 sg13g2_nand3_1 _18808_ (.B(_11976_),
    .C(_11977_),
    .A(_11973_),
    .Y(_11978_));
 sg13g2_buf_1 _18809_ (.A(_11978_),
    .X(\cpu.ex.c_mult[14] ));
 sg13g2_nand2_1 _18810_ (.Y(_11979_),
    .A(\cpu.ex.r_mult[15] ),
    .B(net278));
 sg13g2_nor2_1 _18811_ (.A(_11861_),
    .B(_11877_),
    .Y(_11980_));
 sg13g2_o21ai_1 _18812_ (.B1(net102),
    .Y(_11981_),
    .A1(net175),
    .A2(net116));
 sg13g2_nor2_1 _18813_ (.A(_11970_),
    .B(_11927_),
    .Y(_11982_));
 sg13g2_mux2_1 _18814_ (.A0(_11970_),
    .A1(_11974_),
    .S(net146),
    .X(_11983_));
 sg13g2_a22oi_1 _18815_ (.Y(_11984_),
    .B1(_11983_),
    .B2(_11911_),
    .A2(net116),
    .A1(net490));
 sg13g2_nand4_1 _18816_ (.B(net199),
    .C(net116),
    .A(_11970_),
    .Y(_11985_),
    .D(_11920_));
 sg13g2_o21ai_1 _18817_ (.B1(_11985_),
    .Y(_11986_),
    .A1(net199),
    .A2(_11984_));
 sg13g2_a22oi_1 _18818_ (.Y(_11987_),
    .B1(_11986_),
    .B2(net102),
    .A2(_11982_),
    .A1(_11981_));
 sg13g2_or2_1 _18819_ (.X(_11988_),
    .B(_11987_),
    .A(_11940_));
 sg13g2_nor2_1 _18820_ (.A(_11926_),
    .B(_11919_),
    .Y(_11989_));
 sg13g2_a21oi_1 _18821_ (.A1(net145),
    .A2(_11918_),
    .Y(_11990_),
    .B1(net116));
 sg13g2_a21oi_1 _18822_ (.A1(_11970_),
    .A2(net146),
    .Y(_11991_),
    .B1(_11911_));
 sg13g2_o21ai_1 _18823_ (.B1(_11991_),
    .Y(_11992_),
    .A1(_11914_),
    .A2(_11918_));
 sg13g2_o21ai_1 _18824_ (.B1(_11992_),
    .Y(_11993_),
    .A1(_11970_),
    .A2(_11990_));
 sg13g2_a22oi_1 _18825_ (.Y(_11994_),
    .B1(_11993_),
    .B2(net533),
    .A2(_11989_),
    .A1(net116));
 sg13g2_o21ai_1 _18826_ (.B1(_11994_),
    .Y(_11995_),
    .A1(_11980_),
    .A2(_11988_));
 sg13g2_xnor2_1 _18827_ (.Y(_11996_),
    .A(_11634_),
    .B(_11995_));
 sg13g2_buf_1 _18828_ (.A(_00171_),
    .X(_11997_));
 sg13g2_nor2_1 _18829_ (.A(_11997_),
    .B(net490),
    .Y(_11998_));
 sg13g2_inv_1 _18830_ (.Y(_11999_),
    .A(_11998_));
 sg13g2_nand4_1 _18831_ (.B(_11839_),
    .C(_11996_),
    .A(_11663_),
    .Y(_12000_),
    .D(_11999_));
 sg13g2_or2_1 _18832_ (.X(_12001_),
    .B(_11905_),
    .A(_11997_));
 sg13g2_a21o_1 _18833_ (.A2(_11996_),
    .A1(_11901_),
    .B1(_12001_),
    .X(_12002_));
 sg13g2_nand3_1 _18834_ (.B(_12000_),
    .C(_12002_),
    .A(_11979_),
    .Y(\cpu.ex.c_mult[15] ));
 sg13g2_inv_1 _18835_ (.Y(_00000_),
    .A(net2));
 sg13g2_buf_2 _18836_ (.A(\cpu.qspi.r_state[13] ),
    .X(_12003_));
 sg13g2_buf_1 _18837_ (.A(net803),
    .X(_12004_));
 sg13g2_and2_1 _18838_ (.A(_12003_),
    .B(net667),
    .X(_00006_));
 sg13g2_nor3_1 _18839_ (.A(_09447_),
    .B(_09982_),
    .C(_09983_),
    .Y(_00007_));
 sg13g2_inv_1 _18840_ (.Y(_12005_),
    .A(_09954_));
 sg13g2_nor3_1 _18841_ (.A(_12005_),
    .B(_09447_),
    .C(_09957_),
    .Y(_00008_));
 sg13g2_buf_1 _18842_ (.A(\cpu.qspi.r_state[11] ),
    .X(_12006_));
 sg13g2_inv_1 _18843_ (.Y(_12007_),
    .A(_12006_));
 sg13g2_nor2_1 _18844_ (.A(_12007_),
    .B(net631),
    .Y(_00004_));
 sg13g2_buf_2 _18845_ (.A(\cpu.qspi.r_state[10] ),
    .X(_12008_));
 sg13g2_and2_1 _18846_ (.A(_12008_),
    .B(net706),
    .X(_00003_));
 sg13g2_buf_2 _18847_ (.A(\cpu.qspi.r_state[15] ),
    .X(_12009_));
 sg13g2_and2_1 _18848_ (.A(_12009_),
    .B(net706),
    .X(_00002_));
 sg13g2_inv_1 _18849_ (.Y(_12010_),
    .A(_09950_));
 sg13g2_nor3_1 _18850_ (.A(_12010_),
    .B(net705),
    .C(net788),
    .Y(_00001_));
 sg13g2_and2_1 _18851_ (.A(_11457_),
    .B(_11480_),
    .X(_12011_));
 sg13g2_or4_1 _18852_ (.A(_11427_),
    .B(_11378_),
    .C(_11398_),
    .D(_11557_),
    .X(_12012_));
 sg13g2_nand2b_1 _18853_ (.Y(_12013_),
    .B(_11333_),
    .A_N(_11288_));
 sg13g2_nor4_1 _18854_ (.A(_12011_),
    .B(_11311_),
    .C(_12012_),
    .D(_12013_),
    .Y(_12014_));
 sg13g2_nand4_1 _18855_ (.B(_11237_),
    .C(_11263_),
    .A(_11121_),
    .Y(_12015_),
    .D(_11352_));
 sg13g2_nor4_1 _18856_ (.A(_11452_),
    .B(_11502_),
    .C(_11523_),
    .D(_12015_),
    .Y(_12016_));
 sg13g2_a21oi_1 _18857_ (.A1(_12014_),
    .A2(_12016_),
    .Y(_12017_),
    .B1(\cpu.cond[1] ));
 sg13g2_nor2_1 _18858_ (.A(_11189_),
    .B(_12017_),
    .Y(_12018_));
 sg13g2_xnor2_1 _18859_ (.Y(_12019_),
    .A(_08499_),
    .B(_12018_));
 sg13g2_a21o_1 _18860_ (.A2(_12019_),
    .A1(_11126_),
    .B1(_11137_),
    .X(_12020_));
 sg13g2_nor2b_1 _18861_ (.A(\cpu.dec.jmp ),
    .B_N(_12020_),
    .Y(_12021_));
 sg13g2_buf_1 _18862_ (.A(_09459_),
    .X(_12022_));
 sg13g2_nor2b_1 _18863_ (.A(_12021_),
    .B_N(_12022_),
    .Y(_00053_));
 sg13g2_buf_2 _18864_ (.A(\cpu.qspi.r_state[3] ),
    .X(_12023_));
 sg13g2_and2_1 _18865_ (.A(_12023_),
    .B(net706),
    .X(_00009_));
 sg13g2_buf_2 _18866_ (.A(\cpu.qspi.r_state[6] ),
    .X(_12024_));
 sg13g2_and2_1 _18867_ (.A(_12024_),
    .B(net706),
    .X(_00010_));
 sg13g2_and3_1 _18868_ (.X(_00005_),
    .A(net1047),
    .B(net706),
    .C(_09946_));
 sg13g2_and2_1 _18869_ (.A(net120),
    .B(_09445_),
    .X(_00052_));
 sg13g2_o21ai_1 _18870_ (.B1(net497),
    .Y(_12025_),
    .A1(net1050),
    .A2(net1123));
 sg13g2_inv_1 _18871_ (.Y(_12026_),
    .A(_09377_));
 sg13g2_nor3_1 _18872_ (.A(_09429_),
    .B(_09440_),
    .C(_09436_),
    .Y(_12027_));
 sg13g2_nand2_1 _18873_ (.Y(_12028_),
    .A(_12026_),
    .B(_12027_));
 sg13g2_nand3_1 _18874_ (.B(_12025_),
    .C(_12028_),
    .A(_09387_),
    .Y(_12029_));
 sg13g2_buf_1 _18875_ (.A(_12029_),
    .X(_12030_));
 sg13g2_inv_1 _18876_ (.Y(_12031_),
    .A(_00226_));
 sg13g2_nor3_2 _18877_ (.A(net1123),
    .B(_09436_),
    .C(_12031_),
    .Y(_12032_));
 sg13g2_buf_1 _18878_ (.A(\cpu.spi.r_sel[1] ),
    .X(_12033_));
 sg13g2_buf_1 _18879_ (.A(_12033_),
    .X(_12034_));
 sg13g2_buf_1 _18880_ (.A(\cpu.spi.r_src[2] ),
    .X(_12035_));
 sg13g2_inv_1 _18881_ (.Y(_12036_),
    .A(_00282_));
 sg13g2_buf_1 _18882_ (.A(\cpu.spi.r_sel[0] ),
    .X(_12037_));
 sg13g2_buf_1 _18883_ (.A(_12037_),
    .X(_12038_));
 sg13g2_mux2_1 _18884_ (.A0(_12035_),
    .A1(_12036_),
    .S(_12038_),
    .X(_12039_));
 sg13g2_buf_1 _18885_ (.A(_12033_),
    .X(_12040_));
 sg13g2_buf_1 _18886_ (.A(_12037_),
    .X(_12041_));
 sg13g2_nand2_1 _18887_ (.Y(_12042_),
    .A(_12041_),
    .B(_00283_));
 sg13g2_o21ai_1 _18888_ (.B1(_12042_),
    .Y(_12043_),
    .A1(net1012),
    .A2(_12036_));
 sg13g2_nor2_1 _18889_ (.A(_12040_),
    .B(_12043_),
    .Y(_12044_));
 sg13g2_a21oi_2 _18890_ (.B1(_12044_),
    .Y(_12045_),
    .A2(_12039_),
    .A1(net1015));
 sg13g2_nor2_1 _18891_ (.A(_12032_),
    .B(_12045_),
    .Y(_12046_));
 sg13g2_nor2_1 _18892_ (.A(net1050),
    .B(_09436_),
    .Y(_12047_));
 sg13g2_inv_1 _18893_ (.Y(_12048_),
    .A(_12033_));
 sg13g2_buf_1 _18894_ (.A(\cpu.spi.r_mode[0][1] ),
    .X(_12049_));
 sg13g2_buf_1 _18895_ (.A(\cpu.spi.r_mode[1][1] ),
    .X(_12050_));
 sg13g2_buf_1 _18896_ (.A(_12041_),
    .X(_12051_));
 sg13g2_mux2_1 _18897_ (.A0(_12049_),
    .A1(_12050_),
    .S(net900),
    .X(_12052_));
 sg13g2_nor2_1 _18898_ (.A(_12048_),
    .B(_12037_),
    .Y(_12053_));
 sg13g2_buf_1 _18899_ (.A(\cpu.spi.r_mode[2][1] ),
    .X(_12054_));
 sg13g2_a22oi_1 _18900_ (.Y(_12055_),
    .B1(_12053_),
    .B2(_12054_),
    .A2(_12052_),
    .A1(_12048_));
 sg13g2_xnor2_1 _18901_ (.Y(_12056_),
    .A(_12047_),
    .B(_12055_));
 sg13g2_buf_1 _18902_ (.A(net1042),
    .X(_12057_));
 sg13g2_buf_2 _18903_ (.A(net899),
    .X(_12058_));
 sg13g2_buf_1 _18904_ (.A(net785),
    .X(_12059_));
 sg13g2_nand2_1 _18905_ (.Y(_12060_),
    .A(net785),
    .B(_00283_));
 sg13g2_o21ai_1 _18906_ (.B1(_12060_),
    .Y(_12061_),
    .A1(_12059_),
    .A2(_12036_));
 sg13g2_buf_1 _18907_ (.A(_09495_),
    .X(_12062_));
 sg13g2_nand3_1 _18908_ (.B(net760),
    .C(_12035_),
    .A(net761),
    .Y(_12063_));
 sg13g2_o21ai_1 _18909_ (.B1(_12063_),
    .Y(_12064_),
    .A1(net761),
    .A2(_12061_));
 sg13g2_and2_1 _18910_ (.A(_12032_),
    .B(_12064_),
    .X(_12065_));
 sg13g2_buf_1 _18911_ (.A(net761),
    .X(_12066_));
 sg13g2_buf_1 _18912_ (.A(net665),
    .X(_12067_));
 sg13g2_buf_1 _18913_ (.A(net665),
    .X(_12068_));
 sg13g2_nand2b_1 _18914_ (.Y(_12069_),
    .B(_12068_),
    .A_N(_12049_));
 sg13g2_o21ai_1 _18915_ (.B1(_12069_),
    .Y(_12070_),
    .A1(_12067_),
    .A2(_12054_));
 sg13g2_mux2_1 _18916_ (.A0(_12049_),
    .A1(_12050_),
    .S(_12068_),
    .X(_12071_));
 sg13g2_nor2_1 _18917_ (.A(net664),
    .B(_12071_),
    .Y(_12072_));
 sg13g2_a21oi_1 _18918_ (.A1(net664),
    .A2(_12070_),
    .Y(_12073_),
    .B1(_12072_));
 sg13g2_a22oi_1 _18919_ (.Y(_12074_),
    .B1(_12065_),
    .B2(_12073_),
    .A2(_12056_),
    .A1(_12046_));
 sg13g2_nor2_1 _18920_ (.A(_12046_),
    .B(_12065_),
    .Y(_12075_));
 sg13g2_buf_1 _18921_ (.A(\cpu.gpio.genblk1[3].srcs_o[5] ),
    .X(_12076_));
 sg13g2_o21ai_1 _18922_ (.B1(net1105),
    .Y(_12077_),
    .A1(_12030_),
    .A2(_12075_));
 sg13g2_o21ai_1 _18923_ (.B1(_12077_),
    .Y(_00318_),
    .A1(_12030_),
    .A2(_12074_));
 sg13g2_nor2b_1 _18924_ (.A(_12030_),
    .B_N(_12075_),
    .Y(_12078_));
 sg13g2_or3_1 _18925_ (.A(net1123),
    .B(_09436_),
    .C(_12031_),
    .X(_12079_));
 sg13g2_buf_1 _18926_ (.A(_12079_),
    .X(_12080_));
 sg13g2_and2_1 _18927_ (.A(_12032_),
    .B(_12073_),
    .X(_12081_));
 sg13g2_a21oi_1 _18928_ (.A1(net898),
    .A2(_12056_),
    .Y(_12082_),
    .B1(_12081_));
 sg13g2_buf_1 _18929_ (.A(\cpu.gpio.genblk1[3].srcs_o[4] ),
    .X(_12083_));
 sg13g2_nor2_1 _18930_ (.A(net1104),
    .B(_12078_),
    .Y(_12084_));
 sg13g2_a21oi_1 _18931_ (.A1(_12078_),
    .A2(_12082_),
    .Y(_00319_),
    .B1(_12084_));
 sg13g2_buf_1 _18932_ (.A(\cpu.gpio.genblk1[3].srcs_o[3] ),
    .X(_12085_));
 sg13g2_mux2_1 _18933_ (.A0(\cpu.spi.r_out[7] ),
    .A1(_10229_),
    .S(_09432_),
    .X(_12086_));
 sg13g2_inv_1 _18934_ (.Y(_12087_),
    .A(_00224_));
 sg13g2_mux2_1 _18935_ (.A0(_12087_),
    .A1(\cpu.spi.r_mode[1][0] ),
    .S(_12037_),
    .X(_12088_));
 sg13g2_a22oi_1 _18936_ (.Y(_12089_),
    .B1(_12088_),
    .B2(_12048_),
    .A2(_12053_),
    .A1(\cpu.spi.r_mode[2][0] ));
 sg13g2_buf_1 _18937_ (.A(_12089_),
    .X(_12090_));
 sg13g2_and2_1 _18938_ (.A(_09393_),
    .B(_12090_),
    .X(_12091_));
 sg13g2_a21oi_1 _18939_ (.A1(_00221_),
    .A2(_09397_),
    .Y(_12092_),
    .B1(net1123));
 sg13g2_o21ai_1 _18940_ (.B1(net1123),
    .Y(_12093_),
    .A1(net497),
    .A2(_12090_));
 sg13g2_a22oi_1 _18941_ (.Y(_12094_),
    .B1(_12093_),
    .B2(_09437_),
    .A2(_12092_),
    .A1(_12091_));
 sg13g2_nand2b_1 _18942_ (.Y(_12095_),
    .B(net930),
    .A_N(_12094_));
 sg13g2_buf_1 _18943_ (.A(_12090_),
    .X(_12096_));
 sg13g2_nand3_1 _18944_ (.B(_09434_),
    .C(net608),
    .A(_09365_),
    .Y(_12097_));
 sg13g2_o21ai_1 _18945_ (.B1(_12097_),
    .Y(_12098_),
    .A1(net1124),
    .A2(_12027_));
 sg13g2_nand2b_1 _18946_ (.Y(_12099_),
    .B(_12098_),
    .A_N(_12095_));
 sg13g2_nor2_1 _18947_ (.A(_12045_),
    .B(_12099_),
    .Y(_12100_));
 sg13g2_mux2_1 _18948_ (.A0(net1103),
    .A1(_12086_),
    .S(_12100_),
    .X(_00320_));
 sg13g2_buf_1 _18949_ (.A(\cpu.gpio.genblk1[3].srcs_o[2] ),
    .X(_12101_));
 sg13g2_inv_1 _18950_ (.Y(_12102_),
    .A(_12045_));
 sg13g2_nor2_1 _18951_ (.A(_12102_),
    .B(_12099_),
    .Y(_12103_));
 sg13g2_mux2_1 _18952_ (.A0(net1102),
    .A1(_12086_),
    .S(_12103_),
    .X(_00321_));
 sg13g2_nand2_1 _18953_ (.Y(_12104_),
    .A(net806),
    .B(_09523_));
 sg13g2_buf_2 _18954_ (.A(\cpu.dcache.r_offset[2] ),
    .X(_12105_));
 sg13g2_buf_2 _18955_ (.A(\cpu.dcache.r_offset[1] ),
    .X(_12106_));
 sg13g2_and2_1 _18956_ (.A(_12106_),
    .B(\cpu.dcache.r_offset[0] ),
    .X(_12107_));
 sg13g2_buf_1 _18957_ (.A(_12107_),
    .X(_12108_));
 sg13g2_nand3_1 _18958_ (.B(\cpu.d_wstrobe_d ),
    .C(_12108_),
    .A(_12105_),
    .Y(_12109_));
 sg13g2_buf_1 _18959_ (.A(_12109_),
    .X(_12110_));
 sg13g2_or3_1 _18960_ (.A(_09486_),
    .B(net957),
    .C(_09932_),
    .X(_12111_));
 sg13g2_buf_1 _18961_ (.A(_12111_),
    .X(_12112_));
 sg13g2_a21o_1 _18962_ (.A2(net663),
    .A1(_09924_),
    .B1(_12112_),
    .X(_12113_));
 sg13g2_buf_1 _18963_ (.A(_12113_),
    .X(_12114_));
 sg13g2_or2_1 _18964_ (.X(_12115_),
    .B(_12114_),
    .A(_12104_));
 sg13g2_buf_1 _18965_ (.A(_12115_),
    .X(_12116_));
 sg13g2_buf_1 _18966_ (.A(_08393_),
    .X(_12117_));
 sg13g2_nand2b_1 _18967_ (.Y(_12118_),
    .B(_08389_),
    .A_N(net1011));
 sg13g2_buf_2 _18968_ (.A(_12118_),
    .X(_12119_));
 sg13g2_buf_2 _18969_ (.A(_00275_),
    .X(_12120_));
 sg13g2_o21ai_1 _18970_ (.B1(_12120_),
    .Y(_12121_),
    .A1(_08390_),
    .A2(_12119_));
 sg13g2_nor2_1 _18971_ (.A(_12116_),
    .B(_12121_),
    .Y(_12122_));
 sg13g2_buf_2 _18972_ (.A(_12122_),
    .X(_12123_));
 sg13g2_buf_1 _18973_ (.A(_12123_),
    .X(_12124_));
 sg13g2_buf_1 _18974_ (.A(uio_in[0]),
    .X(_12125_));
 sg13g2_buf_1 _18975_ (.A(_12125_),
    .X(_12126_));
 sg13g2_buf_2 _18976_ (.A(net1101),
    .X(_12127_));
 sg13g2_buf_1 _18977_ (.A(_12104_),
    .X(_12128_));
 sg13g2_buf_1 _18978_ (.A(\cpu.d_wstrobe_d ),
    .X(_12129_));
 sg13g2_buf_1 _18979_ (.A(_00276_),
    .X(_12130_));
 sg13g2_buf_1 _18980_ (.A(_12130_),
    .X(_12131_));
 sg13g2_buf_1 _18981_ (.A(\cpu.dcache.r_offset[0] ),
    .X(_12132_));
 sg13g2_nor2b_1 _18982_ (.A(_12106_),
    .B_N(net1099),
    .Y(_12133_));
 sg13g2_buf_1 _18983_ (.A(_12133_),
    .X(_12134_));
 sg13g2_nand3_1 _18984_ (.B(net1009),
    .C(_12134_),
    .A(net1100),
    .Y(_12135_));
 sg13g2_buf_2 _18985_ (.A(_12135_),
    .X(_12136_));
 sg13g2_nor2_1 _18986_ (.A(net607),
    .B(_12136_),
    .Y(_12137_));
 sg13g2_buf_2 _18987_ (.A(_12137_),
    .X(_12138_));
 sg13g2_nor2b_1 _18988_ (.A(_12138_),
    .B_N(\cpu.dcache.r_data[0][0] ),
    .Y(_12139_));
 sg13g2_a21oi_1 _18989_ (.A1(net1010),
    .A2(_12138_),
    .Y(_12140_),
    .B1(_12139_));
 sg13g2_buf_1 _18990_ (.A(net1041),
    .X(_12141_));
 sg13g2_nand2_1 _18991_ (.Y(_12142_),
    .A(_12141_),
    .B(_12124_));
 sg13g2_o21ai_1 _18992_ (.B1(_12142_),
    .Y(_00322_),
    .A1(net61),
    .A2(_12140_));
 sg13g2_or2_1 _18993_ (.X(_12143_),
    .B(_12119_),
    .A(_08417_));
 sg13g2_buf_2 _18994_ (.A(_12143_),
    .X(_12144_));
 sg13g2_nor2_1 _18995_ (.A(_08417_),
    .B(_12119_),
    .Y(_12145_));
 sg13g2_buf_1 _18996_ (.A(_12145_),
    .X(_12146_));
 sg13g2_and2_1 _18997_ (.A(_10312_),
    .B(_12146_),
    .X(_12147_));
 sg13g2_a21oi_1 _18998_ (.A1(_10200_),
    .A2(_12144_),
    .Y(_12148_),
    .B1(_12147_));
 sg13g2_buf_2 _18999_ (.A(_12148_),
    .X(_12149_));
 sg13g2_buf_1 _19000_ (.A(_12149_),
    .X(_12150_));
 sg13g2_buf_1 _19001_ (.A(net787),
    .X(_12151_));
 sg13g2_inv_2 _19002_ (.Y(_12152_),
    .A(_12120_));
 sg13g2_mux2_1 _19003_ (.A0(net662),
    .A1(_12152_),
    .S(_08417_),
    .X(_12153_));
 sg13g2_or3_1 _19004_ (.A(_12116_),
    .B(_12119_),
    .C(_12153_),
    .X(_12154_));
 sg13g2_buf_1 _19005_ (.A(_12154_),
    .X(_12155_));
 sg13g2_buf_1 _19006_ (.A(_12155_),
    .X(_12156_));
 sg13g2_buf_1 _19007_ (.A(uio_in[2]),
    .X(_12157_));
 sg13g2_buf_1 _19008_ (.A(_12157_),
    .X(_12158_));
 sg13g2_nand3_1 _19009_ (.B(_12131_),
    .C(_12108_),
    .A(_12129_),
    .Y(_12159_));
 sg13g2_buf_4 _19010_ (.X(_12160_),
    .A(_12159_));
 sg13g2_nor2_2 _19011_ (.A(net607),
    .B(_12160_),
    .Y(_12161_));
 sg13g2_mux2_1 _19012_ (.A0(\cpu.dcache.r_data[0][10] ),
    .A1(net1098),
    .S(_12161_),
    .X(_12162_));
 sg13g2_nand2_1 _19013_ (.Y(_12163_),
    .A(net60),
    .B(_12162_));
 sg13g2_o21ai_1 _19014_ (.B1(_12163_),
    .Y(_00323_),
    .A1(net397),
    .A2(net60));
 sg13g2_and2_1 _19015_ (.A(_10319_),
    .B(_12146_),
    .X(_12164_));
 sg13g2_a21oi_1 _19016_ (.A1(net1116),
    .A2(_12144_),
    .Y(_12165_),
    .B1(_12164_));
 sg13g2_buf_2 _19017_ (.A(_12165_),
    .X(_12166_));
 sg13g2_buf_1 _19018_ (.A(_12166_),
    .X(_12167_));
 sg13g2_buf_1 _19019_ (.A(uio_in[3]),
    .X(_12168_));
 sg13g2_buf_1 _19020_ (.A(_12168_),
    .X(_12169_));
 sg13g2_mux2_1 _19021_ (.A0(\cpu.dcache.r_data[0][11] ),
    .A1(net1097),
    .S(_12161_),
    .X(_12170_));
 sg13g2_nand2_1 _19022_ (.Y(_12171_),
    .A(net60),
    .B(_12170_));
 sg13g2_o21ai_1 _19023_ (.B1(_12171_),
    .Y(_00324_),
    .A1(_12156_),
    .A2(net396));
 sg13g2_and2_1 _19024_ (.A(_10324_),
    .B(_12146_),
    .X(_12172_));
 sg13g2_a21oi_1 _19025_ (.A1(_10214_),
    .A2(_12144_),
    .Y(_12173_),
    .B1(_12172_));
 sg13g2_buf_2 _19026_ (.A(_12173_),
    .X(_12174_));
 sg13g2_buf_1 _19027_ (.A(_12174_),
    .X(_12175_));
 sg13g2_buf_1 _19028_ (.A(_12125_),
    .X(_12176_));
 sg13g2_buf_1 _19029_ (.A(_12132_),
    .X(_12177_));
 sg13g2_nor2b_1 _19030_ (.A(_12177_),
    .B_N(_12106_),
    .Y(_12178_));
 sg13g2_nand3_1 _19031_ (.B(net1009),
    .C(_12178_),
    .A(net1100),
    .Y(_12179_));
 sg13g2_buf_4 _19032_ (.X(_12180_),
    .A(_12179_));
 sg13g2_nor2_2 _19033_ (.A(net607),
    .B(_12180_),
    .Y(_12181_));
 sg13g2_mux2_1 _19034_ (.A0(\cpu.dcache.r_data[0][12] ),
    .A1(net1096),
    .S(_12181_),
    .X(_12182_));
 sg13g2_nand2_1 _19035_ (.Y(_12183_),
    .A(_12155_),
    .B(_12182_));
 sg13g2_o21ai_1 _19036_ (.B1(_12183_),
    .Y(_00325_),
    .A1(net60),
    .A2(net395));
 sg13g2_and2_1 _19037_ (.A(_10326_),
    .B(_12146_),
    .X(_12184_));
 sg13g2_a21oi_1 _19038_ (.A1(_10220_),
    .A2(_12144_),
    .Y(_12185_),
    .B1(_12184_));
 sg13g2_buf_2 _19039_ (.A(_12185_),
    .X(_12186_));
 sg13g2_buf_1 _19040_ (.A(_12186_),
    .X(_12187_));
 sg13g2_buf_1 _19041_ (.A(uio_in[1]),
    .X(_12188_));
 sg13g2_buf_1 _19042_ (.A(_12188_),
    .X(_12189_));
 sg13g2_mux2_1 _19043_ (.A0(\cpu.dcache.r_data[0][13] ),
    .A1(net1095),
    .S(_12181_),
    .X(_12190_));
 sg13g2_nand2_1 _19044_ (.Y(_12191_),
    .A(_12155_),
    .B(_12190_));
 sg13g2_o21ai_1 _19045_ (.B1(_12191_),
    .Y(_00326_),
    .A1(net60),
    .A2(net394));
 sg13g2_and2_1 _19046_ (.A(_10339_),
    .B(_12146_),
    .X(_12192_));
 sg13g2_a21oi_1 _19047_ (.A1(_10226_),
    .A2(_12144_),
    .Y(_12193_),
    .B1(_12192_));
 sg13g2_buf_2 _19048_ (.A(_12193_),
    .X(_12194_));
 sg13g2_buf_1 _19049_ (.A(_12194_),
    .X(_12195_));
 sg13g2_mux2_1 _19050_ (.A0(\cpu.dcache.r_data[0][14] ),
    .A1(net1098),
    .S(_12181_),
    .X(_12196_));
 sg13g2_nand2_1 _19051_ (.Y(_12197_),
    .A(_12155_),
    .B(_12196_));
 sg13g2_o21ai_1 _19052_ (.B1(_12197_),
    .Y(_00327_),
    .A1(net60),
    .A2(net393));
 sg13g2_and2_1 _19053_ (.A(_10344_),
    .B(_12146_),
    .X(_12198_));
 sg13g2_a21oi_1 _19054_ (.A1(_10229_),
    .A2(_12144_),
    .Y(_12199_),
    .B1(_12198_));
 sg13g2_buf_2 _19055_ (.A(_12199_),
    .X(_12200_));
 sg13g2_buf_1 _19056_ (.A(_12200_),
    .X(_12201_));
 sg13g2_mux2_1 _19057_ (.A0(\cpu.dcache.r_data[0][15] ),
    .A1(net1097),
    .S(_12181_),
    .X(_12202_));
 sg13g2_nand2_1 _19058_ (.Y(_12203_),
    .A(_12155_),
    .B(_12202_));
 sg13g2_o21ai_1 _19059_ (.B1(_12203_),
    .Y(_00328_),
    .A1(net60),
    .A2(net392));
 sg13g2_o21ai_1 _19060_ (.B1(net662),
    .Y(_12204_),
    .A1(_08390_),
    .A2(_12119_));
 sg13g2_nor2_1 _19061_ (.A(_12116_),
    .B(_12204_),
    .Y(_12205_));
 sg13g2_buf_2 _19062_ (.A(_12205_),
    .X(_12206_));
 sg13g2_buf_1 _19063_ (.A(_12206_),
    .X(_12207_));
 sg13g2_buf_1 _19064_ (.A(_12105_),
    .X(_12208_));
 sg13g2_nand3_1 _19065_ (.B(net1100),
    .C(_12134_),
    .A(net1007),
    .Y(_12209_));
 sg13g2_buf_2 _19066_ (.A(_12209_),
    .X(_12210_));
 sg13g2_nor2_1 _19067_ (.A(_12128_),
    .B(_12210_),
    .Y(_12211_));
 sg13g2_buf_2 _19068_ (.A(_12211_),
    .X(_12212_));
 sg13g2_nor2b_1 _19069_ (.A(_12212_),
    .B_N(\cpu.dcache.r_data[0][16] ),
    .Y(_12213_));
 sg13g2_a21oi_1 _19070_ (.A1(net1010),
    .A2(_12212_),
    .Y(_12214_),
    .B1(_12213_));
 sg13g2_buf_1 _19071_ (.A(_10187_),
    .X(_12215_));
 sg13g2_nand2_1 _19072_ (.Y(_12216_),
    .A(net896),
    .B(_12207_));
 sg13g2_o21ai_1 _19073_ (.B1(_12216_),
    .Y(_00329_),
    .A1(net59),
    .A2(_12214_));
 sg13g2_buf_1 _19074_ (.A(_12188_),
    .X(_12217_));
 sg13g2_buf_2 _19075_ (.A(net1094),
    .X(_12218_));
 sg13g2_nor2b_1 _19076_ (.A(_12212_),
    .B_N(\cpu.dcache.r_data[0][17] ),
    .Y(_12219_));
 sg13g2_a21oi_1 _19077_ (.A1(net1006),
    .A2(_12212_),
    .Y(_12220_),
    .B1(_12219_));
 sg13g2_nand2_1 _19078_ (.Y(_12221_),
    .A(net921),
    .B(net59));
 sg13g2_o21ai_1 _19079_ (.B1(_12221_),
    .Y(_00330_),
    .A1(net59),
    .A2(_12220_));
 sg13g2_buf_1 _19080_ (.A(_12157_),
    .X(_12222_));
 sg13g2_buf_2 _19081_ (.A(net1093),
    .X(_12223_));
 sg13g2_nor2b_1 _19082_ (.A(_12212_),
    .B_N(\cpu.dcache.r_data[0][18] ),
    .Y(_12224_));
 sg13g2_a21oi_1 _19083_ (.A1(net1005),
    .A2(_12212_),
    .Y(_12225_),
    .B1(_12224_));
 sg13g2_buf_1 _19084_ (.A(_10201_),
    .X(_12226_));
 sg13g2_nand2_1 _19085_ (.Y(_12227_),
    .A(_12226_),
    .B(_12206_));
 sg13g2_o21ai_1 _19086_ (.B1(_12227_),
    .Y(_00331_),
    .A1(_12207_),
    .A2(_12225_));
 sg13g2_buf_1 _19087_ (.A(_12168_),
    .X(_12228_));
 sg13g2_buf_2 _19088_ (.A(net1092),
    .X(_12229_));
 sg13g2_nor2b_1 _19089_ (.A(_12212_),
    .B_N(\cpu.dcache.r_data[0][19] ),
    .Y(_12230_));
 sg13g2_a21oi_1 _19090_ (.A1(net1004),
    .A2(_12212_),
    .Y(_12231_),
    .B1(_12230_));
 sg13g2_buf_1 _19091_ (.A(net1116),
    .X(_12232_));
 sg13g2_nand2_1 _19092_ (.Y(_12233_),
    .A(_12232_),
    .B(_12206_));
 sg13g2_o21ai_1 _19093_ (.B1(_12233_),
    .Y(_00332_),
    .A1(net59),
    .A2(_12231_));
 sg13g2_nor2b_1 _19094_ (.A(_12138_),
    .B_N(\cpu.dcache.r_data[0][1] ),
    .Y(_12234_));
 sg13g2_a21oi_1 _19095_ (.A1(net1006),
    .A2(_12138_),
    .Y(_12235_),
    .B1(_12234_));
 sg13g2_nand2_1 _19096_ (.Y(_12236_),
    .A(net921),
    .B(net61));
 sg13g2_o21ai_1 _19097_ (.B1(_12236_),
    .Y(_00333_),
    .A1(net61),
    .A2(_12235_));
 sg13g2_nor2_1 _19098_ (.A(_12106_),
    .B(_12132_),
    .Y(_12237_));
 sg13g2_nand3_1 _19099_ (.B(net1100),
    .C(_12237_),
    .A(net1007),
    .Y(_12238_));
 sg13g2_buf_2 _19100_ (.A(_12238_),
    .X(_12239_));
 sg13g2_nor2_1 _19101_ (.A(_12128_),
    .B(_12239_),
    .Y(_12240_));
 sg13g2_buf_2 _19102_ (.A(_12240_),
    .X(_12241_));
 sg13g2_nor2b_1 _19103_ (.A(_12241_),
    .B_N(\cpu.dcache.r_data[0][20] ),
    .Y(_12242_));
 sg13g2_a21oi_1 _19104_ (.A1(net1010),
    .A2(_12241_),
    .Y(_12243_),
    .B1(_12242_));
 sg13g2_buf_1 _19105_ (.A(_10214_),
    .X(_12244_));
 sg13g2_nand2_1 _19106_ (.Y(_12245_),
    .A(net1002),
    .B(_12206_));
 sg13g2_o21ai_1 _19107_ (.B1(_12245_),
    .Y(_00334_),
    .A1(net59),
    .A2(_12243_));
 sg13g2_nor2b_1 _19108_ (.A(_12241_),
    .B_N(\cpu.dcache.r_data[0][21] ),
    .Y(_12246_));
 sg13g2_a21oi_1 _19109_ (.A1(net1006),
    .A2(_12241_),
    .Y(_12247_),
    .B1(_12246_));
 sg13g2_buf_1 _19110_ (.A(_10220_),
    .X(_12248_));
 sg13g2_nand2_1 _19111_ (.Y(_12249_),
    .A(net1001),
    .B(_12206_));
 sg13g2_o21ai_1 _19112_ (.B1(_12249_),
    .Y(_00335_),
    .A1(net59),
    .A2(_12247_));
 sg13g2_nor2b_1 _19113_ (.A(_12241_),
    .B_N(\cpu.dcache.r_data[0][22] ),
    .Y(_12250_));
 sg13g2_a21oi_1 _19114_ (.A1(net1005),
    .A2(_12241_),
    .Y(_12251_),
    .B1(_12250_));
 sg13g2_buf_1 _19115_ (.A(_10226_),
    .X(_12252_));
 sg13g2_nand2_1 _19116_ (.Y(_12253_),
    .A(net1000),
    .B(_12206_));
 sg13g2_o21ai_1 _19117_ (.B1(_12253_),
    .Y(_00336_),
    .A1(net59),
    .A2(_12251_));
 sg13g2_nor2b_1 _19118_ (.A(_12241_),
    .B_N(\cpu.dcache.r_data[0][23] ),
    .Y(_12254_));
 sg13g2_a21oi_1 _19119_ (.A1(net1004),
    .A2(_12241_),
    .Y(_12255_),
    .B1(_12254_));
 sg13g2_buf_1 _19120_ (.A(_10229_),
    .X(_12256_));
 sg13g2_nand2_1 _19121_ (.Y(_12257_),
    .A(net999),
    .B(_12206_));
 sg13g2_o21ai_1 _19122_ (.B1(_12257_),
    .Y(_00337_),
    .A1(net59),
    .A2(_12255_));
 sg13g2_and2_1 _19123_ (.A(_10302_),
    .B(_12146_),
    .X(_12258_));
 sg13g2_a21oi_1 _19124_ (.A1(_10186_),
    .A2(_12144_),
    .Y(_12259_),
    .B1(_12258_));
 sg13g2_buf_2 _19125_ (.A(_12259_),
    .X(_12260_));
 sg13g2_buf_1 _19126_ (.A(_12260_),
    .X(_12261_));
 sg13g2_nor2_1 _19127_ (.A(_08390_),
    .B(net662),
    .Y(_12262_));
 sg13g2_nor2_1 _19128_ (.A(_08417_),
    .B(_12152_),
    .Y(_12263_));
 sg13g2_or4_1 _19129_ (.A(_12116_),
    .B(_12119_),
    .C(_12262_),
    .D(_12263_),
    .X(_12264_));
 sg13g2_buf_1 _19130_ (.A(_12264_),
    .X(_12265_));
 sg13g2_buf_1 _19131_ (.A(_12265_),
    .X(_12266_));
 sg13g2_or2_1 _19132_ (.X(_12267_),
    .B(net663),
    .A(net607));
 sg13g2_buf_1 _19133_ (.A(_12267_),
    .X(_12268_));
 sg13g2_buf_1 _19134_ (.A(_12268_),
    .X(_12269_));
 sg13g2_mux2_1 _19135_ (.A0(net1096),
    .A1(\cpu.dcache.r_data[0][24] ),
    .S(net440),
    .X(_12270_));
 sg13g2_nand2_1 _19136_ (.Y(_12271_),
    .A(net58),
    .B(_12270_));
 sg13g2_o21ai_1 _19137_ (.B1(_12271_),
    .Y(_00338_),
    .A1(net391),
    .A2(net58));
 sg13g2_and2_1 _19138_ (.A(_10307_),
    .B(_12146_),
    .X(_12272_));
 sg13g2_a21oi_1 _19139_ (.A1(_10194_),
    .A2(_12144_),
    .Y(_12273_),
    .B1(_12272_));
 sg13g2_buf_2 _19140_ (.A(_12273_),
    .X(_12274_));
 sg13g2_buf_1 _19141_ (.A(_12274_),
    .X(_12275_));
 sg13g2_mux2_1 _19142_ (.A0(net1095),
    .A1(\cpu.dcache.r_data[0][25] ),
    .S(net440),
    .X(_12276_));
 sg13g2_nand2_1 _19143_ (.Y(_12277_),
    .A(_12266_),
    .B(_12276_));
 sg13g2_o21ai_1 _19144_ (.B1(_12277_),
    .Y(_00339_),
    .A1(net58),
    .A2(net390));
 sg13g2_mux2_1 _19145_ (.A0(net1098),
    .A1(\cpu.dcache.r_data[0][26] ),
    .S(net440),
    .X(_12278_));
 sg13g2_nand2_1 _19146_ (.Y(_12279_),
    .A(_12265_),
    .B(_12278_));
 sg13g2_o21ai_1 _19147_ (.B1(_12279_),
    .Y(_00340_),
    .A1(net397),
    .A2(net58));
 sg13g2_mux2_1 _19148_ (.A0(net1097),
    .A1(\cpu.dcache.r_data[0][27] ),
    .S(_12268_),
    .X(_12280_));
 sg13g2_nand2_1 _19149_ (.Y(_12281_),
    .A(_12265_),
    .B(_12280_));
 sg13g2_o21ai_1 _19150_ (.B1(_12281_),
    .Y(_00341_),
    .A1(net396),
    .A2(_12266_));
 sg13g2_nand3_1 _19151_ (.B(net1100),
    .C(_12178_),
    .A(net1007),
    .Y(_12282_));
 sg13g2_buf_4 _19152_ (.X(_12283_),
    .A(_12282_));
 sg13g2_nor2_2 _19153_ (.A(net607),
    .B(_12283_),
    .Y(_12284_));
 sg13g2_mux2_1 _19154_ (.A0(\cpu.dcache.r_data[0][28] ),
    .A1(net1096),
    .S(_12284_),
    .X(_12285_));
 sg13g2_nand2_1 _19155_ (.Y(_12286_),
    .A(_12265_),
    .B(_12285_));
 sg13g2_o21ai_1 _19156_ (.B1(_12286_),
    .Y(_00342_),
    .A1(net395),
    .A2(net58));
 sg13g2_mux2_1 _19157_ (.A0(\cpu.dcache.r_data[0][29] ),
    .A1(net1095),
    .S(_12284_),
    .X(_12287_));
 sg13g2_nand2_1 _19158_ (.Y(_12288_),
    .A(_12265_),
    .B(_12287_));
 sg13g2_o21ai_1 _19159_ (.B1(_12288_),
    .Y(_00343_),
    .A1(net394),
    .A2(net58));
 sg13g2_nor2b_1 _19160_ (.A(_12138_),
    .B_N(\cpu.dcache.r_data[0][2] ),
    .Y(_12289_));
 sg13g2_a21oi_1 _19161_ (.A1(net1005),
    .A2(_12138_),
    .Y(_12290_),
    .B1(_12289_));
 sg13g2_nand2_1 _19162_ (.Y(_12291_),
    .A(net895),
    .B(_12123_));
 sg13g2_o21ai_1 _19163_ (.B1(_12291_),
    .Y(_00344_),
    .A1(_12124_),
    .A2(_12290_));
 sg13g2_mux2_1 _19164_ (.A0(\cpu.dcache.r_data[0][30] ),
    .A1(net1098),
    .S(_12284_),
    .X(_12292_));
 sg13g2_nand2_1 _19165_ (.Y(_12293_),
    .A(_12265_),
    .B(_12292_));
 sg13g2_o21ai_1 _19166_ (.B1(_12293_),
    .Y(_00345_),
    .A1(_12195_),
    .A2(net58));
 sg13g2_mux2_1 _19167_ (.A0(\cpu.dcache.r_data[0][31] ),
    .A1(net1097),
    .S(_12284_),
    .X(_12294_));
 sg13g2_nand2_1 _19168_ (.Y(_12295_),
    .A(_12265_),
    .B(_12294_));
 sg13g2_o21ai_1 _19169_ (.B1(_12295_),
    .Y(_00346_),
    .A1(net392),
    .A2(net58));
 sg13g2_nor2b_1 _19170_ (.A(_12138_),
    .B_N(\cpu.dcache.r_data[0][3] ),
    .Y(_12296_));
 sg13g2_a21oi_1 _19171_ (.A1(net1004),
    .A2(_12138_),
    .Y(_12297_),
    .B1(_12296_));
 sg13g2_nand2_1 _19172_ (.Y(_12298_),
    .A(net1003),
    .B(_12123_));
 sg13g2_o21ai_1 _19173_ (.B1(_12298_),
    .Y(_00347_),
    .A1(net61),
    .A2(_12297_));
 sg13g2_nand3_1 _19174_ (.B(net1009),
    .C(_12237_),
    .A(net1100),
    .Y(_12299_));
 sg13g2_buf_2 _19175_ (.A(_12299_),
    .X(_12300_));
 sg13g2_nor2_1 _19176_ (.A(net607),
    .B(_12300_),
    .Y(_12301_));
 sg13g2_buf_2 _19177_ (.A(_12301_),
    .X(_12302_));
 sg13g2_nor2b_1 _19178_ (.A(_12302_),
    .B_N(\cpu.dcache.r_data[0][4] ),
    .Y(_12303_));
 sg13g2_a21oi_1 _19179_ (.A1(net1010),
    .A2(_12302_),
    .Y(_12304_),
    .B1(_12303_));
 sg13g2_nand2_1 _19180_ (.Y(_12305_),
    .A(net1002),
    .B(_12123_));
 sg13g2_o21ai_1 _19181_ (.B1(_12305_),
    .Y(_00348_),
    .A1(net61),
    .A2(_12304_));
 sg13g2_nor2b_1 _19182_ (.A(_12302_),
    .B_N(\cpu.dcache.r_data[0][5] ),
    .Y(_12306_));
 sg13g2_a21oi_1 _19183_ (.A1(net1006),
    .A2(_12302_),
    .Y(_12307_),
    .B1(_12306_));
 sg13g2_nand2_1 _19184_ (.Y(_12308_),
    .A(net1001),
    .B(_12123_));
 sg13g2_o21ai_1 _19185_ (.B1(_12308_),
    .Y(_00349_),
    .A1(net61),
    .A2(_12307_));
 sg13g2_nor2b_1 _19186_ (.A(_12302_),
    .B_N(\cpu.dcache.r_data[0][6] ),
    .Y(_12309_));
 sg13g2_a21oi_1 _19187_ (.A1(net1005),
    .A2(_12302_),
    .Y(_12310_),
    .B1(_12309_));
 sg13g2_nand2_1 _19188_ (.Y(_12311_),
    .A(net1000),
    .B(_12123_));
 sg13g2_o21ai_1 _19189_ (.B1(_12311_),
    .Y(_00350_),
    .A1(net61),
    .A2(_12310_));
 sg13g2_nor2b_1 _19190_ (.A(_12302_),
    .B_N(\cpu.dcache.r_data[0][7] ),
    .Y(_12312_));
 sg13g2_a21oi_1 _19191_ (.A1(net1004),
    .A2(_12302_),
    .Y(_12313_),
    .B1(_12312_));
 sg13g2_nand2_1 _19192_ (.Y(_12314_),
    .A(net999),
    .B(_12123_));
 sg13g2_o21ai_1 _19193_ (.B1(_12314_),
    .Y(_00351_),
    .A1(net61),
    .A2(_12313_));
 sg13g2_mux2_1 _19194_ (.A0(\cpu.dcache.r_data[0][8] ),
    .A1(net1096),
    .S(_12161_),
    .X(_12315_));
 sg13g2_nand2_1 _19195_ (.Y(_12316_),
    .A(_12155_),
    .B(_12315_));
 sg13g2_o21ai_1 _19196_ (.B1(_12316_),
    .Y(_00352_),
    .A1(_12156_),
    .A2(net391));
 sg13g2_mux2_1 _19197_ (.A0(\cpu.dcache.r_data[0][9] ),
    .A1(net1095),
    .S(_12161_),
    .X(_12317_));
 sg13g2_nand2_1 _19198_ (.Y(_12318_),
    .A(_12155_),
    .B(_12317_));
 sg13g2_o21ai_1 _19199_ (.B1(_12318_),
    .Y(_00353_),
    .A1(net60),
    .A2(_12275_));
 sg13g2_buf_1 _19200_ (.A(_09531_),
    .X(_12319_));
 sg13g2_or2_1 _19201_ (.X(_12320_),
    .B(_12121_),
    .A(_12114_));
 sg13g2_buf_2 _19202_ (.A(_12320_),
    .X(_12321_));
 sg13g2_nor2_1 _19203_ (.A(net661),
    .B(_12321_),
    .Y(_12322_));
 sg13g2_buf_2 _19204_ (.A(_12322_),
    .X(_12323_));
 sg13g2_buf_1 _19205_ (.A(_12323_),
    .X(_12324_));
 sg13g2_nor2_1 _19206_ (.A(net661),
    .B(_12136_),
    .Y(_12325_));
 sg13g2_buf_2 _19207_ (.A(_12325_),
    .X(_12326_));
 sg13g2_nor2b_1 _19208_ (.A(_12326_),
    .B_N(\cpu.dcache.r_data[1][0] ),
    .Y(_12327_));
 sg13g2_a21oi_1 _19209_ (.A1(net1010),
    .A2(_12326_),
    .Y(_12328_),
    .B1(_12327_));
 sg13g2_nand2_1 _19210_ (.Y(_12329_),
    .A(net896),
    .B(net57));
 sg13g2_o21ai_1 _19211_ (.B1(_12329_),
    .Y(_00354_),
    .A1(net57),
    .A2(_12328_));
 sg13g2_buf_1 _19212_ (.A(net547),
    .X(_12330_));
 sg13g2_buf_1 _19213_ (.A(net489),
    .X(_12331_));
 sg13g2_buf_1 _19214_ (.A(_12331_),
    .X(_12332_));
 sg13g2_nor3_1 _19215_ (.A(_12114_),
    .B(_12119_),
    .C(_12153_),
    .Y(_12333_));
 sg13g2_buf_2 _19216_ (.A(_12333_),
    .X(_12334_));
 sg13g2_nand2_1 _19217_ (.Y(_12335_),
    .A(net389),
    .B(_12334_));
 sg13g2_buf_1 _19218_ (.A(_12335_),
    .X(_12336_));
 sg13g2_buf_1 _19219_ (.A(_12336_),
    .X(_12337_));
 sg13g2_nor2_2 _19220_ (.A(net661),
    .B(_12160_),
    .Y(_12338_));
 sg13g2_mux2_1 _19221_ (.A0(\cpu.dcache.r_data[1][10] ),
    .A1(net1098),
    .S(_12338_),
    .X(_12339_));
 sg13g2_nand2_1 _19222_ (.Y(_12340_),
    .A(_12337_),
    .B(_12339_));
 sg13g2_o21ai_1 _19223_ (.B1(_12340_),
    .Y(_00355_),
    .A1(_12150_),
    .A2(net56));
 sg13g2_mux2_1 _19224_ (.A0(\cpu.dcache.r_data[1][11] ),
    .A1(net1097),
    .S(_12338_),
    .X(_12341_));
 sg13g2_nand2_1 _19225_ (.Y(_12342_),
    .A(net56),
    .B(_12341_));
 sg13g2_o21ai_1 _19226_ (.B1(_12342_),
    .Y(_00356_),
    .A1(_12167_),
    .A2(_12337_));
 sg13g2_nor2_2 _19227_ (.A(net661),
    .B(_12180_),
    .Y(_12343_));
 sg13g2_mux2_1 _19228_ (.A0(\cpu.dcache.r_data[1][12] ),
    .A1(net1096),
    .S(_12343_),
    .X(_12344_));
 sg13g2_nand2_1 _19229_ (.Y(_12345_),
    .A(_12336_),
    .B(_12344_));
 sg13g2_o21ai_1 _19230_ (.B1(_12345_),
    .Y(_00357_),
    .A1(_12175_),
    .A2(net56));
 sg13g2_mux2_1 _19231_ (.A0(\cpu.dcache.r_data[1][13] ),
    .A1(net1095),
    .S(_12343_),
    .X(_12346_));
 sg13g2_nand2_1 _19232_ (.Y(_12347_),
    .A(_12336_),
    .B(_12346_));
 sg13g2_o21ai_1 _19233_ (.B1(_12347_),
    .Y(_00358_),
    .A1(_12187_),
    .A2(net56));
 sg13g2_buf_1 _19234_ (.A(_12157_),
    .X(_12348_));
 sg13g2_mux2_1 _19235_ (.A0(\cpu.dcache.r_data[1][14] ),
    .A1(_12348_),
    .S(_12343_),
    .X(_12349_));
 sg13g2_nand2_1 _19236_ (.Y(_12350_),
    .A(_12336_),
    .B(_12349_));
 sg13g2_o21ai_1 _19237_ (.B1(_12350_),
    .Y(_00359_),
    .A1(_12195_),
    .A2(net56));
 sg13g2_buf_1 _19238_ (.A(_12168_),
    .X(_12351_));
 sg13g2_mux2_1 _19239_ (.A0(\cpu.dcache.r_data[1][15] ),
    .A1(net1090),
    .S(_12343_),
    .X(_12352_));
 sg13g2_nand2_1 _19240_ (.Y(_12353_),
    .A(_12336_),
    .B(_12352_));
 sg13g2_o21ai_1 _19241_ (.B1(_12353_),
    .Y(_00360_),
    .A1(_12201_),
    .A2(net56));
 sg13g2_or2_1 _19242_ (.X(_12354_),
    .B(_12204_),
    .A(_12114_));
 sg13g2_buf_2 _19243_ (.A(_12354_),
    .X(_12355_));
 sg13g2_nor2_1 _19244_ (.A(net661),
    .B(_12355_),
    .Y(_12356_));
 sg13g2_buf_2 _19245_ (.A(_12356_),
    .X(_12357_));
 sg13g2_buf_1 _19246_ (.A(_12357_),
    .X(_12358_));
 sg13g2_nor2_1 _19247_ (.A(_12319_),
    .B(_12210_),
    .Y(_12359_));
 sg13g2_buf_2 _19248_ (.A(_12359_),
    .X(_12360_));
 sg13g2_nor2b_1 _19249_ (.A(_12360_),
    .B_N(\cpu.dcache.r_data[1][16] ),
    .Y(_12361_));
 sg13g2_a21oi_1 _19250_ (.A1(net1010),
    .A2(_12360_),
    .Y(_12362_),
    .B1(_12361_));
 sg13g2_nand2_1 _19251_ (.Y(_12363_),
    .A(net896),
    .B(net55));
 sg13g2_o21ai_1 _19252_ (.B1(_12363_),
    .Y(_00361_),
    .A1(net55),
    .A2(_12362_));
 sg13g2_nor2b_1 _19253_ (.A(_12360_),
    .B_N(\cpu.dcache.r_data[1][17] ),
    .Y(_12364_));
 sg13g2_a21oi_1 _19254_ (.A1(net1006),
    .A2(_12360_),
    .Y(_12365_),
    .B1(_12364_));
 sg13g2_nand2_1 _19255_ (.Y(_12366_),
    .A(net921),
    .B(net55));
 sg13g2_o21ai_1 _19256_ (.B1(_12366_),
    .Y(_00362_),
    .A1(net55),
    .A2(_12365_));
 sg13g2_nor2b_1 _19257_ (.A(_12360_),
    .B_N(\cpu.dcache.r_data[1][18] ),
    .Y(_12367_));
 sg13g2_a21oi_1 _19258_ (.A1(net1005),
    .A2(_12360_),
    .Y(_12368_),
    .B1(_12367_));
 sg13g2_nand2_1 _19259_ (.Y(_12369_),
    .A(_12226_),
    .B(_12357_));
 sg13g2_o21ai_1 _19260_ (.B1(_12369_),
    .Y(_00363_),
    .A1(net55),
    .A2(_12368_));
 sg13g2_nor2b_1 _19261_ (.A(_12360_),
    .B_N(\cpu.dcache.r_data[1][19] ),
    .Y(_12370_));
 sg13g2_a21oi_1 _19262_ (.A1(net1004),
    .A2(_12360_),
    .Y(_12371_),
    .B1(_12370_));
 sg13g2_nand2_1 _19263_ (.Y(_12372_),
    .A(net1003),
    .B(_12357_));
 sg13g2_o21ai_1 _19264_ (.B1(_12372_),
    .Y(_00364_),
    .A1(_12358_),
    .A2(_12371_));
 sg13g2_nor2b_1 _19265_ (.A(_12326_),
    .B_N(\cpu.dcache.r_data[1][1] ),
    .Y(_12373_));
 sg13g2_a21oi_1 _19266_ (.A1(net1006),
    .A2(_12326_),
    .Y(_12374_),
    .B1(_12373_));
 sg13g2_nand2_1 _19267_ (.Y(_12375_),
    .A(net921),
    .B(net57));
 sg13g2_o21ai_1 _19268_ (.B1(_12375_),
    .Y(_00365_),
    .A1(net57),
    .A2(_12374_));
 sg13g2_buf_1 _19269_ (.A(_12126_),
    .X(_12376_));
 sg13g2_nor2_1 _19270_ (.A(_12319_),
    .B(_12239_),
    .Y(_12377_));
 sg13g2_buf_2 _19271_ (.A(_12377_),
    .X(_12378_));
 sg13g2_nor2b_1 _19272_ (.A(_12378_),
    .B_N(\cpu.dcache.r_data[1][20] ),
    .Y(_12379_));
 sg13g2_a21oi_1 _19273_ (.A1(net998),
    .A2(_12378_),
    .Y(_12380_),
    .B1(_12379_));
 sg13g2_buf_1 _19274_ (.A(_10214_),
    .X(_12381_));
 sg13g2_nand2_1 _19275_ (.Y(_12382_),
    .A(_12381_),
    .B(_12357_));
 sg13g2_o21ai_1 _19276_ (.B1(_12382_),
    .Y(_00366_),
    .A1(_12358_),
    .A2(_12380_));
 sg13g2_buf_1 _19277_ (.A(_12217_),
    .X(_12383_));
 sg13g2_nor2b_1 _19278_ (.A(_12378_),
    .B_N(\cpu.dcache.r_data[1][21] ),
    .Y(_12384_));
 sg13g2_a21oi_1 _19279_ (.A1(net996),
    .A2(_12378_),
    .Y(_12385_),
    .B1(_12384_));
 sg13g2_buf_1 _19280_ (.A(_10220_),
    .X(_12386_));
 sg13g2_nand2_1 _19281_ (.Y(_12387_),
    .A(net995),
    .B(_12357_));
 sg13g2_o21ai_1 _19282_ (.B1(_12387_),
    .Y(_00367_),
    .A1(net55),
    .A2(_12385_));
 sg13g2_nor2b_1 _19283_ (.A(_12378_),
    .B_N(\cpu.dcache.r_data[1][22] ),
    .Y(_12388_));
 sg13g2_a21oi_1 _19284_ (.A1(net1005),
    .A2(_12378_),
    .Y(_12389_),
    .B1(_12388_));
 sg13g2_buf_1 _19285_ (.A(_10226_),
    .X(_12390_));
 sg13g2_nand2_1 _19286_ (.Y(_12391_),
    .A(net994),
    .B(_12357_));
 sg13g2_o21ai_1 _19287_ (.B1(_12391_),
    .Y(_00368_),
    .A1(net55),
    .A2(_12389_));
 sg13g2_nor2b_1 _19288_ (.A(_12378_),
    .B_N(\cpu.dcache.r_data[1][23] ),
    .Y(_12392_));
 sg13g2_a21oi_1 _19289_ (.A1(net1004),
    .A2(_12378_),
    .Y(_12393_),
    .B1(_12392_));
 sg13g2_nand2_1 _19290_ (.Y(_12394_),
    .A(net999),
    .B(_12357_));
 sg13g2_o21ai_1 _19291_ (.B1(_12394_),
    .Y(_00369_),
    .A1(net55),
    .A2(_12393_));
 sg13g2_nor4_1 _19292_ (.A(_12114_),
    .B(_12119_),
    .C(_12262_),
    .D(_12263_),
    .Y(_12395_));
 sg13g2_buf_2 _19293_ (.A(_12395_),
    .X(_12396_));
 sg13g2_nand2_1 _19294_ (.Y(_12397_),
    .A(net389),
    .B(_12396_));
 sg13g2_buf_2 _19295_ (.A(_12397_),
    .X(_12398_));
 sg13g2_buf_1 _19296_ (.A(_12398_),
    .X(_12399_));
 sg13g2_buf_1 _19297_ (.A(_12125_),
    .X(_12400_));
 sg13g2_nor2_1 _19298_ (.A(_09531_),
    .B(net663),
    .Y(_12401_));
 sg13g2_buf_2 _19299_ (.A(_12401_),
    .X(_12402_));
 sg13g2_mux2_1 _19300_ (.A0(\cpu.dcache.r_data[1][24] ),
    .A1(_12400_),
    .S(_12402_),
    .X(_12403_));
 sg13g2_nand2_1 _19301_ (.Y(_12404_),
    .A(net54),
    .B(_12403_));
 sg13g2_o21ai_1 _19302_ (.B1(_12404_),
    .Y(_00370_),
    .A1(net391),
    .A2(net54));
 sg13g2_buf_1 _19303_ (.A(_12188_),
    .X(_12405_));
 sg13g2_mux2_1 _19304_ (.A0(\cpu.dcache.r_data[1][25] ),
    .A1(net1088),
    .S(_12402_),
    .X(_12406_));
 sg13g2_nand2_1 _19305_ (.Y(_12407_),
    .A(net54),
    .B(_12406_));
 sg13g2_o21ai_1 _19306_ (.B1(_12407_),
    .Y(_00371_),
    .A1(_12275_),
    .A2(net54));
 sg13g2_mux2_1 _19307_ (.A0(\cpu.dcache.r_data[1][26] ),
    .A1(_12348_),
    .S(_12402_),
    .X(_12408_));
 sg13g2_nand2_1 _19308_ (.Y(_12409_),
    .A(_12398_),
    .B(_12408_));
 sg13g2_o21ai_1 _19309_ (.B1(_12409_),
    .Y(_00372_),
    .A1(_12150_),
    .A2(_12399_));
 sg13g2_mux2_1 _19310_ (.A0(\cpu.dcache.r_data[1][27] ),
    .A1(net1090),
    .S(_12402_),
    .X(_12410_));
 sg13g2_nand2_1 _19311_ (.Y(_12411_),
    .A(_12398_),
    .B(_12410_));
 sg13g2_o21ai_1 _19312_ (.B1(_12411_),
    .Y(_00373_),
    .A1(_12167_),
    .A2(_12399_));
 sg13g2_nor2_2 _19313_ (.A(net661),
    .B(_12283_),
    .Y(_12412_));
 sg13g2_mux2_1 _19314_ (.A0(\cpu.dcache.r_data[1][28] ),
    .A1(_12400_),
    .S(_12412_),
    .X(_12413_));
 sg13g2_nand2_1 _19315_ (.Y(_12414_),
    .A(_12398_),
    .B(_12413_));
 sg13g2_o21ai_1 _19316_ (.B1(_12414_),
    .Y(_00374_),
    .A1(_12175_),
    .A2(net54));
 sg13g2_mux2_1 _19317_ (.A0(\cpu.dcache.r_data[1][29] ),
    .A1(net1088),
    .S(_12412_),
    .X(_12415_));
 sg13g2_nand2_1 _19318_ (.Y(_12416_),
    .A(_12398_),
    .B(_12415_));
 sg13g2_o21ai_1 _19319_ (.B1(_12416_),
    .Y(_00375_),
    .A1(_12187_),
    .A2(net54));
 sg13g2_buf_1 _19320_ (.A(_12222_),
    .X(_12417_));
 sg13g2_nor2b_1 _19321_ (.A(_12326_),
    .B_N(\cpu.dcache.r_data[1][2] ),
    .Y(_12418_));
 sg13g2_a21oi_1 _19322_ (.A1(net993),
    .A2(_12326_),
    .Y(_12419_),
    .B1(_12418_));
 sg13g2_nand2_1 _19323_ (.Y(_12420_),
    .A(net895),
    .B(_12323_));
 sg13g2_o21ai_1 _19324_ (.B1(_12420_),
    .Y(_00376_),
    .A1(_12324_),
    .A2(_12419_));
 sg13g2_mux2_1 _19325_ (.A0(\cpu.dcache.r_data[1][30] ),
    .A1(net1091),
    .S(_12412_),
    .X(_12421_));
 sg13g2_nand2_1 _19326_ (.Y(_12422_),
    .A(_12398_),
    .B(_12421_));
 sg13g2_o21ai_1 _19327_ (.B1(_12422_),
    .Y(_00377_),
    .A1(net393),
    .A2(net54));
 sg13g2_mux2_1 _19328_ (.A0(\cpu.dcache.r_data[1][31] ),
    .A1(_12351_),
    .S(_12412_),
    .X(_12423_));
 sg13g2_nand2_1 _19329_ (.Y(_12424_),
    .A(_12398_),
    .B(_12423_));
 sg13g2_o21ai_1 _19330_ (.B1(_12424_),
    .Y(_00378_),
    .A1(_12201_),
    .A2(net54));
 sg13g2_buf_1 _19331_ (.A(_12228_),
    .X(_12425_));
 sg13g2_nor2b_1 _19332_ (.A(_12326_),
    .B_N(\cpu.dcache.r_data[1][3] ),
    .Y(_12426_));
 sg13g2_a21oi_1 _19333_ (.A1(net992),
    .A2(_12326_),
    .Y(_12427_),
    .B1(_12426_));
 sg13g2_nand2_1 _19334_ (.Y(_12428_),
    .A(net1003),
    .B(_12323_));
 sg13g2_o21ai_1 _19335_ (.B1(_12428_),
    .Y(_00379_),
    .A1(_12324_),
    .A2(_12427_));
 sg13g2_nor2_1 _19336_ (.A(net661),
    .B(_12300_),
    .Y(_12429_));
 sg13g2_buf_2 _19337_ (.A(_12429_),
    .X(_12430_));
 sg13g2_nor2b_1 _19338_ (.A(_12430_),
    .B_N(\cpu.dcache.r_data[1][4] ),
    .Y(_12431_));
 sg13g2_a21oi_1 _19339_ (.A1(net998),
    .A2(_12430_),
    .Y(_12432_),
    .B1(_12431_));
 sg13g2_nand2_1 _19340_ (.Y(_12433_),
    .A(net997),
    .B(_12323_));
 sg13g2_o21ai_1 _19341_ (.B1(_12433_),
    .Y(_00380_),
    .A1(net57),
    .A2(_12432_));
 sg13g2_nor2b_1 _19342_ (.A(_12430_),
    .B_N(\cpu.dcache.r_data[1][5] ),
    .Y(_12434_));
 sg13g2_a21oi_1 _19343_ (.A1(net996),
    .A2(_12430_),
    .Y(_12435_),
    .B1(_12434_));
 sg13g2_nand2_1 _19344_ (.Y(_12436_),
    .A(net995),
    .B(_12323_));
 sg13g2_o21ai_1 _19345_ (.B1(_12436_),
    .Y(_00381_),
    .A1(net57),
    .A2(_12435_));
 sg13g2_nor2b_1 _19346_ (.A(_12430_),
    .B_N(\cpu.dcache.r_data[1][6] ),
    .Y(_12437_));
 sg13g2_a21oi_1 _19347_ (.A1(net993),
    .A2(_12430_),
    .Y(_12438_),
    .B1(_12437_));
 sg13g2_nand2_1 _19348_ (.Y(_12439_),
    .A(net994),
    .B(_12323_));
 sg13g2_o21ai_1 _19349_ (.B1(_12439_),
    .Y(_00382_),
    .A1(net57),
    .A2(_12438_));
 sg13g2_nor2b_1 _19350_ (.A(_12430_),
    .B_N(\cpu.dcache.r_data[1][7] ),
    .Y(_12440_));
 sg13g2_a21oi_1 _19351_ (.A1(net992),
    .A2(_12430_),
    .Y(_12441_),
    .B1(_12440_));
 sg13g2_nand2_1 _19352_ (.Y(_12442_),
    .A(net999),
    .B(_12323_));
 sg13g2_o21ai_1 _19353_ (.B1(_12442_),
    .Y(_00383_),
    .A1(net57),
    .A2(_12441_));
 sg13g2_mux2_1 _19354_ (.A0(\cpu.dcache.r_data[1][8] ),
    .A1(net1089),
    .S(_12338_),
    .X(_12443_));
 sg13g2_nand2_1 _19355_ (.Y(_12444_),
    .A(_12336_),
    .B(_12443_));
 sg13g2_o21ai_1 _19356_ (.B1(_12444_),
    .Y(_00384_),
    .A1(_12261_),
    .A2(net56));
 sg13g2_mux2_1 _19357_ (.A0(\cpu.dcache.r_data[1][9] ),
    .A1(net1088),
    .S(_12338_),
    .X(_12445_));
 sg13g2_nand2_1 _19358_ (.Y(_12446_),
    .A(_12336_),
    .B(_12445_));
 sg13g2_o21ai_1 _19359_ (.B1(_12446_),
    .Y(_00385_),
    .A1(net390),
    .A2(net56));
 sg13g2_buf_1 _19360_ (.A(net928),
    .X(_12447_));
 sg13g2_nand2_1 _19361_ (.Y(_12448_),
    .A(_09500_),
    .B(net759));
 sg13g2_buf_1 _19362_ (.A(_12448_),
    .X(_12449_));
 sg13g2_nor2_1 _19363_ (.A(net606),
    .B(_12321_),
    .Y(_12450_));
 sg13g2_buf_2 _19364_ (.A(_12450_),
    .X(_12451_));
 sg13g2_buf_1 _19365_ (.A(_12451_),
    .X(_12452_));
 sg13g2_nor2_1 _19366_ (.A(_12449_),
    .B(_12136_),
    .Y(_12453_));
 sg13g2_buf_2 _19367_ (.A(_12453_),
    .X(_12454_));
 sg13g2_nor2b_1 _19368_ (.A(_12454_),
    .B_N(\cpu.dcache.r_data[2][0] ),
    .Y(_12455_));
 sg13g2_a21oi_1 _19369_ (.A1(net998),
    .A2(_12454_),
    .Y(_12456_),
    .B1(_12455_));
 sg13g2_nand2_1 _19370_ (.Y(_12457_),
    .A(net896),
    .B(_12452_));
 sg13g2_o21ai_1 _19371_ (.B1(_12457_),
    .Y(_00386_),
    .A1(net53),
    .A2(_12456_));
 sg13g2_buf_1 _19372_ (.A(net549),
    .X(_12458_));
 sg13g2_buf_1 _19373_ (.A(net488),
    .X(_12459_));
 sg13g2_nand2_1 _19374_ (.Y(_12460_),
    .A(net438),
    .B(_12334_));
 sg13g2_buf_1 _19375_ (.A(_12460_),
    .X(_12461_));
 sg13g2_buf_1 _19376_ (.A(_12461_),
    .X(_12462_));
 sg13g2_nor2_2 _19377_ (.A(net606),
    .B(_12160_),
    .Y(_12463_));
 sg13g2_mux2_1 _19378_ (.A0(\cpu.dcache.r_data[2][10] ),
    .A1(net1091),
    .S(_12463_),
    .X(_12464_));
 sg13g2_nand2_1 _19379_ (.Y(_12465_),
    .A(net52),
    .B(_12464_));
 sg13g2_o21ai_1 _19380_ (.B1(_12465_),
    .Y(_00387_),
    .A1(net397),
    .A2(net52));
 sg13g2_mux2_1 _19381_ (.A0(\cpu.dcache.r_data[2][11] ),
    .A1(net1090),
    .S(_12463_),
    .X(_12466_));
 sg13g2_nand2_1 _19382_ (.Y(_12467_),
    .A(net52),
    .B(_12466_));
 sg13g2_o21ai_1 _19383_ (.B1(_12467_),
    .Y(_00388_),
    .A1(net396),
    .A2(net52));
 sg13g2_nor2_2 _19384_ (.A(net606),
    .B(_12180_),
    .Y(_12468_));
 sg13g2_mux2_1 _19385_ (.A0(\cpu.dcache.r_data[2][12] ),
    .A1(net1089),
    .S(_12468_),
    .X(_12469_));
 sg13g2_nand2_1 _19386_ (.Y(_12470_),
    .A(_12461_),
    .B(_12469_));
 sg13g2_o21ai_1 _19387_ (.B1(_12470_),
    .Y(_00389_),
    .A1(net395),
    .A2(net52));
 sg13g2_mux2_1 _19388_ (.A0(\cpu.dcache.r_data[2][13] ),
    .A1(net1088),
    .S(_12468_),
    .X(_12471_));
 sg13g2_nand2_1 _19389_ (.Y(_12472_),
    .A(_12461_),
    .B(_12471_));
 sg13g2_o21ai_1 _19390_ (.B1(_12472_),
    .Y(_00390_),
    .A1(net394),
    .A2(_12462_));
 sg13g2_mux2_1 _19391_ (.A0(\cpu.dcache.r_data[2][14] ),
    .A1(net1091),
    .S(_12468_),
    .X(_12473_));
 sg13g2_nand2_1 _19392_ (.Y(_12474_),
    .A(_12461_),
    .B(_12473_));
 sg13g2_o21ai_1 _19393_ (.B1(_12474_),
    .Y(_00391_),
    .A1(net393),
    .A2(net52));
 sg13g2_mux2_1 _19394_ (.A0(\cpu.dcache.r_data[2][15] ),
    .A1(net1090),
    .S(_12468_),
    .X(_12475_));
 sg13g2_nand2_1 _19395_ (.Y(_12476_),
    .A(_12461_),
    .B(_12475_));
 sg13g2_o21ai_1 _19396_ (.B1(_12476_),
    .Y(_00392_),
    .A1(net392),
    .A2(net52));
 sg13g2_nor2_1 _19397_ (.A(net606),
    .B(_12355_),
    .Y(_12477_));
 sg13g2_buf_2 _19398_ (.A(_12477_),
    .X(_12478_));
 sg13g2_buf_1 _19399_ (.A(_12478_),
    .X(_12479_));
 sg13g2_nor2_1 _19400_ (.A(_12449_),
    .B(_12210_),
    .Y(_12480_));
 sg13g2_buf_2 _19401_ (.A(_12480_),
    .X(_12481_));
 sg13g2_nor2b_1 _19402_ (.A(_12481_),
    .B_N(\cpu.dcache.r_data[2][16] ),
    .Y(_12482_));
 sg13g2_a21oi_1 _19403_ (.A1(_12376_),
    .A2(_12481_),
    .Y(_12483_),
    .B1(_12482_));
 sg13g2_nand2_1 _19404_ (.Y(_12484_),
    .A(net896),
    .B(net51));
 sg13g2_o21ai_1 _19405_ (.B1(_12484_),
    .Y(_00393_),
    .A1(net51),
    .A2(_12483_));
 sg13g2_nor2b_1 _19406_ (.A(_12481_),
    .B_N(\cpu.dcache.r_data[2][17] ),
    .Y(_12485_));
 sg13g2_a21oi_1 _19407_ (.A1(net996),
    .A2(_12481_),
    .Y(_12486_),
    .B1(_12485_));
 sg13g2_nand2_1 _19408_ (.Y(_12487_),
    .A(_10196_),
    .B(_12479_));
 sg13g2_o21ai_1 _19409_ (.B1(_12487_),
    .Y(_00394_),
    .A1(_12479_),
    .A2(_12486_));
 sg13g2_nor2b_1 _19410_ (.A(_12481_),
    .B_N(\cpu.dcache.r_data[2][18] ),
    .Y(_12488_));
 sg13g2_a21oi_1 _19411_ (.A1(_12417_),
    .A2(_12481_),
    .Y(_12489_),
    .B1(_12488_));
 sg13g2_nand2_1 _19412_ (.Y(_12490_),
    .A(net895),
    .B(_12478_));
 sg13g2_o21ai_1 _19413_ (.B1(_12490_),
    .Y(_00395_),
    .A1(net51),
    .A2(_12489_));
 sg13g2_nor2b_1 _19414_ (.A(_12481_),
    .B_N(\cpu.dcache.r_data[2][19] ),
    .Y(_12491_));
 sg13g2_a21oi_1 _19415_ (.A1(_12425_),
    .A2(_12481_),
    .Y(_12492_),
    .B1(_12491_));
 sg13g2_nand2_1 _19416_ (.Y(_12493_),
    .A(net1003),
    .B(_12478_));
 sg13g2_o21ai_1 _19417_ (.B1(_12493_),
    .Y(_00396_),
    .A1(net51),
    .A2(_12492_));
 sg13g2_nor2b_1 _19418_ (.A(_12454_),
    .B_N(\cpu.dcache.r_data[2][1] ),
    .Y(_12494_));
 sg13g2_a21oi_1 _19419_ (.A1(net996),
    .A2(_12454_),
    .Y(_12495_),
    .B1(_12494_));
 sg13g2_nand2_1 _19420_ (.Y(_12496_),
    .A(net921),
    .B(_12452_));
 sg13g2_o21ai_1 _19421_ (.B1(_12496_),
    .Y(_00397_),
    .A1(net53),
    .A2(_12495_));
 sg13g2_nor2_1 _19422_ (.A(net606),
    .B(_12239_),
    .Y(_12497_));
 sg13g2_buf_2 _19423_ (.A(_12497_),
    .X(_12498_));
 sg13g2_nor2b_1 _19424_ (.A(_12498_),
    .B_N(\cpu.dcache.r_data[2][20] ),
    .Y(_12499_));
 sg13g2_a21oi_1 _19425_ (.A1(net998),
    .A2(_12498_),
    .Y(_12500_),
    .B1(_12499_));
 sg13g2_nand2_1 _19426_ (.Y(_12501_),
    .A(_12381_),
    .B(_12478_));
 sg13g2_o21ai_1 _19427_ (.B1(_12501_),
    .Y(_00398_),
    .A1(net51),
    .A2(_12500_));
 sg13g2_nor2b_1 _19428_ (.A(_12498_),
    .B_N(\cpu.dcache.r_data[2][21] ),
    .Y(_12502_));
 sg13g2_a21oi_1 _19429_ (.A1(net996),
    .A2(_12498_),
    .Y(_12503_),
    .B1(_12502_));
 sg13g2_nand2_1 _19430_ (.Y(_12504_),
    .A(_12386_),
    .B(_12478_));
 sg13g2_o21ai_1 _19431_ (.B1(_12504_),
    .Y(_00399_),
    .A1(net51),
    .A2(_12503_));
 sg13g2_nor2b_1 _19432_ (.A(_12498_),
    .B_N(\cpu.dcache.r_data[2][22] ),
    .Y(_12505_));
 sg13g2_a21oi_1 _19433_ (.A1(net993),
    .A2(_12498_),
    .Y(_12506_),
    .B1(_12505_));
 sg13g2_nand2_1 _19434_ (.Y(_12507_),
    .A(_12390_),
    .B(_12478_));
 sg13g2_o21ai_1 _19435_ (.B1(_12507_),
    .Y(_00400_),
    .A1(net51),
    .A2(_12506_));
 sg13g2_nor2b_1 _19436_ (.A(_12498_),
    .B_N(\cpu.dcache.r_data[2][23] ),
    .Y(_12508_));
 sg13g2_a21oi_1 _19437_ (.A1(net992),
    .A2(_12498_),
    .Y(_12509_),
    .B1(_12508_));
 sg13g2_nand2_1 _19438_ (.Y(_12510_),
    .A(_12256_),
    .B(_12478_));
 sg13g2_o21ai_1 _19439_ (.B1(_12510_),
    .Y(_00401_),
    .A1(net51),
    .A2(_12509_));
 sg13g2_nand2_1 _19440_ (.Y(_12511_),
    .A(net438),
    .B(_12396_));
 sg13g2_buf_2 _19441_ (.A(_12511_),
    .X(_12512_));
 sg13g2_buf_1 _19442_ (.A(_12512_),
    .X(_12513_));
 sg13g2_nor2_1 _19443_ (.A(_12448_),
    .B(net663),
    .Y(_12514_));
 sg13g2_buf_2 _19444_ (.A(_12514_),
    .X(_12515_));
 sg13g2_mux2_1 _19445_ (.A0(\cpu.dcache.r_data[2][24] ),
    .A1(net1089),
    .S(_12515_),
    .X(_12516_));
 sg13g2_nand2_1 _19446_ (.Y(_12517_),
    .A(net50),
    .B(_12516_));
 sg13g2_o21ai_1 _19447_ (.B1(_12517_),
    .Y(_00402_),
    .A1(net391),
    .A2(net50));
 sg13g2_mux2_1 _19448_ (.A0(\cpu.dcache.r_data[2][25] ),
    .A1(_12405_),
    .S(_12515_),
    .X(_12518_));
 sg13g2_nand2_1 _19449_ (.Y(_12519_),
    .A(net50),
    .B(_12518_));
 sg13g2_o21ai_1 _19450_ (.B1(_12519_),
    .Y(_00403_),
    .A1(net390),
    .A2(net50));
 sg13g2_mux2_1 _19451_ (.A0(\cpu.dcache.r_data[2][26] ),
    .A1(net1091),
    .S(_12515_),
    .X(_12520_));
 sg13g2_nand2_1 _19452_ (.Y(_12521_),
    .A(_12512_),
    .B(_12520_));
 sg13g2_o21ai_1 _19453_ (.B1(_12521_),
    .Y(_00404_),
    .A1(net397),
    .A2(_12513_));
 sg13g2_mux2_1 _19454_ (.A0(\cpu.dcache.r_data[2][27] ),
    .A1(_12351_),
    .S(_12515_),
    .X(_12522_));
 sg13g2_nand2_1 _19455_ (.Y(_12523_),
    .A(_12512_),
    .B(_12522_));
 sg13g2_o21ai_1 _19456_ (.B1(_12523_),
    .Y(_00405_),
    .A1(net396),
    .A2(_12513_));
 sg13g2_nor2_2 _19457_ (.A(net606),
    .B(_12283_),
    .Y(_12524_));
 sg13g2_mux2_1 _19458_ (.A0(\cpu.dcache.r_data[2][28] ),
    .A1(net1089),
    .S(_12524_),
    .X(_12525_));
 sg13g2_nand2_1 _19459_ (.Y(_12526_),
    .A(_12512_),
    .B(_12525_));
 sg13g2_o21ai_1 _19460_ (.B1(_12526_),
    .Y(_00406_),
    .A1(net395),
    .A2(net50));
 sg13g2_mux2_1 _19461_ (.A0(\cpu.dcache.r_data[2][29] ),
    .A1(net1088),
    .S(_12524_),
    .X(_12527_));
 sg13g2_nand2_1 _19462_ (.Y(_12528_),
    .A(_12512_),
    .B(_12527_));
 sg13g2_o21ai_1 _19463_ (.B1(_12528_),
    .Y(_00407_),
    .A1(net394),
    .A2(net50));
 sg13g2_nor2b_1 _19464_ (.A(_12454_),
    .B_N(\cpu.dcache.r_data[2][2] ),
    .Y(_12529_));
 sg13g2_a21oi_1 _19465_ (.A1(net993),
    .A2(_12454_),
    .Y(_12530_),
    .B1(_12529_));
 sg13g2_nand2_1 _19466_ (.Y(_12531_),
    .A(net895),
    .B(_12451_));
 sg13g2_o21ai_1 _19467_ (.B1(_12531_),
    .Y(_00408_),
    .A1(net53),
    .A2(_12530_));
 sg13g2_mux2_1 _19468_ (.A0(\cpu.dcache.r_data[2][30] ),
    .A1(net1091),
    .S(_12524_),
    .X(_12532_));
 sg13g2_nand2_1 _19469_ (.Y(_12533_),
    .A(_12512_),
    .B(_12532_));
 sg13g2_o21ai_1 _19470_ (.B1(_12533_),
    .Y(_00409_),
    .A1(net393),
    .A2(net50));
 sg13g2_mux2_1 _19471_ (.A0(\cpu.dcache.r_data[2][31] ),
    .A1(net1090),
    .S(_12524_),
    .X(_12534_));
 sg13g2_nand2_1 _19472_ (.Y(_12535_),
    .A(_12512_),
    .B(_12534_));
 sg13g2_o21ai_1 _19473_ (.B1(_12535_),
    .Y(_00410_),
    .A1(net392),
    .A2(net50));
 sg13g2_nor2b_1 _19474_ (.A(_12454_),
    .B_N(\cpu.dcache.r_data[2][3] ),
    .Y(_12536_));
 sg13g2_a21oi_1 _19475_ (.A1(net992),
    .A2(_12454_),
    .Y(_12537_),
    .B1(_12536_));
 sg13g2_nand2_1 _19476_ (.Y(_12538_),
    .A(net1003),
    .B(_12451_));
 sg13g2_o21ai_1 _19477_ (.B1(_12538_),
    .Y(_00411_),
    .A1(net53),
    .A2(_12537_));
 sg13g2_nor2_1 _19478_ (.A(net606),
    .B(_12300_),
    .Y(_12539_));
 sg13g2_buf_2 _19479_ (.A(_12539_),
    .X(_12540_));
 sg13g2_nor2b_1 _19480_ (.A(_12540_),
    .B_N(\cpu.dcache.r_data[2][4] ),
    .Y(_12541_));
 sg13g2_a21oi_1 _19481_ (.A1(net998),
    .A2(_12540_),
    .Y(_12542_),
    .B1(_12541_));
 sg13g2_nand2_1 _19482_ (.Y(_12543_),
    .A(net997),
    .B(_12451_));
 sg13g2_o21ai_1 _19483_ (.B1(_12543_),
    .Y(_00412_),
    .A1(net53),
    .A2(_12542_));
 sg13g2_nor2b_1 _19484_ (.A(_12540_),
    .B_N(\cpu.dcache.r_data[2][5] ),
    .Y(_12544_));
 sg13g2_a21oi_1 _19485_ (.A1(net996),
    .A2(_12540_),
    .Y(_12545_),
    .B1(_12544_));
 sg13g2_nand2_1 _19486_ (.Y(_12546_),
    .A(net995),
    .B(_12451_));
 sg13g2_o21ai_1 _19487_ (.B1(_12546_),
    .Y(_00413_),
    .A1(net53),
    .A2(_12545_));
 sg13g2_nor2b_1 _19488_ (.A(_12540_),
    .B_N(\cpu.dcache.r_data[2][6] ),
    .Y(_12547_));
 sg13g2_a21oi_1 _19489_ (.A1(net993),
    .A2(_12540_),
    .Y(_12548_),
    .B1(_12547_));
 sg13g2_nand2_1 _19490_ (.Y(_12549_),
    .A(net994),
    .B(_12451_));
 sg13g2_o21ai_1 _19491_ (.B1(_12549_),
    .Y(_00414_),
    .A1(net53),
    .A2(_12548_));
 sg13g2_nor2b_1 _19492_ (.A(_12540_),
    .B_N(\cpu.dcache.r_data[2][7] ),
    .Y(_12550_));
 sg13g2_a21oi_1 _19493_ (.A1(net992),
    .A2(_12540_),
    .Y(_12551_),
    .B1(_12550_));
 sg13g2_nand2_1 _19494_ (.Y(_12552_),
    .A(net999),
    .B(_12451_));
 sg13g2_o21ai_1 _19495_ (.B1(_12552_),
    .Y(_00415_),
    .A1(net53),
    .A2(_12551_));
 sg13g2_mux2_1 _19496_ (.A0(\cpu.dcache.r_data[2][8] ),
    .A1(net1089),
    .S(_12463_),
    .X(_12553_));
 sg13g2_nand2_1 _19497_ (.Y(_12554_),
    .A(_12461_),
    .B(_12553_));
 sg13g2_o21ai_1 _19498_ (.B1(_12554_),
    .Y(_00416_),
    .A1(net391),
    .A2(_12462_));
 sg13g2_mux2_1 _19499_ (.A0(\cpu.dcache.r_data[2][9] ),
    .A1(net1088),
    .S(_12463_),
    .X(_12555_));
 sg13g2_nand2_1 _19500_ (.Y(_12556_),
    .A(_12461_),
    .B(_12555_));
 sg13g2_o21ai_1 _19501_ (.B1(_12556_),
    .Y(_00417_),
    .A1(net390),
    .A2(net52));
 sg13g2_buf_1 _19502_ (.A(net619),
    .X(_12557_));
 sg13g2_buf_2 _19503_ (.A(net496),
    .X(_12558_));
 sg13g2_nand3_1 _19504_ (.B(net437),
    .C(_09500_),
    .A(net531),
    .Y(_12559_));
 sg13g2_buf_1 _19505_ (.A(_12559_),
    .X(_12560_));
 sg13g2_buf_1 _19506_ (.A(_12560_),
    .X(_12561_));
 sg13g2_nor2_1 _19507_ (.A(net271),
    .B(_12321_),
    .Y(_12562_));
 sg13g2_buf_1 _19508_ (.A(_12562_),
    .X(_12563_));
 sg13g2_nor2_1 _19509_ (.A(_12561_),
    .B(_12136_),
    .Y(_12564_));
 sg13g2_buf_2 _19510_ (.A(_12564_),
    .X(_12565_));
 sg13g2_nor2b_1 _19511_ (.A(_12565_),
    .B_N(\cpu.dcache.r_data[3][0] ),
    .Y(_12566_));
 sg13g2_a21oi_1 _19512_ (.A1(net998),
    .A2(_12565_),
    .Y(_12567_),
    .B1(_12566_));
 sg13g2_nand2_1 _19513_ (.Y(_12568_),
    .A(net896),
    .B(net69));
 sg13g2_o21ai_1 _19514_ (.B1(_12568_),
    .Y(_00418_),
    .A1(net69),
    .A2(_12567_));
 sg13g2_buf_1 _19515_ (.A(net627),
    .X(_12569_));
 sg13g2_buf_1 _19516_ (.A(net530),
    .X(_12570_));
 sg13g2_nand2_1 _19517_ (.Y(_12571_),
    .A(net487),
    .B(_12334_));
 sg13g2_buf_1 _19518_ (.A(_12571_),
    .X(_12572_));
 sg13g2_buf_1 _19519_ (.A(_12572_),
    .X(_12573_));
 sg13g2_nor2_2 _19520_ (.A(net271),
    .B(_12160_),
    .Y(_12574_));
 sg13g2_mux2_1 _19521_ (.A0(\cpu.dcache.r_data[3][10] ),
    .A1(net1091),
    .S(_12574_),
    .X(_12575_));
 sg13g2_nand2_1 _19522_ (.Y(_12576_),
    .A(net49),
    .B(_12575_));
 sg13g2_o21ai_1 _19523_ (.B1(_12576_),
    .Y(_00419_),
    .A1(net397),
    .A2(net49));
 sg13g2_mux2_1 _19524_ (.A0(\cpu.dcache.r_data[3][11] ),
    .A1(net1090),
    .S(_12574_),
    .X(_12577_));
 sg13g2_nand2_1 _19525_ (.Y(_12578_),
    .A(net49),
    .B(_12577_));
 sg13g2_o21ai_1 _19526_ (.B1(_12578_),
    .Y(_00420_),
    .A1(net396),
    .A2(net49));
 sg13g2_nor2_2 _19527_ (.A(net271),
    .B(_12180_),
    .Y(_12579_));
 sg13g2_mux2_1 _19528_ (.A0(\cpu.dcache.r_data[3][12] ),
    .A1(net1089),
    .S(_12579_),
    .X(_12580_));
 sg13g2_nand2_1 _19529_ (.Y(_12581_),
    .A(_12572_),
    .B(_12580_));
 sg13g2_o21ai_1 _19530_ (.B1(_12581_),
    .Y(_00421_),
    .A1(net395),
    .A2(net49));
 sg13g2_mux2_1 _19531_ (.A0(\cpu.dcache.r_data[3][13] ),
    .A1(_12405_),
    .S(_12579_),
    .X(_12582_));
 sg13g2_nand2_1 _19532_ (.Y(_12583_),
    .A(_12572_),
    .B(_12582_));
 sg13g2_o21ai_1 _19533_ (.B1(_12583_),
    .Y(_00422_),
    .A1(net394),
    .A2(net49));
 sg13g2_mux2_1 _19534_ (.A0(\cpu.dcache.r_data[3][14] ),
    .A1(net1091),
    .S(_12579_),
    .X(_12584_));
 sg13g2_nand2_1 _19535_ (.Y(_12585_),
    .A(_12572_),
    .B(_12584_));
 sg13g2_o21ai_1 _19536_ (.B1(_12585_),
    .Y(_00423_),
    .A1(net393),
    .A2(_12573_));
 sg13g2_mux2_1 _19537_ (.A0(\cpu.dcache.r_data[3][15] ),
    .A1(net1090),
    .S(_12579_),
    .X(_12586_));
 sg13g2_nand2_1 _19538_ (.Y(_12587_),
    .A(_12572_),
    .B(_12586_));
 sg13g2_o21ai_1 _19539_ (.B1(_12587_),
    .Y(_00424_),
    .A1(net392),
    .A2(_12573_));
 sg13g2_nor2_1 _19540_ (.A(net271),
    .B(_12355_),
    .Y(_12588_));
 sg13g2_buf_1 _19541_ (.A(_12588_),
    .X(_12589_));
 sg13g2_nor2_1 _19542_ (.A(_12561_),
    .B(_12210_),
    .Y(_12590_));
 sg13g2_buf_2 _19543_ (.A(_12590_),
    .X(_12591_));
 sg13g2_nor2b_1 _19544_ (.A(_12591_),
    .B_N(\cpu.dcache.r_data[3][16] ),
    .Y(_12592_));
 sg13g2_a21oi_1 _19545_ (.A1(_12376_),
    .A2(_12591_),
    .Y(_12593_),
    .B1(_12592_));
 sg13g2_nand2_1 _19546_ (.Y(_12594_),
    .A(_12215_),
    .B(net68));
 sg13g2_o21ai_1 _19547_ (.B1(_12594_),
    .Y(_00425_),
    .A1(net68),
    .A2(_12593_));
 sg13g2_nor2b_1 _19548_ (.A(_12591_),
    .B_N(\cpu.dcache.r_data[3][17] ),
    .Y(_12595_));
 sg13g2_a21oi_1 _19549_ (.A1(_12383_),
    .A2(_12591_),
    .Y(_12596_),
    .B1(_12595_));
 sg13g2_nand2_1 _19550_ (.Y(_12597_),
    .A(_10196_),
    .B(_12589_));
 sg13g2_o21ai_1 _19551_ (.B1(_12597_),
    .Y(_00426_),
    .A1(_12589_),
    .A2(_12596_));
 sg13g2_nor2b_1 _19552_ (.A(_12591_),
    .B_N(\cpu.dcache.r_data[3][18] ),
    .Y(_12598_));
 sg13g2_a21oi_1 _19553_ (.A1(_12417_),
    .A2(_12591_),
    .Y(_12599_),
    .B1(_12598_));
 sg13g2_nand2_1 _19554_ (.Y(_12600_),
    .A(net895),
    .B(_12588_));
 sg13g2_o21ai_1 _19555_ (.B1(_12600_),
    .Y(_00427_),
    .A1(net68),
    .A2(_12599_));
 sg13g2_nor2b_1 _19556_ (.A(_12591_),
    .B_N(\cpu.dcache.r_data[3][19] ),
    .Y(_12601_));
 sg13g2_a21oi_1 _19557_ (.A1(_12425_),
    .A2(_12591_),
    .Y(_12602_),
    .B1(_12601_));
 sg13g2_nand2_1 _19558_ (.Y(_12603_),
    .A(net1003),
    .B(_12588_));
 sg13g2_o21ai_1 _19559_ (.B1(_12603_),
    .Y(_00428_),
    .A1(net68),
    .A2(_12602_));
 sg13g2_nor2b_1 _19560_ (.A(_12565_),
    .B_N(\cpu.dcache.r_data[3][1] ),
    .Y(_12604_));
 sg13g2_a21oi_1 _19561_ (.A1(net996),
    .A2(_12565_),
    .Y(_12605_),
    .B1(_12604_));
 sg13g2_nand2_1 _19562_ (.Y(_12606_),
    .A(net921),
    .B(_12563_));
 sg13g2_o21ai_1 _19563_ (.B1(_12606_),
    .Y(_00429_),
    .A1(net69),
    .A2(_12605_));
 sg13g2_or2_1 _19564_ (.X(_12607_),
    .B(_12239_),
    .A(net271));
 sg13g2_buf_1 _19565_ (.A(_12607_),
    .X(_12608_));
 sg13g2_mux2_1 _19566_ (.A0(_12176_),
    .A1(\cpu.dcache.r_data[3][20] ),
    .S(_12608_),
    .X(_12609_));
 sg13g2_mux2_1 _19567_ (.A0(_12609_),
    .A1(net1002),
    .S(net68),
    .X(_00430_));
 sg13g2_mux2_1 _19568_ (.A0(_12189_),
    .A1(\cpu.dcache.r_data[3][21] ),
    .S(_12608_),
    .X(_12610_));
 sg13g2_mux2_1 _19569_ (.A0(_12610_),
    .A1(net1001),
    .S(net68),
    .X(_00431_));
 sg13g2_mux2_1 _19570_ (.A0(_12158_),
    .A1(\cpu.dcache.r_data[3][22] ),
    .S(_12608_),
    .X(_12611_));
 sg13g2_mux2_1 _19571_ (.A0(_12611_),
    .A1(net1000),
    .S(net68),
    .X(_00432_));
 sg13g2_mux2_1 _19572_ (.A0(_12169_),
    .A1(\cpu.dcache.r_data[3][23] ),
    .S(_12608_),
    .X(_12612_));
 sg13g2_buf_1 _19573_ (.A(_10229_),
    .X(_12613_));
 sg13g2_mux2_1 _19574_ (.A0(_12612_),
    .A1(net991),
    .S(net68),
    .X(_00433_));
 sg13g2_nand2_1 _19575_ (.Y(_12614_),
    .A(net487),
    .B(_12396_));
 sg13g2_buf_2 _19576_ (.A(_12614_),
    .X(_12615_));
 sg13g2_buf_1 _19577_ (.A(_12615_),
    .X(_12616_));
 sg13g2_nor2_1 _19578_ (.A(_12560_),
    .B(net663),
    .Y(_12617_));
 sg13g2_buf_2 _19579_ (.A(_12617_),
    .X(_12618_));
 sg13g2_mux2_1 _19580_ (.A0(\cpu.dcache.r_data[3][24] ),
    .A1(net1089),
    .S(_12618_),
    .X(_12619_));
 sg13g2_nand2_1 _19581_ (.Y(_12620_),
    .A(net48),
    .B(_12619_));
 sg13g2_o21ai_1 _19582_ (.B1(_12620_),
    .Y(_00434_),
    .A1(net391),
    .A2(net48));
 sg13g2_mux2_1 _19583_ (.A0(\cpu.dcache.r_data[3][25] ),
    .A1(net1088),
    .S(_12618_),
    .X(_12621_));
 sg13g2_nand2_1 _19584_ (.Y(_12622_),
    .A(net48),
    .B(_12621_));
 sg13g2_o21ai_1 _19585_ (.B1(_12622_),
    .Y(_00435_),
    .A1(net390),
    .A2(net48));
 sg13g2_mux2_1 _19586_ (.A0(\cpu.dcache.r_data[3][26] ),
    .A1(net1091),
    .S(_12618_),
    .X(_12623_));
 sg13g2_nand2_1 _19587_ (.Y(_12624_),
    .A(_12615_),
    .B(_12623_));
 sg13g2_o21ai_1 _19588_ (.B1(_12624_),
    .Y(_00436_),
    .A1(net397),
    .A2(_12616_));
 sg13g2_mux2_1 _19589_ (.A0(\cpu.dcache.r_data[3][27] ),
    .A1(net1090),
    .S(_12618_),
    .X(_12625_));
 sg13g2_nand2_1 _19590_ (.Y(_12626_),
    .A(_12615_),
    .B(_12625_));
 sg13g2_o21ai_1 _19591_ (.B1(_12626_),
    .Y(_00437_),
    .A1(net396),
    .A2(_12616_));
 sg13g2_nor2_2 _19592_ (.A(net271),
    .B(_12283_),
    .Y(_12627_));
 sg13g2_mux2_1 _19593_ (.A0(\cpu.dcache.r_data[3][28] ),
    .A1(net1089),
    .S(_12627_),
    .X(_12628_));
 sg13g2_nand2_1 _19594_ (.Y(_12629_),
    .A(_12615_),
    .B(_12628_));
 sg13g2_o21ai_1 _19595_ (.B1(_12629_),
    .Y(_00438_),
    .A1(net395),
    .A2(net48));
 sg13g2_mux2_1 _19596_ (.A0(\cpu.dcache.r_data[3][29] ),
    .A1(net1088),
    .S(_12627_),
    .X(_12630_));
 sg13g2_nand2_1 _19597_ (.Y(_12631_),
    .A(_12615_),
    .B(_12630_));
 sg13g2_o21ai_1 _19598_ (.B1(_12631_),
    .Y(_00439_),
    .A1(net394),
    .A2(net48));
 sg13g2_nor2b_1 _19599_ (.A(_12565_),
    .B_N(\cpu.dcache.r_data[3][2] ),
    .Y(_12632_));
 sg13g2_a21oi_1 _19600_ (.A1(net993),
    .A2(_12565_),
    .Y(_12633_),
    .B1(_12632_));
 sg13g2_nand2_1 _19601_ (.Y(_12634_),
    .A(net895),
    .B(_12562_));
 sg13g2_o21ai_1 _19602_ (.B1(_12634_),
    .Y(_00440_),
    .A1(_12563_),
    .A2(_12633_));
 sg13g2_buf_1 _19603_ (.A(_12157_),
    .X(_12635_));
 sg13g2_mux2_1 _19604_ (.A0(\cpu.dcache.r_data[3][30] ),
    .A1(net1087),
    .S(_12627_),
    .X(_12636_));
 sg13g2_nand2_1 _19605_ (.Y(_12637_),
    .A(_12615_),
    .B(_12636_));
 sg13g2_o21ai_1 _19606_ (.B1(_12637_),
    .Y(_00441_),
    .A1(net393),
    .A2(net48));
 sg13g2_buf_1 _19607_ (.A(_12168_),
    .X(_12638_));
 sg13g2_mux2_1 _19608_ (.A0(\cpu.dcache.r_data[3][31] ),
    .A1(net1086),
    .S(_12627_),
    .X(_12639_));
 sg13g2_nand2_1 _19609_ (.Y(_12640_),
    .A(_12615_),
    .B(_12639_));
 sg13g2_o21ai_1 _19610_ (.B1(_12640_),
    .Y(_00442_),
    .A1(net392),
    .A2(net48));
 sg13g2_nor2b_1 _19611_ (.A(_12565_),
    .B_N(\cpu.dcache.r_data[3][3] ),
    .Y(_12641_));
 sg13g2_a21oi_1 _19612_ (.A1(net992),
    .A2(_12565_),
    .Y(_12642_),
    .B1(_12641_));
 sg13g2_nand2_1 _19613_ (.Y(_12643_),
    .A(net1003),
    .B(_12562_));
 sg13g2_o21ai_1 _19614_ (.B1(_12643_),
    .Y(_00443_),
    .A1(net69),
    .A2(_12642_));
 sg13g2_or2_1 _19615_ (.X(_12644_),
    .B(_12300_),
    .A(net271));
 sg13g2_buf_1 _19616_ (.A(_12644_),
    .X(_12645_));
 sg13g2_mux2_1 _19617_ (.A0(net1096),
    .A1(\cpu.dcache.r_data[3][4] ),
    .S(_12645_),
    .X(_12646_));
 sg13g2_mux2_1 _19618_ (.A0(_12646_),
    .A1(net1002),
    .S(net69),
    .X(_00444_));
 sg13g2_mux2_1 _19619_ (.A0(net1095),
    .A1(\cpu.dcache.r_data[3][5] ),
    .S(_12645_),
    .X(_12647_));
 sg13g2_mux2_1 _19620_ (.A0(_12647_),
    .A1(net1001),
    .S(net69),
    .X(_00445_));
 sg13g2_mux2_1 _19621_ (.A0(net1098),
    .A1(\cpu.dcache.r_data[3][6] ),
    .S(_12645_),
    .X(_12648_));
 sg13g2_mux2_1 _19622_ (.A0(_12648_),
    .A1(net1000),
    .S(net69),
    .X(_00446_));
 sg13g2_mux2_1 _19623_ (.A0(net1097),
    .A1(\cpu.dcache.r_data[3][7] ),
    .S(_12645_),
    .X(_12649_));
 sg13g2_mux2_1 _19624_ (.A0(_12649_),
    .A1(net991),
    .S(net69),
    .X(_00447_));
 sg13g2_buf_1 _19625_ (.A(_12125_),
    .X(_12650_));
 sg13g2_mux2_1 _19626_ (.A0(\cpu.dcache.r_data[3][8] ),
    .A1(net1085),
    .S(_12574_),
    .X(_12651_));
 sg13g2_nand2_1 _19627_ (.Y(_12652_),
    .A(_12572_),
    .B(_12651_));
 sg13g2_o21ai_1 _19628_ (.B1(_12652_),
    .Y(_00448_),
    .A1(net391),
    .A2(net49));
 sg13g2_buf_1 _19629_ (.A(_12188_),
    .X(_12653_));
 sg13g2_mux2_1 _19630_ (.A0(\cpu.dcache.r_data[3][9] ),
    .A1(net1084),
    .S(_12574_),
    .X(_12654_));
 sg13g2_nand2_1 _19631_ (.Y(_12655_),
    .A(_12572_),
    .B(_12654_));
 sg13g2_o21ai_1 _19632_ (.B1(_12655_),
    .Y(_00449_),
    .A1(net390),
    .A2(net49));
 sg13g2_buf_1 _19633_ (.A(_09519_),
    .X(_12656_));
 sg13g2_nand2_1 _19634_ (.Y(_12657_),
    .A(net758),
    .B(_09839_));
 sg13g2_buf_1 _19635_ (.A(_12657_),
    .X(_12658_));
 sg13g2_nor2_1 _19636_ (.A(net605),
    .B(_12321_),
    .Y(_12659_));
 sg13g2_buf_2 _19637_ (.A(_12659_),
    .X(_12660_));
 sg13g2_buf_1 _19638_ (.A(_12660_),
    .X(_12661_));
 sg13g2_nor2_1 _19639_ (.A(_12658_),
    .B(_12136_),
    .Y(_12662_));
 sg13g2_buf_2 _19640_ (.A(_12662_),
    .X(_12663_));
 sg13g2_nor2b_1 _19641_ (.A(_12663_),
    .B_N(\cpu.dcache.r_data[4][0] ),
    .Y(_12664_));
 sg13g2_a21oi_1 _19642_ (.A1(net998),
    .A2(_12663_),
    .Y(_12665_),
    .B1(_12664_));
 sg13g2_nand2_1 _19643_ (.Y(_12666_),
    .A(net896),
    .B(net47));
 sg13g2_o21ai_1 _19644_ (.B1(_12666_),
    .Y(_00450_),
    .A1(net47),
    .A2(_12665_));
 sg13g2_nand2_1 _19645_ (.Y(_12667_),
    .A(_10236_),
    .B(_12334_));
 sg13g2_buf_1 _19646_ (.A(_12667_),
    .X(_12668_));
 sg13g2_buf_1 _19647_ (.A(_12668_),
    .X(_12669_));
 sg13g2_nor2_2 _19648_ (.A(net605),
    .B(_12160_),
    .Y(_12670_));
 sg13g2_mux2_1 _19649_ (.A0(\cpu.dcache.r_data[4][10] ),
    .A1(net1087),
    .S(_12670_),
    .X(_12671_));
 sg13g2_nand2_1 _19650_ (.Y(_12672_),
    .A(net46),
    .B(_12671_));
 sg13g2_o21ai_1 _19651_ (.B1(_12672_),
    .Y(_00451_),
    .A1(net397),
    .A2(net46));
 sg13g2_mux2_1 _19652_ (.A0(\cpu.dcache.r_data[4][11] ),
    .A1(net1086),
    .S(_12670_),
    .X(_12673_));
 sg13g2_nand2_1 _19653_ (.Y(_12674_),
    .A(net46),
    .B(_12673_));
 sg13g2_o21ai_1 _19654_ (.B1(_12674_),
    .Y(_00452_),
    .A1(net396),
    .A2(net46));
 sg13g2_nor2_2 _19655_ (.A(net605),
    .B(_12180_),
    .Y(_12675_));
 sg13g2_mux2_1 _19656_ (.A0(\cpu.dcache.r_data[4][12] ),
    .A1(net1085),
    .S(_12675_),
    .X(_12676_));
 sg13g2_nand2_1 _19657_ (.Y(_12677_),
    .A(_12668_),
    .B(_12676_));
 sg13g2_o21ai_1 _19658_ (.B1(_12677_),
    .Y(_00453_),
    .A1(net395),
    .A2(net46));
 sg13g2_mux2_1 _19659_ (.A0(\cpu.dcache.r_data[4][13] ),
    .A1(_12653_),
    .S(_12675_),
    .X(_12678_));
 sg13g2_nand2_1 _19660_ (.Y(_12679_),
    .A(_12668_),
    .B(_12678_));
 sg13g2_o21ai_1 _19661_ (.B1(_12679_),
    .Y(_00454_),
    .A1(net394),
    .A2(net46));
 sg13g2_mux2_1 _19662_ (.A0(\cpu.dcache.r_data[4][14] ),
    .A1(net1087),
    .S(_12675_),
    .X(_12680_));
 sg13g2_nand2_1 _19663_ (.Y(_12681_),
    .A(_12668_),
    .B(_12680_));
 sg13g2_o21ai_1 _19664_ (.B1(_12681_),
    .Y(_00455_),
    .A1(net393),
    .A2(_12669_));
 sg13g2_mux2_1 _19665_ (.A0(\cpu.dcache.r_data[4][15] ),
    .A1(net1086),
    .S(_12675_),
    .X(_12682_));
 sg13g2_nand2_1 _19666_ (.Y(_12683_),
    .A(_12668_),
    .B(_12682_));
 sg13g2_o21ai_1 _19667_ (.B1(_12683_),
    .Y(_00456_),
    .A1(net392),
    .A2(net46));
 sg13g2_nor2_1 _19668_ (.A(net605),
    .B(_12355_),
    .Y(_12684_));
 sg13g2_buf_2 _19669_ (.A(_12684_),
    .X(_12685_));
 sg13g2_buf_1 _19670_ (.A(_12685_),
    .X(_12686_));
 sg13g2_nor2_1 _19671_ (.A(_12658_),
    .B(_12210_),
    .Y(_12687_));
 sg13g2_buf_2 _19672_ (.A(_12687_),
    .X(_12688_));
 sg13g2_nor2b_1 _19673_ (.A(_12688_),
    .B_N(\cpu.dcache.r_data[4][16] ),
    .Y(_12689_));
 sg13g2_a21oi_1 _19674_ (.A1(net998),
    .A2(_12688_),
    .Y(_12690_),
    .B1(_12689_));
 sg13g2_nand2_1 _19675_ (.Y(_12691_),
    .A(_12215_),
    .B(_12686_));
 sg13g2_o21ai_1 _19676_ (.B1(_12691_),
    .Y(_00457_),
    .A1(net45),
    .A2(_12690_));
 sg13g2_nor2b_1 _19677_ (.A(_12688_),
    .B_N(\cpu.dcache.r_data[4][17] ),
    .Y(_12692_));
 sg13g2_a21oi_1 _19678_ (.A1(_12383_),
    .A2(_12688_),
    .Y(_12693_),
    .B1(_12692_));
 sg13g2_buf_1 _19679_ (.A(_10195_),
    .X(_12694_));
 sg13g2_nand2_1 _19680_ (.Y(_12695_),
    .A(net894),
    .B(net45));
 sg13g2_o21ai_1 _19681_ (.B1(_12695_),
    .Y(_00458_),
    .A1(net45),
    .A2(_12693_));
 sg13g2_nor2b_1 _19682_ (.A(_12688_),
    .B_N(\cpu.dcache.r_data[4][18] ),
    .Y(_12696_));
 sg13g2_a21oi_1 _19683_ (.A1(net993),
    .A2(_12688_),
    .Y(_12697_),
    .B1(_12696_));
 sg13g2_nand2_1 _19684_ (.Y(_12698_),
    .A(net895),
    .B(_12685_));
 sg13g2_o21ai_1 _19685_ (.B1(_12698_),
    .Y(_00459_),
    .A1(_12686_),
    .A2(_12697_));
 sg13g2_nor2b_1 _19686_ (.A(_12688_),
    .B_N(\cpu.dcache.r_data[4][19] ),
    .Y(_12699_));
 sg13g2_a21oi_1 _19687_ (.A1(net992),
    .A2(_12688_),
    .Y(_12700_),
    .B1(_12699_));
 sg13g2_nand2_1 _19688_ (.Y(_12701_),
    .A(net1003),
    .B(_12685_));
 sg13g2_o21ai_1 _19689_ (.B1(_12701_),
    .Y(_00460_),
    .A1(net45),
    .A2(_12700_));
 sg13g2_nor2b_1 _19690_ (.A(_12663_),
    .B_N(\cpu.dcache.r_data[4][1] ),
    .Y(_12702_));
 sg13g2_a21oi_1 _19691_ (.A1(net996),
    .A2(_12663_),
    .Y(_12703_),
    .B1(_12702_));
 sg13g2_nand2_1 _19692_ (.Y(_12704_),
    .A(net894),
    .B(_12661_));
 sg13g2_o21ai_1 _19693_ (.B1(_12704_),
    .Y(_00461_),
    .A1(net47),
    .A2(_12703_));
 sg13g2_buf_1 _19694_ (.A(_12126_),
    .X(_12705_));
 sg13g2_nor2_1 _19695_ (.A(net605),
    .B(_12239_),
    .Y(_12706_));
 sg13g2_buf_2 _19696_ (.A(_12706_),
    .X(_12707_));
 sg13g2_nor2b_1 _19697_ (.A(_12707_),
    .B_N(\cpu.dcache.r_data[4][20] ),
    .Y(_12708_));
 sg13g2_a21oi_1 _19698_ (.A1(_12705_),
    .A2(_12707_),
    .Y(_12709_),
    .B1(_12708_));
 sg13g2_nand2_1 _19699_ (.Y(_12710_),
    .A(net997),
    .B(_12685_));
 sg13g2_o21ai_1 _19700_ (.B1(_12710_),
    .Y(_00462_),
    .A1(net45),
    .A2(_12709_));
 sg13g2_buf_1 _19701_ (.A(net1094),
    .X(_12711_));
 sg13g2_nor2b_1 _19702_ (.A(_12707_),
    .B_N(\cpu.dcache.r_data[4][21] ),
    .Y(_12712_));
 sg13g2_a21oi_1 _19703_ (.A1(_12711_),
    .A2(_12707_),
    .Y(_12713_),
    .B1(_12712_));
 sg13g2_nand2_1 _19704_ (.Y(_12714_),
    .A(_12386_),
    .B(_12685_));
 sg13g2_o21ai_1 _19705_ (.B1(_12714_),
    .Y(_00463_),
    .A1(net45),
    .A2(_12713_));
 sg13g2_nor2b_1 _19706_ (.A(_12707_),
    .B_N(\cpu.dcache.r_data[4][22] ),
    .Y(_12715_));
 sg13g2_a21oi_1 _19707_ (.A1(net993),
    .A2(_12707_),
    .Y(_12716_),
    .B1(_12715_));
 sg13g2_nand2_1 _19708_ (.Y(_12717_),
    .A(_12390_),
    .B(_12685_));
 sg13g2_o21ai_1 _19709_ (.B1(_12717_),
    .Y(_00464_),
    .A1(net45),
    .A2(_12716_));
 sg13g2_nor2b_1 _19710_ (.A(_12707_),
    .B_N(\cpu.dcache.r_data[4][23] ),
    .Y(_12718_));
 sg13g2_a21oi_1 _19711_ (.A1(net992),
    .A2(_12707_),
    .Y(_12719_),
    .B1(_12718_));
 sg13g2_nand2_1 _19712_ (.Y(_12720_),
    .A(_12256_),
    .B(_12685_));
 sg13g2_o21ai_1 _19713_ (.B1(_12720_),
    .Y(_00465_),
    .A1(net45),
    .A2(_12719_));
 sg13g2_nand2_1 _19714_ (.Y(_12721_),
    .A(net444),
    .B(_12396_));
 sg13g2_buf_2 _19715_ (.A(_12721_),
    .X(_12722_));
 sg13g2_buf_1 _19716_ (.A(_12722_),
    .X(_12723_));
 sg13g2_or2_1 _19717_ (.X(_12724_),
    .B(net663),
    .A(net605));
 sg13g2_buf_1 _19718_ (.A(_12724_),
    .X(_12725_));
 sg13g2_buf_1 _19719_ (.A(_12725_),
    .X(_12726_));
 sg13g2_mux2_1 _19720_ (.A0(net1096),
    .A1(\cpu.dcache.r_data[4][24] ),
    .S(net436),
    .X(_12727_));
 sg13g2_nand2_1 _19721_ (.Y(_12728_),
    .A(_12723_),
    .B(_12727_));
 sg13g2_o21ai_1 _19722_ (.B1(_12728_),
    .Y(_00466_),
    .A1(_12261_),
    .A2(net44));
 sg13g2_mux2_1 _19723_ (.A0(net1095),
    .A1(\cpu.dcache.r_data[4][25] ),
    .S(net436),
    .X(_12729_));
 sg13g2_nand2_1 _19724_ (.Y(_12730_),
    .A(net44),
    .B(_12729_));
 sg13g2_o21ai_1 _19725_ (.B1(_12730_),
    .Y(_00467_),
    .A1(net390),
    .A2(net44));
 sg13g2_mux2_1 _19726_ (.A0(net1098),
    .A1(\cpu.dcache.r_data[4][26] ),
    .S(net436),
    .X(_12731_));
 sg13g2_nand2_1 _19727_ (.Y(_12732_),
    .A(_12722_),
    .B(_12731_));
 sg13g2_o21ai_1 _19728_ (.B1(_12732_),
    .Y(_00468_),
    .A1(net397),
    .A2(net44));
 sg13g2_mux2_1 _19729_ (.A0(net1097),
    .A1(\cpu.dcache.r_data[4][27] ),
    .S(_12725_),
    .X(_12733_));
 sg13g2_nand2_1 _19730_ (.Y(_12734_),
    .A(_12722_),
    .B(_12733_));
 sg13g2_o21ai_1 _19731_ (.B1(_12734_),
    .Y(_00469_),
    .A1(net396),
    .A2(_12723_));
 sg13g2_nor2_2 _19732_ (.A(net605),
    .B(_12283_),
    .Y(_12735_));
 sg13g2_mux2_1 _19733_ (.A0(\cpu.dcache.r_data[4][28] ),
    .A1(_12650_),
    .S(_12735_),
    .X(_12736_));
 sg13g2_nand2_1 _19734_ (.Y(_12737_),
    .A(_12722_),
    .B(_12736_));
 sg13g2_o21ai_1 _19735_ (.B1(_12737_),
    .Y(_00470_),
    .A1(net395),
    .A2(net44));
 sg13g2_mux2_1 _19736_ (.A0(\cpu.dcache.r_data[4][29] ),
    .A1(net1084),
    .S(_12735_),
    .X(_12738_));
 sg13g2_nand2_1 _19737_ (.Y(_12739_),
    .A(_12722_),
    .B(_12738_));
 sg13g2_o21ai_1 _19738_ (.B1(_12739_),
    .Y(_00471_),
    .A1(net394),
    .A2(net44));
 sg13g2_buf_1 _19739_ (.A(_12222_),
    .X(_12740_));
 sg13g2_nor2b_1 _19740_ (.A(_12663_),
    .B_N(\cpu.dcache.r_data[4][2] ),
    .Y(_12741_));
 sg13g2_a21oi_1 _19741_ (.A1(net988),
    .A2(_12663_),
    .Y(_12742_),
    .B1(_12741_));
 sg13g2_nand2_1 _19742_ (.Y(_12743_),
    .A(net895),
    .B(_12660_));
 sg13g2_o21ai_1 _19743_ (.B1(_12743_),
    .Y(_00472_),
    .A1(net47),
    .A2(_12742_));
 sg13g2_mux2_1 _19744_ (.A0(\cpu.dcache.r_data[4][30] ),
    .A1(_12635_),
    .S(_12735_),
    .X(_12744_));
 sg13g2_nand2_1 _19745_ (.Y(_12745_),
    .A(_12722_),
    .B(_12744_));
 sg13g2_o21ai_1 _19746_ (.B1(_12745_),
    .Y(_00473_),
    .A1(net393),
    .A2(net44));
 sg13g2_mux2_1 _19747_ (.A0(\cpu.dcache.r_data[4][31] ),
    .A1(_12638_),
    .S(_12735_),
    .X(_12746_));
 sg13g2_nand2_1 _19748_ (.Y(_12747_),
    .A(_12722_),
    .B(_12746_));
 sg13g2_o21ai_1 _19749_ (.B1(_12747_),
    .Y(_00474_),
    .A1(net392),
    .A2(net44));
 sg13g2_buf_1 _19750_ (.A(net1092),
    .X(_12748_));
 sg13g2_nor2b_1 _19751_ (.A(_12663_),
    .B_N(\cpu.dcache.r_data[4][3] ),
    .Y(_12749_));
 sg13g2_a21oi_1 _19752_ (.A1(net987),
    .A2(_12663_),
    .Y(_12750_),
    .B1(_12749_));
 sg13g2_buf_1 _19753_ (.A(_10208_),
    .X(_12751_));
 sg13g2_nand2_1 _19754_ (.Y(_12752_),
    .A(net986),
    .B(_12660_));
 sg13g2_o21ai_1 _19755_ (.B1(_12752_),
    .Y(_00475_),
    .A1(_12661_),
    .A2(_12750_));
 sg13g2_nor2_1 _19756_ (.A(net605),
    .B(_12300_),
    .Y(_12753_));
 sg13g2_buf_2 _19757_ (.A(_12753_),
    .X(_12754_));
 sg13g2_nor2b_1 _19758_ (.A(_12754_),
    .B_N(\cpu.dcache.r_data[4][4] ),
    .Y(_12755_));
 sg13g2_a21oi_1 _19759_ (.A1(net990),
    .A2(_12754_),
    .Y(_12756_),
    .B1(_12755_));
 sg13g2_nand2_1 _19760_ (.Y(_12757_),
    .A(net997),
    .B(_12660_));
 sg13g2_o21ai_1 _19761_ (.B1(_12757_),
    .Y(_00476_),
    .A1(net47),
    .A2(_12756_));
 sg13g2_nor2b_1 _19762_ (.A(_12754_),
    .B_N(\cpu.dcache.r_data[4][5] ),
    .Y(_12758_));
 sg13g2_a21oi_1 _19763_ (.A1(net989),
    .A2(_12754_),
    .Y(_12759_),
    .B1(_12758_));
 sg13g2_nand2_1 _19764_ (.Y(_12760_),
    .A(net995),
    .B(_12660_));
 sg13g2_o21ai_1 _19765_ (.B1(_12760_),
    .Y(_00477_),
    .A1(net47),
    .A2(_12759_));
 sg13g2_nor2b_1 _19766_ (.A(_12754_),
    .B_N(\cpu.dcache.r_data[4][6] ),
    .Y(_12761_));
 sg13g2_a21oi_1 _19767_ (.A1(net988),
    .A2(_12754_),
    .Y(_12762_),
    .B1(_12761_));
 sg13g2_nand2_1 _19768_ (.Y(_12763_),
    .A(net994),
    .B(_12660_));
 sg13g2_o21ai_1 _19769_ (.B1(_12763_),
    .Y(_00478_),
    .A1(net47),
    .A2(_12762_));
 sg13g2_nor2b_1 _19770_ (.A(_12754_),
    .B_N(\cpu.dcache.r_data[4][7] ),
    .Y(_12764_));
 sg13g2_a21oi_1 _19771_ (.A1(net987),
    .A2(_12754_),
    .Y(_12765_),
    .B1(_12764_));
 sg13g2_nand2_1 _19772_ (.Y(_12766_),
    .A(net999),
    .B(_12660_));
 sg13g2_o21ai_1 _19773_ (.B1(_12766_),
    .Y(_00479_),
    .A1(net47),
    .A2(_12765_));
 sg13g2_mux2_1 _19774_ (.A0(\cpu.dcache.r_data[4][8] ),
    .A1(net1085),
    .S(_12670_),
    .X(_12767_));
 sg13g2_nand2_1 _19775_ (.Y(_12768_),
    .A(_12668_),
    .B(_12767_));
 sg13g2_o21ai_1 _19776_ (.B1(_12768_),
    .Y(_00480_),
    .A1(net391),
    .A2(net46));
 sg13g2_mux2_1 _19777_ (.A0(\cpu.dcache.r_data[4][9] ),
    .A1(_12653_),
    .S(_12670_),
    .X(_12769_));
 sg13g2_nand2_1 _19778_ (.Y(_12770_),
    .A(_12668_),
    .B(_12769_));
 sg13g2_o21ai_1 _19779_ (.B1(_12770_),
    .Y(_00481_),
    .A1(net390),
    .A2(_12669_));
 sg13g2_buf_1 _19780_ (.A(_09836_),
    .X(_12771_));
 sg13g2_nor2_1 _19781_ (.A(net757),
    .B(_12321_),
    .Y(_12772_));
 sg13g2_buf_2 _19782_ (.A(_12772_),
    .X(_12773_));
 sg13g2_buf_1 _19783_ (.A(_12773_),
    .X(_12774_));
 sg13g2_nor2_1 _19784_ (.A(net757),
    .B(_12136_),
    .Y(_12775_));
 sg13g2_buf_2 _19785_ (.A(_12775_),
    .X(_12776_));
 sg13g2_nor2b_1 _19786_ (.A(_12776_),
    .B_N(\cpu.dcache.r_data[5][0] ),
    .Y(_12777_));
 sg13g2_a21oi_1 _19787_ (.A1(net990),
    .A2(_12776_),
    .Y(_12778_),
    .B1(_12777_));
 sg13g2_nand2_1 _19788_ (.Y(_12779_),
    .A(net896),
    .B(net43));
 sg13g2_o21ai_1 _19789_ (.B1(_12779_),
    .Y(_00482_),
    .A1(net43),
    .A2(_12778_));
 sg13g2_buf_1 _19790_ (.A(net702),
    .X(_12780_));
 sg13g2_buf_1 _19791_ (.A(net604),
    .X(_12781_));
 sg13g2_buf_1 _19792_ (.A(_12781_),
    .X(_12782_));
 sg13g2_nand2_1 _19793_ (.Y(_12783_),
    .A(net486),
    .B(_12334_));
 sg13g2_buf_1 _19794_ (.A(_12783_),
    .X(_12784_));
 sg13g2_buf_1 _19795_ (.A(_12784_),
    .X(_12785_));
 sg13g2_nor2_2 _19796_ (.A(net757),
    .B(_12160_),
    .Y(_12786_));
 sg13g2_mux2_1 _19797_ (.A0(\cpu.dcache.r_data[5][10] ),
    .A1(net1087),
    .S(_12786_),
    .X(_12787_));
 sg13g2_nand2_1 _19798_ (.Y(_12788_),
    .A(net42),
    .B(_12787_));
 sg13g2_o21ai_1 _19799_ (.B1(_12788_),
    .Y(_00483_),
    .A1(_12149_),
    .A2(net42));
 sg13g2_mux2_1 _19800_ (.A0(\cpu.dcache.r_data[5][11] ),
    .A1(net1086),
    .S(_12786_),
    .X(_12789_));
 sg13g2_nand2_1 _19801_ (.Y(_12790_),
    .A(net42),
    .B(_12789_));
 sg13g2_o21ai_1 _19802_ (.B1(_12790_),
    .Y(_00484_),
    .A1(_12166_),
    .A2(net42));
 sg13g2_nor2_2 _19803_ (.A(net757),
    .B(_12180_),
    .Y(_12791_));
 sg13g2_mux2_1 _19804_ (.A0(\cpu.dcache.r_data[5][12] ),
    .A1(net1085),
    .S(_12791_),
    .X(_12792_));
 sg13g2_nand2_1 _19805_ (.Y(_12793_),
    .A(_12784_),
    .B(_12792_));
 sg13g2_o21ai_1 _19806_ (.B1(_12793_),
    .Y(_00485_),
    .A1(_12174_),
    .A2(_12785_));
 sg13g2_mux2_1 _19807_ (.A0(\cpu.dcache.r_data[5][13] ),
    .A1(net1084),
    .S(_12791_),
    .X(_12794_));
 sg13g2_nand2_1 _19808_ (.Y(_12795_),
    .A(_12784_),
    .B(_12794_));
 sg13g2_o21ai_1 _19809_ (.B1(_12795_),
    .Y(_00486_),
    .A1(_12186_),
    .A2(_12785_));
 sg13g2_mux2_1 _19810_ (.A0(\cpu.dcache.r_data[5][14] ),
    .A1(net1087),
    .S(_12791_),
    .X(_12796_));
 sg13g2_nand2_1 _19811_ (.Y(_12797_),
    .A(_12784_),
    .B(_12796_));
 sg13g2_o21ai_1 _19812_ (.B1(_12797_),
    .Y(_00487_),
    .A1(_12194_),
    .A2(net42));
 sg13g2_mux2_1 _19813_ (.A0(\cpu.dcache.r_data[5][15] ),
    .A1(net1086),
    .S(_12791_),
    .X(_12798_));
 sg13g2_nand2_1 _19814_ (.Y(_12799_),
    .A(_12784_),
    .B(_12798_));
 sg13g2_o21ai_1 _19815_ (.B1(_12799_),
    .Y(_00488_),
    .A1(_12200_),
    .A2(net42));
 sg13g2_nor2_1 _19816_ (.A(net757),
    .B(_12355_),
    .Y(_12800_));
 sg13g2_buf_2 _19817_ (.A(_12800_),
    .X(_12801_));
 sg13g2_buf_1 _19818_ (.A(_12801_),
    .X(_12802_));
 sg13g2_nor2_1 _19819_ (.A(net757),
    .B(_12210_),
    .Y(_12803_));
 sg13g2_buf_2 _19820_ (.A(_12803_),
    .X(_12804_));
 sg13g2_nor2b_1 _19821_ (.A(_12804_),
    .B_N(\cpu.dcache.r_data[5][16] ),
    .Y(_12805_));
 sg13g2_a21oi_1 _19822_ (.A1(_12705_),
    .A2(_12804_),
    .Y(_12806_),
    .B1(_12805_));
 sg13g2_buf_1 _19823_ (.A(net1041),
    .X(_12807_));
 sg13g2_nand2_1 _19824_ (.Y(_12808_),
    .A(net893),
    .B(net41));
 sg13g2_o21ai_1 _19825_ (.B1(_12808_),
    .Y(_00489_),
    .A1(net41),
    .A2(_12806_));
 sg13g2_nor2b_1 _19826_ (.A(_12804_),
    .B_N(\cpu.dcache.r_data[5][17] ),
    .Y(_12809_));
 sg13g2_a21oi_1 _19827_ (.A1(net989),
    .A2(_12804_),
    .Y(_12810_),
    .B1(_12809_));
 sg13g2_nand2_1 _19828_ (.Y(_12811_),
    .A(net894),
    .B(net41));
 sg13g2_o21ai_1 _19829_ (.B1(_12811_),
    .Y(_00490_),
    .A1(net41),
    .A2(_12810_));
 sg13g2_nor2b_1 _19830_ (.A(_12804_),
    .B_N(\cpu.dcache.r_data[5][18] ),
    .Y(_12812_));
 sg13g2_a21oi_1 _19831_ (.A1(_12740_),
    .A2(_12804_),
    .Y(_12813_),
    .B1(_12812_));
 sg13g2_buf_1 _19832_ (.A(_10201_),
    .X(_12814_));
 sg13g2_nand2_1 _19833_ (.Y(_12815_),
    .A(net892),
    .B(_12801_));
 sg13g2_o21ai_1 _19834_ (.B1(_12815_),
    .Y(_00491_),
    .A1(net41),
    .A2(_12813_));
 sg13g2_nor2b_1 _19835_ (.A(_12804_),
    .B_N(\cpu.dcache.r_data[5][19] ),
    .Y(_12816_));
 sg13g2_a21oi_1 _19836_ (.A1(net987),
    .A2(_12804_),
    .Y(_12817_),
    .B1(_12816_));
 sg13g2_nand2_1 _19837_ (.Y(_12818_),
    .A(net986),
    .B(_12801_));
 sg13g2_o21ai_1 _19838_ (.B1(_12818_),
    .Y(_00492_),
    .A1(net41),
    .A2(_12817_));
 sg13g2_nor2b_1 _19839_ (.A(_12776_),
    .B_N(\cpu.dcache.r_data[5][1] ),
    .Y(_12819_));
 sg13g2_a21oi_1 _19840_ (.A1(net989),
    .A2(_12776_),
    .Y(_12820_),
    .B1(_12819_));
 sg13g2_nand2_1 _19841_ (.Y(_12821_),
    .A(net894),
    .B(net43));
 sg13g2_o21ai_1 _19842_ (.B1(_12821_),
    .Y(_00493_),
    .A1(net43),
    .A2(_12820_));
 sg13g2_nor2_1 _19843_ (.A(_12771_),
    .B(_12239_),
    .Y(_12822_));
 sg13g2_buf_2 _19844_ (.A(_12822_),
    .X(_12823_));
 sg13g2_nor2b_1 _19845_ (.A(_12823_),
    .B_N(\cpu.dcache.r_data[5][20] ),
    .Y(_12824_));
 sg13g2_a21oi_1 _19846_ (.A1(net990),
    .A2(_12823_),
    .Y(_12825_),
    .B1(_12824_));
 sg13g2_nand2_1 _19847_ (.Y(_12826_),
    .A(net997),
    .B(_12801_));
 sg13g2_o21ai_1 _19848_ (.B1(_12826_),
    .Y(_00494_),
    .A1(net41),
    .A2(_12825_));
 sg13g2_nor2b_1 _19849_ (.A(_12823_),
    .B_N(\cpu.dcache.r_data[5][21] ),
    .Y(_12827_));
 sg13g2_a21oi_1 _19850_ (.A1(_12711_),
    .A2(_12823_),
    .Y(_12828_),
    .B1(_12827_));
 sg13g2_nand2_1 _19851_ (.Y(_12829_),
    .A(net995),
    .B(_12801_));
 sg13g2_o21ai_1 _19852_ (.B1(_12829_),
    .Y(_00495_),
    .A1(_12802_),
    .A2(_12828_));
 sg13g2_nor2b_1 _19853_ (.A(_12823_),
    .B_N(\cpu.dcache.r_data[5][22] ),
    .Y(_12830_));
 sg13g2_a21oi_1 _19854_ (.A1(_12740_),
    .A2(_12823_),
    .Y(_12831_),
    .B1(_12830_));
 sg13g2_nand2_1 _19855_ (.Y(_12832_),
    .A(net994),
    .B(_12801_));
 sg13g2_o21ai_1 _19856_ (.B1(_12832_),
    .Y(_00496_),
    .A1(net41),
    .A2(_12831_));
 sg13g2_nor2b_1 _19857_ (.A(_12823_),
    .B_N(\cpu.dcache.r_data[5][23] ),
    .Y(_12833_));
 sg13g2_a21oi_1 _19858_ (.A1(_12748_),
    .A2(_12823_),
    .Y(_12834_),
    .B1(_12833_));
 sg13g2_nand2_1 _19859_ (.Y(_12835_),
    .A(net999),
    .B(_12801_));
 sg13g2_o21ai_1 _19860_ (.B1(_12835_),
    .Y(_00497_),
    .A1(_12802_),
    .A2(_12834_));
 sg13g2_nand2_1 _19861_ (.Y(_12836_),
    .A(net486),
    .B(_12396_));
 sg13g2_buf_2 _19862_ (.A(_12836_),
    .X(_12837_));
 sg13g2_buf_1 _19863_ (.A(_12837_),
    .X(_12838_));
 sg13g2_nor2_1 _19864_ (.A(_09836_),
    .B(_12110_),
    .Y(_12839_));
 sg13g2_buf_2 _19865_ (.A(_12839_),
    .X(_12840_));
 sg13g2_mux2_1 _19866_ (.A0(\cpu.dcache.r_data[5][24] ),
    .A1(net1085),
    .S(_12840_),
    .X(_12841_));
 sg13g2_nand2_1 _19867_ (.Y(_12842_),
    .A(_12838_),
    .B(_12841_));
 sg13g2_o21ai_1 _19868_ (.B1(_12842_),
    .Y(_00498_),
    .A1(_12260_),
    .A2(_12838_));
 sg13g2_mux2_1 _19869_ (.A0(\cpu.dcache.r_data[5][25] ),
    .A1(net1084),
    .S(_12840_),
    .X(_12843_));
 sg13g2_nand2_1 _19870_ (.Y(_02684_),
    .A(net40),
    .B(_12843_));
 sg13g2_o21ai_1 _19871_ (.B1(_02684_),
    .Y(_00499_),
    .A1(_12274_),
    .A2(net40));
 sg13g2_mux2_1 _19872_ (.A0(\cpu.dcache.r_data[5][26] ),
    .A1(_12635_),
    .S(_12840_),
    .X(_02685_));
 sg13g2_nand2_1 _19873_ (.Y(_02686_),
    .A(_12837_),
    .B(_02685_));
 sg13g2_o21ai_1 _19874_ (.B1(_02686_),
    .Y(_00500_),
    .A1(_12149_),
    .A2(net40));
 sg13g2_mux2_1 _19875_ (.A0(\cpu.dcache.r_data[5][27] ),
    .A1(_12638_),
    .S(_12840_),
    .X(_02687_));
 sg13g2_nand2_1 _19876_ (.Y(_02688_),
    .A(_12837_),
    .B(_02687_));
 sg13g2_o21ai_1 _19877_ (.B1(_02688_),
    .Y(_00501_),
    .A1(_12166_),
    .A2(net40));
 sg13g2_nor2_2 _19878_ (.A(net757),
    .B(_12283_),
    .Y(_02689_));
 sg13g2_mux2_1 _19879_ (.A0(\cpu.dcache.r_data[5][28] ),
    .A1(net1085),
    .S(_02689_),
    .X(_02690_));
 sg13g2_nand2_1 _19880_ (.Y(_02691_),
    .A(_12837_),
    .B(_02690_));
 sg13g2_o21ai_1 _19881_ (.B1(_02691_),
    .Y(_00502_),
    .A1(_12174_),
    .A2(net40));
 sg13g2_mux2_1 _19882_ (.A0(\cpu.dcache.r_data[5][29] ),
    .A1(net1084),
    .S(_02689_),
    .X(_02692_));
 sg13g2_nand2_1 _19883_ (.Y(_02693_),
    .A(_12837_),
    .B(_02692_));
 sg13g2_o21ai_1 _19884_ (.B1(_02693_),
    .Y(_00503_),
    .A1(_12186_),
    .A2(net40));
 sg13g2_nor2b_1 _19885_ (.A(_12776_),
    .B_N(\cpu.dcache.r_data[5][2] ),
    .Y(_02694_));
 sg13g2_a21oi_1 _19886_ (.A1(net988),
    .A2(_12776_),
    .Y(_02695_),
    .B1(_02694_));
 sg13g2_nand2_1 _19887_ (.Y(_02696_),
    .A(net892),
    .B(_12773_));
 sg13g2_o21ai_1 _19888_ (.B1(_02696_),
    .Y(_00504_),
    .A1(_12774_),
    .A2(_02695_));
 sg13g2_mux2_1 _19889_ (.A0(\cpu.dcache.r_data[5][30] ),
    .A1(net1087),
    .S(_02689_),
    .X(_02697_));
 sg13g2_nand2_1 _19890_ (.Y(_02698_),
    .A(_12837_),
    .B(_02697_));
 sg13g2_o21ai_1 _19891_ (.B1(_02698_),
    .Y(_00505_),
    .A1(_12194_),
    .A2(net40));
 sg13g2_mux2_1 _19892_ (.A0(\cpu.dcache.r_data[5][31] ),
    .A1(net1086),
    .S(_02689_),
    .X(_02699_));
 sg13g2_nand2_1 _19893_ (.Y(_02700_),
    .A(_12837_),
    .B(_02699_));
 sg13g2_o21ai_1 _19894_ (.B1(_02700_),
    .Y(_00506_),
    .A1(_12200_),
    .A2(net40));
 sg13g2_nor2b_1 _19895_ (.A(_12776_),
    .B_N(\cpu.dcache.r_data[5][3] ),
    .Y(_02701_));
 sg13g2_a21oi_1 _19896_ (.A1(net987),
    .A2(_12776_),
    .Y(_02702_),
    .B1(_02701_));
 sg13g2_nand2_1 _19897_ (.Y(_02703_),
    .A(net986),
    .B(_12773_));
 sg13g2_o21ai_1 _19898_ (.B1(_02703_),
    .Y(_00507_),
    .A1(_12774_),
    .A2(_02702_));
 sg13g2_nor2_1 _19899_ (.A(net757),
    .B(_12300_),
    .Y(_02704_));
 sg13g2_buf_2 _19900_ (.A(_02704_),
    .X(_02705_));
 sg13g2_nor2b_1 _19901_ (.A(_02705_),
    .B_N(\cpu.dcache.r_data[5][4] ),
    .Y(_02706_));
 sg13g2_a21oi_1 _19902_ (.A1(net990),
    .A2(_02705_),
    .Y(_02707_),
    .B1(_02706_));
 sg13g2_nand2_1 _19903_ (.Y(_02708_),
    .A(net997),
    .B(_12773_));
 sg13g2_o21ai_1 _19904_ (.B1(_02708_),
    .Y(_00508_),
    .A1(net43),
    .A2(_02707_));
 sg13g2_nor2b_1 _19905_ (.A(_02705_),
    .B_N(\cpu.dcache.r_data[5][5] ),
    .Y(_02709_));
 sg13g2_a21oi_1 _19906_ (.A1(net989),
    .A2(_02705_),
    .Y(_02710_),
    .B1(_02709_));
 sg13g2_nand2_1 _19907_ (.Y(_02711_),
    .A(net995),
    .B(_12773_));
 sg13g2_o21ai_1 _19908_ (.B1(_02711_),
    .Y(_00509_),
    .A1(net43),
    .A2(_02710_));
 sg13g2_nor2b_1 _19909_ (.A(_02705_),
    .B_N(\cpu.dcache.r_data[5][6] ),
    .Y(_02712_));
 sg13g2_a21oi_1 _19910_ (.A1(net988),
    .A2(_02705_),
    .Y(_02713_),
    .B1(_02712_));
 sg13g2_nand2_1 _19911_ (.Y(_02714_),
    .A(net994),
    .B(_12773_));
 sg13g2_o21ai_1 _19912_ (.B1(_02714_),
    .Y(_00510_),
    .A1(net43),
    .A2(_02713_));
 sg13g2_nor2b_1 _19913_ (.A(_02705_),
    .B_N(\cpu.dcache.r_data[5][7] ),
    .Y(_02715_));
 sg13g2_a21oi_1 _19914_ (.A1(net987),
    .A2(_02705_),
    .Y(_02716_),
    .B1(_02715_));
 sg13g2_nand2_1 _19915_ (.Y(_02717_),
    .A(net999),
    .B(_12773_));
 sg13g2_o21ai_1 _19916_ (.B1(_02717_),
    .Y(_00511_),
    .A1(net43),
    .A2(_02716_));
 sg13g2_mux2_1 _19917_ (.A0(\cpu.dcache.r_data[5][8] ),
    .A1(net1085),
    .S(_12786_),
    .X(_02718_));
 sg13g2_nand2_1 _19918_ (.Y(_02719_),
    .A(_12784_),
    .B(_02718_));
 sg13g2_o21ai_1 _19919_ (.B1(_02719_),
    .Y(_00512_),
    .A1(_12260_),
    .A2(net42));
 sg13g2_mux2_1 _19920_ (.A0(\cpu.dcache.r_data[5][9] ),
    .A1(net1084),
    .S(_12786_),
    .X(_02720_));
 sg13g2_nand2_1 _19921_ (.Y(_02721_),
    .A(_12784_),
    .B(_02720_));
 sg13g2_o21ai_1 _19922_ (.B1(_02721_),
    .Y(_00513_),
    .A1(_12274_),
    .A2(net42));
 sg13g2_buf_1 _19923_ (.A(_09831_),
    .X(_02722_));
 sg13g2_nor2_1 _19924_ (.A(net660),
    .B(_12321_),
    .Y(_02723_));
 sg13g2_buf_2 _19925_ (.A(_02723_),
    .X(_02724_));
 sg13g2_buf_1 _19926_ (.A(_02724_),
    .X(_02725_));
 sg13g2_nor2_1 _19927_ (.A(net660),
    .B(_12136_),
    .Y(_02726_));
 sg13g2_buf_2 _19928_ (.A(_02726_),
    .X(_02727_));
 sg13g2_nor2b_1 _19929_ (.A(_02727_),
    .B_N(\cpu.dcache.r_data[6][0] ),
    .Y(_02728_));
 sg13g2_a21oi_1 _19930_ (.A1(net990),
    .A2(_02727_),
    .Y(_02729_),
    .B1(_02728_));
 sg13g2_nand2_1 _19931_ (.Y(_02730_),
    .A(net893),
    .B(net39));
 sg13g2_o21ai_1 _19932_ (.B1(_02730_),
    .Y(_00514_),
    .A1(net39),
    .A2(_02729_));
 sg13g2_buf_1 _19933_ (.A(net701),
    .X(_02731_));
 sg13g2_buf_1 _19934_ (.A(net603),
    .X(_02732_));
 sg13g2_buf_1 _19935_ (.A(net528),
    .X(_02733_));
 sg13g2_buf_1 _19936_ (.A(net485),
    .X(_02734_));
 sg13g2_nand2_1 _19937_ (.Y(_02735_),
    .A(net435),
    .B(_12334_));
 sg13g2_buf_2 _19938_ (.A(_02735_),
    .X(_02736_));
 sg13g2_buf_1 _19939_ (.A(_02736_),
    .X(_02737_));
 sg13g2_nor2_2 _19940_ (.A(net660),
    .B(_12160_),
    .Y(_02738_));
 sg13g2_mux2_1 _19941_ (.A0(\cpu.dcache.r_data[6][10] ),
    .A1(net1087),
    .S(_02738_),
    .X(_02739_));
 sg13g2_nand2_1 _19942_ (.Y(_02740_),
    .A(net38),
    .B(_02739_));
 sg13g2_o21ai_1 _19943_ (.B1(_02740_),
    .Y(_00515_),
    .A1(_12149_),
    .A2(net38));
 sg13g2_mux2_1 _19944_ (.A0(\cpu.dcache.r_data[6][11] ),
    .A1(net1086),
    .S(_02738_),
    .X(_02741_));
 sg13g2_nand2_1 _19945_ (.Y(_02742_),
    .A(net38),
    .B(_02741_));
 sg13g2_o21ai_1 _19946_ (.B1(_02742_),
    .Y(_00516_),
    .A1(_12166_),
    .A2(net38));
 sg13g2_nor2_2 _19947_ (.A(net660),
    .B(_12180_),
    .Y(_02743_));
 sg13g2_mux2_1 _19948_ (.A0(\cpu.dcache.r_data[6][12] ),
    .A1(net1085),
    .S(_02743_),
    .X(_02744_));
 sg13g2_nand2_1 _19949_ (.Y(_02745_),
    .A(_02736_),
    .B(_02744_));
 sg13g2_o21ai_1 _19950_ (.B1(_02745_),
    .Y(_00517_),
    .A1(_12174_),
    .A2(net38));
 sg13g2_mux2_1 _19951_ (.A0(\cpu.dcache.r_data[6][13] ),
    .A1(net1084),
    .S(_02743_),
    .X(_02746_));
 sg13g2_nand2_1 _19952_ (.Y(_02747_),
    .A(_02736_),
    .B(_02746_));
 sg13g2_o21ai_1 _19953_ (.B1(_02747_),
    .Y(_00518_),
    .A1(_12186_),
    .A2(_02737_));
 sg13g2_mux2_1 _19954_ (.A0(\cpu.dcache.r_data[6][14] ),
    .A1(net1087),
    .S(_02743_),
    .X(_02748_));
 sg13g2_nand2_1 _19955_ (.Y(_02749_),
    .A(_02736_),
    .B(_02748_));
 sg13g2_o21ai_1 _19956_ (.B1(_02749_),
    .Y(_00519_),
    .A1(_12194_),
    .A2(net38));
 sg13g2_mux2_1 _19957_ (.A0(\cpu.dcache.r_data[6][15] ),
    .A1(net1086),
    .S(_02743_),
    .X(_02750_));
 sg13g2_nand2_1 _19958_ (.Y(_02751_),
    .A(_02736_),
    .B(_02750_));
 sg13g2_o21ai_1 _19959_ (.B1(_02751_),
    .Y(_00520_),
    .A1(_12200_),
    .A2(net38));
 sg13g2_nor2_1 _19960_ (.A(net660),
    .B(_12355_),
    .Y(_02752_));
 sg13g2_buf_2 _19961_ (.A(_02752_),
    .X(_02753_));
 sg13g2_buf_1 _19962_ (.A(_02753_),
    .X(_02754_));
 sg13g2_nor2_1 _19963_ (.A(_02722_),
    .B(_12210_),
    .Y(_02755_));
 sg13g2_buf_2 _19964_ (.A(_02755_),
    .X(_02756_));
 sg13g2_nor2b_1 _19965_ (.A(_02756_),
    .B_N(\cpu.dcache.r_data[6][16] ),
    .Y(_02757_));
 sg13g2_a21oi_1 _19966_ (.A1(net990),
    .A2(_02756_),
    .Y(_02758_),
    .B1(_02757_));
 sg13g2_nand2_1 _19967_ (.Y(_02759_),
    .A(net893),
    .B(net37));
 sg13g2_o21ai_1 _19968_ (.B1(_02759_),
    .Y(_00521_),
    .A1(net37),
    .A2(_02758_));
 sg13g2_nor2b_1 _19969_ (.A(_02756_),
    .B_N(\cpu.dcache.r_data[6][17] ),
    .Y(_02760_));
 sg13g2_a21oi_1 _19970_ (.A1(net989),
    .A2(_02756_),
    .Y(_02761_),
    .B1(_02760_));
 sg13g2_nand2_1 _19971_ (.Y(_02762_),
    .A(net894),
    .B(net37));
 sg13g2_o21ai_1 _19972_ (.B1(_02762_),
    .Y(_00522_),
    .A1(net37),
    .A2(_02761_));
 sg13g2_nor2b_1 _19973_ (.A(_02756_),
    .B_N(\cpu.dcache.r_data[6][18] ),
    .Y(_02763_));
 sg13g2_a21oi_1 _19974_ (.A1(net988),
    .A2(_02756_),
    .Y(_02764_),
    .B1(_02763_));
 sg13g2_nand2_1 _19975_ (.Y(_02765_),
    .A(net892),
    .B(_02753_));
 sg13g2_o21ai_1 _19976_ (.B1(_02765_),
    .Y(_00523_),
    .A1(net37),
    .A2(_02764_));
 sg13g2_nor2b_1 _19977_ (.A(_02756_),
    .B_N(\cpu.dcache.r_data[6][19] ),
    .Y(_02766_));
 sg13g2_a21oi_1 _19978_ (.A1(net987),
    .A2(_02756_),
    .Y(_02767_),
    .B1(_02766_));
 sg13g2_nand2_1 _19979_ (.Y(_02768_),
    .A(net986),
    .B(_02753_));
 sg13g2_o21ai_1 _19980_ (.B1(_02768_),
    .Y(_00524_),
    .A1(net37),
    .A2(_02767_));
 sg13g2_nor2b_1 _19981_ (.A(_02727_),
    .B_N(\cpu.dcache.r_data[6][1] ),
    .Y(_02769_));
 sg13g2_a21oi_1 _19982_ (.A1(net989),
    .A2(_02727_),
    .Y(_02770_),
    .B1(_02769_));
 sg13g2_nand2_1 _19983_ (.Y(_02771_),
    .A(net894),
    .B(net39));
 sg13g2_o21ai_1 _19984_ (.B1(_02771_),
    .Y(_00525_),
    .A1(net39),
    .A2(_02770_));
 sg13g2_nor2_1 _19985_ (.A(net660),
    .B(_12239_),
    .Y(_02772_));
 sg13g2_buf_2 _19986_ (.A(_02772_),
    .X(_02773_));
 sg13g2_nor2b_1 _19987_ (.A(_02773_),
    .B_N(\cpu.dcache.r_data[6][20] ),
    .Y(_02774_));
 sg13g2_a21oi_1 _19988_ (.A1(net990),
    .A2(_02773_),
    .Y(_02775_),
    .B1(_02774_));
 sg13g2_nand2_1 _19989_ (.Y(_02776_),
    .A(net997),
    .B(_02753_));
 sg13g2_o21ai_1 _19990_ (.B1(_02776_),
    .Y(_00526_),
    .A1(_02754_),
    .A2(_02775_));
 sg13g2_nor2b_1 _19991_ (.A(_02773_),
    .B_N(\cpu.dcache.r_data[6][21] ),
    .Y(_02777_));
 sg13g2_a21oi_1 _19992_ (.A1(net989),
    .A2(_02773_),
    .Y(_02778_),
    .B1(_02777_));
 sg13g2_nand2_1 _19993_ (.Y(_02779_),
    .A(net995),
    .B(_02753_));
 sg13g2_o21ai_1 _19994_ (.B1(_02779_),
    .Y(_00527_),
    .A1(_02754_),
    .A2(_02778_));
 sg13g2_nor2b_1 _19995_ (.A(_02773_),
    .B_N(\cpu.dcache.r_data[6][22] ),
    .Y(_02780_));
 sg13g2_a21oi_1 _19996_ (.A1(net988),
    .A2(_02773_),
    .Y(_02781_),
    .B1(_02780_));
 sg13g2_nand2_1 _19997_ (.Y(_02782_),
    .A(net994),
    .B(_02753_));
 sg13g2_o21ai_1 _19998_ (.B1(_02782_),
    .Y(_00528_),
    .A1(net37),
    .A2(_02781_));
 sg13g2_nor2b_1 _19999_ (.A(_02773_),
    .B_N(\cpu.dcache.r_data[6][23] ),
    .Y(_02783_));
 sg13g2_a21oi_1 _20000_ (.A1(_12748_),
    .A2(_02773_),
    .Y(_02784_),
    .B1(_02783_));
 sg13g2_buf_1 _20001_ (.A(_10229_),
    .X(_02785_));
 sg13g2_nand2_1 _20002_ (.Y(_02786_),
    .A(net985),
    .B(_02753_));
 sg13g2_o21ai_1 _20003_ (.B1(_02786_),
    .Y(_00529_),
    .A1(net37),
    .A2(_02784_));
 sg13g2_nand2_1 _20004_ (.Y(_02787_),
    .A(net435),
    .B(_12396_));
 sg13g2_buf_2 _20005_ (.A(_02787_),
    .X(_02788_));
 sg13g2_buf_1 _20006_ (.A(_02788_),
    .X(_02789_));
 sg13g2_nor2_1 _20007_ (.A(_09831_),
    .B(_12110_),
    .Y(_02790_));
 sg13g2_buf_2 _20008_ (.A(_02790_),
    .X(_02791_));
 sg13g2_mux2_1 _20009_ (.A0(\cpu.dcache.r_data[6][24] ),
    .A1(_12650_),
    .S(_02791_),
    .X(_02792_));
 sg13g2_nand2_1 _20010_ (.Y(_02793_),
    .A(net36),
    .B(_02792_));
 sg13g2_o21ai_1 _20011_ (.B1(_02793_),
    .Y(_00530_),
    .A1(_12260_),
    .A2(net36));
 sg13g2_mux2_1 _20012_ (.A0(\cpu.dcache.r_data[6][25] ),
    .A1(net1084),
    .S(_02791_),
    .X(_02794_));
 sg13g2_nand2_1 _20013_ (.Y(_02795_),
    .A(_02789_),
    .B(_02794_));
 sg13g2_o21ai_1 _20014_ (.B1(_02795_),
    .Y(_00531_),
    .A1(_12274_),
    .A2(net36));
 sg13g2_mux2_1 _20015_ (.A0(\cpu.dcache.r_data[6][26] ),
    .A1(net1093),
    .S(_02791_),
    .X(_02796_));
 sg13g2_nand2_1 _20016_ (.Y(_02797_),
    .A(_02788_),
    .B(_02796_));
 sg13g2_o21ai_1 _20017_ (.B1(_02797_),
    .Y(_00532_),
    .A1(_12149_),
    .A2(net36));
 sg13g2_mux2_1 _20018_ (.A0(\cpu.dcache.r_data[6][27] ),
    .A1(net1092),
    .S(_02791_),
    .X(_02798_));
 sg13g2_nand2_1 _20019_ (.Y(_02799_),
    .A(_02788_),
    .B(_02798_));
 sg13g2_o21ai_1 _20020_ (.B1(_02799_),
    .Y(_00533_),
    .A1(_12166_),
    .A2(_02789_));
 sg13g2_nor2_2 _20021_ (.A(net660),
    .B(_12283_),
    .Y(_02800_));
 sg13g2_mux2_1 _20022_ (.A0(\cpu.dcache.r_data[6][28] ),
    .A1(net1101),
    .S(_02800_),
    .X(_02801_));
 sg13g2_nand2_1 _20023_ (.Y(_02802_),
    .A(_02788_),
    .B(_02801_));
 sg13g2_o21ai_1 _20024_ (.B1(_02802_),
    .Y(_00534_),
    .A1(_12174_),
    .A2(net36));
 sg13g2_mux2_1 _20025_ (.A0(\cpu.dcache.r_data[6][29] ),
    .A1(net1094),
    .S(_02800_),
    .X(_02803_));
 sg13g2_nand2_1 _20026_ (.Y(_02804_),
    .A(_02788_),
    .B(_02803_));
 sg13g2_o21ai_1 _20027_ (.B1(_02804_),
    .Y(_00535_),
    .A1(_12186_),
    .A2(net36));
 sg13g2_nor2b_1 _20028_ (.A(_02727_),
    .B_N(\cpu.dcache.r_data[6][2] ),
    .Y(_02805_));
 sg13g2_a21oi_1 _20029_ (.A1(net988),
    .A2(_02727_),
    .Y(_02806_),
    .B1(_02805_));
 sg13g2_nand2_1 _20030_ (.Y(_02807_),
    .A(net892),
    .B(_02724_));
 sg13g2_o21ai_1 _20031_ (.B1(_02807_),
    .Y(_00536_),
    .A1(_02725_),
    .A2(_02806_));
 sg13g2_mux2_1 _20032_ (.A0(\cpu.dcache.r_data[6][30] ),
    .A1(net1093),
    .S(_02800_),
    .X(_02808_));
 sg13g2_nand2_1 _20033_ (.Y(_02809_),
    .A(_02788_),
    .B(_02808_));
 sg13g2_o21ai_1 _20034_ (.B1(_02809_),
    .Y(_00537_),
    .A1(_12194_),
    .A2(net36));
 sg13g2_mux2_1 _20035_ (.A0(\cpu.dcache.r_data[6][31] ),
    .A1(net1092),
    .S(_02800_),
    .X(_02810_));
 sg13g2_nand2_1 _20036_ (.Y(_02811_),
    .A(_02788_),
    .B(_02810_));
 sg13g2_o21ai_1 _20037_ (.B1(_02811_),
    .Y(_00538_),
    .A1(_12200_),
    .A2(net36));
 sg13g2_nor2b_1 _20038_ (.A(_02727_),
    .B_N(\cpu.dcache.r_data[6][3] ),
    .Y(_02812_));
 sg13g2_a21oi_1 _20039_ (.A1(net987),
    .A2(_02727_),
    .Y(_02813_),
    .B1(_02812_));
 sg13g2_nand2_1 _20040_ (.Y(_02814_),
    .A(net986),
    .B(_02724_));
 sg13g2_o21ai_1 _20041_ (.B1(_02814_),
    .Y(_00539_),
    .A1(_02725_),
    .A2(_02813_));
 sg13g2_nor2_1 _20042_ (.A(net660),
    .B(_12300_),
    .Y(_02815_));
 sg13g2_buf_2 _20043_ (.A(_02815_),
    .X(_02816_));
 sg13g2_nor2b_1 _20044_ (.A(_02816_),
    .B_N(\cpu.dcache.r_data[6][4] ),
    .Y(_02817_));
 sg13g2_a21oi_1 _20045_ (.A1(net990),
    .A2(_02816_),
    .Y(_02818_),
    .B1(_02817_));
 sg13g2_nand2_1 _20046_ (.Y(_02819_),
    .A(net997),
    .B(_02724_));
 sg13g2_o21ai_1 _20047_ (.B1(_02819_),
    .Y(_00540_),
    .A1(net39),
    .A2(_02818_));
 sg13g2_nor2b_1 _20048_ (.A(_02816_),
    .B_N(\cpu.dcache.r_data[6][5] ),
    .Y(_02820_));
 sg13g2_a21oi_1 _20049_ (.A1(net989),
    .A2(_02816_),
    .Y(_02821_),
    .B1(_02820_));
 sg13g2_nand2_1 _20050_ (.Y(_02822_),
    .A(net995),
    .B(_02724_));
 sg13g2_o21ai_1 _20051_ (.B1(_02822_),
    .Y(_00541_),
    .A1(net39),
    .A2(_02821_));
 sg13g2_nor2b_1 _20052_ (.A(_02816_),
    .B_N(\cpu.dcache.r_data[6][6] ),
    .Y(_02823_));
 sg13g2_a21oi_1 _20053_ (.A1(net988),
    .A2(_02816_),
    .Y(_02824_),
    .B1(_02823_));
 sg13g2_nand2_1 _20054_ (.Y(_02825_),
    .A(net994),
    .B(_02724_));
 sg13g2_o21ai_1 _20055_ (.B1(_02825_),
    .Y(_00542_),
    .A1(net39),
    .A2(_02824_));
 sg13g2_nor2b_1 _20056_ (.A(_02816_),
    .B_N(\cpu.dcache.r_data[6][7] ),
    .Y(_02826_));
 sg13g2_a21oi_1 _20057_ (.A1(net987),
    .A2(_02816_),
    .Y(_02827_),
    .B1(_02826_));
 sg13g2_nand2_1 _20058_ (.Y(_02828_),
    .A(net985),
    .B(_02724_));
 sg13g2_o21ai_1 _20059_ (.B1(_02828_),
    .Y(_00543_),
    .A1(net39),
    .A2(_02827_));
 sg13g2_mux2_1 _20060_ (.A0(\cpu.dcache.r_data[6][8] ),
    .A1(net1101),
    .S(_02738_),
    .X(_02829_));
 sg13g2_nand2_1 _20061_ (.Y(_02830_),
    .A(_02736_),
    .B(_02829_));
 sg13g2_o21ai_1 _20062_ (.B1(_02830_),
    .Y(_00544_),
    .A1(_12260_),
    .A2(net38));
 sg13g2_mux2_1 _20063_ (.A0(\cpu.dcache.r_data[6][9] ),
    .A1(net1094),
    .S(_02738_),
    .X(_02831_));
 sg13g2_nand2_1 _20064_ (.Y(_02832_),
    .A(_02736_),
    .B(_02831_));
 sg13g2_o21ai_1 _20065_ (.B1(_02832_),
    .Y(_00545_),
    .A1(_12274_),
    .A2(_02737_));
 sg13g2_buf_1 _20066_ (.A(_10178_),
    .X(_02833_));
 sg13g2_nor2_1 _20067_ (.A(net345),
    .B(_12321_),
    .Y(_02834_));
 sg13g2_buf_1 _20068_ (.A(_02834_),
    .X(_02835_));
 sg13g2_buf_2 _20069_ (.A(net1101),
    .X(_02836_));
 sg13g2_nor2_1 _20070_ (.A(net345),
    .B(_12136_),
    .Y(_02837_));
 sg13g2_buf_2 _20071_ (.A(_02837_),
    .X(_02838_));
 sg13g2_nor2b_1 _20072_ (.A(_02838_),
    .B_N(\cpu.dcache.r_data[7][0] ),
    .Y(_02839_));
 sg13g2_a21oi_1 _20073_ (.A1(_02836_),
    .A2(_02838_),
    .Y(_02840_),
    .B1(_02839_));
 sg13g2_nand2_1 _20074_ (.Y(_02841_),
    .A(net893),
    .B(net67));
 sg13g2_o21ai_1 _20075_ (.B1(_02841_),
    .Y(_00546_),
    .A1(net67),
    .A2(_02840_));
 sg13g2_nand2_1 _20076_ (.Y(_02842_),
    .A(net445),
    .B(_12334_));
 sg13g2_buf_1 _20077_ (.A(_02842_),
    .X(_02843_));
 sg13g2_buf_1 _20078_ (.A(_02843_),
    .X(_02844_));
 sg13g2_nor2_2 _20079_ (.A(net345),
    .B(_12160_),
    .Y(_02845_));
 sg13g2_mux2_1 _20080_ (.A0(\cpu.dcache.r_data[7][10] ),
    .A1(net1093),
    .S(_02845_),
    .X(_02846_));
 sg13g2_nand2_1 _20081_ (.Y(_02847_),
    .A(net35),
    .B(_02846_));
 sg13g2_o21ai_1 _20082_ (.B1(_02847_),
    .Y(_00547_),
    .A1(_12149_),
    .A2(net35));
 sg13g2_mux2_1 _20083_ (.A0(\cpu.dcache.r_data[7][11] ),
    .A1(net1092),
    .S(_02845_),
    .X(_02848_));
 sg13g2_nand2_1 _20084_ (.Y(_02849_),
    .A(net35),
    .B(_02848_));
 sg13g2_o21ai_1 _20085_ (.B1(_02849_),
    .Y(_00548_),
    .A1(_12166_),
    .A2(net35));
 sg13g2_nor2_2 _20086_ (.A(net345),
    .B(_12180_),
    .Y(_02850_));
 sg13g2_mux2_1 _20087_ (.A0(\cpu.dcache.r_data[7][12] ),
    .A1(net1101),
    .S(_02850_),
    .X(_02851_));
 sg13g2_nand2_1 _20088_ (.Y(_02852_),
    .A(_02843_),
    .B(_02851_));
 sg13g2_o21ai_1 _20089_ (.B1(_02852_),
    .Y(_00549_),
    .A1(_12174_),
    .A2(net35));
 sg13g2_mux2_1 _20090_ (.A0(\cpu.dcache.r_data[7][13] ),
    .A1(net1094),
    .S(_02850_),
    .X(_02853_));
 sg13g2_nand2_1 _20091_ (.Y(_02854_),
    .A(_02843_),
    .B(_02853_));
 sg13g2_o21ai_1 _20092_ (.B1(_02854_),
    .Y(_00550_),
    .A1(_12186_),
    .A2(net35));
 sg13g2_mux2_1 _20093_ (.A0(\cpu.dcache.r_data[7][14] ),
    .A1(net1093),
    .S(_02850_),
    .X(_02855_));
 sg13g2_nand2_1 _20094_ (.Y(_02856_),
    .A(_02843_),
    .B(_02855_));
 sg13g2_o21ai_1 _20095_ (.B1(_02856_),
    .Y(_00551_),
    .A1(_12194_),
    .A2(_02844_));
 sg13g2_mux2_1 _20096_ (.A0(\cpu.dcache.r_data[7][15] ),
    .A1(net1092),
    .S(_02850_),
    .X(_02857_));
 sg13g2_nand2_1 _20097_ (.Y(_02858_),
    .A(_02843_),
    .B(_02857_));
 sg13g2_o21ai_1 _20098_ (.B1(_02858_),
    .Y(_00552_),
    .A1(_12200_),
    .A2(net35));
 sg13g2_nor2_1 _20099_ (.A(net345),
    .B(_12355_),
    .Y(_02859_));
 sg13g2_buf_1 _20100_ (.A(_02859_),
    .X(_02860_));
 sg13g2_nor2_1 _20101_ (.A(_02833_),
    .B(_12210_),
    .Y(_02861_));
 sg13g2_buf_2 _20102_ (.A(_02861_),
    .X(_02862_));
 sg13g2_nor2b_1 _20103_ (.A(_02862_),
    .B_N(\cpu.dcache.r_data[7][16] ),
    .Y(_02863_));
 sg13g2_a21oi_1 _20104_ (.A1(_02836_),
    .A2(_02862_),
    .Y(_02864_),
    .B1(_02863_));
 sg13g2_nand2_1 _20105_ (.Y(_02865_),
    .A(net893),
    .B(net66));
 sg13g2_o21ai_1 _20106_ (.B1(_02865_),
    .Y(_00553_),
    .A1(net66),
    .A2(_02864_));
 sg13g2_buf_2 _20107_ (.A(net1094),
    .X(_02866_));
 sg13g2_nor2b_1 _20108_ (.A(_02862_),
    .B_N(\cpu.dcache.r_data[7][17] ),
    .Y(_02867_));
 sg13g2_a21oi_1 _20109_ (.A1(_02866_),
    .A2(_02862_),
    .Y(_02868_),
    .B1(_02867_));
 sg13g2_nand2_1 _20110_ (.Y(_02869_),
    .A(net894),
    .B(net66));
 sg13g2_o21ai_1 _20111_ (.B1(_02869_),
    .Y(_00554_),
    .A1(net66),
    .A2(_02868_));
 sg13g2_buf_2 _20112_ (.A(net1093),
    .X(_02870_));
 sg13g2_nor2b_1 _20113_ (.A(_02862_),
    .B_N(\cpu.dcache.r_data[7][18] ),
    .Y(_02871_));
 sg13g2_a21oi_1 _20114_ (.A1(_02870_),
    .A2(_02862_),
    .Y(_02872_),
    .B1(_02871_));
 sg13g2_nand2_1 _20115_ (.Y(_02873_),
    .A(net892),
    .B(_02859_));
 sg13g2_o21ai_1 _20116_ (.B1(_02873_),
    .Y(_00555_),
    .A1(net66),
    .A2(_02872_));
 sg13g2_buf_2 _20117_ (.A(_12228_),
    .X(_02874_));
 sg13g2_nor2b_1 _20118_ (.A(_02862_),
    .B_N(\cpu.dcache.r_data[7][19] ),
    .Y(_02875_));
 sg13g2_a21oi_1 _20119_ (.A1(_02874_),
    .A2(_02862_),
    .Y(_02876_),
    .B1(_02875_));
 sg13g2_nand2_1 _20120_ (.Y(_02877_),
    .A(net986),
    .B(_02859_));
 sg13g2_o21ai_1 _20121_ (.B1(_02877_),
    .Y(_00556_),
    .A1(net66),
    .A2(_02876_));
 sg13g2_nor2b_1 _20122_ (.A(_02838_),
    .B_N(\cpu.dcache.r_data[7][1] ),
    .Y(_02878_));
 sg13g2_a21oi_1 _20123_ (.A1(_02866_),
    .A2(_02838_),
    .Y(_02879_),
    .B1(_02878_));
 sg13g2_nand2_1 _20124_ (.Y(_02880_),
    .A(net894),
    .B(net67));
 sg13g2_o21ai_1 _20125_ (.B1(_02880_),
    .Y(_00557_),
    .A1(net67),
    .A2(_02879_));
 sg13g2_or2_1 _20126_ (.X(_02881_),
    .B(_12239_),
    .A(net345));
 sg13g2_buf_1 _20127_ (.A(_02881_),
    .X(_02882_));
 sg13g2_mux2_1 _20128_ (.A0(_12176_),
    .A1(\cpu.dcache.r_data[7][20] ),
    .S(_02882_),
    .X(_02883_));
 sg13g2_mux2_1 _20129_ (.A0(_02883_),
    .A1(_12244_),
    .S(_02860_),
    .X(_00558_));
 sg13g2_mux2_1 _20130_ (.A0(_12189_),
    .A1(\cpu.dcache.r_data[7][21] ),
    .S(_02882_),
    .X(_02884_));
 sg13g2_mux2_1 _20131_ (.A0(_02884_),
    .A1(_12248_),
    .S(_02860_),
    .X(_00559_));
 sg13g2_mux2_1 _20132_ (.A0(_12158_),
    .A1(\cpu.dcache.r_data[7][22] ),
    .S(_02882_),
    .X(_02885_));
 sg13g2_mux2_1 _20133_ (.A0(_02885_),
    .A1(_12252_),
    .S(net66),
    .X(_00560_));
 sg13g2_mux2_1 _20134_ (.A0(_12169_),
    .A1(\cpu.dcache.r_data[7][23] ),
    .S(_02882_),
    .X(_02886_));
 sg13g2_mux2_1 _20135_ (.A0(_02886_),
    .A1(_12613_),
    .S(net66),
    .X(_00561_));
 sg13g2_nand2_1 _20136_ (.Y(_02887_),
    .A(net445),
    .B(_12396_));
 sg13g2_buf_2 _20137_ (.A(_02887_),
    .X(_02888_));
 sg13g2_buf_1 _20138_ (.A(_02888_),
    .X(_02889_));
 sg13g2_nor2_1 _20139_ (.A(_10178_),
    .B(net663),
    .Y(_02890_));
 sg13g2_buf_2 _20140_ (.A(_02890_),
    .X(_02891_));
 sg13g2_mux2_1 _20141_ (.A0(\cpu.dcache.r_data[7][24] ),
    .A1(net1101),
    .S(_02891_),
    .X(_02892_));
 sg13g2_nand2_1 _20142_ (.Y(_02893_),
    .A(_02889_),
    .B(_02892_));
 sg13g2_o21ai_1 _20143_ (.B1(_02893_),
    .Y(_00562_),
    .A1(_12260_),
    .A2(_02889_));
 sg13g2_mux2_1 _20144_ (.A0(\cpu.dcache.r_data[7][25] ),
    .A1(_12217_),
    .S(_02891_),
    .X(_02894_));
 sg13g2_nand2_1 _20145_ (.Y(_02895_),
    .A(net34),
    .B(_02894_));
 sg13g2_o21ai_1 _20146_ (.B1(_02895_),
    .Y(_00563_),
    .A1(_12274_),
    .A2(net34));
 sg13g2_mux2_1 _20147_ (.A0(\cpu.dcache.r_data[7][26] ),
    .A1(net1093),
    .S(_02891_),
    .X(_02896_));
 sg13g2_nand2_1 _20148_ (.Y(_02897_),
    .A(_02888_),
    .B(_02896_));
 sg13g2_o21ai_1 _20149_ (.B1(_02897_),
    .Y(_00564_),
    .A1(_12149_),
    .A2(net34));
 sg13g2_mux2_1 _20150_ (.A0(\cpu.dcache.r_data[7][27] ),
    .A1(net1092),
    .S(_02891_),
    .X(_02898_));
 sg13g2_nand2_1 _20151_ (.Y(_02899_),
    .A(_02888_),
    .B(_02898_));
 sg13g2_o21ai_1 _20152_ (.B1(_02899_),
    .Y(_00565_),
    .A1(_12166_),
    .A2(net34));
 sg13g2_nor2_2 _20153_ (.A(net345),
    .B(_12283_),
    .Y(_02900_));
 sg13g2_mux2_1 _20154_ (.A0(\cpu.dcache.r_data[7][28] ),
    .A1(net1101),
    .S(_02900_),
    .X(_02901_));
 sg13g2_nand2_1 _20155_ (.Y(_02902_),
    .A(_02888_),
    .B(_02901_));
 sg13g2_o21ai_1 _20156_ (.B1(_02902_),
    .Y(_00566_),
    .A1(_12174_),
    .A2(net34));
 sg13g2_mux2_1 _20157_ (.A0(\cpu.dcache.r_data[7][29] ),
    .A1(net1094),
    .S(_02900_),
    .X(_02903_));
 sg13g2_nand2_1 _20158_ (.Y(_02904_),
    .A(_02888_),
    .B(_02903_));
 sg13g2_o21ai_1 _20159_ (.B1(_02904_),
    .Y(_00567_),
    .A1(_12186_),
    .A2(net34));
 sg13g2_nor2b_1 _20160_ (.A(_02838_),
    .B_N(\cpu.dcache.r_data[7][2] ),
    .Y(_02905_));
 sg13g2_a21oi_1 _20161_ (.A1(_02870_),
    .A2(_02838_),
    .Y(_02906_),
    .B1(_02905_));
 sg13g2_nand2_1 _20162_ (.Y(_02907_),
    .A(net892),
    .B(_02834_));
 sg13g2_o21ai_1 _20163_ (.B1(_02907_),
    .Y(_00568_),
    .A1(_02835_),
    .A2(_02906_));
 sg13g2_mux2_1 _20164_ (.A0(\cpu.dcache.r_data[7][30] ),
    .A1(net1093),
    .S(_02900_),
    .X(_02908_));
 sg13g2_nand2_1 _20165_ (.Y(_02909_),
    .A(_02888_),
    .B(_02908_));
 sg13g2_o21ai_1 _20166_ (.B1(_02909_),
    .Y(_00569_),
    .A1(_12194_),
    .A2(net34));
 sg13g2_mux2_1 _20167_ (.A0(\cpu.dcache.r_data[7][31] ),
    .A1(net1092),
    .S(_02900_),
    .X(_02910_));
 sg13g2_nand2_1 _20168_ (.Y(_02911_),
    .A(_02888_),
    .B(_02910_));
 sg13g2_o21ai_1 _20169_ (.B1(_02911_),
    .Y(_00570_),
    .A1(_12200_),
    .A2(net34));
 sg13g2_nor2b_1 _20170_ (.A(_02838_),
    .B_N(\cpu.dcache.r_data[7][3] ),
    .Y(_02912_));
 sg13g2_a21oi_1 _20171_ (.A1(_02874_),
    .A2(_02838_),
    .Y(_02913_),
    .B1(_02912_));
 sg13g2_nand2_1 _20172_ (.Y(_02914_),
    .A(net986),
    .B(_02834_));
 sg13g2_o21ai_1 _20173_ (.B1(_02914_),
    .Y(_00571_),
    .A1(_02835_),
    .A2(_02913_));
 sg13g2_or2_1 _20174_ (.X(_02915_),
    .B(_12300_),
    .A(net345));
 sg13g2_buf_1 _20175_ (.A(_02915_),
    .X(_02916_));
 sg13g2_mux2_1 _20176_ (.A0(net1096),
    .A1(\cpu.dcache.r_data[7][4] ),
    .S(_02916_),
    .X(_02917_));
 sg13g2_mux2_1 _20177_ (.A0(_02917_),
    .A1(_12244_),
    .S(net67),
    .X(_00572_));
 sg13g2_mux2_1 _20178_ (.A0(net1095),
    .A1(\cpu.dcache.r_data[7][5] ),
    .S(_02916_),
    .X(_02918_));
 sg13g2_mux2_1 _20179_ (.A0(_02918_),
    .A1(_12248_),
    .S(net67),
    .X(_00573_));
 sg13g2_mux2_1 _20180_ (.A0(net1098),
    .A1(\cpu.dcache.r_data[7][6] ),
    .S(_02916_),
    .X(_02919_));
 sg13g2_mux2_1 _20181_ (.A0(_02919_),
    .A1(_12252_),
    .S(net67),
    .X(_00574_));
 sg13g2_mux2_1 _20182_ (.A0(net1097),
    .A1(\cpu.dcache.r_data[7][7] ),
    .S(_02916_),
    .X(_02920_));
 sg13g2_mux2_1 _20183_ (.A0(_02920_),
    .A1(_12613_),
    .S(net67),
    .X(_00575_));
 sg13g2_mux2_1 _20184_ (.A0(\cpu.dcache.r_data[7][8] ),
    .A1(net1101),
    .S(_02845_),
    .X(_02921_));
 sg13g2_nand2_1 _20185_ (.Y(_02922_),
    .A(_02843_),
    .B(_02921_));
 sg13g2_o21ai_1 _20186_ (.B1(_02922_),
    .Y(_00576_),
    .A1(_12260_),
    .A2(net35));
 sg13g2_mux2_1 _20187_ (.A0(\cpu.dcache.r_data[7][9] ),
    .A1(net1094),
    .S(_02845_),
    .X(_02923_));
 sg13g2_nand2_1 _20188_ (.Y(_02924_),
    .A(_02843_),
    .B(_02923_));
 sg13g2_o21ai_1 _20189_ (.B1(_02924_),
    .Y(_00577_),
    .A1(_12274_),
    .A2(_02844_));
 sg13g2_buf_1 _20190_ (.A(net1011),
    .X(_02925_));
 sg13g2_buf_1 _20191_ (.A(\cpu.d_rstrobe_d ),
    .X(_02926_));
 sg13g2_nand2b_1 _20192_ (.Y(_02927_),
    .B(net1100),
    .A_N(_02926_));
 sg13g2_or4_1 _20193_ (.A(_02925_),
    .B(_09486_),
    .C(net957),
    .D(_02927_),
    .X(_02928_));
 sg13g2_o21ai_1 _20194_ (.B1(_02928_),
    .Y(_02929_),
    .A1(_09924_),
    .A2(_12112_));
 sg13g2_buf_2 _20195_ (.A(_02929_),
    .X(_02930_));
 sg13g2_xor2_1 _20196_ (.B(_12129_),
    .A(_02926_),
    .X(_02931_));
 sg13g2_nand3_1 _20197_ (.B(_12108_),
    .C(_02931_),
    .A(_12208_),
    .Y(_02932_));
 sg13g2_o21ai_1 _20198_ (.B1(_02932_),
    .Y(_02933_),
    .A1(_09924_),
    .A2(_12112_));
 sg13g2_buf_2 _20199_ (.A(_02933_),
    .X(_02934_));
 sg13g2_nor2b_1 _20200_ (.A(net607),
    .B_N(_02934_),
    .Y(_02935_));
 sg13g2_mux2_1 _20201_ (.A0(\cpu.dcache.r_dirty[0] ),
    .A1(_02930_),
    .S(_02935_),
    .X(_00578_));
 sg13g2_nand2_1 _20202_ (.Y(_02936_),
    .A(net389),
    .B(_02934_));
 sg13g2_mux2_1 _20203_ (.A0(_02930_),
    .A1(\cpu.dcache.r_dirty[1] ),
    .S(_02936_),
    .X(_00579_));
 sg13g2_nand2_1 _20204_ (.Y(_02937_),
    .A(_12459_),
    .B(_02934_));
 sg13g2_mux2_1 _20205_ (.A0(_02930_),
    .A1(\cpu.dcache.r_dirty[2] ),
    .S(_02937_),
    .X(_00580_));
 sg13g2_nand2_1 _20206_ (.Y(_02938_),
    .A(_12570_),
    .B(_02934_));
 sg13g2_mux2_1 _20207_ (.A0(_02930_),
    .A1(\cpu.dcache.r_dirty[3] ),
    .S(_02938_),
    .X(_00581_));
 sg13g2_nand2_1 _20208_ (.Y(_02939_),
    .A(net444),
    .B(_02934_));
 sg13g2_mux2_1 _20209_ (.A0(_02930_),
    .A1(\cpu.dcache.r_dirty[4] ),
    .S(_02939_),
    .X(_00582_));
 sg13g2_nand2_1 _20210_ (.Y(_02940_),
    .A(net486),
    .B(_02934_));
 sg13g2_mux2_1 _20211_ (.A0(_02930_),
    .A1(\cpu.dcache.r_dirty[5] ),
    .S(_02940_),
    .X(_00583_));
 sg13g2_nand2_1 _20212_ (.Y(_02941_),
    .A(_02734_),
    .B(_02934_));
 sg13g2_mux2_1 _20213_ (.A0(_02930_),
    .A1(\cpu.dcache.r_dirty[6] ),
    .S(_02941_),
    .X(_00584_));
 sg13g2_nand2_1 _20214_ (.Y(_02942_),
    .A(_10121_),
    .B(_02934_));
 sg13g2_mux2_1 _20215_ (.A0(_02930_),
    .A1(\cpu.dcache.r_dirty[7] ),
    .S(_02942_),
    .X(_00585_));
 sg13g2_buf_1 _20216_ (.A(_11383_),
    .X(_02943_));
 sg13g2_buf_1 _20217_ (.A(net890),
    .X(_02944_));
 sg13g2_buf_1 _20218_ (.A(net440),
    .X(_02945_));
 sg13g2_buf_1 _20219_ (.A(net440),
    .X(_02946_));
 sg13g2_nand2_1 _20220_ (.Y(_02947_),
    .A(\cpu.dcache.r_tag[0][5] ),
    .B(net387));
 sg13g2_o21ai_1 _20221_ (.B1(_02947_),
    .Y(_00589_),
    .A1(net756),
    .A2(_02945_));
 sg13g2_mux2_1 _20222_ (.A0(net407),
    .A1(\cpu.dcache.r_tag[0][15] ),
    .S(net388),
    .X(_00590_));
 sg13g2_mux2_1 _20223_ (.A0(net406),
    .A1(\cpu.dcache.r_tag[0][16] ),
    .S(net388),
    .X(_00591_));
 sg13g2_mux2_1 _20224_ (.A0(net408),
    .A1(\cpu.dcache.r_tag[0][17] ),
    .S(net388),
    .X(_00592_));
 sg13g2_mux2_1 _20225_ (.A0(_09722_),
    .A1(\cpu.dcache.r_tag[0][18] ),
    .S(net388),
    .X(_00593_));
 sg13g2_nand2_1 _20226_ (.Y(_02948_),
    .A(\cpu.dcache.r_tag[0][19] ),
    .B(net440));
 sg13g2_o21ai_1 _20227_ (.B1(_02948_),
    .Y(_00594_),
    .A1(_09667_),
    .A2(net388));
 sg13g2_mux2_1 _20228_ (.A0(net404),
    .A1(\cpu.dcache.r_tag[0][20] ),
    .S(net388),
    .X(_00595_));
 sg13g2_mux2_1 _20229_ (.A0(net401),
    .A1(\cpu.dcache.r_tag[0][21] ),
    .S(net387),
    .X(_00596_));
 sg13g2_mux2_1 _20230_ (.A0(net400),
    .A1(\cpu.dcache.r_tag[0][22] ),
    .S(net387),
    .X(_00597_));
 sg13g2_nand2_1 _20231_ (.Y(_02949_),
    .A(\cpu.dcache.r_tag[0][23] ),
    .B(net440));
 sg13g2_o21ai_1 _20232_ (.B1(_02949_),
    .Y(_00598_),
    .A1(_09968_),
    .A2(net388));
 sg13g2_buf_2 _20233_ (.A(_09277_),
    .X(_02950_));
 sg13g2_buf_1 _20234_ (.A(net984),
    .X(_02951_));
 sg13g2_buf_1 _20235_ (.A(net889),
    .X(_02952_));
 sg13g2_mux2_1 _20236_ (.A0(net755),
    .A1(\cpu.dcache.r_tag[0][6] ),
    .S(net387),
    .X(_00599_));
 sg13g2_buf_1 _20237_ (.A(_09280_),
    .X(_02953_));
 sg13g2_buf_1 _20238_ (.A(net983),
    .X(_02954_));
 sg13g2_buf_1 _20239_ (.A(net888),
    .X(_02955_));
 sg13g2_mux2_1 _20240_ (.A0(_02955_),
    .A1(\cpu.dcache.r_tag[0][7] ),
    .S(_02946_),
    .X(_00600_));
 sg13g2_buf_1 _20241_ (.A(net1056),
    .X(_02956_));
 sg13g2_buf_1 _20242_ (.A(net887),
    .X(_02957_));
 sg13g2_mux2_1 _20243_ (.A0(_02957_),
    .A1(\cpu.dcache.r_tag[0][8] ),
    .S(_02946_),
    .X(_00601_));
 sg13g2_inv_2 _20244_ (.Y(_02958_),
    .A(_10716_));
 sg13g2_nand2_1 _20245_ (.Y(_02959_),
    .A(\cpu.dcache.r_tag[0][9] ),
    .B(_12269_));
 sg13g2_o21ai_1 _20246_ (.B1(_02959_),
    .Y(_00602_),
    .A1(_02958_),
    .A2(_02945_));
 sg13g2_buf_1 _20247_ (.A(net1107),
    .X(_02960_));
 sg13g2_buf_1 _20248_ (.A(net982),
    .X(_02961_));
 sg13g2_mux2_1 _20249_ (.A0(net886),
    .A1(\cpu.dcache.r_tag[0][10] ),
    .S(net387),
    .X(_00603_));
 sg13g2_buf_1 _20250_ (.A(_11274_),
    .X(_02962_));
 sg13g2_buf_1 _20251_ (.A(net885),
    .X(_02963_));
 sg13g2_nand2_1 _20252_ (.Y(_02964_),
    .A(\cpu.dcache.r_tag[0][11] ),
    .B(_12269_));
 sg13g2_o21ai_1 _20253_ (.B1(_02964_),
    .Y(_00604_),
    .A1(net752),
    .A2(net388));
 sg13g2_mux2_1 _20254_ (.A0(net403),
    .A1(\cpu.dcache.r_tag[0][12] ),
    .S(net387),
    .X(_00605_));
 sg13g2_mux2_1 _20255_ (.A0(net402),
    .A1(\cpu.dcache.r_tag[0][13] ),
    .S(net387),
    .X(_00606_));
 sg13g2_mux2_1 _20256_ (.A0(_09565_),
    .A1(\cpu.dcache.r_tag[0][14] ),
    .S(net387),
    .X(_00607_));
 sg13g2_buf_2 _20257_ (.A(net761),
    .X(_02965_));
 sg13g2_buf_1 _20258_ (.A(net659),
    .X(_02966_));
 sg13g2_buf_1 _20259_ (.A(net602),
    .X(_02967_));
 sg13g2_buf_1 _20260_ (.A(_12402_),
    .X(_02968_));
 sg13g2_mux2_1 _20261_ (.A0(\cpu.dcache.r_tag[1][5] ),
    .A1(net527),
    .S(_02968_),
    .X(_00608_));
 sg13g2_mux2_1 _20262_ (.A0(\cpu.dcache.r_tag[1][15] ),
    .A1(net407),
    .S(net484),
    .X(_00609_));
 sg13g2_mux2_1 _20263_ (.A0(\cpu.dcache.r_tag[1][16] ),
    .A1(net406),
    .S(net484),
    .X(_00610_));
 sg13g2_mux2_1 _20264_ (.A0(\cpu.dcache.r_tag[1][17] ),
    .A1(net408),
    .S(_02968_),
    .X(_00611_));
 sg13g2_mux2_1 _20265_ (.A0(\cpu.dcache.r_tag[1][18] ),
    .A1(net405),
    .S(net484),
    .X(_00612_));
 sg13g2_mux2_1 _20266_ (.A0(\cpu.dcache.r_tag[1][19] ),
    .A1(_09666_),
    .S(net484),
    .X(_00613_));
 sg13g2_mux2_1 _20267_ (.A0(\cpu.dcache.r_tag[1][20] ),
    .A1(_09743_),
    .S(net484),
    .X(_00614_));
 sg13g2_mux2_1 _20268_ (.A0(\cpu.dcache.r_tag[1][21] ),
    .A1(net401),
    .S(net484),
    .X(_00615_));
 sg13g2_mux2_1 _20269_ (.A0(\cpu.dcache.r_tag[1][22] ),
    .A1(net400),
    .S(net484),
    .X(_00616_));
 sg13g2_mux2_1 _20270_ (.A0(\cpu.dcache.r_tag[1][23] ),
    .A1(_09609_),
    .S(net484),
    .X(_00617_));
 sg13g2_buf_1 _20271_ (.A(net889),
    .X(_02969_));
 sg13g2_buf_1 _20272_ (.A(_12402_),
    .X(_02970_));
 sg13g2_mux2_1 _20273_ (.A0(\cpu.dcache.r_tag[1][6] ),
    .A1(net751),
    .S(net483),
    .X(_00618_));
 sg13g2_buf_1 _20274_ (.A(net888),
    .X(_02971_));
 sg13g2_mux2_1 _20275_ (.A0(\cpu.dcache.r_tag[1][7] ),
    .A1(net750),
    .S(net483),
    .X(_00619_));
 sg13g2_buf_1 _20276_ (.A(net887),
    .X(_02972_));
 sg13g2_mux2_1 _20277_ (.A0(\cpu.dcache.r_tag[1][8] ),
    .A1(_02972_),
    .S(net483),
    .X(_00620_));
 sg13g2_buf_2 _20278_ (.A(_10716_),
    .X(_02973_));
 sg13g2_buf_1 _20279_ (.A(_02973_),
    .X(_02974_));
 sg13g2_mux2_1 _20280_ (.A0(\cpu.dcache.r_tag[1][9] ),
    .A1(net884),
    .S(net483),
    .X(_00621_));
 sg13g2_buf_1 _20281_ (.A(net982),
    .X(_02975_));
 sg13g2_mux2_1 _20282_ (.A0(\cpu.dcache.r_tag[1][10] ),
    .A1(net883),
    .S(net483),
    .X(_00622_));
 sg13g2_buf_1 _20283_ (.A(_10680_),
    .X(_02976_));
 sg13g2_buf_1 _20284_ (.A(net981),
    .X(_02977_));
 sg13g2_mux2_1 _20285_ (.A0(\cpu.dcache.r_tag[1][11] ),
    .A1(net882),
    .S(_02970_),
    .X(_00623_));
 sg13g2_mux2_1 _20286_ (.A0(\cpu.dcache.r_tag[1][12] ),
    .A1(net403),
    .S(_02970_),
    .X(_00624_));
 sg13g2_mux2_1 _20287_ (.A0(\cpu.dcache.r_tag[1][13] ),
    .A1(net402),
    .S(net483),
    .X(_00625_));
 sg13g2_mux2_1 _20288_ (.A0(\cpu.dcache.r_tag[1][14] ),
    .A1(net409),
    .S(net483),
    .X(_00626_));
 sg13g2_buf_1 _20289_ (.A(_12515_),
    .X(_02978_));
 sg13g2_mux2_1 _20290_ (.A0(\cpu.dcache.r_tag[2][5] ),
    .A1(net527),
    .S(net482),
    .X(_00627_));
 sg13g2_mux2_1 _20291_ (.A0(\cpu.dcache.r_tag[2][15] ),
    .A1(net407),
    .S(net482),
    .X(_00628_));
 sg13g2_mux2_1 _20292_ (.A0(\cpu.dcache.r_tag[2][16] ),
    .A1(net406),
    .S(net482),
    .X(_00629_));
 sg13g2_mux2_1 _20293_ (.A0(\cpu.dcache.r_tag[2][17] ),
    .A1(net408),
    .S(net482),
    .X(_00630_));
 sg13g2_mux2_1 _20294_ (.A0(\cpu.dcache.r_tag[2][18] ),
    .A1(net405),
    .S(net482),
    .X(_00631_));
 sg13g2_mux2_1 _20295_ (.A0(\cpu.dcache.r_tag[2][19] ),
    .A1(_09666_),
    .S(net482),
    .X(_00632_));
 sg13g2_mux2_1 _20296_ (.A0(\cpu.dcache.r_tag[2][20] ),
    .A1(net404),
    .S(net482),
    .X(_00633_));
 sg13g2_mux2_1 _20297_ (.A0(\cpu.dcache.r_tag[2][21] ),
    .A1(net401),
    .S(_02978_),
    .X(_00634_));
 sg13g2_mux2_1 _20298_ (.A0(\cpu.dcache.r_tag[2][22] ),
    .A1(net400),
    .S(net482),
    .X(_00635_));
 sg13g2_mux2_1 _20299_ (.A0(\cpu.dcache.r_tag[2][23] ),
    .A1(_09609_),
    .S(_02978_),
    .X(_00636_));
 sg13g2_buf_1 _20300_ (.A(_12515_),
    .X(_02979_));
 sg13g2_mux2_1 _20301_ (.A0(\cpu.dcache.r_tag[2][6] ),
    .A1(net751),
    .S(net481),
    .X(_00637_));
 sg13g2_mux2_1 _20302_ (.A0(\cpu.dcache.r_tag[2][7] ),
    .A1(net750),
    .S(net481),
    .X(_00638_));
 sg13g2_mux2_1 _20303_ (.A0(\cpu.dcache.r_tag[2][8] ),
    .A1(net749),
    .S(net481),
    .X(_00639_));
 sg13g2_mux2_1 _20304_ (.A0(\cpu.dcache.r_tag[2][9] ),
    .A1(net884),
    .S(net481),
    .X(_00640_));
 sg13g2_mux2_1 _20305_ (.A0(\cpu.dcache.r_tag[2][10] ),
    .A1(net883),
    .S(net481),
    .X(_00641_));
 sg13g2_mux2_1 _20306_ (.A0(\cpu.dcache.r_tag[2][11] ),
    .A1(net882),
    .S(_02979_),
    .X(_00642_));
 sg13g2_mux2_1 _20307_ (.A0(\cpu.dcache.r_tag[2][12] ),
    .A1(net403),
    .S(_02979_),
    .X(_00643_));
 sg13g2_mux2_1 _20308_ (.A0(\cpu.dcache.r_tag[2][13] ),
    .A1(net402),
    .S(net481),
    .X(_00644_));
 sg13g2_mux2_1 _20309_ (.A0(\cpu.dcache.r_tag[2][14] ),
    .A1(net409),
    .S(net481),
    .X(_00645_));
 sg13g2_buf_1 _20310_ (.A(_12618_),
    .X(_02980_));
 sg13g2_mux2_1 _20311_ (.A0(\cpu.dcache.r_tag[3][5] ),
    .A1(net527),
    .S(net198),
    .X(_00646_));
 sg13g2_mux2_1 _20312_ (.A0(\cpu.dcache.r_tag[3][15] ),
    .A1(net407),
    .S(net198),
    .X(_00647_));
 sg13g2_mux2_1 _20313_ (.A0(\cpu.dcache.r_tag[3][16] ),
    .A1(net406),
    .S(_02980_),
    .X(_00648_));
 sg13g2_mux2_1 _20314_ (.A0(\cpu.dcache.r_tag[3][17] ),
    .A1(net408),
    .S(_02980_),
    .X(_00649_));
 sg13g2_mux2_1 _20315_ (.A0(\cpu.dcache.r_tag[3][18] ),
    .A1(net405),
    .S(net198),
    .X(_00650_));
 sg13g2_mux2_1 _20316_ (.A0(\cpu.dcache.r_tag[3][19] ),
    .A1(_09666_),
    .S(net198),
    .X(_00651_));
 sg13g2_mux2_1 _20317_ (.A0(\cpu.dcache.r_tag[3][20] ),
    .A1(net404),
    .S(net198),
    .X(_00652_));
 sg13g2_mux2_1 _20318_ (.A0(\cpu.dcache.r_tag[3][21] ),
    .A1(net401),
    .S(net198),
    .X(_00653_));
 sg13g2_mux2_1 _20319_ (.A0(\cpu.dcache.r_tag[3][22] ),
    .A1(net400),
    .S(net198),
    .X(_00654_));
 sg13g2_mux2_1 _20320_ (.A0(\cpu.dcache.r_tag[3][23] ),
    .A1(_09609_),
    .S(net198),
    .X(_00655_));
 sg13g2_buf_1 _20321_ (.A(_12618_),
    .X(_02981_));
 sg13g2_mux2_1 _20322_ (.A0(\cpu.dcache.r_tag[3][6] ),
    .A1(_02969_),
    .S(net197),
    .X(_00656_));
 sg13g2_mux2_1 _20323_ (.A0(\cpu.dcache.r_tag[3][7] ),
    .A1(_02971_),
    .S(net197),
    .X(_00657_));
 sg13g2_mux2_1 _20324_ (.A0(\cpu.dcache.r_tag[3][8] ),
    .A1(net749),
    .S(net197),
    .X(_00658_));
 sg13g2_mux2_1 _20325_ (.A0(\cpu.dcache.r_tag[3][9] ),
    .A1(net884),
    .S(net197),
    .X(_00659_));
 sg13g2_mux2_1 _20326_ (.A0(\cpu.dcache.r_tag[3][10] ),
    .A1(_02975_),
    .S(net197),
    .X(_00660_));
 sg13g2_mux2_1 _20327_ (.A0(\cpu.dcache.r_tag[3][11] ),
    .A1(net882),
    .S(_02981_),
    .X(_00661_));
 sg13g2_mux2_1 _20328_ (.A0(\cpu.dcache.r_tag[3][12] ),
    .A1(_09768_),
    .S(_02981_),
    .X(_00662_));
 sg13g2_mux2_1 _20329_ (.A0(\cpu.dcache.r_tag[3][13] ),
    .A1(net402),
    .S(net197),
    .X(_00663_));
 sg13g2_mux2_1 _20330_ (.A0(\cpu.dcache.r_tag[3][14] ),
    .A1(net409),
    .S(net197),
    .X(_00664_));
 sg13g2_buf_1 _20331_ (.A(net436),
    .X(_02982_));
 sg13g2_nand2_1 _20332_ (.Y(_02983_),
    .A(\cpu.dcache.r_tag[4][5] ),
    .B(net436));
 sg13g2_o21ai_1 _20333_ (.B1(_02983_),
    .Y(_00665_),
    .A1(net756),
    .A2(net386));
 sg13g2_mux2_1 _20334_ (.A0(net407),
    .A1(\cpu.dcache.r_tag[4][15] ),
    .S(net386),
    .X(_00666_));
 sg13g2_mux2_1 _20335_ (.A0(net406),
    .A1(\cpu.dcache.r_tag[4][16] ),
    .S(net386),
    .X(_00667_));
 sg13g2_mux2_1 _20336_ (.A0(net408),
    .A1(\cpu.dcache.r_tag[4][17] ),
    .S(net386),
    .X(_00668_));
 sg13g2_mux2_1 _20337_ (.A0(net405),
    .A1(\cpu.dcache.r_tag[4][18] ),
    .S(net386),
    .X(_00669_));
 sg13g2_nand2_1 _20338_ (.Y(_02984_),
    .A(\cpu.dcache.r_tag[4][19] ),
    .B(net436));
 sg13g2_o21ai_1 _20339_ (.B1(_02984_),
    .Y(_00670_),
    .A1(_09667_),
    .A2(net386));
 sg13g2_buf_1 _20340_ (.A(net436),
    .X(_02985_));
 sg13g2_mux2_1 _20341_ (.A0(net404),
    .A1(\cpu.dcache.r_tag[4][20] ),
    .S(net385),
    .X(_00671_));
 sg13g2_mux2_1 _20342_ (.A0(net401),
    .A1(\cpu.dcache.r_tag[4][21] ),
    .S(net385),
    .X(_00672_));
 sg13g2_mux2_1 _20343_ (.A0(net400),
    .A1(\cpu.dcache.r_tag[4][22] ),
    .S(net385),
    .X(_00673_));
 sg13g2_nand2_1 _20344_ (.Y(_02986_),
    .A(\cpu.dcache.r_tag[4][23] ),
    .B(net436));
 sg13g2_o21ai_1 _20345_ (.B1(_02986_),
    .Y(_00674_),
    .A1(_09968_),
    .A2(net386));
 sg13g2_mux2_1 _20346_ (.A0(net755),
    .A1(\cpu.dcache.r_tag[4][6] ),
    .S(net385),
    .X(_00675_));
 sg13g2_mux2_1 _20347_ (.A0(_02955_),
    .A1(\cpu.dcache.r_tag[4][7] ),
    .S(_02985_),
    .X(_00676_));
 sg13g2_mux2_1 _20348_ (.A0(_02957_),
    .A1(\cpu.dcache.r_tag[4][8] ),
    .S(_02985_),
    .X(_00677_));
 sg13g2_nand2_1 _20349_ (.Y(_02987_),
    .A(\cpu.dcache.r_tag[4][9] ),
    .B(_12726_));
 sg13g2_o21ai_1 _20350_ (.B1(_02987_),
    .Y(_00678_),
    .A1(_02958_),
    .A2(_02982_));
 sg13g2_mux2_1 _20351_ (.A0(_02961_),
    .A1(\cpu.dcache.r_tag[4][10] ),
    .S(net385),
    .X(_00679_));
 sg13g2_nand2_1 _20352_ (.Y(_02988_),
    .A(\cpu.dcache.r_tag[4][11] ),
    .B(_12726_));
 sg13g2_o21ai_1 _20353_ (.B1(_02988_),
    .Y(_00680_),
    .A1(net752),
    .A2(_02982_));
 sg13g2_mux2_1 _20354_ (.A0(net403),
    .A1(\cpu.dcache.r_tag[4][12] ),
    .S(net385),
    .X(_00681_));
 sg13g2_mux2_1 _20355_ (.A0(net402),
    .A1(\cpu.dcache.r_tag[4][13] ),
    .S(net385),
    .X(_00682_));
 sg13g2_mux2_1 _20356_ (.A0(net409),
    .A1(\cpu.dcache.r_tag[4][14] ),
    .S(net385),
    .X(_00683_));
 sg13g2_buf_1 _20357_ (.A(_12840_),
    .X(_02989_));
 sg13g2_buf_1 _20358_ (.A(_12840_),
    .X(_02990_));
 sg13g2_nand2_1 _20359_ (.Y(_02991_),
    .A(net602),
    .B(_02990_));
 sg13g2_o21ai_1 _20360_ (.B1(_02991_),
    .Y(_00684_),
    .A1(_09834_),
    .A2(_02989_));
 sg13g2_mux2_1 _20361_ (.A0(\cpu.dcache.r_tag[5][15] ),
    .A1(net407),
    .S(net480),
    .X(_00685_));
 sg13g2_mux2_1 _20362_ (.A0(\cpu.dcache.r_tag[5][16] ),
    .A1(net406),
    .S(_02989_),
    .X(_00686_));
 sg13g2_mux2_1 _20363_ (.A0(\cpu.dcache.r_tag[5][17] ),
    .A1(net408),
    .S(net480),
    .X(_00687_));
 sg13g2_mux2_1 _20364_ (.A0(\cpu.dcache.r_tag[5][18] ),
    .A1(net405),
    .S(net480),
    .X(_00688_));
 sg13g2_mux2_1 _20365_ (.A0(\cpu.dcache.r_tag[5][19] ),
    .A1(_09666_),
    .S(net480),
    .X(_00689_));
 sg13g2_mux2_1 _20366_ (.A0(\cpu.dcache.r_tag[5][20] ),
    .A1(net404),
    .S(net480),
    .X(_00690_));
 sg13g2_mux2_1 _20367_ (.A0(\cpu.dcache.r_tag[5][21] ),
    .A1(net401),
    .S(net480),
    .X(_00691_));
 sg13g2_mux2_1 _20368_ (.A0(\cpu.dcache.r_tag[5][22] ),
    .A1(net400),
    .S(net480),
    .X(_00692_));
 sg13g2_mux2_1 _20369_ (.A0(\cpu.dcache.r_tag[5][23] ),
    .A1(_09609_),
    .S(net480),
    .X(_00693_));
 sg13g2_mux2_1 _20370_ (.A0(\cpu.dcache.r_tag[5][6] ),
    .A1(_02969_),
    .S(_02990_),
    .X(_00694_));
 sg13g2_mux2_1 _20371_ (.A0(\cpu.dcache.r_tag[5][7] ),
    .A1(_02971_),
    .S(net479),
    .X(_00695_));
 sg13g2_mux2_1 _20372_ (.A0(\cpu.dcache.r_tag[5][8] ),
    .A1(_02972_),
    .S(net479),
    .X(_00696_));
 sg13g2_mux2_1 _20373_ (.A0(\cpu.dcache.r_tag[5][9] ),
    .A1(net884),
    .S(net479),
    .X(_00697_));
 sg13g2_mux2_1 _20374_ (.A0(\cpu.dcache.r_tag[5][10] ),
    .A1(_02975_),
    .S(net479),
    .X(_00698_));
 sg13g2_mux2_1 _20375_ (.A0(\cpu.dcache.r_tag[5][11] ),
    .A1(net882),
    .S(net479),
    .X(_00699_));
 sg13g2_mux2_1 _20376_ (.A0(\cpu.dcache.r_tag[5][12] ),
    .A1(_09768_),
    .S(net479),
    .X(_00700_));
 sg13g2_mux2_1 _20377_ (.A0(\cpu.dcache.r_tag[5][13] ),
    .A1(net402),
    .S(net479),
    .X(_00701_));
 sg13g2_mux2_1 _20378_ (.A0(\cpu.dcache.r_tag[5][14] ),
    .A1(net409),
    .S(net479),
    .X(_00702_));
 sg13g2_buf_1 _20379_ (.A(_02791_),
    .X(_02992_));
 sg13g2_buf_1 _20380_ (.A(_02791_),
    .X(_02993_));
 sg13g2_nand2_1 _20381_ (.Y(_02994_),
    .A(net602),
    .B(net477));
 sg13g2_o21ai_1 _20382_ (.B1(_02994_),
    .Y(_00703_),
    .A1(_09829_),
    .A2(_02992_));
 sg13g2_mux2_1 _20383_ (.A0(\cpu.dcache.r_tag[6][15] ),
    .A1(net407),
    .S(net478),
    .X(_00704_));
 sg13g2_mux2_1 _20384_ (.A0(\cpu.dcache.r_tag[6][16] ),
    .A1(_09696_),
    .S(_02992_),
    .X(_00705_));
 sg13g2_mux2_1 _20385_ (.A0(\cpu.dcache.r_tag[6][17] ),
    .A1(_09588_),
    .S(net478),
    .X(_00706_));
 sg13g2_mux2_1 _20386_ (.A0(\cpu.dcache.r_tag[6][18] ),
    .A1(net405),
    .S(net478),
    .X(_00707_));
 sg13g2_mux2_1 _20387_ (.A0(\cpu.dcache.r_tag[6][19] ),
    .A1(_09666_),
    .S(net478),
    .X(_00708_));
 sg13g2_mux2_1 _20388_ (.A0(\cpu.dcache.r_tag[6][20] ),
    .A1(net404),
    .S(net478),
    .X(_00709_));
 sg13g2_mux2_1 _20389_ (.A0(\cpu.dcache.r_tag[6][21] ),
    .A1(net401),
    .S(net478),
    .X(_00710_));
 sg13g2_mux2_1 _20390_ (.A0(\cpu.dcache.r_tag[6][22] ),
    .A1(_09913_),
    .S(net478),
    .X(_00711_));
 sg13g2_mux2_1 _20391_ (.A0(\cpu.dcache.r_tag[6][23] ),
    .A1(_09609_),
    .S(net478),
    .X(_00712_));
 sg13g2_buf_1 _20392_ (.A(net889),
    .X(_02995_));
 sg13g2_mux2_1 _20393_ (.A0(\cpu.dcache.r_tag[6][6] ),
    .A1(net748),
    .S(net477),
    .X(_00713_));
 sg13g2_buf_1 _20394_ (.A(net888),
    .X(_02996_));
 sg13g2_mux2_1 _20395_ (.A0(\cpu.dcache.r_tag[6][7] ),
    .A1(net747),
    .S(net477),
    .X(_00714_));
 sg13g2_buf_1 _20396_ (.A(net887),
    .X(_02997_));
 sg13g2_mux2_1 _20397_ (.A0(\cpu.dcache.r_tag[6][8] ),
    .A1(net746),
    .S(net477),
    .X(_00715_));
 sg13g2_mux2_1 _20398_ (.A0(\cpu.dcache.r_tag[6][9] ),
    .A1(_02974_),
    .S(net477),
    .X(_00716_));
 sg13g2_buf_1 _20399_ (.A(net982),
    .X(_02998_));
 sg13g2_mux2_1 _20400_ (.A0(\cpu.dcache.r_tag[6][10] ),
    .A1(net881),
    .S(net477),
    .X(_00717_));
 sg13g2_mux2_1 _20401_ (.A0(\cpu.dcache.r_tag[6][11] ),
    .A1(net882),
    .S(_02993_),
    .X(_00718_));
 sg13g2_mux2_1 _20402_ (.A0(\cpu.dcache.r_tag[6][12] ),
    .A1(net403),
    .S(_02993_),
    .X(_00719_));
 sg13g2_mux2_1 _20403_ (.A0(\cpu.dcache.r_tag[6][13] ),
    .A1(_09797_),
    .S(net477),
    .X(_00720_));
 sg13g2_mux2_1 _20404_ (.A0(\cpu.dcache.r_tag[6][14] ),
    .A1(net409),
    .S(net477),
    .X(_00721_));
 sg13g2_buf_1 _20405_ (.A(_02891_),
    .X(_02999_));
 sg13g2_mux2_1 _20406_ (.A0(\cpu.dcache.r_tag[7][5] ),
    .A1(net527),
    .S(net228),
    .X(_00722_));
 sg13g2_mux2_1 _20407_ (.A0(\cpu.dcache.r_tag[7][15] ),
    .A1(net407),
    .S(net228),
    .X(_00723_));
 sg13g2_mux2_1 _20408_ (.A0(\cpu.dcache.r_tag[7][16] ),
    .A1(_09696_),
    .S(_02999_),
    .X(_00724_));
 sg13g2_mux2_1 _20409_ (.A0(\cpu.dcache.r_tag[7][17] ),
    .A1(_09588_),
    .S(_02999_),
    .X(_00725_));
 sg13g2_mux2_1 _20410_ (.A0(\cpu.dcache.r_tag[7][18] ),
    .A1(_09722_),
    .S(net228),
    .X(_00726_));
 sg13g2_mux2_1 _20411_ (.A0(\cpu.dcache.r_tag[7][19] ),
    .A1(_09666_),
    .S(net228),
    .X(_00727_));
 sg13g2_mux2_1 _20412_ (.A0(\cpu.dcache.r_tag[7][20] ),
    .A1(net404),
    .S(net228),
    .X(_00728_));
 sg13g2_mux2_1 _20413_ (.A0(\cpu.dcache.r_tag[7][21] ),
    .A1(_09890_),
    .S(net228),
    .X(_00729_));
 sg13g2_mux2_1 _20414_ (.A0(\cpu.dcache.r_tag[7][22] ),
    .A1(net400),
    .S(net228),
    .X(_00730_));
 sg13g2_mux2_1 _20415_ (.A0(\cpu.dcache.r_tag[7][23] ),
    .A1(_09609_),
    .S(net228),
    .X(_00731_));
 sg13g2_buf_1 _20416_ (.A(_02891_),
    .X(_03000_));
 sg13g2_mux2_1 _20417_ (.A0(\cpu.dcache.r_tag[7][6] ),
    .A1(net748),
    .S(net227),
    .X(_00732_));
 sg13g2_mux2_1 _20418_ (.A0(\cpu.dcache.r_tag[7][7] ),
    .A1(net747),
    .S(net227),
    .X(_00733_));
 sg13g2_mux2_1 _20419_ (.A0(\cpu.dcache.r_tag[7][8] ),
    .A1(net746),
    .S(net227),
    .X(_00734_));
 sg13g2_mux2_1 _20420_ (.A0(\cpu.dcache.r_tag[7][9] ),
    .A1(_02974_),
    .S(_03000_),
    .X(_00735_));
 sg13g2_mux2_1 _20421_ (.A0(\cpu.dcache.r_tag[7][10] ),
    .A1(net881),
    .S(_03000_),
    .X(_00736_));
 sg13g2_mux2_1 _20422_ (.A0(\cpu.dcache.r_tag[7][11] ),
    .A1(net882),
    .S(net227),
    .X(_00737_));
 sg13g2_mux2_1 _20423_ (.A0(\cpu.dcache.r_tag[7][12] ),
    .A1(net403),
    .S(net227),
    .X(_00738_));
 sg13g2_mux2_1 _20424_ (.A0(\cpu.dcache.r_tag[7][13] ),
    .A1(_09797_),
    .S(net227),
    .X(_00739_));
 sg13g2_mux2_1 _20425_ (.A0(\cpu.dcache.r_tag[7][14] ),
    .A1(_09565_),
    .S(net227),
    .X(_00740_));
 sg13g2_nor2_1 _20426_ (.A(_09058_),
    .B(_10026_),
    .Y(_03001_));
 sg13g2_buf_1 _20427_ (.A(_03001_),
    .X(_03002_));
 sg13g2_a21o_1 _20428_ (.A2(_09048_),
    .A1(_08976_),
    .B1(_09056_),
    .X(_03003_));
 sg13g2_buf_1 _20429_ (.A(_03003_),
    .X(_03004_));
 sg13g2_nor2_1 _20430_ (.A(net280),
    .B(_03004_),
    .Y(_03005_));
 sg13g2_buf_2 _20431_ (.A(_03005_),
    .X(_03006_));
 sg13g2_a21oi_1 _20432_ (.A1(net240),
    .A2(net226),
    .Y(_03007_),
    .B1(_03006_));
 sg13g2_nor2_1 _20433_ (.A(_10003_),
    .B(_03007_),
    .Y(_03008_));
 sg13g2_nand2_1 _20434_ (.Y(_03009_),
    .A(_10003_),
    .B(net240));
 sg13g2_buf_2 _20435_ (.A(_03009_),
    .X(_03010_));
 sg13g2_nor2_1 _20436_ (.A(net152),
    .B(_03010_),
    .Y(_03011_));
 sg13g2_buf_1 _20437_ (.A(_08972_),
    .X(_03012_));
 sg13g2_o21ai_1 _20438_ (.B1(_03012_),
    .Y(_03013_),
    .A1(_03008_),
    .A2(_03011_));
 sg13g2_o21ai_1 _20439_ (.B1(_03013_),
    .Y(_00749_),
    .A1(_11137_),
    .A2(net118));
 sg13g2_buf_1 _20440_ (.A(net279),
    .X(_03014_));
 sg13g2_buf_1 _20441_ (.A(_10026_),
    .X(_03015_));
 sg13g2_buf_1 _20442_ (.A(_09199_),
    .X(_03016_));
 sg13g2_nand2_1 _20443_ (.Y(_03017_),
    .A(net168),
    .B(net180));
 sg13g2_buf_1 _20444_ (.A(_10003_),
    .X(_03018_));
 sg13g2_a22oi_1 _20445_ (.Y(_03019_),
    .B1(_03017_),
    .B2(net167),
    .A2(net270),
    .A1(net177));
 sg13g2_nor2_1 _20446_ (.A(net225),
    .B(_03019_),
    .Y(_03020_));
 sg13g2_buf_1 _20447_ (.A(net280),
    .X(_03021_));
 sg13g2_nand2_1 _20448_ (.Y(_03022_),
    .A(net207),
    .B(net224));
 sg13g2_buf_1 _20449_ (.A(_09079_),
    .X(_03023_));
 sg13g2_nand2_1 _20450_ (.Y(_03024_),
    .A(net212),
    .B(net280));
 sg13g2_nand3_1 _20451_ (.B(net223),
    .C(_03024_),
    .A(net225),
    .Y(_03025_));
 sg13g2_o21ai_1 _20452_ (.B1(_03025_),
    .Y(_03026_),
    .A1(net167),
    .A2(_03022_));
 sg13g2_o21ai_1 _20453_ (.B1(net115),
    .Y(_03027_),
    .A1(_03020_),
    .A2(_03026_));
 sg13g2_o21ai_1 _20454_ (.B1(_03027_),
    .Y(_00750_),
    .A1(_11680_),
    .A2(net118));
 sg13g2_buf_1 _20455_ (.A(net108),
    .X(_03028_));
 sg13g2_nand2_1 _20456_ (.Y(_03029_),
    .A(net239),
    .B(net225));
 sg13g2_nor3_1 _20457_ (.A(_09998_),
    .B(net151),
    .C(_03029_),
    .Y(_03030_));
 sg13g2_a21o_1 _20458_ (.A2(net87),
    .A1(\cpu.cond[1] ),
    .B1(_03030_),
    .X(_00751_));
 sg13g2_a21oi_1 _20459_ (.A1(net225),
    .A2(_03024_),
    .Y(_03031_),
    .B1(net168));
 sg13g2_buf_1 _20460_ (.A(_08972_),
    .X(_03032_));
 sg13g2_mux2_1 _20461_ (.A0(\cpu.cond[2] ),
    .A1(_03031_),
    .S(net114),
    .X(_00752_));
 sg13g2_nor4_1 _20462_ (.A(net108),
    .B(_09136_),
    .C(_09203_),
    .D(_09205_),
    .Y(_03033_));
 sg13g2_a21o_1 _20463_ (.A2(net87),
    .A1(\cpu.dec.div ),
    .B1(_03033_),
    .X(_00753_));
 sg13g2_nand2_1 _20464_ (.Y(_03034_),
    .A(net150),
    .B(net149));
 sg13g2_mux4_1 _20465_ (.S0(net1061),
    .A0(\cpu.icache.r_data[4][8] ),
    .A1(\cpu.icache.r_data[5][8] ),
    .A2(\cpu.icache.r_data[6][8] ),
    .A3(\cpu.icache.r_data[7][8] ),
    .S1(net942),
    .X(_03035_));
 sg13g2_nand2_1 _20466_ (.Y(_03036_),
    .A(net935),
    .B(_03035_));
 sg13g2_a22oi_1 _20467_ (.Y(_03037_),
    .B1(net638),
    .B2(\cpu.icache.r_data[3][8] ),
    .A2(net717),
    .A1(\cpu.icache.r_data[2][8] ));
 sg13g2_nand2_1 _20468_ (.Y(_03038_),
    .A(\cpu.icache.r_data[1][8] ),
    .B(_08589_));
 sg13g2_and4_1 _20469_ (.A(net560),
    .B(_03036_),
    .C(_03037_),
    .D(_03038_),
    .X(_03039_));
 sg13g2_a21oi_1 _20470_ (.A1(_00174_),
    .A2(_08981_),
    .Y(_03040_),
    .B1(_03039_));
 sg13g2_nor2_1 _20471_ (.A(_00175_),
    .B(_08570_),
    .Y(_03041_));
 sg13g2_mux2_1 _20472_ (.A0(\cpu.icache.r_data[7][24] ),
    .A1(\cpu.icache.r_data[3][24] ),
    .S(net1064),
    .X(_03042_));
 sg13g2_a22oi_1 _20473_ (.Y(_03043_),
    .B1(_03042_),
    .B2(_08801_),
    .A2(_08582_),
    .A1(\cpu.icache.r_data[5][24] ));
 sg13g2_nor2_1 _20474_ (.A(_08608_),
    .B(_03043_),
    .Y(_03044_));
 sg13g2_a22oi_1 _20475_ (.Y(_03045_),
    .B1(net811),
    .B2(\cpu.icache.r_data[4][24] ),
    .A2(net717),
    .A1(\cpu.icache.r_data[2][24] ));
 sg13g2_a22oi_1 _20476_ (.Y(_03046_),
    .B1(_08665_),
    .B2(\cpu.icache.r_data[6][24] ),
    .A2(net639),
    .A1(\cpu.icache.r_data[1][24] ));
 sg13g2_nand2_1 _20477_ (.Y(_03047_),
    .A(_03045_),
    .B(_03046_));
 sg13g2_or4_1 _20478_ (.A(net936),
    .B(_03041_),
    .C(_03044_),
    .D(_03047_),
    .X(_03048_));
 sg13g2_o21ai_1 _20479_ (.B1(_03048_),
    .Y(_03049_),
    .A1(net1060),
    .A2(_03040_));
 sg13g2_buf_1 _20480_ (.A(_03049_),
    .X(_03050_));
 sg13g2_mux4_1 _20481_ (.S0(net1061),
    .A0(\cpu.icache.r_data[4][25] ),
    .A1(\cpu.icache.r_data[5][25] ),
    .A2(\cpu.icache.r_data[6][25] ),
    .A3(\cpu.icache.r_data[7][25] ),
    .S1(net942),
    .X(_03051_));
 sg13g2_and2_1 _20482_ (.A(\cpu.icache.r_data[1][25] ),
    .B(_08588_),
    .X(_03052_));
 sg13g2_a221oi_1 _20483_ (.B2(\cpu.icache.r_data[3][25] ),
    .C1(_03052_),
    .B1(_08595_),
    .A1(\cpu.icache.r_data[2][25] ),
    .Y(_03053_),
    .A2(_08577_));
 sg13g2_o21ai_1 _20484_ (.B1(_03053_),
    .Y(_03054_),
    .A1(_00177_),
    .A2(_08569_));
 sg13g2_a21oi_1 _20485_ (.A1(net935),
    .A2(_03051_),
    .Y(_03055_),
    .B1(_03054_));
 sg13g2_nand2_1 _20486_ (.Y(_03056_),
    .A(_00176_),
    .B(_08980_));
 sg13g2_mux4_1 _20487_ (.S0(_08564_),
    .A0(\cpu.icache.r_data[4][9] ),
    .A1(\cpu.icache.r_data[5][9] ),
    .A2(\cpu.icache.r_data[6][9] ),
    .A3(\cpu.icache.r_data[7][9] ),
    .S1(net1063),
    .X(_03057_));
 sg13g2_nand2_1 _20488_ (.Y(_03058_),
    .A(net935),
    .B(_03057_));
 sg13g2_a22oi_1 _20489_ (.Y(_03059_),
    .B1(_08595_),
    .B2(\cpu.icache.r_data[3][9] ),
    .A2(_08577_),
    .A1(\cpu.icache.r_data[2][9] ));
 sg13g2_nand2_1 _20490_ (.Y(_03060_),
    .A(\cpu.icache.r_data[1][9] ),
    .B(_08588_));
 sg13g2_nand4_1 _20491_ (.B(_03058_),
    .C(_03059_),
    .A(_08570_),
    .Y(_03061_),
    .D(_03060_));
 sg13g2_nand3_1 _20492_ (.B(_03056_),
    .C(_03061_),
    .A(_09012_),
    .Y(_03062_));
 sg13g2_o21ai_1 _20493_ (.B1(_03062_),
    .Y(_03063_),
    .A1(_09012_),
    .A2(_03055_));
 sg13g2_buf_1 _20494_ (.A(_03063_),
    .X(_03064_));
 sg13g2_mux4_1 _20495_ (.S0(net1061),
    .A0(\cpu.icache.r_data[4][23] ),
    .A1(\cpu.icache.r_data[5][23] ),
    .A2(\cpu.icache.r_data[6][23] ),
    .A3(\cpu.icache.r_data[7][23] ),
    .S1(net946),
    .X(_03065_));
 sg13g2_and2_1 _20496_ (.A(\cpu.icache.r_data[1][23] ),
    .B(_08588_),
    .X(_03066_));
 sg13g2_a221oi_1 _20497_ (.B2(\cpu.icache.r_data[3][23] ),
    .C1(_03066_),
    .B1(_08595_),
    .A1(\cpu.icache.r_data[2][23] ),
    .Y(_03067_),
    .A2(_08577_));
 sg13g2_o21ai_1 _20498_ (.B1(_03067_),
    .Y(_03068_),
    .A1(_00173_),
    .A2(net560));
 sg13g2_a21oi_1 _20499_ (.A1(net935),
    .A2(_03065_),
    .Y(_03069_),
    .B1(_03068_));
 sg13g2_nand2_1 _20500_ (.Y(_03070_),
    .A(_00172_),
    .B(_08980_));
 sg13g2_mux4_1 _20501_ (.S0(net1126),
    .A0(\cpu.icache.r_data[4][7] ),
    .A1(\cpu.icache.r_data[5][7] ),
    .A2(\cpu.icache.r_data[6][7] ),
    .A3(\cpu.icache.r_data[7][7] ),
    .S1(net1063),
    .X(_03071_));
 sg13g2_nand2_1 _20502_ (.Y(_03072_),
    .A(_09064_),
    .B(_03071_));
 sg13g2_a22oi_1 _20503_ (.Y(_03073_),
    .B1(_08595_),
    .B2(\cpu.icache.r_data[3][7] ),
    .A2(_08577_),
    .A1(\cpu.icache.r_data[2][7] ));
 sg13g2_nand2_1 _20504_ (.Y(_03074_),
    .A(\cpu.icache.r_data[1][7] ),
    .B(_08588_));
 sg13g2_nand4_1 _20505_ (.B(_03072_),
    .C(_03073_),
    .A(net560),
    .Y(_03075_),
    .D(_03074_));
 sg13g2_nand3_1 _20506_ (.B(_03070_),
    .C(_03075_),
    .A(_09012_),
    .Y(_03076_));
 sg13g2_o21ai_1 _20507_ (.B1(_03076_),
    .Y(_03077_),
    .A1(_09013_),
    .A2(_03069_));
 sg13g2_buf_1 _20508_ (.A(_03077_),
    .X(_03078_));
 sg13g2_nor2_1 _20509_ (.A(_03064_),
    .B(_03078_),
    .Y(_03079_));
 sg13g2_and2_1 _20510_ (.A(_03050_),
    .B(_03079_),
    .X(_03080_));
 sg13g2_buf_1 _20511_ (.A(_03080_),
    .X(_03081_));
 sg13g2_nand3_1 _20512_ (.B(_09995_),
    .C(_03081_),
    .A(_09192_),
    .Y(_03082_));
 sg13g2_buf_1 _20513_ (.A(_03082_),
    .X(_03083_));
 sg13g2_nor4_1 _20514_ (.A(net108),
    .B(_09258_),
    .C(_03034_),
    .D(_03083_),
    .Y(_03084_));
 sg13g2_a21o_1 _20515_ (.A2(net87),
    .A1(\cpu.dec.do_flush_all ),
    .B1(_03084_),
    .X(_00754_));
 sg13g2_nand2_1 _20516_ (.Y(_03085_),
    .A(net239),
    .B(net226));
 sg13g2_nor3_1 _20517_ (.A(net106),
    .B(net151),
    .C(_03085_),
    .Y(_03086_));
 sg13g2_a21o_1 _20518_ (.A2(net87),
    .A1(\cpu.dec.do_flush_write ),
    .B1(_03086_),
    .X(_00755_));
 sg13g2_nor2_1 _20519_ (.A(net212),
    .B(_03016_),
    .Y(_03087_));
 sg13g2_buf_1 _20520_ (.A(_03087_),
    .X(_03088_));
 sg13g2_inv_1 _20521_ (.Y(_03089_),
    .A(_10006_));
 sg13g2_nor2_1 _20522_ (.A(net280),
    .B(net223),
    .Y(_03090_));
 sg13g2_buf_1 _20523_ (.A(_03004_),
    .X(_03091_));
 sg13g2_o21ai_1 _20524_ (.B1(net269),
    .Y(_03092_),
    .A1(net167),
    .A2(_03090_));
 sg13g2_o21ai_1 _20525_ (.B1(_03092_),
    .Y(_03093_),
    .A1(_09020_),
    .A2(net206));
 sg13g2_a22oi_1 _20526_ (.Y(_03094_),
    .B1(_03093_),
    .B2(net211),
    .A2(net149),
    .A1(_03089_));
 sg13g2_buf_1 _20527_ (.A(_09256_),
    .X(_03095_));
 sg13g2_nand2_1 _20528_ (.Y(_03096_),
    .A(_10003_),
    .B(_09199_));
 sg13g2_buf_2 _20529_ (.A(_03096_),
    .X(_03097_));
 sg13g2_nor2_1 _20530_ (.A(net222),
    .B(_03097_),
    .Y(_03098_));
 sg13g2_nor2_1 _20531_ (.A(_09174_),
    .B(_03010_),
    .Y(_03099_));
 sg13g2_nor2_2 _20532_ (.A(net269),
    .B(net270),
    .Y(_03100_));
 sg13g2_o21ai_1 _20533_ (.B1(_03100_),
    .Y(_03101_),
    .A1(_03098_),
    .A2(_03099_));
 sg13g2_o21ai_1 _20534_ (.B1(_03101_),
    .Y(_03102_),
    .A1(_03088_),
    .A2(_03094_));
 sg13g2_mux2_1 _20535_ (.A0(_10962_),
    .A1(_03102_),
    .S(net114),
    .X(_00756_));
 sg13g2_nand2_1 _20536_ (.Y(_03103_),
    .A(net280),
    .B(net226));
 sg13g2_buf_2 _20537_ (.A(_03103_),
    .X(_03104_));
 sg13g2_nor2_1 _20538_ (.A(net240),
    .B(_03104_),
    .Y(_03105_));
 sg13g2_a21oi_1 _20539_ (.A1(net240),
    .A2(_09197_),
    .Y(_03106_),
    .B1(_03105_));
 sg13g2_nor3_1 _20540_ (.A(net212),
    .B(net222),
    .C(_03106_),
    .Y(_03107_));
 sg13g2_buf_2 _20541_ (.A(_03107_),
    .X(_03108_));
 sg13g2_a21oi_2 _20542_ (.B1(_10003_),
    .Y(_03109_),
    .A2(net270),
    .A1(net280));
 sg13g2_nand2_1 _20543_ (.Y(_03110_),
    .A(net240),
    .B(_03109_));
 sg13g2_o21ai_1 _20544_ (.B1(_03110_),
    .Y(_03111_),
    .A1(_09020_),
    .A2(net222));
 sg13g2_buf_2 _20545_ (.A(_03111_),
    .X(_03112_));
 sg13g2_nor2_1 _20546_ (.A(net151),
    .B(net149),
    .Y(_03113_));
 sg13g2_buf_1 _20547_ (.A(_03113_),
    .X(_03114_));
 sg13g2_nor2_1 _20548_ (.A(_03112_),
    .B(net113),
    .Y(_03115_));
 sg13g2_nand2_2 _20549_ (.Y(_03116_),
    .A(_03091_),
    .B(_03023_));
 sg13g2_buf_1 _20550_ (.A(_03050_),
    .X(_03117_));
 sg13g2_o21ai_1 _20551_ (.B1(net206),
    .Y(_03118_),
    .A1(_03116_),
    .A2(net268));
 sg13g2_nor2_1 _20552_ (.A(_09040_),
    .B(_03004_),
    .Y(_03119_));
 sg13g2_buf_1 _20553_ (.A(_03119_),
    .X(_03120_));
 sg13g2_nand2_1 _20554_ (.Y(_03121_),
    .A(_09079_),
    .B(_03120_));
 sg13g2_buf_1 _20555_ (.A(_03121_),
    .X(_03122_));
 sg13g2_buf_1 _20556_ (.A(_03122_),
    .X(_03123_));
 sg13g2_nand2_1 _20557_ (.Y(_03124_),
    .A(_10008_),
    .B(_03006_));
 sg13g2_buf_2 _20558_ (.A(_03124_),
    .X(_03125_));
 sg13g2_o21ai_1 _20559_ (.B1(_03125_),
    .Y(_03126_),
    .A1(net222),
    .A2(net112));
 sg13g2_a21oi_1 _20560_ (.A1(_03112_),
    .A2(_03118_),
    .Y(_03127_),
    .B1(_03126_));
 sg13g2_nor2_1 _20561_ (.A(_03115_),
    .B(_03127_),
    .Y(_03128_));
 sg13g2_o21ai_1 _20562_ (.B1(net115),
    .Y(_03129_),
    .A1(_03108_),
    .A2(_03128_));
 sg13g2_o21ai_1 _20563_ (.B1(_03129_),
    .Y(_00757_),
    .A1(_10649_),
    .A2(_09994_));
 sg13g2_o21ai_1 _20564_ (.B1(_03125_),
    .Y(_03130_),
    .A1(_09174_),
    .A2(net112));
 sg13g2_nand2_1 _20565_ (.Y(_03131_),
    .A(_09153_),
    .B(_03079_));
 sg13g2_nor2_1 _20566_ (.A(net268),
    .B(_03131_),
    .Y(_03132_));
 sg13g2_buf_1 _20567_ (.A(_03132_),
    .X(_03133_));
 sg13g2_a21o_1 _20568_ (.A2(net144),
    .A1(net222),
    .B1(_03122_),
    .X(_03134_));
 sg13g2_buf_1 _20569_ (.A(_03134_),
    .X(_03135_));
 sg13g2_nor2_1 _20570_ (.A(net211),
    .B(_03133_),
    .Y(_03136_));
 sg13g2_o21ai_1 _20571_ (.B1(net223),
    .Y(_03137_),
    .A1(net210),
    .A2(net166));
 sg13g2_o21ai_1 _20572_ (.B1(net239),
    .Y(_03138_),
    .A1(_09081_),
    .A2(net210));
 sg13g2_nand2_1 _20573_ (.Y(_03139_),
    .A(_03137_),
    .B(_03138_));
 sg13g2_o21ai_1 _20574_ (.B1(_03139_),
    .Y(_03140_),
    .A1(_03135_),
    .A2(_03136_));
 sg13g2_a221oi_1 _20575_ (.B2(_03112_),
    .C1(_03108_),
    .B1(_03140_),
    .A1(net113),
    .Y(_03141_),
    .A2(_03130_));
 sg13g2_nor2_1 _20576_ (.A(\cpu.dec.imm[11] ),
    .B(net114),
    .Y(_03142_));
 sg13g2_a21oi_1 _20577_ (.A1(net120),
    .A2(_03141_),
    .Y(_00758_),
    .B1(_03142_));
 sg13g2_o21ai_1 _20578_ (.B1(_03125_),
    .Y(_03143_),
    .A1(net281),
    .A2(net112));
 sg13g2_nor2_1 _20579_ (.A(_09136_),
    .B(net144),
    .Y(_03144_));
 sg13g2_o21ai_1 _20580_ (.B1(_03139_),
    .Y(_03145_),
    .A1(_03135_),
    .A2(_03144_));
 sg13g2_a221oi_1 _20581_ (.B2(_03112_),
    .C1(_03108_),
    .B1(_03145_),
    .A1(net113),
    .Y(_03146_),
    .A2(_03143_));
 sg13g2_nor2_1 _20582_ (.A(\cpu.dec.imm[12] ),
    .B(net114),
    .Y(_03147_));
 sg13g2_a21oi_1 _20583_ (.A1(net120),
    .A2(_03146_),
    .Y(_00759_),
    .B1(_03147_));
 sg13g2_nor3_1 _20584_ (.A(net269),
    .B(net180),
    .C(net151),
    .Y(_03148_));
 sg13g2_nor2_1 _20585_ (.A(_10008_),
    .B(net144),
    .Y(_03149_));
 sg13g2_o21ai_1 _20586_ (.B1(_03139_),
    .Y(_03150_),
    .A1(_03135_),
    .A2(_03149_));
 sg13g2_a221oi_1 _20587_ (.B2(_03112_),
    .C1(_03108_),
    .B1(_03150_),
    .A1(net206),
    .Y(_03151_),
    .A2(_03148_));
 sg13g2_nor2_1 _20588_ (.A(\cpu.dec.imm[13] ),
    .B(net115),
    .Y(_03152_));
 sg13g2_a21oi_1 _20589_ (.A1(net120),
    .A2(_03151_),
    .Y(_00760_),
    .B1(_03152_));
 sg13g2_nor2_1 _20590_ (.A(net208),
    .B(net144),
    .Y(_03153_));
 sg13g2_o21ai_1 _20591_ (.B1(_03139_),
    .Y(_03154_),
    .A1(_03135_),
    .A2(_03153_));
 sg13g2_a21oi_1 _20592_ (.A1(_03112_),
    .A2(_03154_),
    .Y(_03155_),
    .B1(_03108_));
 sg13g2_o21ai_1 _20593_ (.B1(_03125_),
    .Y(_03156_),
    .A1(_09117_),
    .A2(net112));
 sg13g2_nand2_1 _20594_ (.Y(_03157_),
    .A(net113),
    .B(_03156_));
 sg13g2_a21oi_1 _20595_ (.A1(_03155_),
    .A2(_03157_),
    .Y(_03158_),
    .B1(net106));
 sg13g2_a21o_1 _20596_ (.A2(_03028_),
    .A1(\cpu.dec.imm[14] ),
    .B1(_03158_),
    .X(_00761_));
 sg13g2_o21ai_1 _20597_ (.B1(_03125_),
    .Y(_03159_),
    .A1(net208),
    .A2(net112));
 sg13g2_nand2_1 _20598_ (.Y(_03160_),
    .A(net113),
    .B(_03159_));
 sg13g2_a21oi_1 _20599_ (.A1(_03155_),
    .A2(_03160_),
    .Y(_03161_),
    .B1(net106));
 sg13g2_a21o_1 _20600_ (.A2(_03028_),
    .A1(\cpu.dec.imm[15] ),
    .B1(_03161_),
    .X(_00762_));
 sg13g2_nor3_2 _20601_ (.A(net279),
    .B(net151),
    .C(net206),
    .Y(_03162_));
 sg13g2_nor2_1 _20602_ (.A(_03008_),
    .B(_03162_),
    .Y(_03163_));
 sg13g2_nand2_1 _20603_ (.Y(_03164_),
    .A(_10001_),
    .B(_03010_));
 sg13g2_or3_1 _20604_ (.A(_09040_),
    .B(_09081_),
    .C(_03100_),
    .X(_03165_));
 sg13g2_buf_1 _20605_ (.A(_03165_),
    .X(_03166_));
 sg13g2_nand2_1 _20606_ (.Y(_03167_),
    .A(net212),
    .B(net206));
 sg13g2_nor3_2 _20607_ (.A(_03117_),
    .B(_03122_),
    .C(_03131_),
    .Y(_03168_));
 sg13g2_nor3_1 _20608_ (.A(net150),
    .B(_03167_),
    .C(_03168_),
    .Y(_03169_));
 sg13g2_a21oi_1 _20609_ (.A1(net150),
    .A2(_03166_),
    .Y(_03170_),
    .B1(_03169_));
 sg13g2_o21ai_1 _20610_ (.B1(_09136_),
    .Y(_03171_),
    .A1(net179),
    .A2(_03170_));
 sg13g2_o21ai_1 _20611_ (.B1(_03171_),
    .Y(_03172_),
    .A1(_03163_),
    .A2(_03164_));
 sg13g2_mux2_1 _20612_ (.A0(_03172_),
    .A1(_10796_),
    .S(net91),
    .X(_00763_));
 sg13g2_inv_1 _20613_ (.Y(_03173_),
    .A(_10805_));
 sg13g2_nor2_1 _20614_ (.A(_09083_),
    .B(_09222_),
    .Y(_03174_));
 sg13g2_a21oi_1 _20615_ (.A1(net211),
    .A2(_03168_),
    .Y(_03175_),
    .B1(_03174_));
 sg13g2_o21ai_1 _20616_ (.B1(net177),
    .Y(_03176_),
    .A1(net238),
    .A2(_03109_));
 sg13g2_a21oi_1 _20617_ (.A1(_03109_),
    .A2(_03175_),
    .Y(_03177_),
    .B1(_03176_));
 sg13g2_nand2_1 _20618_ (.Y(_03178_),
    .A(_10025_),
    .B(_09150_));
 sg13g2_o21ai_1 _20619_ (.B1(_03178_),
    .Y(_03179_),
    .A1(_10025_),
    .A2(_09222_));
 sg13g2_nand2_1 _20620_ (.Y(_03180_),
    .A(_03104_),
    .B(_03179_));
 sg13g2_o21ai_1 _20621_ (.B1(_03180_),
    .Y(_03181_),
    .A1(_09153_),
    .A2(_03104_));
 sg13g2_inv_1 _20622_ (.Y(_03182_),
    .A(_03166_));
 sg13g2_a21o_1 _20623_ (.A2(_03182_),
    .A1(_09101_),
    .B1(_03174_),
    .X(_03183_));
 sg13g2_a22oi_1 _20624_ (.Y(_03184_),
    .B1(_03183_),
    .B2(net113),
    .A2(_03181_),
    .A1(_10032_));
 sg13g2_o21ai_1 _20625_ (.B1(_03184_),
    .Y(_03185_),
    .A1(net222),
    .A2(_03163_));
 sg13g2_o21ai_1 _20626_ (.B1(net115),
    .Y(_03186_),
    .A1(_03177_),
    .A2(_03185_));
 sg13g2_o21ai_1 _20627_ (.B1(_03186_),
    .Y(_00764_),
    .A1(_03173_),
    .A2(net118));
 sg13g2_o21ai_1 _20628_ (.B1(net208),
    .Y(_03187_),
    .A1(_03167_),
    .A2(_03168_));
 sg13g2_nand3_1 _20629_ (.B(_03002_),
    .C(_03109_),
    .A(net211),
    .Y(_03188_));
 sg13g2_a21oi_1 _20630_ (.A1(_03187_),
    .A2(_03188_),
    .Y(_03189_),
    .B1(net168));
 sg13g2_nand2_1 _20631_ (.Y(_03190_),
    .A(net269),
    .B(_03104_));
 sg13g2_nor2_1 _20632_ (.A(net222),
    .B(_03190_),
    .Y(_03191_));
 sg13g2_a21oi_1 _20633_ (.A1(net208),
    .A2(_03190_),
    .Y(_03192_),
    .B1(_03191_));
 sg13g2_nor2_1 _20634_ (.A(_03097_),
    .B(_03192_),
    .Y(_03193_));
 sg13g2_a22oi_1 _20635_ (.Y(_03194_),
    .B1(_03182_),
    .B2(net208),
    .A2(net149),
    .A1(net211));
 sg13g2_nor2_1 _20636_ (.A(_09201_),
    .B(_03194_),
    .Y(_03195_));
 sg13g2_a21oi_1 _20637_ (.A1(_10015_),
    .A2(_03109_),
    .Y(_03196_),
    .B1(_03114_));
 sg13g2_inv_1 _20638_ (.Y(_03197_),
    .A(_09256_));
 sg13g2_a22oi_1 _20639_ (.Y(_03198_),
    .B1(_03006_),
    .B2(_09102_),
    .A2(_03197_),
    .A1(_09198_));
 sg13g2_nor2_1 _20640_ (.A(_03196_),
    .B(_03198_),
    .Y(_03199_));
 sg13g2_nor4_1 _20641_ (.A(_03189_),
    .B(_03193_),
    .C(_03195_),
    .D(_03199_),
    .Y(_03200_));
 sg13g2_nand2_1 _20642_ (.Y(_03201_),
    .A(_10937_),
    .B(net89));
 sg13g2_o21ai_1 _20643_ (.B1(_03201_),
    .Y(_00765_),
    .A1(net92),
    .A2(_03200_));
 sg13g2_a21oi_1 _20644_ (.A1(net225),
    .A2(net144),
    .Y(_03202_),
    .B1(net270));
 sg13g2_nor2_1 _20645_ (.A(_03022_),
    .B(_03202_),
    .Y(_03203_));
 sg13g2_nor3_1 _20646_ (.A(net167),
    .B(net179),
    .C(_03203_),
    .Y(_03204_));
 sg13g2_nand4_1 _20647_ (.B(net206),
    .C(_03008_),
    .A(net208),
    .Y(_03205_),
    .D(_03010_));
 sg13g2_o21ai_1 _20648_ (.B1(_03205_),
    .Y(_03206_),
    .A1(net180),
    .A2(_03204_));
 sg13g2_mux2_1 _20649_ (.A0(_03206_),
    .A1(\cpu.dec.imm[4] ),
    .S(net91),
    .X(_00766_));
 sg13g2_o21ai_1 _20650_ (.B1(net209),
    .Y(_03207_),
    .A1(net168),
    .A2(net179));
 sg13g2_or4_1 _20651_ (.A(net168),
    .B(_09197_),
    .C(_09174_),
    .D(_03100_),
    .X(_03208_));
 sg13g2_a21oi_1 _20652_ (.A1(_03207_),
    .A2(_03208_),
    .Y(_03209_),
    .B1(net178));
 sg13g2_o21ai_1 _20653_ (.B1(net207),
    .Y(_03210_),
    .A1(net112),
    .A2(net144));
 sg13g2_o21ai_1 _20654_ (.B1(_03210_),
    .Y(_03211_),
    .A1(net224),
    .A2(net226));
 sg13g2_nand3_1 _20655_ (.B(net209),
    .C(_03211_),
    .A(net178),
    .Y(_03212_));
 sg13g2_nand2b_1 _20656_ (.Y(_03213_),
    .B(_03212_),
    .A_N(_03209_));
 sg13g2_mux2_1 _20657_ (.A0(_03213_),
    .A1(\cpu.dec.imm[5] ),
    .S(_09264_),
    .X(_00767_));
 sg13g2_buf_1 _20658_ (.A(_03078_),
    .X(_03214_));
 sg13g2_nor2_1 _20659_ (.A(net279),
    .B(_09197_),
    .Y(_03215_));
 sg13g2_a21oi_1 _20660_ (.A1(net267),
    .A2(_03215_),
    .Y(_03216_),
    .B1(_03174_));
 sg13g2_nand2_1 _20661_ (.Y(_03217_),
    .A(net226),
    .B(net267));
 sg13g2_nand3_1 _20662_ (.B(net211),
    .C(_03006_),
    .A(net178),
    .Y(_03218_));
 sg13g2_o21ai_1 _20663_ (.B1(_03218_),
    .Y(_03219_),
    .A1(_03110_),
    .A2(_03217_));
 sg13g2_inv_1 _20664_ (.Y(_03220_),
    .A(_03168_));
 sg13g2_a21oi_1 _20665_ (.A1(net206),
    .A2(_03220_),
    .Y(_03221_),
    .B1(_09020_));
 sg13g2_a21oi_1 _20666_ (.A1(_10032_),
    .A2(_03190_),
    .Y(_03222_),
    .B1(_03221_));
 sg13g2_nor2_1 _20667_ (.A(_09222_),
    .B(_03222_),
    .Y(_03223_));
 sg13g2_nor3_1 _20668_ (.A(_03088_),
    .B(_03219_),
    .C(_03223_),
    .Y(_03224_));
 sg13g2_a21oi_1 _20669_ (.A1(_03088_),
    .A2(_03216_),
    .Y(_03225_),
    .B1(_03224_));
 sg13g2_mux2_1 _20670_ (.A0(_03225_),
    .A1(\cpu.dec.imm[6] ),
    .S(net91),
    .X(_00768_));
 sg13g2_nand2_1 _20671_ (.Y(_03226_),
    .A(_03197_),
    .B(_03221_));
 sg13g2_nand3_1 _20672_ (.B(net270),
    .C(_03098_),
    .A(net225),
    .Y(_03227_));
 sg13g2_nor2_1 _20673_ (.A(net279),
    .B(net268),
    .Y(_03228_));
 sg13g2_nand3b_1 _20674_ (.B(_03228_),
    .C(_03088_),
    .Y(_03229_),
    .A_N(_03090_));
 sg13g2_a21oi_1 _20675_ (.A1(_09136_),
    .A2(_03008_),
    .Y(_03230_),
    .B1(_03108_));
 sg13g2_nand4_1 _20676_ (.B(_03227_),
    .C(_03229_),
    .A(_03226_),
    .Y(_03231_),
    .D(_03230_));
 sg13g2_mux2_1 _20677_ (.A0(_03231_),
    .A1(\cpu.dec.imm[7] ),
    .S(_09264_),
    .X(_00769_));
 sg13g2_nor2_1 _20678_ (.A(net209),
    .B(net144),
    .Y(_03232_));
 sg13g2_nand2_1 _20679_ (.Y(_03233_),
    .A(net206),
    .B(_03125_));
 sg13g2_a21oi_1 _20680_ (.A1(net226),
    .A2(net344),
    .Y(_03234_),
    .B1(_03233_));
 sg13g2_o21ai_1 _20681_ (.B1(_03234_),
    .Y(_03235_),
    .A1(_03135_),
    .A2(_03232_));
 sg13g2_o21ai_1 _20682_ (.B1(_03125_),
    .Y(_03236_),
    .A1(_09240_),
    .A2(net112));
 sg13g2_nand3_1 _20683_ (.B(net344),
    .C(_03215_),
    .A(_03088_),
    .Y(_03237_));
 sg13g2_nand2b_1 _20684_ (.Y(_03238_),
    .B(_03237_),
    .A_N(_03108_));
 sg13g2_a221oi_1 _20685_ (.B2(net113),
    .C1(_03238_),
    .B1(_03236_),
    .A1(_03112_),
    .Y(_03239_),
    .A2(_03235_));
 sg13g2_nor2_1 _20686_ (.A(\cpu.dec.imm[8] ),
    .B(net115),
    .Y(_03240_));
 sg13g2_a21oi_1 _20687_ (.A1(net120),
    .A2(_03239_),
    .Y(_00770_),
    .B1(_03240_));
 sg13g2_o21ai_1 _20688_ (.B1(_03125_),
    .Y(_03241_),
    .A1(_09222_),
    .A2(net112));
 sg13g2_nor2_1 _20689_ (.A(_10001_),
    .B(net144),
    .Y(_03242_));
 sg13g2_a21oi_1 _20690_ (.A1(net238),
    .A2(net226),
    .Y(_03243_),
    .B1(_03233_));
 sg13g2_o21ai_1 _20691_ (.B1(_03243_),
    .Y(_03244_),
    .A1(_03135_),
    .A2(_03242_));
 sg13g2_a221oi_1 _20692_ (.B2(_03112_),
    .C1(_03108_),
    .B1(_03244_),
    .A1(net113),
    .Y(_03245_),
    .A2(_03241_));
 sg13g2_nor2_1 _20693_ (.A(\cpu.dec.imm[9] ),
    .B(_03012_),
    .Y(_03246_));
 sg13g2_a21oi_1 _20694_ (.A1(net120),
    .A2(_03245_),
    .Y(_00771_),
    .B1(_03246_));
 sg13g2_buf_1 _20695_ (.A(_08533_),
    .X(_03247_));
 sg13g2_nand2_1 _20696_ (.Y(_03248_),
    .A(_03247_),
    .B(_09136_));
 sg13g2_nor4_1 _20697_ (.A(_09170_),
    .B(_03034_),
    .C(_03083_),
    .D(_03248_),
    .Y(_03249_));
 sg13g2_a21o_1 _20698_ (.A2(net87),
    .A1(\cpu.dec.do_inv_mmu ),
    .B1(_03249_),
    .X(_00772_));
 sg13g2_nor3_1 _20699_ (.A(net106),
    .B(_09201_),
    .C(_03166_),
    .Y(_03250_));
 sg13g2_a21o_1 _20700_ (.A2(net87),
    .A1(\cpu.dec.io ),
    .B1(_03250_),
    .X(_00773_));
 sg13g2_nor2_1 _20701_ (.A(_10001_),
    .B(_09238_),
    .Y(_03251_));
 sg13g2_nand4_1 _20702_ (.B(_09174_),
    .C(_09256_),
    .A(net281),
    .Y(_03252_),
    .D(_03251_));
 sg13g2_buf_2 _20703_ (.A(_03252_),
    .X(_03253_));
 sg13g2_nor4_1 _20704_ (.A(_09170_),
    .B(net152),
    .C(_03097_),
    .D(_03253_),
    .Y(_03254_));
 sg13g2_a21o_1 _20705_ (.A2(net87),
    .A1(\cpu.dec.jmp ),
    .B1(_03254_),
    .X(_00774_));
 sg13g2_inv_1 _20706_ (.Y(_03255_),
    .A(_11669_));
 sg13g2_o21ai_1 _20707_ (.B1(net212),
    .Y(_03256_),
    .A1(net207),
    .A2(net223));
 sg13g2_nand3_1 _20708_ (.B(net166),
    .C(_03256_),
    .A(net119),
    .Y(_03257_));
 sg13g2_o21ai_1 _20709_ (.B1(_03257_),
    .Y(_00775_),
    .A1(_03255_),
    .A2(net118));
 sg13g2_nor4_1 _20710_ (.A(net108),
    .B(_09175_),
    .C(_10008_),
    .D(_09203_),
    .Y(_03258_));
 sg13g2_a21o_1 _20711_ (.A2(net87),
    .A1(_09455_),
    .B1(_03258_),
    .X(_00776_));
 sg13g2_nor2_1 _20712_ (.A(_10013_),
    .B(net180),
    .Y(_03259_));
 sg13g2_o21ai_1 _20713_ (.B1(_10014_),
    .Y(_03260_),
    .A1(_09154_),
    .A2(_03259_));
 sg13g2_a21oi_1 _20714_ (.A1(net224),
    .A2(_09194_),
    .Y(_03261_),
    .B1(_03097_));
 sg13g2_buf_1 _20715_ (.A(_09081_),
    .X(_03262_));
 sg13g2_o21ai_1 _20716_ (.B1(_03262_),
    .Y(_03263_),
    .A1(_09202_),
    .A2(_03261_));
 sg13g2_o21ai_1 _20717_ (.B1(_03263_),
    .Y(_03264_),
    .A1(net152),
    .A2(_03260_));
 sg13g2_o21ai_1 _20718_ (.B1(_03010_),
    .Y(_03265_),
    .A1(_03162_),
    .A2(_03264_));
 sg13g2_nand2_1 _20719_ (.Y(_03266_),
    .A(net915),
    .B(net89));
 sg13g2_o21ai_1 _20720_ (.B1(_03266_),
    .Y(_00777_),
    .A1(net92),
    .A2(_03265_));
 sg13g2_nor3_1 _20721_ (.A(_09195_),
    .B(_09194_),
    .C(_03253_),
    .Y(_03267_));
 sg13g2_a21o_1 _20722_ (.A2(_03253_),
    .A1(net267),
    .B1(_03267_),
    .X(_03268_));
 sg13g2_a22oi_1 _20723_ (.Y(_03269_),
    .B1(_03268_),
    .B2(net165),
    .A2(_03214_),
    .A1(_03021_));
 sg13g2_nand2_1 _20724_ (.Y(_03270_),
    .A(_03023_),
    .B(_03214_));
 sg13g2_o21ai_1 _20725_ (.B1(_03270_),
    .Y(_03271_),
    .A1(net223),
    .A2(_09240_));
 sg13g2_a22oi_1 _20726_ (.Y(_03272_),
    .B1(net166),
    .B2(_03271_),
    .A2(net267),
    .A1(_09197_));
 sg13g2_inv_1 _20727_ (.Y(_03273_),
    .A(_03272_));
 sg13g2_inv_1 _20728_ (.Y(_03274_),
    .A(_03104_));
 sg13g2_a21oi_1 _20729_ (.A1(_03116_),
    .A2(net267),
    .Y(_03275_),
    .B1(_03274_));
 sg13g2_nor2_1 _20730_ (.A(net226),
    .B(_03010_),
    .Y(_03276_));
 sg13g2_o21ai_1 _20731_ (.B1(_03276_),
    .Y(_03277_),
    .A1(net239),
    .A2(_09239_));
 sg13g2_o21ai_1 _20732_ (.B1(_03277_),
    .Y(_03278_),
    .A1(_09020_),
    .A2(_03275_));
 sg13g2_a22oi_1 _20733_ (.Y(_03279_),
    .B1(_03278_),
    .B2(_03029_),
    .A2(_03273_),
    .A1(_10005_));
 sg13g2_o21ai_1 _20734_ (.B1(_03279_),
    .Y(_03280_),
    .A1(_03097_),
    .A2(_03269_));
 sg13g2_mux2_1 _20735_ (.A0(_03280_),
    .A1(\cpu.dec.r_rd[0] ),
    .S(net91),
    .X(_00778_));
 sg13g2_a21oi_1 _20736_ (.A1(net165),
    .A2(_03253_),
    .Y(_03281_),
    .B1(net224));
 sg13g2_inv_1 _20737_ (.Y(_03282_),
    .A(_09020_));
 sg13g2_o21ai_1 _20738_ (.B1(_03282_),
    .Y(_03283_),
    .A1(net165),
    .A2(net166));
 sg13g2_o21ai_1 _20739_ (.B1(_03283_),
    .Y(_03284_),
    .A1(_03097_),
    .A2(_03281_));
 sg13g2_nand2b_1 _20740_ (.Y(_03285_),
    .B(_03284_),
    .A_N(_03117_));
 sg13g2_a21oi_1 _20741_ (.A1(net279),
    .A2(_09222_),
    .Y(_03286_),
    .B1(net239));
 sg13g2_o21ai_1 _20742_ (.B1(net270),
    .Y(_03287_),
    .A1(_03228_),
    .A2(_03286_));
 sg13g2_o21ai_1 _20743_ (.B1(_03287_),
    .Y(_03288_),
    .A1(net268),
    .A2(_03123_));
 sg13g2_nor3_1 _20744_ (.A(_09175_),
    .B(_03095_),
    .C(_03083_),
    .Y(_03289_));
 sg13g2_and2_1 _20745_ (.A(_10042_),
    .B(_03289_),
    .X(_03290_));
 sg13g2_buf_1 _20746_ (.A(_03290_),
    .X(_03291_));
 sg13g2_nand2b_1 _20747_ (.Y(_03292_),
    .B(net149),
    .A_N(_03291_));
 sg13g2_nand3_1 _20748_ (.B(_03288_),
    .C(_03292_),
    .A(net150),
    .Y(_03293_));
 sg13g2_nand3_1 _20749_ (.B(_10001_),
    .C(_03276_),
    .A(net224),
    .Y(_03294_));
 sg13g2_nand3_1 _20750_ (.B(_03293_),
    .C(_03294_),
    .A(_03285_),
    .Y(_03295_));
 sg13g2_mux2_1 _20751_ (.A0(_03295_),
    .A1(\cpu.dec.r_rd[1] ),
    .S(net89),
    .X(_00779_));
 sg13g2_nand2_1 _20752_ (.Y(_03296_),
    .A(net223),
    .B(net344));
 sg13g2_o21ai_1 _20753_ (.B1(_03296_),
    .Y(_03297_),
    .A1(net223),
    .A2(_03095_));
 sg13g2_a22oi_1 _20754_ (.Y(_03298_),
    .B1(net166),
    .B2(_03297_),
    .A2(net344),
    .A1(net179));
 sg13g2_nand3_1 _20755_ (.B(_03197_),
    .C(_03276_),
    .A(_03021_),
    .Y(_03299_));
 sg13g2_o21ai_1 _20756_ (.B1(_03299_),
    .Y(_03300_),
    .A1(net151),
    .A2(_03298_));
 sg13g2_a21oi_1 _20757_ (.A1(net344),
    .A2(_03284_),
    .Y(_03301_),
    .B1(_03300_));
 sg13g2_nor2_1 _20758_ (.A(\cpu.dec.r_rd[2] ),
    .B(net115),
    .Y(_03302_));
 sg13g2_a21oi_1 _20759_ (.A1(net120),
    .A2(_03301_),
    .Y(_00780_),
    .B1(_03302_));
 sg13g2_nand3_1 _20760_ (.B(net239),
    .C(_03253_),
    .A(_03018_),
    .Y(_03303_));
 sg13g2_nand2_1 _20761_ (.Y(_03304_),
    .A(net168),
    .B(_03303_));
 sg13g2_a21oi_1 _20762_ (.A1(net165),
    .A2(_03304_),
    .Y(_03305_),
    .B1(net166));
 sg13g2_nand2_1 _20763_ (.Y(_03306_),
    .A(net238),
    .B(_03010_));
 sg13g2_a21oi_1 _20764_ (.A1(net207),
    .A2(net225),
    .Y(_03307_),
    .B1(net165));
 sg13g2_a21oi_1 _20765_ (.A1(net212),
    .A2(net279),
    .Y(_03308_),
    .B1(net207));
 sg13g2_nand2b_1 _20766_ (.Y(_03309_),
    .B(net270),
    .A_N(_03308_));
 sg13g2_o21ai_1 _20767_ (.B1(_03309_),
    .Y(_03310_),
    .A1(net178),
    .A2(_03307_));
 sg13g2_a22oi_1 _20768_ (.Y(_03311_),
    .B1(_03310_),
    .B2(net224),
    .A2(net179),
    .A1(net178));
 sg13g2_o21ai_1 _20769_ (.B1(_03311_),
    .Y(_03312_),
    .A1(_03305_),
    .A2(_03306_));
 sg13g2_mux2_1 _20770_ (.A0(_03312_),
    .A1(\cpu.dec.r_rd[3] ),
    .S(net89),
    .X(_00781_));
 sg13g2_o21ai_1 _20771_ (.B1(_03116_),
    .Y(_03313_),
    .A1(net269),
    .A2(_03024_));
 sg13g2_a21oi_1 _20772_ (.A1(_09193_),
    .A2(_03253_),
    .Y(_03314_),
    .B1(net152));
 sg13g2_or2_1 _20773_ (.X(_03315_),
    .B(_03314_),
    .A(_03215_));
 sg13g2_nand2_1 _20774_ (.Y(_03316_),
    .A(net207),
    .B(net269));
 sg13g2_o21ai_1 _20775_ (.B1(_03316_),
    .Y(_03317_),
    .A1(net207),
    .A2(_03315_));
 sg13g2_a21oi_1 _20776_ (.A1(net168),
    .A2(net165),
    .Y(_03318_),
    .B1(_03100_));
 sg13g2_o21ai_1 _20777_ (.B1(net267),
    .Y(_03319_),
    .A1(_03024_),
    .A2(_03318_));
 sg13g2_a221oi_1 _20778_ (.B2(net167),
    .C1(_03319_),
    .B1(_03317_),
    .A1(net177),
    .Y(_03320_),
    .A2(_03313_));
 sg13g2_o21ai_1 _20779_ (.B1(net115),
    .Y(_03321_),
    .A1(_03011_),
    .A2(_03320_));
 sg13g2_o21ai_1 _20780_ (.B1(_03321_),
    .Y(_00782_),
    .A1(_11152_),
    .A2(net118));
 sg13g2_a21oi_1 _20781_ (.A1(_03014_),
    .A2(net268),
    .Y(_03322_),
    .B1(_09197_));
 sg13g2_nand2_1 _20782_ (.Y(_03323_),
    .A(net207),
    .B(_03322_));
 sg13g2_o21ai_1 _20783_ (.B1(_03323_),
    .Y(_03324_),
    .A1(net177),
    .A2(net269));
 sg13g2_o21ai_1 _20784_ (.B1(net224),
    .Y(_03325_),
    .A1(_03015_),
    .A2(_03131_));
 sg13g2_a21o_1 _20785_ (.A2(_03325_),
    .A1(_03014_),
    .B1(net165),
    .X(_03326_));
 sg13g2_nor2_1 _20786_ (.A(_09020_),
    .B(net268),
    .Y(_03327_));
 sg13g2_a22oi_1 _20787_ (.Y(_03328_),
    .B1(_03315_),
    .B2(_10032_),
    .A2(_03123_),
    .A1(net150));
 sg13g2_a21oi_1 _20788_ (.A1(_03034_),
    .A2(net268),
    .Y(_03329_),
    .B1(_03328_));
 sg13g2_a221oi_1 _20789_ (.B2(_03327_),
    .C1(_03329_),
    .B1(_03326_),
    .A1(net167),
    .Y(_03330_),
    .A2(_03324_));
 sg13g2_nand2_1 _20790_ (.Y(_03331_),
    .A(_11069_),
    .B(net89));
 sg13g2_o21ai_1 _20791_ (.B1(_03331_),
    .Y(_00783_),
    .A1(net92),
    .A2(_03330_));
 sg13g2_and3_1 _20792_ (.X(_03332_),
    .A(net225),
    .B(_03088_),
    .C(net344));
 sg13g2_nand3b_1 _20793_ (.B(_03282_),
    .C(_03116_),
    .Y(_03333_),
    .A_N(net166));
 sg13g2_o21ai_1 _20794_ (.B1(_03010_),
    .Y(_03334_),
    .A1(_03162_),
    .A2(net344));
 sg13g2_a21oi_1 _20795_ (.A1(_03328_),
    .A2(_03333_),
    .Y(_03335_),
    .B1(_03334_));
 sg13g2_o21ai_1 _20796_ (.B1(net119),
    .Y(_03336_),
    .A1(_03332_),
    .A2(_03335_));
 sg13g2_o21ai_1 _20797_ (.B1(_03336_),
    .Y(_00784_),
    .A1(net673),
    .A2(net118));
 sg13g2_nand2_1 _20798_ (.Y(_03337_),
    .A(net238),
    .B(_03314_));
 sg13g2_nor2_1 _20799_ (.A(net178),
    .B(_03215_),
    .Y(_03338_));
 sg13g2_mux2_1 _20800_ (.A0(net223),
    .A1(net165),
    .S(net178),
    .X(_03339_));
 sg13g2_a22oi_1 _20801_ (.Y(_03340_),
    .B1(_03339_),
    .B2(net224),
    .A2(_03338_),
    .A1(_03337_));
 sg13g2_inv_1 _20802_ (.Y(_03341_),
    .A(_03256_));
 sg13g2_a21oi_1 _20803_ (.A1(net178),
    .A2(net270),
    .Y(_03342_),
    .B1(_03316_));
 sg13g2_a21oi_1 _20804_ (.A1(net166),
    .A2(_03341_),
    .Y(_03343_),
    .B1(_03342_));
 sg13g2_o21ai_1 _20805_ (.B1(_03343_),
    .Y(_03344_),
    .A1(net177),
    .A2(_03340_));
 sg13g2_nand2_1 _20806_ (.Y(_03345_),
    .A(_11222_),
    .B(net89));
 sg13g2_o21ai_1 _20807_ (.B1(_03345_),
    .Y(_00785_),
    .A1(net92),
    .A2(_03344_));
 sg13g2_o21ai_1 _20808_ (.B1(_09197_),
    .Y(_03346_),
    .A1(_09999_),
    .A2(_03251_));
 sg13g2_nand3_1 _20809_ (.B(_03104_),
    .C(_03346_),
    .A(net150),
    .Y(_03347_));
 sg13g2_inv_1 _20810_ (.Y(_03348_),
    .A(_03347_));
 sg13g2_a21oi_1 _20811_ (.A1(_10032_),
    .A2(_03006_),
    .Y(_03349_),
    .B1(_03348_));
 sg13g2_a22oi_1 _20812_ (.Y(_03350_),
    .B1(_03006_),
    .B2(net267),
    .A2(net209),
    .A1(net179));
 sg13g2_nor2_1 _20813_ (.A(_03097_),
    .B(_03350_),
    .Y(_03351_));
 sg13g2_a21oi_1 _20814_ (.A1(net209),
    .A2(_03349_),
    .Y(_03352_),
    .B1(_03351_));
 sg13g2_nand2_1 _20815_ (.Y(_03353_),
    .A(_10445_),
    .B(net89));
 sg13g2_o21ai_1 _20816_ (.B1(_03353_),
    .Y(_00786_),
    .A1(net92),
    .A2(_03352_));
 sg13g2_nor2_1 _20817_ (.A(_03029_),
    .B(net268),
    .Y(_03354_));
 sg13g2_o21ai_1 _20818_ (.B1(_10032_),
    .Y(_03355_),
    .A1(_03174_),
    .A2(_03354_));
 sg13g2_nand2_1 _20819_ (.Y(_03356_),
    .A(_10001_),
    .B(_03349_));
 sg13g2_a21oi_1 _20820_ (.A1(_03355_),
    .A2(_03356_),
    .Y(_03357_),
    .B1(net106));
 sg13g2_a21o_1 _20821_ (.A2(net91),
    .A1(_10412_),
    .B1(_03357_),
    .X(_00787_));
 sg13g2_nand3_1 _20822_ (.B(_03006_),
    .C(net344),
    .A(_10032_),
    .Y(_03358_));
 sg13g2_o21ai_1 _20823_ (.B1(net269),
    .Y(_03359_),
    .A1(_10003_),
    .A2(_03015_));
 sg13g2_a21oi_1 _20824_ (.A1(_03091_),
    .A2(_10028_),
    .Y(_03360_),
    .B1(_03018_));
 sg13g2_a21oi_1 _20825_ (.A1(net239),
    .A2(_03359_),
    .Y(_03361_),
    .B1(_03360_));
 sg13g2_o21ai_1 _20826_ (.B1(_03197_),
    .Y(_03362_),
    .A1(_10015_),
    .A2(_03361_));
 sg13g2_a21oi_1 _20827_ (.A1(_03358_),
    .A2(_03362_),
    .Y(_03363_),
    .B1(net106));
 sg13g2_a21o_1 _20828_ (.A2(net91),
    .A1(_10420_),
    .B1(_03363_),
    .X(_00788_));
 sg13g2_nor2_1 _20829_ (.A(net152),
    .B(net211),
    .Y(_03364_));
 sg13g2_nor2_1 _20830_ (.A(net238),
    .B(_03029_),
    .Y(_03365_));
 sg13g2_o21ai_1 _20831_ (.B1(_10032_),
    .Y(_03366_),
    .A1(_03364_),
    .A2(_03365_));
 sg13g2_nand3_1 _20832_ (.B(_03347_),
    .C(_03366_),
    .A(net119),
    .Y(_03367_));
 sg13g2_o21ai_1 _20833_ (.B1(_03367_),
    .Y(_00789_),
    .A1(_10548_),
    .A2(net114));
 sg13g2_nand2_1 _20834_ (.Y(_03368_),
    .A(_10371_),
    .B(_10021_));
 sg13g2_o21ai_1 _20835_ (.B1(_03368_),
    .Y(_00790_),
    .A1(_09171_),
    .A2(_09260_));
 sg13g2_nand3_1 _20836_ (.B(_10041_),
    .C(_03251_),
    .A(net119),
    .Y(_03369_));
 sg13g2_o21ai_1 _20837_ (.B1(_03369_),
    .Y(_00791_),
    .A1(net906),
    .A2(_03032_));
 sg13g2_nor3_1 _20838_ (.A(net106),
    .B(net180),
    .C(_09206_),
    .Y(_03370_));
 sg13g2_a21o_1 _20839_ (.A2(net91),
    .A1(\cpu.dec.r_set_cc ),
    .B1(_03370_),
    .X(_00792_));
 sg13g2_nor3_1 _20840_ (.A(net167),
    .B(net177),
    .C(_03116_),
    .Y(_03371_));
 sg13g2_a21oi_1 _20841_ (.A1(net167),
    .A2(_03006_),
    .Y(_03372_),
    .B1(_03371_));
 sg13g2_buf_1 _20842_ (.A(\cpu.dec.r_store ),
    .X(_03373_));
 sg13g2_nor2_1 _20843_ (.A(_03373_),
    .B(net115),
    .Y(_03374_));
 sg13g2_a21oi_1 _20844_ (.A1(net120),
    .A2(_03372_),
    .Y(_00793_),
    .B1(_03374_));
 sg13g2_inv_1 _20845_ (.Y(_03375_),
    .A(\cpu.dec.r_swapsp ));
 sg13g2_nand3_1 _20846_ (.B(_03162_),
    .C(_03291_),
    .A(net119),
    .Y(_03376_));
 sg13g2_o21ai_1 _20847_ (.B1(_03376_),
    .Y(_00794_),
    .A1(_03375_),
    .A2(_03032_));
 sg13g2_inv_1 _20848_ (.Y(_03377_),
    .A(\cpu.dec.r_sys_call ));
 sg13g2_nand4_1 _20849_ (.B(_10007_),
    .C(net149),
    .A(_08972_),
    .Y(_03378_),
    .D(_03289_));
 sg13g2_o21ai_1 _20850_ (.B1(_03378_),
    .Y(_00795_),
    .A1(_03377_),
    .A2(net114));
 sg13g2_a21oi_1 _20851_ (.A1(_09174_),
    .A2(_03081_),
    .Y(_03379_),
    .B1(_09083_));
 sg13g2_nor2b_1 _20852_ (.A(_03379_),
    .B_N(_03276_),
    .Y(_03380_));
 sg13g2_nor3_1 _20853_ (.A(_09101_),
    .B(_09116_),
    .C(_03253_),
    .Y(_03381_));
 sg13g2_nand3_1 _20854_ (.B(_03081_),
    .C(_03381_),
    .A(net149),
    .Y(_03382_));
 sg13g2_o21ai_1 _20855_ (.B1(_09153_),
    .Y(_03383_),
    .A1(net279),
    .A2(_03314_));
 sg13g2_nand2b_1 _20856_ (.Y(_03384_),
    .B(net267),
    .A_N(_03050_));
 sg13g2_xnor2_1 _20857_ (.Y(_03385_),
    .A(_03064_),
    .B(_03384_));
 sg13g2_nand2b_1 _20858_ (.Y(_03386_),
    .B(_03385_),
    .A_N(net955));
 sg13g2_a21oi_1 _20859_ (.A1(_03104_),
    .A2(_03383_),
    .Y(_03387_),
    .B1(_03386_));
 sg13g2_xnor2_1 _20860_ (.Y(_03388_),
    .A(_09241_),
    .B(net222));
 sg13g2_nand2_1 _20861_ (.Y(_03389_),
    .A(_08388_),
    .B(net210));
 sg13g2_o21ai_1 _20862_ (.B1(_03389_),
    .Y(_03390_),
    .A1(net955),
    .A2(net210));
 sg13g2_nand3_1 _20863_ (.B(_03388_),
    .C(_03390_),
    .A(_03364_),
    .Y(_03391_));
 sg13g2_nand2_1 _20864_ (.Y(_03392_),
    .A(_09175_),
    .B(_10008_));
 sg13g2_o21ai_1 _20865_ (.B1(_03392_),
    .Y(_03393_),
    .A1(_10008_),
    .A2(_09240_));
 sg13g2_nand2_1 _20866_ (.Y(_03394_),
    .A(net149),
    .B(_03393_));
 sg13g2_nand4_1 _20867_ (.B(_03085_),
    .C(_03391_),
    .A(_03016_),
    .Y(_03395_),
    .D(_03394_));
 sg13g2_a22oi_1 _20868_ (.Y(_03396_),
    .B1(_09175_),
    .B2(_09117_),
    .A2(_09136_),
    .A1(_09101_));
 sg13g2_nand3_1 _20869_ (.B(net210),
    .C(_09239_),
    .A(_09117_),
    .Y(_03397_));
 sg13g2_o21ai_1 _20870_ (.B1(_03397_),
    .Y(_03398_),
    .A1(net210),
    .A2(_03396_));
 sg13g2_nor3_1 _20871_ (.A(_09101_),
    .B(_03122_),
    .C(_03386_),
    .Y(_03399_));
 sg13g2_a21oi_1 _20872_ (.A1(_09197_),
    .A2(_03398_),
    .Y(_03400_),
    .B1(_03399_));
 sg13g2_o21ai_1 _20873_ (.B1(_10012_),
    .Y(_03401_),
    .A1(net168),
    .A2(_03400_));
 sg13g2_o21ai_1 _20874_ (.B1(_03401_),
    .Y(_03402_),
    .A1(_03387_),
    .A2(_03395_));
 sg13g2_nand3_1 _20875_ (.B(net180),
    .C(_03381_),
    .A(_03247_),
    .Y(_03403_));
 sg13g2_nand2b_1 _20876_ (.Y(_03404_),
    .B(_03403_),
    .A_N(_03085_));
 sg13g2_nor3_1 _20877_ (.A(_08533_),
    .B(_11029_),
    .C(_03100_),
    .Y(_03405_));
 sg13g2_o21ai_1 _20878_ (.B1(_09195_),
    .Y(_03406_),
    .A1(_09081_),
    .A2(_03405_));
 sg13g2_nand2_1 _20879_ (.Y(_03407_),
    .A(_09101_),
    .B(_10008_));
 sg13g2_a21oi_1 _20880_ (.A1(_09150_),
    .A2(_03197_),
    .Y(_03408_),
    .B1(_09136_));
 sg13g2_o21ai_1 _20881_ (.B1(net208),
    .Y(_03409_),
    .A1(_03407_),
    .A2(_03408_));
 sg13g2_a21oi_1 _20882_ (.A1(_03262_),
    .A2(_03409_),
    .Y(_03410_),
    .B1(_03399_));
 sg13g2_nand3_1 _20883_ (.B(_03406_),
    .C(_03410_),
    .A(_03404_),
    .Y(_03411_));
 sg13g2_a21oi_1 _20884_ (.A1(_09173_),
    .A2(_09258_),
    .Y(_03412_),
    .B1(_03083_));
 sg13g2_and2_1 _20885_ (.A(net745),
    .B(_10030_),
    .X(_03413_));
 sg13g2_o21ai_1 _20886_ (.B1(_03413_),
    .Y(_03414_),
    .A1(_03291_),
    .A2(_03412_));
 sg13g2_nand3_1 _20887_ (.B(_03411_),
    .C(_03414_),
    .A(net150),
    .Y(_03415_));
 sg13g2_a22oi_1 _20888_ (.Y(_03416_),
    .B1(_03402_),
    .B2(_03415_),
    .A2(_03382_),
    .A1(_03380_));
 sg13g2_nand2_1 _20889_ (.Y(_03417_),
    .A(net114),
    .B(_03416_));
 sg13g2_o21ai_1 _20890_ (.B1(_03417_),
    .Y(_00796_),
    .A1(_11536_),
    .A2(net114));
 sg13g2_buf_1 _20891_ (.A(net1052),
    .X(_03418_));
 sg13g2_buf_1 _20892_ (.A(_03418_),
    .X(_03419_));
 sg13g2_nand2b_1 _20893_ (.Y(_03420_),
    .B(net1114),
    .A_N(net1113));
 sg13g2_buf_1 _20894_ (.A(_03420_),
    .X(_03421_));
 sg13g2_nand3_1 _20895_ (.B(_10354_),
    .C(net1115),
    .A(net1112),
    .Y(_03422_));
 sg13g2_buf_1 _20896_ (.A(_03422_),
    .X(_03423_));
 sg13g2_nor2_1 _20897_ (.A(_03421_),
    .B(_03423_),
    .Y(_03424_));
 sg13g2_buf_2 _20898_ (.A(_03424_),
    .X(_03425_));
 sg13g2_buf_1 _20899_ (.A(_03425_),
    .X(_03426_));
 sg13g2_mux2_1 _20900_ (.A0(\cpu.ex.r_10[0] ),
    .A1(net744),
    .S(_03426_),
    .X(_00801_));
 sg13g2_mux2_1 _20901_ (.A0(\cpu.ex.r_10[10] ),
    .A1(net881),
    .S(net526),
    .X(_00802_));
 sg13g2_mux2_1 _20902_ (.A0(\cpu.ex.r_10[11] ),
    .A1(net882),
    .S(net526),
    .X(_00803_));
 sg13g2_buf_1 _20903_ (.A(net687),
    .X(_03427_));
 sg13g2_mux2_1 _20904_ (.A0(\cpu.ex.r_10[12] ),
    .A1(net601),
    .S(net526),
    .X(_00804_));
 sg13g2_buf_1 _20905_ (.A(net791),
    .X(_03428_));
 sg13g2_mux2_1 _20906_ (.A0(\cpu.ex.r_10[13] ),
    .A1(net658),
    .S(net526),
    .X(_00805_));
 sg13g2_buf_1 _20907_ (.A(net622),
    .X(_03429_));
 sg13g2_mux2_1 _20908_ (.A0(\cpu.ex.r_10[14] ),
    .A1(net525),
    .S(net526),
    .X(_00806_));
 sg13g2_buf_1 _20909_ (.A(net926),
    .X(_03430_));
 sg13g2_mux2_1 _20910_ (.A0(\cpu.ex.r_10[15] ),
    .A1(net743),
    .S(net526),
    .X(_00807_));
 sg13g2_buf_1 _20911_ (.A(net542),
    .X(_03431_));
 sg13g2_mux2_1 _20912_ (.A0(\cpu.ex.r_10[1] ),
    .A1(net476),
    .S(net526),
    .X(_00808_));
 sg13g2_buf_1 _20913_ (.A(_12557_),
    .X(_03432_));
 sg13g2_buf_1 _20914_ (.A(net475),
    .X(_03433_));
 sg13g2_mux2_1 _20915_ (.A0(\cpu.ex.r_10[2] ),
    .A1(net434),
    .S(net526),
    .X(_00809_));
 sg13g2_buf_1 _20916_ (.A(_12558_),
    .X(_03434_));
 sg13g2_mux2_1 _20917_ (.A0(\cpu.ex.r_10[3] ),
    .A1(net384),
    .S(_03426_),
    .X(_00810_));
 sg13g2_buf_2 _20918_ (.A(net610),
    .X(_03435_));
 sg13g2_buf_1 _20919_ (.A(net524),
    .X(_03436_));
 sg13g2_mux2_1 _20920_ (.A0(\cpu.ex.r_10[4] ),
    .A1(net474),
    .S(_03425_),
    .X(_00811_));
 sg13g2_mux2_1 _20921_ (.A0(\cpu.ex.r_10[5] ),
    .A1(net527),
    .S(_03425_),
    .X(_00812_));
 sg13g2_mux2_1 _20922_ (.A0(\cpu.ex.r_10[6] ),
    .A1(net748),
    .S(_03425_),
    .X(_00813_));
 sg13g2_mux2_1 _20923_ (.A0(\cpu.ex.r_10[7] ),
    .A1(net747),
    .S(_03425_),
    .X(_00814_));
 sg13g2_mux2_1 _20924_ (.A0(\cpu.ex.r_10[8] ),
    .A1(net746),
    .S(_03425_),
    .X(_00815_));
 sg13g2_mux2_1 _20925_ (.A0(\cpu.ex.r_10[9] ),
    .A1(net884),
    .S(_03425_),
    .X(_00816_));
 sg13g2_nor2_1 _20926_ (.A(_10351_),
    .B(_03423_),
    .Y(_03437_));
 sg13g2_buf_2 _20927_ (.A(_03437_),
    .X(_03438_));
 sg13g2_buf_1 _20928_ (.A(_03438_),
    .X(_03439_));
 sg13g2_mux2_1 _20929_ (.A0(\cpu.ex.r_11[0] ),
    .A1(net744),
    .S(net523),
    .X(_00817_));
 sg13g2_mux2_1 _20930_ (.A0(\cpu.ex.r_11[10] ),
    .A1(net881),
    .S(net523),
    .X(_00818_));
 sg13g2_mux2_1 _20931_ (.A0(\cpu.ex.r_11[11] ),
    .A1(_02977_),
    .S(_03439_),
    .X(_00819_));
 sg13g2_mux2_1 _20932_ (.A0(\cpu.ex.r_11[12] ),
    .A1(net601),
    .S(net523),
    .X(_00820_));
 sg13g2_mux2_1 _20933_ (.A0(\cpu.ex.r_11[13] ),
    .A1(net658),
    .S(net523),
    .X(_00821_));
 sg13g2_mux2_1 _20934_ (.A0(\cpu.ex.r_11[14] ),
    .A1(net525),
    .S(net523),
    .X(_00822_));
 sg13g2_mux2_1 _20935_ (.A0(\cpu.ex.r_11[15] ),
    .A1(net743),
    .S(net523),
    .X(_00823_));
 sg13g2_mux2_1 _20936_ (.A0(\cpu.ex.r_11[1] ),
    .A1(net476),
    .S(net523),
    .X(_00824_));
 sg13g2_mux2_1 _20937_ (.A0(\cpu.ex.r_11[2] ),
    .A1(net434),
    .S(_03439_),
    .X(_00825_));
 sg13g2_mux2_1 _20938_ (.A0(\cpu.ex.r_11[3] ),
    .A1(net384),
    .S(net523),
    .X(_00826_));
 sg13g2_mux2_1 _20939_ (.A0(\cpu.ex.r_11[4] ),
    .A1(net474),
    .S(_03438_),
    .X(_00827_));
 sg13g2_mux2_1 _20940_ (.A0(\cpu.ex.r_11[5] ),
    .A1(net527),
    .S(_03438_),
    .X(_00828_));
 sg13g2_mux2_1 _20941_ (.A0(\cpu.ex.r_11[6] ),
    .A1(net748),
    .S(_03438_),
    .X(_00829_));
 sg13g2_mux2_1 _20942_ (.A0(\cpu.ex.r_11[7] ),
    .A1(net747),
    .S(_03438_),
    .X(_00830_));
 sg13g2_mux2_1 _20943_ (.A0(\cpu.ex.r_11[8] ),
    .A1(net746),
    .S(_03438_),
    .X(_00831_));
 sg13g2_mux2_1 _20944_ (.A0(\cpu.ex.r_11[9] ),
    .A1(net884),
    .S(_03438_),
    .X(_00832_));
 sg13g2_nand3_1 _20945_ (.B(net1111),
    .C(net1115),
    .A(net1112),
    .Y(_03440_));
 sg13g2_buf_1 _20946_ (.A(_03440_),
    .X(_03441_));
 sg13g2_nor3_1 _20947_ (.A(net1114),
    .B(net1113),
    .C(_03441_),
    .Y(_03442_));
 sg13g2_buf_4 _20948_ (.X(_03443_),
    .A(_03442_));
 sg13g2_buf_1 _20949_ (.A(_03443_),
    .X(_03444_));
 sg13g2_mux2_1 _20950_ (.A0(\cpu.ex.r_12[0] ),
    .A1(_03419_),
    .S(_03444_),
    .X(_00833_));
 sg13g2_mux2_1 _20951_ (.A0(\cpu.ex.r_12[10] ),
    .A1(_02998_),
    .S(net600),
    .X(_00834_));
 sg13g2_mux2_1 _20952_ (.A0(\cpu.ex.r_12[11] ),
    .A1(net882),
    .S(net600),
    .X(_00835_));
 sg13g2_mux2_1 _20953_ (.A0(\cpu.ex.r_12[12] ),
    .A1(net601),
    .S(net600),
    .X(_00836_));
 sg13g2_mux2_1 _20954_ (.A0(\cpu.ex.r_12[13] ),
    .A1(net658),
    .S(net600),
    .X(_00837_));
 sg13g2_mux2_1 _20955_ (.A0(\cpu.ex.r_12[14] ),
    .A1(net525),
    .S(net600),
    .X(_00838_));
 sg13g2_nand2_1 _20956_ (.Y(_03445_),
    .A(net926),
    .B(_03443_));
 sg13g2_o21ai_1 _20957_ (.B1(_03445_),
    .Y(_00839_),
    .A1(_10403_),
    .A2(net600));
 sg13g2_mux2_1 _20958_ (.A0(\cpu.ex.r_12[1] ),
    .A1(net476),
    .S(net600),
    .X(_00840_));
 sg13g2_mux2_1 _20959_ (.A0(\cpu.ex.r_12[2] ),
    .A1(net434),
    .S(net600),
    .X(_00841_));
 sg13g2_mux2_1 _20960_ (.A0(\cpu.ex.r_12[3] ),
    .A1(net384),
    .S(_03444_),
    .X(_00842_));
 sg13g2_mux2_1 _20961_ (.A0(\cpu.ex.r_12[4] ),
    .A1(net474),
    .S(_03443_),
    .X(_00843_));
 sg13g2_mux2_1 _20962_ (.A0(\cpu.ex.r_12[5] ),
    .A1(net527),
    .S(_03443_),
    .X(_00844_));
 sg13g2_mux2_1 _20963_ (.A0(\cpu.ex.r_12[6] ),
    .A1(net748),
    .S(_03443_),
    .X(_00845_));
 sg13g2_mux2_1 _20964_ (.A0(\cpu.ex.r_12[7] ),
    .A1(_02996_),
    .S(_03443_),
    .X(_00846_));
 sg13g2_mux2_1 _20965_ (.A0(\cpu.ex.r_12[8] ),
    .A1(net746),
    .S(_03443_),
    .X(_00847_));
 sg13g2_buf_1 _20966_ (.A(_02973_),
    .X(_03446_));
 sg13g2_mux2_1 _20967_ (.A0(\cpu.ex.r_12[9] ),
    .A1(net879),
    .S(_03443_),
    .X(_00848_));
 sg13g2_nand2b_1 _20968_ (.Y(_03447_),
    .B(_10350_),
    .A_N(_10349_));
 sg13g2_buf_1 _20969_ (.A(_03447_),
    .X(_03448_));
 sg13g2_nor2_1 _20970_ (.A(_03441_),
    .B(_03448_),
    .Y(_03449_));
 sg13g2_buf_2 _20971_ (.A(_03449_),
    .X(_03450_));
 sg13g2_buf_1 _20972_ (.A(_03450_),
    .X(_03451_));
 sg13g2_mux2_1 _20973_ (.A0(\cpu.ex.r_13[0] ),
    .A1(net744),
    .S(net599),
    .X(_00849_));
 sg13g2_mux2_1 _20974_ (.A0(\cpu.ex.r_13[10] ),
    .A1(net881),
    .S(net599),
    .X(_00850_));
 sg13g2_mux2_1 _20975_ (.A0(\cpu.ex.r_13[11] ),
    .A1(_02977_),
    .S(net599),
    .X(_00851_));
 sg13g2_mux2_1 _20976_ (.A0(\cpu.ex.r_13[12] ),
    .A1(net601),
    .S(net599),
    .X(_00852_));
 sg13g2_mux2_1 _20977_ (.A0(\cpu.ex.r_13[13] ),
    .A1(net658),
    .S(net599),
    .X(_00853_));
 sg13g2_mux2_1 _20978_ (.A0(\cpu.ex.r_13[14] ),
    .A1(net525),
    .S(net599),
    .X(_00854_));
 sg13g2_mux2_1 _20979_ (.A0(\cpu.ex.r_13[15] ),
    .A1(net743),
    .S(_03451_),
    .X(_00855_));
 sg13g2_mux2_1 _20980_ (.A0(\cpu.ex.r_13[1] ),
    .A1(net476),
    .S(net599),
    .X(_00856_));
 sg13g2_mux2_1 _20981_ (.A0(\cpu.ex.r_13[2] ),
    .A1(net434),
    .S(_03451_),
    .X(_00857_));
 sg13g2_mux2_1 _20982_ (.A0(\cpu.ex.r_13[3] ),
    .A1(net384),
    .S(net599),
    .X(_00858_));
 sg13g2_mux2_1 _20983_ (.A0(\cpu.ex.r_13[4] ),
    .A1(net474),
    .S(_03450_),
    .X(_00859_));
 sg13g2_mux2_1 _20984_ (.A0(\cpu.ex.r_13[5] ),
    .A1(net527),
    .S(_03450_),
    .X(_00860_));
 sg13g2_mux2_1 _20985_ (.A0(\cpu.ex.r_13[6] ),
    .A1(net748),
    .S(_03450_),
    .X(_00861_));
 sg13g2_mux2_1 _20986_ (.A0(\cpu.ex.r_13[7] ),
    .A1(net747),
    .S(_03450_),
    .X(_00862_));
 sg13g2_mux2_1 _20987_ (.A0(\cpu.ex.r_13[8] ),
    .A1(_02997_),
    .S(_03450_),
    .X(_00863_));
 sg13g2_mux2_1 _20988_ (.A0(\cpu.ex.r_13[9] ),
    .A1(net879),
    .S(_03450_),
    .X(_00864_));
 sg13g2_nor2_1 _20989_ (.A(_03421_),
    .B(_03441_),
    .Y(_03452_));
 sg13g2_buf_4 _20990_ (.X(_03453_),
    .A(_03452_));
 sg13g2_buf_1 _20991_ (.A(_03453_),
    .X(_03454_));
 sg13g2_mux2_1 _20992_ (.A0(\cpu.ex.r_14[0] ),
    .A1(net744),
    .S(net598),
    .X(_00865_));
 sg13g2_mux2_1 _20993_ (.A0(\cpu.ex.r_14[10] ),
    .A1(net881),
    .S(net598),
    .X(_00866_));
 sg13g2_buf_1 _20994_ (.A(net981),
    .X(_03455_));
 sg13g2_mux2_1 _20995_ (.A0(\cpu.ex.r_14[11] ),
    .A1(net878),
    .S(net598),
    .X(_00867_));
 sg13g2_mux2_1 _20996_ (.A0(\cpu.ex.r_14[12] ),
    .A1(net601),
    .S(net598),
    .X(_00868_));
 sg13g2_mux2_1 _20997_ (.A0(\cpu.ex.r_14[13] ),
    .A1(net658),
    .S(net598),
    .X(_00869_));
 sg13g2_mux2_1 _20998_ (.A0(\cpu.ex.r_14[14] ),
    .A1(net525),
    .S(net598),
    .X(_00870_));
 sg13g2_mux2_1 _20999_ (.A0(\cpu.ex.r_14[15] ),
    .A1(net743),
    .S(net598),
    .X(_00871_));
 sg13g2_nand2_1 _21000_ (.Y(_03456_),
    .A(net476),
    .B(_03453_));
 sg13g2_o21ai_1 _21001_ (.B1(_03456_),
    .Y(_00872_),
    .A1(_10775_),
    .A2(_03454_));
 sg13g2_mux2_1 _21002_ (.A0(\cpu.ex.r_14[2] ),
    .A1(net434),
    .S(_03454_),
    .X(_00873_));
 sg13g2_mux2_1 _21003_ (.A0(\cpu.ex.r_14[3] ),
    .A1(net384),
    .S(net598),
    .X(_00874_));
 sg13g2_mux2_1 _21004_ (.A0(\cpu.ex.r_14[4] ),
    .A1(net474),
    .S(_03453_),
    .X(_00875_));
 sg13g2_mux2_1 _21005_ (.A0(\cpu.ex.r_14[5] ),
    .A1(_02967_),
    .S(_03453_),
    .X(_00876_));
 sg13g2_mux2_1 _21006_ (.A0(\cpu.ex.r_14[6] ),
    .A1(net748),
    .S(_03453_),
    .X(_00877_));
 sg13g2_mux2_1 _21007_ (.A0(\cpu.ex.r_14[7] ),
    .A1(net747),
    .S(_03453_),
    .X(_00878_));
 sg13g2_mux2_1 _21008_ (.A0(\cpu.ex.r_14[8] ),
    .A1(net746),
    .S(_03453_),
    .X(_00879_));
 sg13g2_mux2_1 _21009_ (.A0(\cpu.ex.r_14[9] ),
    .A1(net879),
    .S(_03453_),
    .X(_00880_));
 sg13g2_nor2_1 _21010_ (.A(_10351_),
    .B(_03441_),
    .Y(_03457_));
 sg13g2_buf_2 _21011_ (.A(_03457_),
    .X(_03458_));
 sg13g2_buf_1 _21012_ (.A(_03458_),
    .X(_03459_));
 sg13g2_mux2_1 _21013_ (.A0(\cpu.ex.r_15[0] ),
    .A1(net744),
    .S(net597),
    .X(_00881_));
 sg13g2_mux2_1 _21014_ (.A0(\cpu.ex.r_15[10] ),
    .A1(net881),
    .S(net597),
    .X(_00882_));
 sg13g2_mux2_1 _21015_ (.A0(\cpu.ex.r_15[11] ),
    .A1(net878),
    .S(_03459_),
    .X(_00883_));
 sg13g2_mux2_1 _21016_ (.A0(\cpu.ex.r_15[12] ),
    .A1(_03427_),
    .S(net597),
    .X(_00884_));
 sg13g2_mux2_1 _21017_ (.A0(\cpu.ex.r_15[13] ),
    .A1(net658),
    .S(net597),
    .X(_00885_));
 sg13g2_mux2_1 _21018_ (.A0(\cpu.ex.r_15[14] ),
    .A1(net525),
    .S(net597),
    .X(_00886_));
 sg13g2_mux2_1 _21019_ (.A0(\cpu.ex.r_15[15] ),
    .A1(net743),
    .S(net597),
    .X(_00887_));
 sg13g2_mux2_1 _21020_ (.A0(\cpu.ex.r_15[1] ),
    .A1(net476),
    .S(net597),
    .X(_00888_));
 sg13g2_mux2_1 _21021_ (.A0(\cpu.ex.r_15[2] ),
    .A1(_03433_),
    .S(_03459_),
    .X(_00889_));
 sg13g2_mux2_1 _21022_ (.A0(\cpu.ex.r_15[3] ),
    .A1(net384),
    .S(net597),
    .X(_00890_));
 sg13g2_mux2_1 _21023_ (.A0(\cpu.ex.r_15[4] ),
    .A1(net474),
    .S(_03458_),
    .X(_00891_));
 sg13g2_mux2_1 _21024_ (.A0(\cpu.ex.r_15[5] ),
    .A1(_02967_),
    .S(_03458_),
    .X(_00892_));
 sg13g2_mux2_1 _21025_ (.A0(\cpu.ex.r_15[6] ),
    .A1(_02995_),
    .S(_03458_),
    .X(_00893_));
 sg13g2_mux2_1 _21026_ (.A0(\cpu.ex.r_15[7] ),
    .A1(_02996_),
    .S(_03458_),
    .X(_00894_));
 sg13g2_mux2_1 _21027_ (.A0(\cpu.ex.r_15[8] ),
    .A1(_02997_),
    .S(_03458_),
    .X(_00895_));
 sg13g2_mux2_1 _21028_ (.A0(\cpu.ex.r_15[9] ),
    .A1(net879),
    .S(_03458_),
    .X(_00896_));
 sg13g2_nor3_1 _21029_ (.A(net1114),
    .B(net1113),
    .C(_03423_),
    .Y(_03460_));
 sg13g2_buf_1 _21030_ (.A(_03460_),
    .X(_03461_));
 sg13g2_buf_1 _21031_ (.A(net596),
    .X(_03462_));
 sg13g2_mux2_1 _21032_ (.A0(\cpu.ex.r_8[0] ),
    .A1(net744),
    .S(net522),
    .X(_00897_));
 sg13g2_mux2_1 _21033_ (.A0(\cpu.ex.r_8[10] ),
    .A1(_02998_),
    .S(net522),
    .X(_00898_));
 sg13g2_mux2_1 _21034_ (.A0(\cpu.ex.r_8[11] ),
    .A1(net878),
    .S(net522),
    .X(_00899_));
 sg13g2_mux2_1 _21035_ (.A0(\cpu.ex.r_8[12] ),
    .A1(net601),
    .S(net522),
    .X(_00900_));
 sg13g2_mux2_1 _21036_ (.A0(\cpu.ex.r_8[13] ),
    .A1(net658),
    .S(net522),
    .X(_00901_));
 sg13g2_mux2_1 _21037_ (.A0(\cpu.ex.r_8[14] ),
    .A1(net525),
    .S(net522),
    .X(_00902_));
 sg13g2_mux2_1 _21038_ (.A0(\cpu.ex.r_8[15] ),
    .A1(net743),
    .S(net522),
    .X(_00903_));
 sg13g2_mux2_1 _21039_ (.A0(\cpu.ex.r_8[1] ),
    .A1(net476),
    .S(_03462_),
    .X(_00904_));
 sg13g2_mux2_1 _21040_ (.A0(\cpu.ex.r_8[2] ),
    .A1(net434),
    .S(net596),
    .X(_00905_));
 sg13g2_mux2_1 _21041_ (.A0(\cpu.ex.r_8[3] ),
    .A1(net384),
    .S(net596),
    .X(_00906_));
 sg13g2_buf_1 _21042_ (.A(net524),
    .X(_03463_));
 sg13g2_nand2_1 _21043_ (.Y(_03464_),
    .A(_03463_),
    .B(_03461_));
 sg13g2_o21ai_1 _21044_ (.B1(_03464_),
    .Y(_00907_),
    .A1(_10889_),
    .A2(net522));
 sg13g2_buf_1 _21045_ (.A(net602),
    .X(_03465_));
 sg13g2_mux2_1 _21046_ (.A0(\cpu.ex.r_8[5] ),
    .A1(net521),
    .S(net596),
    .X(_00908_));
 sg13g2_inv_1 _21047_ (.Y(_03466_),
    .A(\cpu.ex.r_8[6] ));
 sg13g2_nand2_1 _21048_ (.Y(_03467_),
    .A(net889),
    .B(net596));
 sg13g2_o21ai_1 _21049_ (.B1(_03467_),
    .Y(_00909_),
    .A1(_03466_),
    .A2(_03462_));
 sg13g2_mux2_1 _21050_ (.A0(\cpu.ex.r_8[7] ),
    .A1(net747),
    .S(net596),
    .X(_00910_));
 sg13g2_mux2_1 _21051_ (.A0(\cpu.ex.r_8[8] ),
    .A1(net746),
    .S(net596),
    .X(_00911_));
 sg13g2_mux2_1 _21052_ (.A0(\cpu.ex.r_8[9] ),
    .A1(net879),
    .S(net596),
    .X(_00912_));
 sg13g2_nor2_1 _21053_ (.A(_03423_),
    .B(_03448_),
    .Y(_03468_));
 sg13g2_buf_4 _21054_ (.X(_03469_),
    .A(_03468_));
 sg13g2_buf_1 _21055_ (.A(_03469_),
    .X(_03470_));
 sg13g2_mux2_1 _21056_ (.A0(\cpu.ex.r_9[0] ),
    .A1(net744),
    .S(net520),
    .X(_00913_));
 sg13g2_mux2_1 _21057_ (.A0(\cpu.ex.r_9[10] ),
    .A1(net881),
    .S(net520),
    .X(_00914_));
 sg13g2_mux2_1 _21058_ (.A0(\cpu.ex.r_9[11] ),
    .A1(net878),
    .S(net520),
    .X(_00915_));
 sg13g2_mux2_1 _21059_ (.A0(\cpu.ex.r_9[12] ),
    .A1(net601),
    .S(net520),
    .X(_00916_));
 sg13g2_mux2_1 _21060_ (.A0(\cpu.ex.r_9[13] ),
    .A1(net658),
    .S(net520),
    .X(_00917_));
 sg13g2_mux2_1 _21061_ (.A0(\cpu.ex.r_9[14] ),
    .A1(_03429_),
    .S(net520),
    .X(_00918_));
 sg13g2_mux2_1 _21062_ (.A0(\cpu.ex.r_9[15] ),
    .A1(net743),
    .S(net520),
    .X(_00919_));
 sg13g2_mux2_1 _21063_ (.A0(\cpu.ex.r_9[1] ),
    .A1(net476),
    .S(_03470_),
    .X(_00920_));
 sg13g2_mux2_1 _21064_ (.A0(\cpu.ex.r_9[2] ),
    .A1(_03433_),
    .S(net520),
    .X(_00921_));
 sg13g2_mux2_1 _21065_ (.A0(\cpu.ex.r_9[3] ),
    .A1(net384),
    .S(_03469_),
    .X(_00922_));
 sg13g2_nand2_1 _21066_ (.Y(_03471_),
    .A(net524),
    .B(_03469_));
 sg13g2_o21ai_1 _21067_ (.B1(_03471_),
    .Y(_00923_),
    .A1(_10880_),
    .A2(_03470_));
 sg13g2_mux2_1 _21068_ (.A0(\cpu.ex.r_9[5] ),
    .A1(net521),
    .S(_03469_),
    .X(_00924_));
 sg13g2_mux2_1 _21069_ (.A0(\cpu.ex.r_9[6] ),
    .A1(net748),
    .S(_03469_),
    .X(_00925_));
 sg13g2_mux2_1 _21070_ (.A0(\cpu.ex.r_9[7] ),
    .A1(net747),
    .S(_03469_),
    .X(_00926_));
 sg13g2_mux2_1 _21071_ (.A0(\cpu.ex.r_9[8] ),
    .A1(net746),
    .S(_03469_),
    .X(_00927_));
 sg13g2_mux2_1 _21072_ (.A0(\cpu.ex.r_9[9] ),
    .A1(net879),
    .S(_03469_),
    .X(_00928_));
 sg13g2_buf_1 _21073_ (.A(_11194_),
    .X(_03472_));
 sg13g2_buf_1 _21074_ (.A(net196),
    .X(_03473_));
 sg13g2_buf_1 _21075_ (.A(_11267_),
    .X(_03474_));
 sg13g2_nor2_1 _21076_ (.A(_00195_),
    .B(net221),
    .Y(_03475_));
 sg13g2_nand2b_1 _21077_ (.Y(_03476_),
    .B(net221),
    .A_N(_11121_));
 sg13g2_nand2b_1 _21078_ (.Y(_03477_),
    .B(_03476_),
    .A_N(_03475_));
 sg13g2_buf_1 _21079_ (.A(_03477_),
    .X(_03478_));
 sg13g2_buf_1 _21080_ (.A(_03478_),
    .X(_03479_));
 sg13g2_nand2_1 _21081_ (.Y(_03480_),
    .A(net146),
    .B(net131));
 sg13g2_a21oi_1 _21082_ (.A1(_08404_),
    .A2(_11150_),
    .Y(_03481_),
    .B1(_11236_));
 sg13g2_nor2_1 _21083_ (.A(_00196_),
    .B(net221),
    .Y(_03482_));
 sg13g2_a21o_1 _21084_ (.A2(_03481_),
    .A1(net221),
    .B1(_03482_),
    .X(_03483_));
 sg13g2_buf_1 _21085_ (.A(_03483_),
    .X(_03484_));
 sg13g2_buf_1 _21086_ (.A(_03484_),
    .X(_03485_));
 sg13g2_nor2_1 _21087_ (.A(net169),
    .B(net130),
    .Y(_03486_));
 sg13g2_buf_1 _21088_ (.A(net176),
    .X(_03487_));
 sg13g2_nor2_1 _21089_ (.A(_00289_),
    .B(net221),
    .Y(_03488_));
 sg13g2_nand2b_1 _21090_ (.Y(_03489_),
    .B(net221),
    .A_N(_11263_));
 sg13g2_nand2b_1 _21091_ (.Y(_03490_),
    .B(_03489_),
    .A_N(_03488_));
 sg13g2_buf_1 _21092_ (.A(_03490_),
    .X(_03491_));
 sg13g2_buf_1 _21093_ (.A(net142),
    .X(_03492_));
 sg13g2_nor2_1 _21094_ (.A(net143),
    .B(net129),
    .Y(_03493_));
 sg13g2_nor2_1 _21095_ (.A(_03486_),
    .B(_03493_),
    .Y(_03494_));
 sg13g2_a21oi_1 _21096_ (.A1(_10474_),
    .A2(_10800_),
    .Y(_03495_),
    .B1(_10801_));
 sg13g2_buf_2 _21097_ (.A(_03495_),
    .X(_03496_));
 sg13g2_or4_1 _21098_ (.A(_08388_),
    .B(_11137_),
    .C(_08434_),
    .D(net505),
    .X(_03497_));
 sg13g2_nand2_1 _21099_ (.Y(_03498_),
    .A(_11536_),
    .B(_11537_));
 sg13g2_o21ai_1 _21100_ (.B1(_11535_),
    .Y(_03499_),
    .A1(_08431_),
    .A2(_03498_));
 sg13g2_and4_1 _21101_ (.A(_10983_),
    .B(_03496_),
    .C(_03497_),
    .D(_03499_),
    .X(_03500_));
 sg13g2_nand3_1 _21102_ (.B(_11557_),
    .C(_11523_),
    .A(net275),
    .Y(_03501_));
 sg13g2_o21ai_1 _21103_ (.B1(_03501_),
    .Y(_03502_),
    .A1(_11528_),
    .A2(_03500_));
 sg13g2_buf_1 _21104_ (.A(_03496_),
    .X(_03503_));
 sg13g2_a21oi_1 _21105_ (.A1(_10983_),
    .A2(_11559_),
    .Y(_03504_),
    .B1(net220));
 sg13g2_and4_1 _21106_ (.A(_11360_),
    .B(_11361_),
    .C(_11379_),
    .D(_11380_),
    .X(_03505_));
 sg13g2_buf_2 _21107_ (.A(_03505_),
    .X(_03506_));
 sg13g2_buf_1 _21108_ (.A(_03506_),
    .X(_03507_));
 sg13g2_mux2_1 _21109_ (.A0(_00297_),
    .A1(_11481_),
    .S(_11192_),
    .X(_03508_));
 sg13g2_buf_2 _21110_ (.A(_03508_),
    .X(_03509_));
 sg13g2_buf_8 _21111_ (.A(_03509_),
    .X(_03510_));
 sg13g2_nor3_1 _21112_ (.A(_10936_),
    .B(_10941_),
    .C(_11502_),
    .Y(_03511_));
 sg13g2_inv_1 _21113_ (.Y(_03512_),
    .A(_00191_));
 sg13g2_nor3_1 _21114_ (.A(_03512_),
    .B(_10936_),
    .C(_10941_),
    .Y(_03513_));
 sg13g2_mux2_1 _21115_ (.A0(_03511_),
    .A1(_03513_),
    .S(_11141_),
    .X(_03514_));
 sg13g2_a221oi_1 _21116_ (.B2(_10959_),
    .C1(_03514_),
    .B1(net195),
    .A1(_11652_),
    .Y(_03515_),
    .A2(net219));
 sg13g2_o21ai_1 _21117_ (.B1(_03515_),
    .Y(_03516_),
    .A1(_03502_),
    .A2(_03504_));
 sg13g2_nand2_1 _21118_ (.Y(_03517_),
    .A(net277),
    .B(net235));
 sg13g2_inv_1 _21119_ (.Y(_03518_),
    .A(_11502_));
 sg13g2_mux2_1 _21120_ (.A0(_00191_),
    .A1(_03518_),
    .S(_11191_),
    .X(_03519_));
 sg13g2_buf_1 _21121_ (.A(_03519_),
    .X(_03520_));
 sg13g2_o21ai_1 _21122_ (.B1(net219),
    .Y(_03521_),
    .A1(_03517_),
    .A2(net266));
 sg13g2_o21ai_1 _21123_ (.B1(_11653_),
    .Y(_03522_),
    .A1(_10943_),
    .A2(net266));
 sg13g2_nor2_1 _21124_ (.A(net272),
    .B(_03514_),
    .Y(_03523_));
 sg13g2_a21oi_1 _21125_ (.A1(_11652_),
    .A2(net219),
    .Y(_03524_),
    .B1(net195));
 sg13g2_a22oi_1 _21126_ (.Y(_03525_),
    .B1(_03523_),
    .B2(_03524_),
    .A2(_03522_),
    .A1(_03521_));
 sg13g2_nand2b_1 _21127_ (.Y(_03526_),
    .B(_11426_),
    .A_N(_11408_));
 sg13g2_mux2_1 _21128_ (.A0(_00295_),
    .A1(_03526_),
    .S(net347),
    .X(_03527_));
 sg13g2_buf_2 _21129_ (.A(_03527_),
    .X(_03528_));
 sg13g2_buf_8 _21130_ (.A(_03528_),
    .X(_03529_));
 sg13g2_nor2_1 _21131_ (.A(net202),
    .B(net194),
    .Y(_03530_));
 sg13g2_a22oi_1 _21132_ (.Y(_03531_),
    .B1(_11402_),
    .B2(_11526_),
    .A2(_11398_),
    .A1(net347));
 sg13g2_buf_2 _21133_ (.A(_03531_),
    .X(_03532_));
 sg13g2_nor2_1 _21134_ (.A(_11645_),
    .B(_03532_),
    .Y(_03533_));
 sg13g2_nor3_1 _21135_ (.A(net276),
    .B(_03530_),
    .C(_03533_),
    .Y(_03534_));
 sg13g2_and3_1 _21136_ (.X(_03535_),
    .A(_03516_),
    .B(_03525_),
    .C(_03534_));
 sg13g2_nand2_1 _21137_ (.Y(_03536_),
    .A(net202),
    .B(net194));
 sg13g2_buf_1 _21138_ (.A(_11406_),
    .X(_03537_));
 sg13g2_nor2_1 _21139_ (.A(net236),
    .B(net193),
    .Y(_03538_));
 sg13g2_nand2b_1 _21140_ (.Y(_03539_),
    .B(_03538_),
    .A_N(_03530_));
 sg13g2_a21oi_1 _21141_ (.A1(_03536_),
    .A2(_03539_),
    .Y(_03540_),
    .B1(net276));
 sg13g2_mux2_1 _21142_ (.A0(_11317_),
    .A1(_11333_),
    .S(net275),
    .X(_03541_));
 sg13g2_buf_2 _21143_ (.A(_03541_),
    .X(_03542_));
 sg13g2_nor2_1 _21144_ (.A(_10757_),
    .B(_03542_),
    .Y(_03543_));
 sg13g2_inv_1 _21145_ (.Y(_03544_),
    .A(_03543_));
 sg13g2_o21ai_1 _21146_ (.B1(_03544_),
    .Y(_03545_),
    .A1(_03535_),
    .A2(_03540_));
 sg13g2_nand3b_1 _21147_ (.B(_11038_),
    .C(_03536_),
    .Y(_03546_),
    .A_N(_03538_));
 sg13g2_a21oi_1 _21148_ (.A1(_03516_),
    .A2(_03525_),
    .Y(_03547_),
    .B1(_03546_));
 sg13g2_a21oi_1 _21149_ (.A1(_03536_),
    .A2(_03533_),
    .Y(_03548_),
    .B1(_03530_));
 sg13g2_nor2_1 _21150_ (.A(net273),
    .B(_03548_),
    .Y(_03549_));
 sg13g2_or4_1 _21151_ (.A(_11454_),
    .B(_03547_),
    .C(_03549_),
    .D(_03543_),
    .X(_03550_));
 sg13g2_buf_1 _21152_ (.A(_03550_),
    .X(_03551_));
 sg13g2_inv_1 _21153_ (.Y(_03552_),
    .A(_11311_));
 sg13g2_mux2_1 _21154_ (.A0(_00291_),
    .A1(_03552_),
    .S(net275),
    .X(_03553_));
 sg13g2_buf_1 _21155_ (.A(_03553_),
    .X(_03554_));
 sg13g2_a22oi_1 _21156_ (.Y(_03555_),
    .B1(_03542_),
    .B2(_11806_),
    .A2(_03554_),
    .A1(net200));
 sg13g2_and2_1 _21157_ (.A(net172),
    .B(_03555_),
    .X(_03556_));
 sg13g2_nand3_1 _21158_ (.B(_03551_),
    .C(_03556_),
    .A(_03545_),
    .Y(_03557_));
 sg13g2_buf_1 _21159_ (.A(_03554_),
    .X(_03558_));
 sg13g2_inv_1 _21160_ (.Y(_03559_),
    .A(_11352_));
 sg13g2_nor2_1 _21161_ (.A(_11316_),
    .B(net275),
    .Y(_03560_));
 sg13g2_a21o_1 _21162_ (.A2(_03559_),
    .A1(_11267_),
    .B1(_03560_),
    .X(_03561_));
 sg13g2_buf_1 _21163_ (.A(_03561_),
    .X(_03562_));
 sg13g2_nand2_1 _21164_ (.Y(_03563_),
    .A(net172),
    .B(_03562_));
 sg13g2_a21oi_1 _21165_ (.A1(net200),
    .A2(net163),
    .Y(_03564_),
    .B1(_03563_));
 sg13g2_a21oi_1 _21166_ (.A1(net174),
    .A2(_11313_),
    .Y(_03565_),
    .B1(_03564_));
 sg13g2_buf_1 _21167_ (.A(_03562_),
    .X(_03566_));
 sg13g2_nand4_1 _21168_ (.B(_03545_),
    .C(_03551_),
    .A(net141),
    .Y(_03567_),
    .D(_03555_));
 sg13g2_nand3_1 _21169_ (.B(_03565_),
    .C(_03567_),
    .A(_03557_),
    .Y(_03568_));
 sg13g2_buf_1 _21170_ (.A(net233),
    .X(_03569_));
 sg13g2_nand2b_1 _21171_ (.Y(_03570_),
    .B(net170),
    .A_N(net192));
 sg13g2_and2_1 _21172_ (.A(net147),
    .B(net192),
    .X(_03571_));
 sg13g2_a21o_1 _21173_ (.A2(_03570_),
    .A1(_03568_),
    .B1(_03571_),
    .X(_03572_));
 sg13g2_buf_2 _21174_ (.A(_03572_),
    .X(_03573_));
 sg13g2_a22oi_1 _21175_ (.Y(_03574_),
    .B1(net129),
    .B2(net143),
    .A2(net130),
    .A1(net169));
 sg13g2_nor2_1 _21176_ (.A(_03486_),
    .B(_03574_),
    .Y(_03575_));
 sg13g2_a21oi_1 _21177_ (.A1(_03494_),
    .A2(_03573_),
    .Y(_03576_),
    .B1(_03575_));
 sg13g2_nand2_1 _21178_ (.Y(_03577_),
    .A(_03480_),
    .B(_03576_));
 sg13g2_nor2b_1 _21179_ (.A(_03475_),
    .B_N(_03476_),
    .Y(_03578_));
 sg13g2_buf_2 _21180_ (.A(_03578_),
    .X(_03579_));
 sg13g2_nand2_1 _21181_ (.Y(_03580_),
    .A(_11954_),
    .B(_03579_));
 sg13g2_a22oi_1 _21182_ (.Y(_03581_),
    .B1(_03577_),
    .B2(_03580_),
    .A2(net164),
    .A1(net132));
 sg13g2_nor2_1 _21183_ (.A(_11634_),
    .B(net164),
    .Y(_03582_));
 sg13g2_a21oi_2 _21184_ (.B1(_11688_),
    .Y(_03583_),
    .A2(_11694_),
    .A1(net1053));
 sg13g2_nor2_1 _21185_ (.A(_09121_),
    .B(_03583_),
    .Y(_03584_));
 sg13g2_o21ai_1 _21186_ (.B1(_03584_),
    .Y(_03585_),
    .A1(_03581_),
    .A2(_03582_));
 sg13g2_buf_1 _21187_ (.A(net1059),
    .X(_03586_));
 sg13g2_nor2_1 _21188_ (.A(_10461_),
    .B(_11194_),
    .Y(_03587_));
 sg13g2_nor3_1 _21189_ (.A(net877),
    .B(_03583_),
    .C(_03587_),
    .Y(_03588_));
 sg13g2_nand2_2 _21190_ (.Y(_03589_),
    .A(net146),
    .B(_03579_));
 sg13g2_a21oi_1 _21191_ (.A1(net221),
    .A2(_03481_),
    .Y(_03590_),
    .B1(_03482_));
 sg13g2_buf_1 _21192_ (.A(_03590_),
    .X(_03591_));
 sg13g2_buf_1 _21193_ (.A(_03591_),
    .X(_03592_));
 sg13g2_nand2b_1 _21194_ (.Y(_03593_),
    .B(_11451_),
    .A_N(_11431_));
 sg13g2_mux2_1 _21195_ (.A0(_00294_),
    .A1(_03593_),
    .S(net347),
    .X(_03594_));
 sg13g2_buf_1 _21196_ (.A(_03594_),
    .X(_03595_));
 sg13g2_nand2_2 _21197_ (.Y(_03596_),
    .A(net276),
    .B(net218));
 sg13g2_nand2_1 _21198_ (.Y(_03597_),
    .A(_10757_),
    .B(_03596_));
 sg13g2_nand2_1 _21199_ (.Y(_03598_),
    .A(_11587_),
    .B(_11454_));
 sg13g2_and2_1 _21200_ (.A(_03542_),
    .B(_03598_),
    .X(_03599_));
 sg13g2_nor3_1 _21201_ (.A(_11652_),
    .B(net274),
    .C(_11406_),
    .Y(_03600_));
 sg13g2_o21ai_1 _21202_ (.B1(net193),
    .Y(_03601_),
    .A1(_11652_),
    .A2(net274));
 sg13g2_o21ai_1 _21203_ (.B1(_03601_),
    .Y(_03602_),
    .A1(net236),
    .A2(_03600_));
 sg13g2_a21oi_1 _21204_ (.A1(_11429_),
    .A2(_03602_),
    .Y(_03603_),
    .B1(_11584_));
 sg13g2_a22oi_1 _21205_ (.Y(_03604_),
    .B1(_03599_),
    .B2(_03603_),
    .A2(_03597_),
    .A1(_03542_));
 sg13g2_buf_1 _21206_ (.A(_03604_),
    .X(_03605_));
 sg13g2_nand2_2 _21207_ (.Y(_03606_),
    .A(net236),
    .B(_03532_));
 sg13g2_inv_1 _21208_ (.Y(_03607_),
    .A(_03606_));
 sg13g2_nor2_2 _21209_ (.A(_10983_),
    .B(_03496_),
    .Y(_03608_));
 sg13g2_a221oi_1 _21210_ (.B2(net347),
    .C1(_03496_),
    .B1(_11557_),
    .A1(_11535_),
    .Y(_03609_),
    .A2(net398));
 sg13g2_nor3_1 _21211_ (.A(_03608_),
    .B(_11528_),
    .C(_03609_),
    .Y(_03610_));
 sg13g2_nand2_1 _21212_ (.Y(_03611_),
    .A(_10983_),
    .B(_03496_));
 sg13g2_buf_8 _21213_ (.A(_03611_),
    .X(_03612_));
 sg13g2_nand4_1 _21214_ (.B(_10836_),
    .C(_11457_),
    .A(_10807_),
    .Y(_03613_),
    .D(_11480_));
 sg13g2_nand3b_1 _21215_ (.B(_10807_),
    .C(_10836_),
    .Y(_03614_),
    .A_N(_00297_));
 sg13g2_mux2_1 _21216_ (.A0(_03613_),
    .A1(_03614_),
    .S(_11141_),
    .X(_03615_));
 sg13g2_buf_2 _21217_ (.A(_03615_),
    .X(_03616_));
 sg13g2_o21ai_1 _21218_ (.B1(_03616_),
    .Y(_03617_),
    .A1(_11559_),
    .A2(_03612_));
 sg13g2_a22oi_1 _21219_ (.Y(_03618_),
    .B1(_03509_),
    .B2(_10838_),
    .A2(net266),
    .A1(net277));
 sg13g2_o21ai_1 _21220_ (.B1(_03618_),
    .Y(_03619_),
    .A1(_03610_),
    .A2(_03617_));
 sg13g2_buf_1 _21221_ (.A(_03619_),
    .X(_03620_));
 sg13g2_nand3_1 _21222_ (.B(net274),
    .C(_11406_),
    .A(_11652_),
    .Y(_03621_));
 sg13g2_nand2_2 _21223_ (.Y(_03622_),
    .A(_11645_),
    .B(_11406_));
 sg13g2_nand3_1 _21224_ (.B(_11652_),
    .C(net274),
    .A(_11645_),
    .Y(_03623_));
 sg13g2_nand3_1 _21225_ (.B(_10940_),
    .C(_11502_),
    .A(_10946_),
    .Y(_03624_));
 sg13g2_nand3_1 _21226_ (.B(_10946_),
    .C(_10940_),
    .A(_03512_),
    .Y(_03625_));
 sg13g2_mux2_1 _21227_ (.A0(_03624_),
    .A1(_03625_),
    .S(_11141_),
    .X(_03626_));
 sg13g2_buf_2 _21228_ (.A(_03626_),
    .X(_03627_));
 sg13g2_and2_1 _21229_ (.A(_11010_),
    .B(_03627_),
    .X(_03628_));
 sg13g2_and4_1 _21230_ (.A(_03621_),
    .B(_03622_),
    .C(_03623_),
    .D(_03628_),
    .X(_03629_));
 sg13g2_nand2_1 _21231_ (.Y(_03630_),
    .A(net235),
    .B(_03627_));
 sg13g2_o21ai_1 _21232_ (.B1(_03506_),
    .Y(_03631_),
    .A1(net235),
    .A2(_03627_));
 sg13g2_a221oi_1 _21233_ (.B2(_03631_),
    .C1(_11429_),
    .B1(_03630_),
    .A1(_11645_),
    .Y(_03632_),
    .A2(net193));
 sg13g2_a221oi_1 _21234_ (.B2(_03629_),
    .C1(_03632_),
    .B1(_03620_),
    .A1(_03528_),
    .Y(_03633_),
    .A2(_03607_));
 sg13g2_nand2_2 _21235_ (.Y(_03634_),
    .A(net235),
    .B(_03506_));
 sg13g2_nand2_1 _21236_ (.Y(_03635_),
    .A(_03634_),
    .B(_03606_));
 sg13g2_o21ai_1 _21237_ (.B1(_03599_),
    .Y(_03636_),
    .A1(_03620_),
    .A2(_03635_));
 sg13g2_or2_1 _21238_ (.X(_03637_),
    .B(_03636_),
    .A(_03633_));
 sg13g2_buf_8 _21239_ (.A(_03637_),
    .X(_03638_));
 sg13g2_and3_1 _21240_ (.X(_03639_),
    .A(_03621_),
    .B(_03622_),
    .C(_03623_));
 sg13g2_nand2_1 _21241_ (.Y(_03640_),
    .A(_11583_),
    .B(_11429_));
 sg13g2_and2_1 _21242_ (.A(_03598_),
    .B(_03640_),
    .X(_03641_));
 sg13g2_nor2_1 _21243_ (.A(_11038_),
    .B(net218),
    .Y(_03642_));
 sg13g2_nand2_1 _21244_ (.Y(_03643_),
    .A(_11011_),
    .B(_03528_));
 sg13g2_o21ai_1 _21245_ (.B1(_03596_),
    .Y(_03644_),
    .A1(_03642_),
    .A2(_03643_));
 sg13g2_a21oi_1 _21246_ (.A1(_03639_),
    .A2(_03641_),
    .Y(_03645_),
    .B1(_03644_));
 sg13g2_nand4_1 _21247_ (.B(_03596_),
    .C(_03606_),
    .A(_03634_),
    .Y(_03646_),
    .D(_03643_));
 sg13g2_a21oi_1 _21248_ (.A1(_03627_),
    .A2(_03620_),
    .Y(_03647_),
    .B1(_03646_));
 sg13g2_or3_1 _21249_ (.A(_10757_),
    .B(_03645_),
    .C(_03647_),
    .X(_03648_));
 sg13g2_buf_1 _21250_ (.A(_03648_),
    .X(_03649_));
 sg13g2_a21oi_1 _21251_ (.A1(_03474_),
    .A2(_03559_),
    .Y(_03650_),
    .B1(_03560_));
 sg13g2_nor2_1 _21252_ (.A(net204),
    .B(_03650_),
    .Y(_03651_));
 sg13g2_nand4_1 _21253_ (.B(_03638_),
    .C(_03649_),
    .A(_03605_),
    .Y(_03652_),
    .D(_03651_));
 sg13g2_nor2_1 _21254_ (.A(net174),
    .B(net172),
    .Y(_03653_));
 sg13g2_nand4_1 _21255_ (.B(_03638_),
    .C(_03649_),
    .A(_03605_),
    .Y(_03654_),
    .D(_03653_));
 sg13g2_a21oi_1 _21256_ (.A1(net173),
    .A2(_03651_),
    .Y(_03655_),
    .B1(_11313_));
 sg13g2_nand3_1 _21257_ (.B(_03654_),
    .C(_03655_),
    .A(_03652_),
    .Y(_03656_));
 sg13g2_nand4_1 _21258_ (.B(_03605_),
    .C(_03638_),
    .A(_03562_),
    .Y(_03657_),
    .D(_03649_));
 sg13g2_nor2_1 _21259_ (.A(_11840_),
    .B(net141),
    .Y(_03658_));
 sg13g2_nand3_1 _21260_ (.B(_03638_),
    .C(_03649_),
    .A(_03605_),
    .Y(_03659_));
 sg13g2_buf_1 _21261_ (.A(_03659_),
    .X(_03660_));
 sg13g2_a22oi_1 _21262_ (.Y(_03661_),
    .B1(_03658_),
    .B2(_03660_),
    .A2(_03657_),
    .A1(_11862_));
 sg13g2_and2_1 _21263_ (.A(net170),
    .B(net233),
    .X(_03662_));
 sg13g2_buf_2 _21264_ (.A(_03662_),
    .X(_03663_));
 sg13g2_a21o_1 _21265_ (.A2(_03661_),
    .A1(_03656_),
    .B1(_03663_),
    .X(_03664_));
 sg13g2_buf_8 _21266_ (.A(_03664_),
    .X(_03665_));
 sg13g2_nor2b_1 _21267_ (.A(_03488_),
    .B_N(_03489_),
    .Y(_03666_));
 sg13g2_buf_2 _21268_ (.A(_03666_),
    .X(_03667_));
 sg13g2_nor2_1 _21269_ (.A(net170),
    .B(net192),
    .Y(_03668_));
 sg13g2_nor2_1 _21270_ (.A(_03667_),
    .B(_03668_),
    .Y(_03669_));
 sg13g2_nor2_1 _21271_ (.A(net143),
    .B(_03668_),
    .Y(_03670_));
 sg13g2_and2_1 _21272_ (.A(_03656_),
    .B(_03661_),
    .X(_03671_));
 sg13g2_buf_8 _21273_ (.A(_03671_),
    .X(_03672_));
 sg13g2_nor2_1 _21274_ (.A(net176),
    .B(_03667_),
    .Y(_03673_));
 sg13g2_buf_1 _21275_ (.A(_03673_),
    .X(_03674_));
 sg13g2_a21o_1 _21276_ (.A2(_03663_),
    .A1(net171),
    .B1(_03674_),
    .X(_03675_));
 sg13g2_a221oi_1 _21277_ (.B2(_03672_),
    .C1(_03675_),
    .B1(_03670_),
    .A1(_03665_),
    .Y(_03676_),
    .A2(_03669_));
 sg13g2_buf_1 _21278_ (.A(_03676_),
    .X(_03677_));
 sg13g2_nand2_1 _21279_ (.Y(_03678_),
    .A(net128),
    .B(_03677_));
 sg13g2_o21ai_1 _21280_ (.B1(net169),
    .Y(_03679_),
    .A1(net128),
    .A2(_03677_));
 sg13g2_nor2_1 _21281_ (.A(_11650_),
    .B(_03579_),
    .Y(_03680_));
 sg13g2_buf_1 _21282_ (.A(_03680_),
    .X(_03681_));
 sg13g2_a21o_1 _21283_ (.A2(_03679_),
    .A1(_03678_),
    .B1(_03681_),
    .X(_03682_));
 sg13g2_nand3_1 _21284_ (.B(_03589_),
    .C(_03682_),
    .A(_03588_),
    .Y(_03683_));
 sg13g2_inv_2 _21285_ (.Y(_03684_),
    .A(_11194_));
 sg13g2_nor2_1 _21286_ (.A(_11633_),
    .B(_03684_),
    .Y(_03685_));
 sg13g2_a22oi_1 _21287_ (.Y(_03686_),
    .B1(_03588_),
    .B2(_03685_),
    .A2(_03583_),
    .A1(\cpu.ex.r_cc ));
 sg13g2_nand3_1 _21288_ (.B(_03683_),
    .C(_03686_),
    .A(_03585_),
    .Y(_00929_));
 sg13g2_or4_1 _21289_ (.A(_10352_),
    .B(net1111),
    .C(_10348_),
    .D(_10351_),
    .X(_03687_));
 sg13g2_nand2b_1 _21290_ (.Y(_03688_),
    .B(_08418_),
    .A_N(_03687_));
 sg13g2_buf_2 _21291_ (.A(_03688_),
    .X(_03689_));
 sg13g2_buf_1 _21292_ (.A(_03689_),
    .X(_03690_));
 sg13g2_buf_1 _21293_ (.A(_03689_),
    .X(_03691_));
 sg13g2_nand2_1 _21294_ (.Y(_03692_),
    .A(\cpu.ex.r_epc[1] ),
    .B(net594));
 sg13g2_o21ai_1 _21295_ (.B1(_03692_),
    .Y(_00931_),
    .A1(_10240_),
    .A2(net595));
 sg13g2_nand2_1 _21296_ (.Y(_03693_),
    .A(\cpu.ex.r_epc[11] ),
    .B(net594));
 sg13g2_o21ai_1 _21297_ (.B1(_03693_),
    .Y(_00932_),
    .A1(_02963_),
    .A2(_03690_));
 sg13g2_buf_1 _21298_ (.A(_08400_),
    .X(_03694_));
 sg13g2_buf_1 _21299_ (.A(net876),
    .X(_03695_));
 sg13g2_nand2_1 _21300_ (.Y(_03696_),
    .A(\cpu.ex.r_epc[12] ),
    .B(net594));
 sg13g2_o21ai_1 _21301_ (.B1(_03696_),
    .Y(_00933_),
    .A1(net742),
    .A2(net595));
 sg13g2_buf_1 _21302_ (.A(_08404_),
    .X(_03697_));
 sg13g2_buf_1 _21303_ (.A(net875),
    .X(_03698_));
 sg13g2_nand2_1 _21304_ (.Y(_03699_),
    .A(\cpu.ex.r_epc[13] ),
    .B(net594));
 sg13g2_o21ai_1 _21305_ (.B1(_03699_),
    .Y(_00934_),
    .A1(net741),
    .A2(net595));
 sg13g2_buf_1 _21306_ (.A(_08512_),
    .X(_03700_));
 sg13g2_buf_1 _21307_ (.A(net740),
    .X(_03701_));
 sg13g2_nand2_1 _21308_ (.Y(_03702_),
    .A(\cpu.ex.r_epc[14] ),
    .B(net594));
 sg13g2_o21ai_1 _21309_ (.B1(_03702_),
    .Y(_00935_),
    .A1(_03701_),
    .A2(net595));
 sg13g2_buf_1 _21310_ (.A(net670),
    .X(_03703_));
 sg13g2_nand2_1 _21311_ (.Y(_03704_),
    .A(\cpu.ex.r_epc[15] ),
    .B(_03689_));
 sg13g2_o21ai_1 _21312_ (.B1(_03704_),
    .Y(_00936_),
    .A1(net593),
    .A2(net595));
 sg13g2_nand2_1 _21313_ (.Y(_03705_),
    .A(\cpu.ex.r_epc[2] ),
    .B(_03689_));
 sg13g2_o21ai_1 _21314_ (.B1(_03705_),
    .Y(_00937_),
    .A1(net806),
    .A2(net595));
 sg13g2_nand2_1 _21315_ (.Y(_03706_),
    .A(\cpu.ex.r_epc[3] ),
    .B(_03689_));
 sg13g2_o21ai_1 _21316_ (.B1(_03706_),
    .Y(_00938_),
    .A1(net758),
    .A2(_03690_));
 sg13g2_buf_1 _21317_ (.A(net760),
    .X(_03707_));
 sg13g2_buf_1 _21318_ (.A(_03707_),
    .X(_03708_));
 sg13g2_nand2_1 _21319_ (.Y(_03709_),
    .A(\cpu.ex.r_epc[4] ),
    .B(_03689_));
 sg13g2_o21ai_1 _21320_ (.B1(_03709_),
    .Y(_00939_),
    .A1(net592),
    .A2(net595));
 sg13g2_nand2_1 _21321_ (.Y(_03710_),
    .A(\cpu.ex.r_epc[5] ),
    .B(_03689_));
 sg13g2_o21ai_1 _21322_ (.B1(_03710_),
    .Y(_00940_),
    .A1(_02944_),
    .A2(net595));
 sg13g2_mux2_1 _21323_ (.A0(_02952_),
    .A1(\cpu.ex.r_epc[6] ),
    .S(net594),
    .X(_00941_));
 sg13g2_mux2_1 _21324_ (.A0(net754),
    .A1(\cpu.ex.r_epc[7] ),
    .S(_03691_),
    .X(_00942_));
 sg13g2_mux2_1 _21325_ (.A0(net753),
    .A1(\cpu.ex.r_epc[8] ),
    .S(_03691_),
    .X(_00943_));
 sg13g2_nand2_1 _21326_ (.Y(_03711_),
    .A(\cpu.ex.r_epc[9] ),
    .B(_03689_));
 sg13g2_o21ai_1 _21327_ (.B1(_03711_),
    .Y(_00944_),
    .A1(_02958_),
    .A2(net594));
 sg13g2_mux2_1 _21328_ (.A0(_02961_),
    .A1(\cpu.ex.r_epc[10] ),
    .S(net594),
    .X(_00945_));
 sg13g2_or4_1 _21329_ (.A(_10352_),
    .B(_10353_),
    .C(_10348_),
    .D(_03448_),
    .X(_03712_));
 sg13g2_buf_2 _21330_ (.A(_03712_),
    .X(_03713_));
 sg13g2_buf_1 _21331_ (.A(_03713_),
    .X(_03714_));
 sg13g2_buf_1 _21332_ (.A(_03713_),
    .X(_03715_));
 sg13g2_nand2_1 _21333_ (.Y(_03716_),
    .A(\cpu.ex.r_lr[1] ),
    .B(net590));
 sg13g2_o21ai_1 _21334_ (.B1(_03716_),
    .Y(_00951_),
    .A1(_10240_),
    .A2(net591));
 sg13g2_nand2_1 _21335_ (.Y(_03717_),
    .A(\cpu.ex.r_lr[11] ),
    .B(net590));
 sg13g2_o21ai_1 _21336_ (.B1(_03717_),
    .Y(_00952_),
    .A1(_02963_),
    .A2(net591));
 sg13g2_nand2_1 _21337_ (.Y(_03718_),
    .A(\cpu.ex.r_lr[12] ),
    .B(net590));
 sg13g2_o21ai_1 _21338_ (.B1(_03718_),
    .Y(_00953_),
    .A1(net742),
    .A2(net591));
 sg13g2_nand2_1 _21339_ (.Y(_03719_),
    .A(\cpu.ex.r_lr[13] ),
    .B(net590));
 sg13g2_o21ai_1 _21340_ (.B1(_03719_),
    .Y(_00954_),
    .A1(net741),
    .A2(net591));
 sg13g2_nand2_1 _21341_ (.Y(_03720_),
    .A(\cpu.ex.r_lr[14] ),
    .B(net590));
 sg13g2_o21ai_1 _21342_ (.B1(_03720_),
    .Y(_00955_),
    .A1(_03701_),
    .A2(net591));
 sg13g2_nand2_1 _21343_ (.Y(_03721_),
    .A(\cpu.ex.r_lr[15] ),
    .B(_03713_));
 sg13g2_o21ai_1 _21344_ (.B1(_03721_),
    .Y(_00956_),
    .A1(net593),
    .A2(net591));
 sg13g2_nand2_1 _21345_ (.Y(_03722_),
    .A(\cpu.ex.r_lr[2] ),
    .B(_03713_));
 sg13g2_o21ai_1 _21346_ (.B1(_03722_),
    .Y(_00957_),
    .A1(net806),
    .A2(_03714_));
 sg13g2_nand2_1 _21347_ (.Y(_03723_),
    .A(\cpu.ex.r_lr[3] ),
    .B(_03713_));
 sg13g2_o21ai_1 _21348_ (.B1(_03723_),
    .Y(_00958_),
    .A1(net758),
    .A2(_03714_));
 sg13g2_nand2_1 _21349_ (.Y(_03724_),
    .A(\cpu.ex.r_lr[4] ),
    .B(_03713_));
 sg13g2_o21ai_1 _21350_ (.B1(_03724_),
    .Y(_00959_),
    .A1(net592),
    .A2(net591));
 sg13g2_nand2_1 _21351_ (.Y(_03725_),
    .A(\cpu.ex.r_lr[5] ),
    .B(_03713_));
 sg13g2_o21ai_1 _21352_ (.B1(_03725_),
    .Y(_00960_),
    .A1(_02944_),
    .A2(net591));
 sg13g2_mux2_1 _21353_ (.A0(net755),
    .A1(\cpu.ex.r_lr[6] ),
    .S(net590),
    .X(_00961_));
 sg13g2_mux2_1 _21354_ (.A0(net754),
    .A1(\cpu.ex.r_lr[7] ),
    .S(_03715_),
    .X(_00962_));
 sg13g2_mux2_1 _21355_ (.A0(net753),
    .A1(\cpu.ex.r_lr[8] ),
    .S(_03715_),
    .X(_00963_));
 sg13g2_nand2_1 _21356_ (.Y(_03726_),
    .A(\cpu.ex.r_lr[9] ),
    .B(_03713_));
 sg13g2_o21ai_1 _21357_ (.B1(_03726_),
    .Y(_00964_),
    .A1(_02958_),
    .A2(net590));
 sg13g2_mux2_1 _21358_ (.A0(net886),
    .A1(\cpu.ex.r_lr[10] ),
    .S(net590),
    .X(_00965_));
 sg13g2_nor2_1 _21359_ (.A(_10467_),
    .B(_11636_),
    .Y(_03727_));
 sg13g2_buf_8 _21360_ (.A(_03727_),
    .X(_03728_));
 sg13g2_buf_8 _21361_ (.A(_03728_),
    .X(_03729_));
 sg13g2_nor2_1 _21362_ (.A(_10984_),
    .B(net29),
    .Y(_03730_));
 sg13g2_xnor2_1 _21363_ (.Y(_03731_),
    .A(net70),
    .B(_03730_));
 sg13g2_buf_1 _21364_ (.A(_10358_),
    .X(_03732_));
 sg13g2_buf_1 _21365_ (.A(net519),
    .X(_03733_));
 sg13g2_nand3_1 _21366_ (.B(_11967_),
    .C(_11998_),
    .A(_11971_),
    .Y(_03734_));
 sg13g2_nand2_1 _21367_ (.Y(_03735_),
    .A(_11564_),
    .B(_11974_));
 sg13g2_a22oi_1 _21368_ (.Y(_03736_),
    .B1(_03735_),
    .B2(net146),
    .A2(_11966_),
    .A1(_11963_));
 sg13g2_o21ai_1 _21369_ (.B1(_10461_),
    .Y(_03737_),
    .A1(_11998_),
    .A2(_03736_));
 sg13g2_nand2_1 _21370_ (.Y(_03738_),
    .A(_10461_),
    .B(_11564_));
 sg13g2_a21oi_1 _21371_ (.A1(_11997_),
    .A2(_03738_),
    .Y(_03739_),
    .B1(_11970_));
 sg13g2_a21oi_1 _21372_ (.A1(_11963_),
    .A2(_11966_),
    .Y(_03740_),
    .B1(_11997_));
 sg13g2_nor2_1 _21373_ (.A(net532),
    .B(net146),
    .Y(_03741_));
 sg13g2_o21ai_1 _21374_ (.B1(_03741_),
    .Y(_03742_),
    .A1(_03739_),
    .A2(_03740_));
 sg13g2_a21oi_1 _21375_ (.A1(_11564_),
    .A2(_03741_),
    .Y(_03743_),
    .B1(_11974_));
 sg13g2_nand2_1 _21376_ (.Y(_03744_),
    .A(net146),
    .B(_11972_));
 sg13g2_nand3_1 _21377_ (.B(_11564_),
    .C(_03744_),
    .A(_10461_),
    .Y(_03745_));
 sg13g2_o21ai_1 _21378_ (.B1(_03745_),
    .Y(_03746_),
    .A1(_11997_),
    .A2(_03743_));
 sg13g2_nand3_1 _21379_ (.B(_11961_),
    .C(_03746_),
    .A(_11844_),
    .Y(_03747_));
 sg13g2_nand4_1 _21380_ (.B(_03737_),
    .C(_03742_),
    .A(_03734_),
    .Y(_03748_),
    .D(_03747_));
 sg13g2_buf_1 _21381_ (.A(_03748_),
    .X(_03749_));
 sg13g2_nand2_1 _21382_ (.Y(_03750_),
    .A(net70),
    .B(_03749_));
 sg13g2_and2_1 _21383_ (.A(\cpu.ex.r_mult[15] ),
    .B(net533),
    .X(_03751_));
 sg13g2_buf_1 _21384_ (.A(_03751_),
    .X(_03752_));
 sg13g2_xnor2_1 _21385_ (.Y(_03753_),
    .A(_03750_),
    .B(_03752_));
 sg13g2_nand3_1 _21386_ (.B(_10359_),
    .C(\cpu.ex.r_cc ),
    .A(_10347_),
    .Y(_03754_));
 sg13g2_and2_1 _21387_ (.A(_09465_),
    .B(_10363_),
    .X(_03755_));
 sg13g2_buf_1 _21388_ (.A(_03755_),
    .X(_03756_));
 sg13g2_nand3_1 _21389_ (.B(_10360_),
    .C(_03756_),
    .A(\cpu.ex.r_mult[16] ),
    .Y(_03757_));
 sg13g2_a21oi_1 _21390_ (.A1(_03754_),
    .A2(_03757_),
    .Y(_03758_),
    .B1(net519));
 sg13g2_a221oi_1 _21391_ (.B2(_03753_),
    .C1(_03758_),
    .B1(_11839_),
    .A1(_03419_),
    .Y(_03759_),
    .A2(net472));
 sg13g2_o21ai_1 _21392_ (.B1(_03759_),
    .Y(_00966_),
    .A1(_11853_),
    .A2(_03731_));
 sg13g2_nand2_1 _21393_ (.Y(_03760_),
    .A(net346),
    .B(_11740_));
 sg13g2_xnor2_1 _21394_ (.Y(_03761_),
    .A(net231),
    .B(_03760_));
 sg13g2_nor2_1 _21395_ (.A(_11635_),
    .B(_03761_),
    .Y(_03762_));
 sg13g2_nor2_2 _21396_ (.A(_10840_),
    .B(_09474_),
    .Y(_03763_));
 sg13g2_nor2b_1 _21397_ (.A(_03762_),
    .B_N(_03763_),
    .Y(_03764_));
 sg13g2_nor3_1 _21398_ (.A(_03729_),
    .B(_03761_),
    .C(_03763_),
    .Y(_03765_));
 sg13g2_o21ai_1 _21399_ (.B1(_11658_),
    .Y(_03766_),
    .A1(_03764_),
    .A2(_03765_));
 sg13g2_nor2_1 _21400_ (.A(_09477_),
    .B(net441),
    .Y(_03767_));
 sg13g2_buf_2 _21401_ (.A(_03767_),
    .X(_03768_));
 sg13g2_nand3_1 _21402_ (.B(_03749_),
    .C(_03752_),
    .A(net70),
    .Y(_03769_));
 sg13g2_nor2_1 _21403_ (.A(net491),
    .B(_11786_),
    .Y(_03770_));
 sg13g2_nor3_1 _21404_ (.A(_11614_),
    .B(_11629_),
    .C(_11631_),
    .Y(_03771_));
 sg13g2_buf_2 _21405_ (.A(_03771_),
    .X(_03772_));
 sg13g2_nor2_1 _21406_ (.A(_03772_),
    .B(_10467_),
    .Y(_03773_));
 sg13g2_a221oi_1 _21407_ (.B2(_03773_),
    .C1(_10840_),
    .B1(_03770_),
    .A1(_03768_),
    .Y(_03774_),
    .A2(_03769_));
 sg13g2_nand2_1 _21408_ (.Y(_03775_),
    .A(net1122),
    .B(net533));
 sg13g2_o21ai_1 _21409_ (.B1(_10840_),
    .Y(_03776_),
    .A1(_03775_),
    .A2(_03769_));
 sg13g2_nand2b_1 _21410_ (.Y(_03777_),
    .B(_03776_),
    .A_N(_03774_));
 sg13g2_nand2_1 _21411_ (.Y(_03778_),
    .A(_10360_),
    .B(_03756_));
 sg13g2_buf_1 _21412_ (.A(_03778_),
    .X(_03779_));
 sg13g2_nand4_1 _21413_ (.B(_10347_),
    .C(_10359_),
    .A(_09120_),
    .Y(_03780_),
    .D(\cpu.ex.r_cc ));
 sg13g2_a21oi_1 _21414_ (.A1(_03779_),
    .A2(_03780_),
    .Y(_03781_),
    .B1(_10358_));
 sg13g2_buf_2 _21415_ (.A(_03781_),
    .X(_03782_));
 sg13g2_inv_1 _21416_ (.Y(_03783_),
    .A(_03782_));
 sg13g2_and3_1 _21417_ (.X(_03784_),
    .A(_03766_),
    .B(_03777_),
    .C(_03783_));
 sg13g2_nor2_1 _21418_ (.A(_10360_),
    .B(_03782_),
    .Y(_03785_));
 sg13g2_nor2_2 _21419_ (.A(_03732_),
    .B(_03785_),
    .Y(_03786_));
 sg13g2_o21ai_1 _21420_ (.B1(_03786_),
    .Y(_03787_),
    .A1(\cpu.ex.r_mult[17] ),
    .A2(_03779_));
 sg13g2_nand2_1 _21421_ (.Y(_03788_),
    .A(_03431_),
    .B(net472));
 sg13g2_o21ai_1 _21422_ (.B1(_03788_),
    .Y(_00967_),
    .A1(_03784_),
    .A2(_03787_));
 sg13g2_buf_1 _21423_ (.A(_03782_),
    .X(_03789_));
 sg13g2_a21oi_1 _21424_ (.A1(net475),
    .A2(net472),
    .Y(_03790_),
    .B1(net162));
 sg13g2_nand2b_1 _21425_ (.Y(_03791_),
    .B(net220),
    .A_N(_03763_));
 sg13g2_and2_1 _21426_ (.A(net231),
    .B(_03763_),
    .X(_03792_));
 sg13g2_buf_1 _21427_ (.A(_03792_),
    .X(_03793_));
 sg13g2_a21oi_1 _21428_ (.A1(_03760_),
    .A2(_03791_),
    .Y(_03794_),
    .B1(_03793_));
 sg13g2_xnor2_1 _21429_ (.Y(_03795_),
    .A(net272),
    .B(_03794_));
 sg13g2_nor2_1 _21430_ (.A(_10844_),
    .B(net491),
    .Y(_03796_));
 sg13g2_o21ai_1 _21431_ (.B1(_03796_),
    .Y(_03797_),
    .A1(_03729_),
    .A2(_03795_));
 sg13g2_or3_1 _21432_ (.A(_03728_),
    .B(_03796_),
    .C(_03795_),
    .X(_03798_));
 sg13g2_a21o_1 _21433_ (.A2(_03798_),
    .A1(_03797_),
    .B1(_11786_),
    .X(_03799_));
 sg13g2_nand4_1 _21434_ (.B(net88),
    .C(_03749_),
    .A(_10841_),
    .Y(_03800_),
    .D(_03752_));
 sg13g2_buf_8 _21435_ (.A(_03800_),
    .X(_03801_));
 sg13g2_nor2_1 _21436_ (.A(_10844_),
    .B(net27),
    .Y(_03802_));
 sg13g2_nand2_1 _21437_ (.Y(_03803_),
    .A(_10844_),
    .B(net27));
 sg13g2_nand3b_1 _21438_ (.B(_03803_),
    .C(_03768_),
    .Y(_03804_),
    .A_N(_03802_));
 sg13g2_a21o_1 _21439_ (.A2(_03804_),
    .A1(_03799_),
    .B1(net442),
    .X(_03805_));
 sg13g2_nand2_1 _21440_ (.Y(_03806_),
    .A(net492),
    .B(_03756_));
 sg13g2_buf_2 _21441_ (.A(_03806_),
    .X(_03807_));
 sg13g2_nor2_1 _21442_ (.A(\cpu.ex.r_mult[18] ),
    .B(_03807_),
    .Y(_03808_));
 sg13g2_a21oi_1 _21443_ (.A1(_03790_),
    .A2(_03805_),
    .Y(_00968_),
    .B1(_03808_));
 sg13g2_o21ai_1 _21444_ (.B1(_03786_),
    .Y(_03809_),
    .A1(\cpu.ex.r_mult[19] ),
    .A2(_03779_));
 sg13g2_nand2_1 _21445_ (.Y(_03810_),
    .A(_10843_),
    .B(_10846_));
 sg13g2_a21oi_1 _21446_ (.A1(_10985_),
    .A2(_11740_),
    .Y(_03811_),
    .B1(_03810_));
 sg13g2_xnor2_1 _21447_ (.Y(_03812_),
    .A(net230),
    .B(_03811_));
 sg13g2_nor2_1 _21448_ (.A(net29),
    .B(_03812_),
    .Y(_03813_));
 sg13g2_xnor2_1 _21449_ (.Y(_03814_),
    .A(_11571_),
    .B(_03813_));
 sg13g2_xnor2_1 _21450_ (.Y(_03815_),
    .A(_10913_),
    .B(_03802_));
 sg13g2_a221oi_1 _21451_ (.B2(_03768_),
    .C1(_03789_),
    .B1(_03815_),
    .A1(net71),
    .Y(_03816_),
    .A2(_03814_));
 sg13g2_nand2_1 _21452_ (.Y(_03817_),
    .A(_03434_),
    .B(net472));
 sg13g2_o21ai_1 _21453_ (.B1(_03817_),
    .Y(_00969_),
    .A1(_03809_),
    .A2(_03816_));
 sg13g2_nand2_1 _21454_ (.Y(_03818_),
    .A(net524),
    .B(net472));
 sg13g2_o21ai_1 _21455_ (.B1(_03786_),
    .Y(_03819_),
    .A1(\cpu.ex.r_mult[20] ),
    .A2(_03779_));
 sg13g2_or2_1 _21456_ (.X(_03820_),
    .B(_10844_),
    .A(_10913_));
 sg13g2_buf_1 _21457_ (.A(_03820_),
    .X(_03821_));
 sg13g2_nor2_1 _21458_ (.A(net27),
    .B(_03821_),
    .Y(_03822_));
 sg13g2_nor3_1 _21459_ (.A(_10909_),
    .B(_11707_),
    .C(_03822_),
    .Y(_03823_));
 sg13g2_nor3_1 _21460_ (.A(_10910_),
    .B(net27),
    .C(_03821_),
    .Y(_03824_));
 sg13g2_o21ai_1 _21461_ (.B1(net1122),
    .Y(_03825_),
    .A1(_03823_),
    .A2(_03824_));
 sg13g2_nand2_1 _21462_ (.Y(_03826_),
    .A(net229),
    .B(_11571_));
 sg13g2_a21oi_1 _21463_ (.A1(_03811_),
    .A2(_03826_),
    .Y(_03827_),
    .B1(_11572_));
 sg13g2_xnor2_1 _21464_ (.Y(_03828_),
    .A(net235),
    .B(_03827_));
 sg13g2_and2_1 _21465_ (.A(_03772_),
    .B(_10465_),
    .X(_03829_));
 sg13g2_or2_1 _21466_ (.X(_03830_),
    .B(_10465_),
    .A(_03772_));
 sg13g2_and2_1 _21467_ (.A(net132),
    .B(_03828_),
    .X(_03831_));
 sg13g2_a22oi_1 _21468_ (.Y(_03832_),
    .B1(_03830_),
    .B2(_03831_),
    .A2(_03829_),
    .A1(_03828_));
 sg13g2_xnor2_1 _21469_ (.Y(_03833_),
    .A(_11566_),
    .B(_03832_));
 sg13g2_a221oi_1 _21470_ (.B2(_03833_),
    .C1(_03789_),
    .B1(net71),
    .A1(net524),
    .Y(_03834_),
    .A2(net472));
 sg13g2_a22oi_1 _21471_ (.Y(_00970_),
    .B1(_03825_),
    .B2(_03834_),
    .A2(_03819_),
    .A1(_03818_));
 sg13g2_or2_1 _21472_ (.X(_03835_),
    .B(_03779_),
    .A(\cpu.ex.r_mult[21] ));
 sg13g2_a22oi_1 _21473_ (.Y(_03836_),
    .B1(_03786_),
    .B2(_03835_),
    .A2(_03733_),
    .A1(_02965_));
 sg13g2_xnor2_1 _21474_ (.Y(_03837_),
    .A(_10841_),
    .B(net220));
 sg13g2_nand2_1 _21475_ (.Y(_03838_),
    .A(_03796_),
    .B(_03837_));
 sg13g2_nand2_1 _21476_ (.Y(_03839_),
    .A(_10913_),
    .B(net230));
 sg13g2_o21ai_1 _21477_ (.B1(_03839_),
    .Y(_03840_),
    .A1(net230),
    .A2(_11571_));
 sg13g2_a22oi_1 _21478_ (.Y(_03841_),
    .B1(_03840_),
    .B2(_10909_),
    .A2(net230),
    .A1(net491));
 sg13g2_or2_1 _21479_ (.X(_03842_),
    .B(_03841_),
    .A(net232));
 sg13g2_xnor2_1 _21480_ (.Y(_03843_),
    .A(_10913_),
    .B(net230));
 sg13g2_nand3_1 _21481_ (.B(_11566_),
    .C(_03843_),
    .A(net232),
    .Y(_03844_));
 sg13g2_nand2_1 _21482_ (.Y(_03845_),
    .A(net220),
    .B(_03763_));
 sg13g2_o21ai_1 _21483_ (.B1(_03845_),
    .Y(_03846_),
    .A1(_10841_),
    .A2(net220));
 sg13g2_a221oi_1 _21484_ (.B2(_10844_),
    .C1(net272),
    .B1(_03846_),
    .A1(_10463_),
    .Y(_03847_),
    .A2(net231));
 sg13g2_a221oi_1 _21485_ (.B2(_03844_),
    .C1(_03847_),
    .B1(_03842_),
    .A1(net272),
    .Y(_03848_),
    .A2(_03838_));
 sg13g2_buf_1 _21486_ (.A(_10838_),
    .X(_03849_));
 sg13g2_o21ai_1 _21487_ (.B1(_03796_),
    .Y(_03850_),
    .A1(net265),
    .A2(_03793_));
 sg13g2_nand2_1 _21488_ (.Y(_03851_),
    .A(net265),
    .B(_03793_));
 sg13g2_and2_1 _21489_ (.A(_03850_),
    .B(_03851_),
    .X(_03852_));
 sg13g2_buf_1 _21490_ (.A(_03852_),
    .X(_03853_));
 sg13g2_nor2_1 _21491_ (.A(net229),
    .B(_03853_),
    .Y(_03854_));
 sg13g2_o21ai_1 _21492_ (.B1(net232),
    .Y(_03855_),
    .A1(net229),
    .A2(_03853_));
 sg13g2_a221oi_1 _21493_ (.B2(net229),
    .C1(_10913_),
    .B1(_03853_),
    .A1(_10909_),
    .Y(_03856_),
    .A2(net232));
 sg13g2_a21oi_1 _21494_ (.A1(_10910_),
    .A2(_03855_),
    .Y(_03857_),
    .B1(_03856_));
 sg13g2_nor2_1 _21495_ (.A(net491),
    .B(_03857_),
    .Y(_03858_));
 sg13g2_a221oi_1 _21496_ (.B2(net235),
    .C1(_03858_),
    .B1(_03854_),
    .A1(_03760_),
    .Y(_03859_),
    .A2(_03848_));
 sg13g2_xnor2_1 _21497_ (.Y(_03860_),
    .A(_11645_),
    .B(_03859_));
 sg13g2_nor3_1 _21498_ (.A(_11786_),
    .B(_03728_),
    .C(_03860_),
    .Y(_03861_));
 sg13g2_a21oi_1 _21499_ (.A1(_12058_),
    .A2(_10358_),
    .Y(_03862_),
    .B1(_03782_));
 sg13g2_nand2_1 _21500_ (.Y(_03863_),
    .A(_10847_),
    .B(_03862_));
 sg13g2_nor2_1 _21501_ (.A(_03861_),
    .B(_03863_),
    .Y(_03864_));
 sg13g2_o21ai_1 _21502_ (.B1(_03770_),
    .Y(_03865_),
    .A1(_03728_),
    .A2(_03860_));
 sg13g2_and3_1 _21503_ (.X(_03866_),
    .A(_10848_),
    .B(_03865_),
    .C(_03862_));
 sg13g2_nand2b_1 _21504_ (.Y(_03867_),
    .B(_10910_),
    .A_N(_03821_));
 sg13g2_buf_2 _21505_ (.A(_03867_),
    .X(_03868_));
 sg13g2_nor2_1 _21506_ (.A(_03801_),
    .B(_03868_),
    .Y(_03869_));
 sg13g2_mux2_1 _21507_ (.A0(_03864_),
    .A1(_03866_),
    .S(_03869_),
    .X(_03870_));
 sg13g2_and2_1 _21508_ (.A(_03775_),
    .B(_03866_),
    .X(_03871_));
 sg13g2_nor3_1 _21509_ (.A(_03768_),
    .B(_03861_),
    .C(_03863_),
    .Y(_03872_));
 sg13g2_nor4_1 _21510_ (.A(_03836_),
    .B(_03870_),
    .C(_03871_),
    .D(_03872_),
    .Y(_00971_));
 sg13g2_a21o_1 _21511_ (.A2(_11577_),
    .A1(net537),
    .B1(_11626_),
    .X(_03873_));
 sg13g2_xnor2_1 _21512_ (.Y(_03874_),
    .A(net202),
    .B(_03873_));
 sg13g2_o21ai_1 _21513_ (.B1(_03874_),
    .Y(_03875_),
    .A1(_10467_),
    .A2(_11636_));
 sg13g2_xnor2_1 _21514_ (.Y(_03876_),
    .A(_11041_),
    .B(_03875_));
 sg13g2_a221oi_1 _21515_ (.B2(_03876_),
    .C1(net162),
    .B1(net62),
    .A1(net984),
    .Y(_03877_),
    .A2(_03733_));
 sg13g2_nor3_1 _21516_ (.A(_10847_),
    .B(net27),
    .C(_03868_),
    .Y(_03878_));
 sg13g2_nor2_1 _21517_ (.A(_11013_),
    .B(_11707_),
    .Y(_03879_));
 sg13g2_xor2_1 _21518_ (.B(_03879_),
    .A(_03878_),
    .X(_03880_));
 sg13g2_nand2_1 _21519_ (.Y(_03881_),
    .A(_11839_),
    .B(_03880_));
 sg13g2_nor2_1 _21520_ (.A(_10997_),
    .B(_03807_),
    .Y(_03882_));
 sg13g2_a21oi_1 _21521_ (.A1(_03877_),
    .A2(_03881_),
    .Y(_00972_),
    .B1(_03882_));
 sg13g2_nor4_1 _21522_ (.A(_11013_),
    .B(_10847_),
    .C(_03801_),
    .D(_03868_),
    .Y(_03883_));
 sg13g2_xnor2_1 _21523_ (.Y(_03884_),
    .A(_11012_),
    .B(_03883_));
 sg13g2_nand2_1 _21524_ (.Y(_03885_),
    .A(_10470_),
    .B(_11616_));
 sg13g2_nand2_1 _21525_ (.Y(_03886_),
    .A(_11618_),
    .B(_03885_));
 sg13g2_xnor2_1 _21526_ (.Y(_03887_),
    .A(net273),
    .B(_03886_));
 sg13g2_o21ai_1 _21527_ (.B1(_03887_),
    .Y(_03888_),
    .A1(_10467_),
    .A2(_11636_));
 sg13g2_xnor2_1 _21528_ (.Y(_03889_),
    .A(_11040_),
    .B(_03888_));
 sg13g2_a221oi_1 _21529_ (.B2(net71),
    .C1(net162),
    .B1(_03889_),
    .A1(_03768_),
    .Y(_03890_),
    .A2(_03884_));
 sg13g2_o21ai_1 _21530_ (.B1(_03786_),
    .Y(_03891_),
    .A1(\cpu.ex.r_mult[23] ),
    .A2(_03779_));
 sg13g2_nand2_1 _21531_ (.Y(_03892_),
    .A(_02954_),
    .B(net472));
 sg13g2_o21ai_1 _21532_ (.B1(_03892_),
    .Y(_00973_),
    .A1(_03890_),
    .A2(_03891_));
 sg13g2_a21oi_1 _21533_ (.A1(net1056),
    .A2(net519),
    .Y(_03893_),
    .B1(_03782_));
 sg13g2_nand3_1 _21534_ (.B(_11578_),
    .C(_10848_),
    .A(_10997_),
    .Y(_03894_));
 sg13g2_nor3_1 _21535_ (.A(net27),
    .B(_03868_),
    .C(_03894_),
    .Y(_03895_));
 sg13g2_xnor2_1 _21536_ (.Y(_03896_),
    .A(net1106),
    .B(_03895_));
 sg13g2_nand2_1 _21537_ (.Y(_03897_),
    .A(_03768_),
    .B(_03896_));
 sg13g2_nor2_1 _21538_ (.A(net132),
    .B(_03772_),
    .Y(_03898_));
 sg13g2_xnor2_1 _21539_ (.Y(_03899_),
    .A(net201),
    .B(_11592_));
 sg13g2_nor2_1 _21540_ (.A(_10462_),
    .B(net1106),
    .Y(_03900_));
 sg13g2_a21oi_1 _21541_ (.A1(_10462_),
    .A2(net132),
    .Y(_03901_),
    .B1(_03900_));
 sg13g2_nor2_1 _21542_ (.A(_03899_),
    .B(_03901_),
    .Y(_03902_));
 sg13g2_nand3b_1 _21543_ (.B(_03900_),
    .C(net132),
    .Y(_03903_),
    .A_N(_03899_));
 sg13g2_o21ai_1 _21544_ (.B1(net1106),
    .Y(_03904_),
    .A1(_10462_),
    .A2(_03899_));
 sg13g2_nand3_1 _21545_ (.B(_03903_),
    .C(_03904_),
    .A(_10470_),
    .Y(_03905_));
 sg13g2_a221oi_1 _21546_ (.B2(_03772_),
    .C1(_03905_),
    .B1(_03902_),
    .A1(_10754_),
    .Y(_03906_),
    .A2(_03898_));
 sg13g2_nand2_1 _21547_ (.Y(_03907_),
    .A(net132),
    .B(_03772_));
 sg13g2_nor3_1 _21548_ (.A(_10755_),
    .B(_03907_),
    .C(_03899_),
    .Y(_03908_));
 sg13g2_o21ai_1 _21549_ (.B1(net71),
    .Y(_03909_),
    .A1(_03906_),
    .A2(_03908_));
 sg13g2_and2_1 _21550_ (.A(_03893_),
    .B(_03909_),
    .X(_03910_));
 sg13g2_nor2_1 _21551_ (.A(\cpu.ex.r_mult[24] ),
    .B(_03807_),
    .Y(_03911_));
 sg13g2_a221oi_1 _21552_ (.B2(_03910_),
    .C1(_03911_),
    .B1(_03897_),
    .A1(net442),
    .Y(_00974_),
    .A2(_03893_));
 sg13g2_or2_1 _21553_ (.X(_03912_),
    .B(_03894_),
    .A(net1106));
 sg13g2_nor3_1 _21554_ (.A(net27),
    .B(_03868_),
    .C(_03912_),
    .Y(_03913_));
 sg13g2_xnor2_1 _21555_ (.Y(_03914_),
    .A(_10759_),
    .B(_03913_));
 sg13g2_nand2_1 _21556_ (.Y(_03915_),
    .A(_11904_),
    .B(_03914_));
 sg13g2_nor2_1 _21557_ (.A(net203),
    .B(_10755_),
    .Y(_03916_));
 sg13g2_nand2_1 _21558_ (.Y(_03917_),
    .A(net203),
    .B(_10755_));
 sg13g2_o21ai_1 _21559_ (.B1(_03917_),
    .Y(_03918_),
    .A1(_11592_),
    .A2(_03916_));
 sg13g2_xnor2_1 _21560_ (.Y(_03919_),
    .A(net173),
    .B(_03918_));
 sg13g2_o21ai_1 _21561_ (.B1(_03919_),
    .Y(_03920_),
    .A1(_03772_),
    .A2(_10467_));
 sg13g2_nand2_1 _21562_ (.Y(_03921_),
    .A(_10762_),
    .B(_03920_));
 sg13g2_nor2b_1 _21563_ (.A(_10762_),
    .B_N(_03919_),
    .Y(_03922_));
 sg13g2_nor2b_1 _21564_ (.A(_10465_),
    .B_N(_10762_),
    .Y(_03923_));
 sg13g2_a22oi_1 _21565_ (.Y(_03924_),
    .B1(_03923_),
    .B2(_03907_),
    .A2(_03922_),
    .A1(_03829_));
 sg13g2_nand3_1 _21566_ (.B(_03830_),
    .C(_03922_),
    .A(net132),
    .Y(_03925_));
 sg13g2_nand3_1 _21567_ (.B(_03924_),
    .C(_03925_),
    .A(_03921_),
    .Y(_03926_));
 sg13g2_a221oi_1 _21568_ (.B2(_03926_),
    .C1(net162),
    .B1(net62),
    .A1(_02973_),
    .Y(_03927_),
    .A2(_03732_));
 sg13g2_nor2_1 _21569_ (.A(\cpu.ex.r_mult[25] ),
    .B(_03807_),
    .Y(_03928_));
 sg13g2_a21oi_1 _21570_ (.A1(_03915_),
    .A2(_03927_),
    .Y(_00975_),
    .B1(_03928_));
 sg13g2_a21oi_1 _21571_ (.A1(net1107),
    .A2(net519),
    .Y(_03929_),
    .B1(net162));
 sg13g2_nor2_1 _21572_ (.A(_10759_),
    .B(_03912_),
    .Y(_03930_));
 sg13g2_nand2_1 _21573_ (.Y(_03931_),
    .A(_10690_),
    .B(_03930_));
 sg13g2_nor3_1 _21574_ (.A(net27),
    .B(_03868_),
    .C(_03931_),
    .Y(_03932_));
 sg13g2_a21oi_1 _21575_ (.A1(_03869_),
    .A2(_03930_),
    .Y(_03933_),
    .B1(_10690_));
 sg13g2_or3_1 _21576_ (.A(_03775_),
    .B(_03932_),
    .C(_03933_),
    .X(_03934_));
 sg13g2_nand2_1 _21577_ (.Y(_03935_),
    .A(net172),
    .B(net203));
 sg13g2_nand2_1 _21578_ (.Y(_03936_),
    .A(net537),
    .B(_11597_));
 sg13g2_a21oi_1 _21579_ (.A1(_03935_),
    .A2(_03936_),
    .Y(_03937_),
    .B1(_11592_));
 sg13g2_nand2_1 _21580_ (.Y(_03938_),
    .A(net203),
    .B(_10762_));
 sg13g2_o21ai_1 _21581_ (.B1(_11601_),
    .Y(_03939_),
    .A1(_11592_),
    .A2(_03938_));
 sg13g2_nor2_1 _21582_ (.A(_03937_),
    .B(_03939_),
    .Y(_03940_));
 sg13g2_xnor2_1 _21583_ (.Y(_03941_),
    .A(net200),
    .B(_03940_));
 sg13g2_nor2_1 _21584_ (.A(_03728_),
    .B(_03941_),
    .Y(_03942_));
 sg13g2_xnor2_1 _21585_ (.Y(_03943_),
    .A(_11608_),
    .B(_03942_));
 sg13g2_a221oi_1 _21586_ (.B2(_03943_),
    .C1(net162),
    .B1(net71),
    .A1(net1107),
    .Y(_03944_),
    .A2(net519));
 sg13g2_nor3_1 _21587_ (.A(net1108),
    .B(net442),
    .C(_10364_),
    .Y(_03945_));
 sg13g2_a221oi_1 _21588_ (.B2(_03944_),
    .C1(_03945_),
    .B1(_03934_),
    .A1(net442),
    .Y(_00976_),
    .A2(_03929_));
 sg13g2_a21oi_1 _21589_ (.A1(_10680_),
    .A2(_10358_),
    .Y(_03946_),
    .B1(_03782_));
 sg13g2_nor2_1 _21590_ (.A(\cpu.ex.r_mult[27] ),
    .B(net442),
    .Y(_03947_));
 sg13g2_nand2_1 _21591_ (.Y(_03948_),
    .A(net200),
    .B(_11608_));
 sg13g2_o21ai_1 _21592_ (.B1(_03948_),
    .Y(_03949_),
    .A1(_03937_),
    .A2(_03939_));
 sg13g2_buf_1 _21593_ (.A(_03949_),
    .X(_03950_));
 sg13g2_nand2_1 _21594_ (.Y(_03951_),
    .A(net174),
    .B(_11595_));
 sg13g2_nand2_1 _21595_ (.Y(_03952_),
    .A(_03950_),
    .B(_03951_));
 sg13g2_xnor2_1 _21596_ (.Y(_03953_),
    .A(net147),
    .B(_03952_));
 sg13g2_nor2_1 _21597_ (.A(net29),
    .B(_03953_),
    .Y(_03954_));
 sg13g2_xnor2_1 _21598_ (.Y(_03955_),
    .A(_10688_),
    .B(_03954_));
 sg13g2_xnor2_1 _21599_ (.Y(_03956_),
    .A(_11603_),
    .B(_03932_));
 sg13g2_inv_1 _21600_ (.Y(_03957_),
    .A(_03946_));
 sg13g2_a221oi_1 _21601_ (.B2(_03768_),
    .C1(_03957_),
    .B1(_03956_),
    .A1(net71),
    .Y(_03958_),
    .A2(_03955_));
 sg13g2_a221oi_1 _21602_ (.B2(_03756_),
    .C1(_03958_),
    .B1(_03947_),
    .A1(net442),
    .Y(_00977_),
    .A2(_03946_));
 sg13g2_a21oi_1 _21603_ (.A1(net687),
    .A2(net472),
    .Y(_03959_),
    .B1(net162));
 sg13g2_o21ai_1 _21604_ (.B1(_11619_),
    .Y(_03960_),
    .A1(_10767_),
    .A2(_11592_));
 sg13g2_buf_1 _21605_ (.A(_03960_),
    .X(_03961_));
 sg13g2_xnor2_1 _21606_ (.Y(_03962_),
    .A(net143),
    .B(_03961_));
 sg13g2_nor2_1 _21607_ (.A(net1023),
    .B(net491),
    .Y(_03963_));
 sg13g2_o21ai_1 _21608_ (.B1(_03963_),
    .Y(_03964_),
    .A1(net29),
    .A2(_03962_));
 sg13g2_or3_1 _21609_ (.A(_03728_),
    .B(_03963_),
    .C(_03962_),
    .X(_03965_));
 sg13g2_a21o_1 _21610_ (.A2(_03965_),
    .A1(_03964_),
    .B1(_11786_),
    .X(_03966_));
 sg13g2_nor2_1 _21611_ (.A(net1023),
    .B(net441),
    .Y(_03967_));
 sg13g2_nor4_1 _21612_ (.A(_11603_),
    .B(_10840_),
    .C(_03868_),
    .D(_03931_),
    .Y(_03968_));
 sg13g2_nand4_1 _21613_ (.B(_03749_),
    .C(_03752_),
    .A(net70),
    .Y(_03969_),
    .D(_03968_));
 sg13g2_buf_2 _21614_ (.A(_03969_),
    .X(_03970_));
 sg13g2_mux2_1 _21615_ (.A0(net1023),
    .A1(_03967_),
    .S(_03970_),
    .X(_03971_));
 sg13g2_nand2_1 _21616_ (.Y(_03972_),
    .A(net1122),
    .B(_03971_));
 sg13g2_a21o_1 _21617_ (.A2(_03972_),
    .A1(_03966_),
    .B1(net442),
    .X(_03973_));
 sg13g2_nor2_1 _21618_ (.A(net1022),
    .B(_03807_),
    .Y(_03974_));
 sg13g2_a21oi_1 _21619_ (.A1(_03959_),
    .A2(_03973_),
    .Y(_00978_),
    .B1(_03974_));
 sg13g2_a22oi_1 _21620_ (.Y(_03975_),
    .B1(_03950_),
    .B2(_03951_),
    .A2(net170),
    .A1(_11603_));
 sg13g2_nor2_1 _21621_ (.A(_11603_),
    .B(net170),
    .Y(_03976_));
 sg13g2_o21ai_1 _21622_ (.B1(_10472_),
    .Y(_03977_),
    .A1(_03975_),
    .A2(_03976_));
 sg13g2_nand3_1 _21623_ (.B(_03950_),
    .C(_03951_),
    .A(net170),
    .Y(_03978_));
 sg13g2_a221oi_1 _21624_ (.B2(_10637_),
    .C1(_10472_),
    .B1(_03978_),
    .A1(_11933_),
    .Y(_03979_),
    .A2(_03952_));
 sg13g2_a21o_1 _21625_ (.A2(_03977_),
    .A1(net171),
    .B1(_03979_),
    .X(_03980_));
 sg13g2_nand2_1 _21626_ (.Y(_03981_),
    .A(_10637_),
    .B(_03978_));
 sg13g2_a221oi_1 _21627_ (.B2(net1023),
    .C1(net491),
    .B1(_03981_),
    .A1(net171),
    .Y(_03982_),
    .A2(_03977_));
 sg13g2_mux2_1 _21628_ (.A0(_03980_),
    .A1(_03982_),
    .S(net145),
    .X(_03983_));
 sg13g2_nor2_1 _21629_ (.A(net1022),
    .B(net29),
    .Y(_03984_));
 sg13g2_and2_1 _21630_ (.A(net1022),
    .B(net537),
    .X(_03985_));
 sg13g2_xnor2_1 _21631_ (.Y(_03986_),
    .A(net145),
    .B(_03980_));
 sg13g2_nand2_1 _21632_ (.Y(_03987_),
    .A(_11933_),
    .B(_03952_));
 sg13g2_nor4_1 _21633_ (.A(_10572_),
    .B(net169),
    .C(net29),
    .D(_03987_),
    .Y(_03988_));
 sg13g2_a21o_1 _21634_ (.A2(_03985_),
    .A1(net29),
    .B1(_03988_),
    .X(_03989_));
 sg13g2_a221oi_1 _21635_ (.B2(_03986_),
    .C1(_03989_),
    .B1(_03985_),
    .A1(_03983_),
    .Y(_03990_),
    .A2(_03984_));
 sg13g2_a21o_1 _21636_ (.A2(net519),
    .A1(net791),
    .B1(_03782_),
    .X(_03991_));
 sg13g2_o21ai_1 _21637_ (.B1(net1022),
    .Y(_03992_),
    .A1(net1023),
    .A2(_03970_));
 sg13g2_or3_1 _21638_ (.A(net1022),
    .B(net1023),
    .C(_03970_),
    .X(_03993_));
 sg13g2_a221oi_1 _21639_ (.B2(_03993_),
    .C1(_11792_),
    .B1(_03992_),
    .A1(_09455_),
    .Y(_03994_),
    .A2(_12022_));
 sg13g2_inv_1 _21640_ (.Y(_03995_),
    .A(_10540_));
 sg13g2_nand3_1 _21641_ (.B(net492),
    .C(_03756_),
    .A(_03995_),
    .Y(_03996_));
 sg13g2_o21ai_1 _21642_ (.B1(_03996_),
    .Y(_03997_),
    .A1(_03991_),
    .A2(_03994_));
 sg13g2_o21ai_1 _21643_ (.B1(_03997_),
    .Y(_00979_),
    .A1(_11853_),
    .A2(_03990_));
 sg13g2_nor2_1 _21644_ (.A(\cpu.ex.r_mult[30] ),
    .B(_03807_),
    .Y(_03998_));
 sg13g2_nand2_1 _21645_ (.Y(_03999_),
    .A(net1022),
    .B(_10472_));
 sg13g2_nor2_1 _21646_ (.A(_03970_),
    .B(_03999_),
    .Y(_04000_));
 sg13g2_xnor2_1 _21647_ (.Y(_04001_),
    .A(_03995_),
    .B(_04000_));
 sg13g2_o21ai_1 _21648_ (.B1(_10472_),
    .Y(_04002_),
    .A1(net143),
    .A2(_03961_));
 sg13g2_a21oi_1 _21649_ (.A1(net143),
    .A2(_03961_),
    .Y(_04003_),
    .B1(net169));
 sg13g2_nand2_1 _21650_ (.Y(_04004_),
    .A(_10572_),
    .B(net537));
 sg13g2_a21oi_1 _21651_ (.A1(_04002_),
    .A2(_04003_),
    .Y(_04005_),
    .B1(_04004_));
 sg13g2_nor2_1 _21652_ (.A(net1023),
    .B(net145),
    .Y(_04006_));
 sg13g2_o21ai_1 _21653_ (.B1(_04006_),
    .Y(_04007_),
    .A1(net143),
    .A2(_03961_));
 sg13g2_nand2_1 _21654_ (.Y(_04008_),
    .A(_10576_),
    .B(_03961_));
 sg13g2_o21ai_1 _21655_ (.B1(_04008_),
    .Y(_04009_),
    .A1(net491),
    .A2(_04007_));
 sg13g2_o21ai_1 _21656_ (.B1(net116),
    .Y(_04010_),
    .A1(_04005_),
    .A2(_04009_));
 sg13g2_or3_1 _21657_ (.A(net116),
    .B(_04005_),
    .C(_04009_),
    .X(_04011_));
 sg13g2_a21oi_1 _21658_ (.A1(_04010_),
    .A2(_04011_),
    .Y(_04012_),
    .B1(net29));
 sg13g2_nand2_1 _21659_ (.Y(_04013_),
    .A(_10540_),
    .B(net537));
 sg13g2_xnor2_1 _21660_ (.Y(_04014_),
    .A(_04012_),
    .B(_04013_));
 sg13g2_a21o_1 _21661_ (.A2(net519),
    .A1(net622),
    .B1(_03782_),
    .X(_04015_));
 sg13g2_a221oi_1 _21662_ (.B2(net62),
    .C1(_04015_),
    .B1(_04014_),
    .A1(_11904_),
    .Y(_04016_),
    .A2(_04001_));
 sg13g2_nor2_1 _21663_ (.A(_03998_),
    .B(_04016_),
    .Y(_00980_));
 sg13g2_nor3_1 _21664_ (.A(_03995_),
    .B(_03970_),
    .C(_03999_),
    .Y(_04017_));
 sg13g2_xnor2_1 _21665_ (.Y(_04018_),
    .A(_10462_),
    .B(_04017_));
 sg13g2_nand2_1 _21666_ (.Y(_04019_),
    .A(_11904_),
    .B(_04018_));
 sg13g2_nand2b_1 _21667_ (.Y(_04020_),
    .B(_03907_),
    .A_N(_03898_));
 sg13g2_and2_1 _21668_ (.A(_10465_),
    .B(net62),
    .X(_04021_));
 sg13g2_a221oi_1 _21669_ (.B2(_04021_),
    .C1(net162),
    .B1(_04020_),
    .A1(net926),
    .Y(_04022_),
    .A2(net519));
 sg13g2_nor2_1 _21670_ (.A(\cpu.ex.r_mult[31] ),
    .B(_03807_),
    .Y(_04023_));
 sg13g2_a21oi_1 _21671_ (.A1(_04019_),
    .A2(_04022_),
    .Y(_00981_),
    .B1(_04023_));
 sg13g2_nor2b_1 _21672_ (.A(_08525_),
    .B_N(_11538_),
    .Y(_04024_));
 sg13g2_buf_1 _21673_ (.A(_04024_),
    .X(_04025_));
 sg13g2_inv_1 _21674_ (.Y(_04026_),
    .A(net1053));
 sg13g2_nor2_1 _21675_ (.A(_09356_),
    .B(_11678_),
    .Y(_04027_));
 sg13g2_mux2_1 _21676_ (.A0(_04026_),
    .A1(_04027_),
    .S(_12020_),
    .X(_04028_));
 sg13g2_nand3_1 _21677_ (.B(_04025_),
    .C(_04028_),
    .A(net666),
    .Y(_04029_));
 sg13g2_buf_1 _21678_ (.A(_04029_),
    .X(_04030_));
 sg13g2_buf_1 _21679_ (.A(_04030_),
    .X(_04031_));
 sg13g2_buf_1 _21680_ (.A(_03542_),
    .X(_04032_));
 sg13g2_nand2_1 _21681_ (.Y(_04033_),
    .A(net272),
    .B(net277));
 sg13g2_buf_2 _21682_ (.A(_04033_),
    .X(_04034_));
 sg13g2_nor2_1 _21683_ (.A(_03612_),
    .B(_04034_),
    .Y(_04035_));
 sg13g2_buf_1 _21684_ (.A(_04035_),
    .X(_04036_));
 sg13g2_nand2b_1 _21685_ (.Y(_04037_),
    .B(net140),
    .A_N(net161));
 sg13g2_nand2_1 _21686_ (.Y(_04038_),
    .A(net272),
    .B(net229));
 sg13g2_buf_2 _21687_ (.A(_04038_),
    .X(_04039_));
 sg13g2_or2_1 _21688_ (.X(_04040_),
    .B(_10981_),
    .A(_10963_));
 sg13g2_nor2_1 _21689_ (.A(_10370_),
    .B(_10800_),
    .Y(_04041_));
 sg13g2_a22oi_1 _21690_ (.Y(_04042_),
    .B1(_04040_),
    .B2(_04041_),
    .A2(net1030),
    .A1(net1060));
 sg13g2_buf_1 _21691_ (.A(_04042_),
    .X(_04043_));
 sg13g2_nor2_1 _21692_ (.A(_04039_),
    .B(net217),
    .Y(_04044_));
 sg13g2_nor2_1 _21693_ (.A(net265),
    .B(net230),
    .Y(_04045_));
 sg13g2_nor2_1 _21694_ (.A(_10984_),
    .B(net231),
    .Y(_04046_));
 sg13g2_a21oi_1 _21695_ (.A1(_04045_),
    .A2(_04046_),
    .Y(_04047_),
    .B1(_11643_));
 sg13g2_nor2_1 _21696_ (.A(_08373_),
    .B(_04047_),
    .Y(_04048_));
 sg13g2_o21ai_1 _21697_ (.B1(net164),
    .Y(_04049_),
    .A1(_04044_),
    .A2(_04048_));
 sg13g2_nand2_1 _21698_ (.Y(_04050_),
    .A(_03608_),
    .B(_04045_));
 sg13g2_nor2_1 _21699_ (.A(_03591_),
    .B(_04050_),
    .Y(_04051_));
 sg13g2_or2_1 _21700_ (.X(_04052_),
    .B(net217),
    .A(_04034_));
 sg13g2_buf_1 _21701_ (.A(_04052_),
    .X(_04053_));
 sg13g2_nor2_1 _21702_ (.A(net218),
    .B(_04053_),
    .Y(_04054_));
 sg13g2_or2_1 _21703_ (.X(_04055_),
    .B(net217),
    .A(_11642_));
 sg13g2_buf_2 _21704_ (.A(_04055_),
    .X(_04056_));
 sg13g2_nor2_1 _21705_ (.A(net266),
    .B(_04056_),
    .Y(_04057_));
 sg13g2_nand4_1 _21706_ (.B(net220),
    .C(net265),
    .A(net346),
    .Y(_04058_),
    .D(net277));
 sg13g2_buf_2 _21707_ (.A(_04058_),
    .X(_04059_));
 sg13g2_nand4_1 _21708_ (.B(net231),
    .C(_03849_),
    .A(net346),
    .Y(_04060_),
    .D(net277));
 sg13g2_buf_1 _21709_ (.A(_04060_),
    .X(_04061_));
 sg13g2_buf_1 _21710_ (.A(_04061_),
    .X(_04062_));
 sg13g2_o21ai_1 _21711_ (.B1(net139),
    .Y(_04063_),
    .A1(net219),
    .A2(_04059_));
 sg13g2_nor4_1 _21712_ (.A(_04051_),
    .B(_04054_),
    .C(_04057_),
    .D(_04063_),
    .Y(_04064_));
 sg13g2_or4_1 _21713_ (.A(net346),
    .B(net220),
    .C(_03849_),
    .D(_10943_),
    .X(_04065_));
 sg13g2_buf_1 _21714_ (.A(_04065_),
    .X(_04066_));
 sg13g2_buf_1 _21715_ (.A(_04066_),
    .X(_04067_));
 sg13g2_nor2_1 _21716_ (.A(_03532_),
    .B(net138),
    .Y(_04068_));
 sg13g2_nand2_1 _21717_ (.Y(_04069_),
    .A(_10838_),
    .B(_10943_));
 sg13g2_buf_1 _21718_ (.A(_04069_),
    .X(_04070_));
 sg13g2_nand2_1 _21719_ (.Y(_04071_),
    .A(_10983_),
    .B(net231));
 sg13g2_buf_1 _21720_ (.A(_04071_),
    .X(_04072_));
 sg13g2_or2_1 _21721_ (.X(_04073_),
    .B(_04072_),
    .A(net191));
 sg13g2_buf_1 _21722_ (.A(_04073_),
    .X(_04074_));
 sg13g2_nor2_1 _21723_ (.A(net163),
    .B(_04074_),
    .Y(_04075_));
 sg13g2_buf_1 _21724_ (.A(_03650_),
    .X(_04076_));
 sg13g2_nand2b_1 _21725_ (.Y(_04077_),
    .B(_03608_),
    .A_N(net191));
 sg13g2_buf_1 _21726_ (.A(_04077_),
    .X(_04078_));
 sg13g2_nor2_1 _21727_ (.A(net217),
    .B(net191),
    .Y(_04079_));
 sg13g2_buf_1 _21728_ (.A(_04079_),
    .X(_04080_));
 sg13g2_nor2_1 _21729_ (.A(_03612_),
    .B(net191),
    .Y(_04081_));
 sg13g2_buf_2 _21730_ (.A(_04081_),
    .X(_04082_));
 sg13g2_a22oi_1 _21731_ (.Y(_04083_),
    .B1(_04082_),
    .B2(net142),
    .A2(_04080_),
    .A1(net233));
 sg13g2_o21ai_1 _21732_ (.B1(_04083_),
    .Y(_04084_),
    .A1(_04076_),
    .A2(_04078_));
 sg13g2_or2_1 _21733_ (.X(_04085_),
    .B(_04072_),
    .A(_04039_));
 sg13g2_buf_1 _21734_ (.A(_04085_),
    .X(_04086_));
 sg13g2_nor2_1 _21735_ (.A(_04034_),
    .B(_04072_),
    .Y(_04087_));
 sg13g2_buf_2 _21736_ (.A(_04087_),
    .X(_04088_));
 sg13g2_nand2_1 _21737_ (.Y(_04089_),
    .A(_11429_),
    .B(_04088_));
 sg13g2_o21ai_1 _21738_ (.B1(_04089_),
    .Y(_04090_),
    .A1(_03579_),
    .A2(_04086_));
 sg13g2_nor4_1 _21739_ (.A(_04068_),
    .B(_04075_),
    .C(_04084_),
    .D(_04090_),
    .Y(_04091_));
 sg13g2_nand4_1 _21740_ (.B(_04049_),
    .C(_04064_),
    .A(_04037_),
    .Y(_04092_),
    .D(_04091_));
 sg13g2_buf_1 _21741_ (.A(net195),
    .X(_04093_));
 sg13g2_nor2_1 _21742_ (.A(_11642_),
    .B(_04072_),
    .Y(_04094_));
 sg13g2_buf_1 _21743_ (.A(_04094_),
    .X(_04095_));
 sg13g2_buf_1 _21744_ (.A(net127),
    .X(_04096_));
 sg13g2_buf_1 _21745_ (.A(net111),
    .X(_04097_));
 sg13g2_nor2_1 _21746_ (.A(net1135),
    .B(_09991_),
    .Y(_04098_));
 sg13g2_buf_2 _21747_ (.A(_04098_),
    .X(_04099_));
 sg13g2_a21oi_1 _21748_ (.A1(net159),
    .A2(_04097_),
    .Y(_04100_),
    .B1(_04099_));
 sg13g2_nand2_1 _21749_ (.Y(_04101_),
    .A(_04092_),
    .B(_04100_));
 sg13g2_nor2_1 _21750_ (.A(net231),
    .B(_11528_),
    .Y(_04102_));
 sg13g2_nand2_1 _21751_ (.Y(_04103_),
    .A(_11700_),
    .B(_11528_));
 sg13g2_nor2b_1 _21752_ (.A(_04102_),
    .B_N(_04103_),
    .Y(_04104_));
 sg13g2_buf_1 _21753_ (.A(_04104_),
    .X(_04105_));
 sg13g2_buf_1 _21754_ (.A(_11559_),
    .X(_04106_));
 sg13g2_buf_1 _21755_ (.A(net190),
    .X(_04107_));
 sg13g2_o21ai_1 _21756_ (.B1(net346),
    .Y(_04108_),
    .A1(_09997_),
    .A2(net158));
 sg13g2_nand2b_1 _21757_ (.Y(_04109_),
    .B(_04108_),
    .A_N(_04105_));
 sg13g2_nand3b_1 _21758_ (.B(net346),
    .C(_04105_),
    .Y(_04110_),
    .A_N(_09997_));
 sg13g2_o21ai_1 _21759_ (.B1(_04110_),
    .Y(_04111_),
    .A1(net1059),
    .A2(_04105_));
 sg13g2_nor2_1 _21760_ (.A(_10984_),
    .B(net190),
    .Y(_04112_));
 sg13g2_nand2_1 _21761_ (.Y(_04113_),
    .A(_04112_),
    .B(_04105_));
 sg13g2_nand2_1 _21762_ (.Y(_04114_),
    .A(_09997_),
    .B(_04113_));
 sg13g2_a22oi_1 _21763_ (.Y(_04115_),
    .B1(_04114_),
    .B2(_09121_),
    .A2(_04111_),
    .A1(net158));
 sg13g2_nor4_1 _21764_ (.A(_09156_),
    .B(_10019_),
    .C(net1118),
    .D(net1117),
    .Y(_04116_));
 sg13g2_nor4_1 _21765_ (.A(_09119_),
    .B(net1125),
    .C(_09997_),
    .D(_10045_),
    .Y(_04117_));
 sg13g2_and2_1 _21766_ (.A(_04116_),
    .B(_04117_),
    .X(_04118_));
 sg13g2_and2_1 _21767_ (.A(_04099_),
    .B(_04118_),
    .X(_04119_));
 sg13g2_buf_1 _21768_ (.A(_04119_),
    .X(_04120_));
 sg13g2_xor2_1 _21769_ (.B(_04105_),
    .A(_04112_),
    .X(_04121_));
 sg13g2_o21ai_1 _21770_ (.B1(_04121_),
    .Y(_04122_),
    .A1(_10045_),
    .A2(_04120_));
 sg13g2_nor2_1 _21771_ (.A(net1044),
    .B(net190),
    .Y(_04123_));
 sg13g2_nor2_1 _21772_ (.A(_10363_),
    .B(_11672_),
    .Y(_04124_));
 sg13g2_buf_2 _21773_ (.A(_04124_),
    .X(_04125_));
 sg13g2_a221oi_1 _21774_ (.B2(_04123_),
    .C1(_04125_),
    .B1(_04096_),
    .A1(_09156_),
    .Y(_04126_),
    .A2(net173));
 sg13g2_mux2_1 _21775_ (.A0(net1125),
    .A1(net1117),
    .S(_04102_),
    .X(_04127_));
 sg13g2_o21ai_1 _21776_ (.B1(_04103_),
    .Y(_04128_),
    .A1(_10019_),
    .A2(_04127_));
 sg13g2_nand3_1 _21777_ (.B(_04126_),
    .C(_04128_),
    .A(_04122_),
    .Y(_04129_));
 sg13g2_a21oi_1 _21778_ (.A1(_04109_),
    .A2(_04115_),
    .Y(_04130_),
    .B1(_04129_));
 sg13g2_nand2_1 _21779_ (.Y(_04131_),
    .A(_04101_),
    .B(_04130_));
 sg13g2_o21ai_1 _21780_ (.B1(_04131_),
    .Y(_04132_),
    .A1(_11674_),
    .A2(\cpu.ex.c_mult[1] ));
 sg13g2_nor3_1 _21781_ (.A(_09356_),
    .B(_09385_),
    .C(_09457_),
    .Y(_04133_));
 sg13g2_and3_1 _21782_ (.X(_04134_),
    .A(_04025_),
    .B(_12021_),
    .C(_04133_));
 sg13g2_buf_1 _21783_ (.A(_04134_),
    .X(_04135_));
 sg13g2_inv_1 _21784_ (.Y(_04136_),
    .A(_04030_));
 sg13g2_nand2_1 _21785_ (.Y(_04137_),
    .A(\cpu.dec.iready ),
    .B(_00199_));
 sg13g2_nor2_1 _21786_ (.A(\cpu.ex.r_branch_stall ),
    .B(_04137_),
    .Y(_04138_));
 sg13g2_buf_1 _21787_ (.A(_04138_),
    .X(_04139_));
 sg13g2_nand3_1 _21788_ (.B(net282),
    .C(_04139_),
    .A(_09284_),
    .Y(_04140_));
 sg13g2_o21ai_1 _21789_ (.B1(_09457_),
    .Y(_04141_),
    .A1(_08431_),
    .A2(_08525_));
 sg13g2_a21oi_1 _21790_ (.A1(_04140_),
    .A2(_04141_),
    .Y(_04142_),
    .B1(_09357_));
 sg13g2_nand4_1 _21791_ (.B(_08526_),
    .C(_09334_),
    .A(_11536_),
    .Y(_04143_),
    .D(_04133_));
 sg13g2_nand2_1 _21792_ (.Y(_04144_),
    .A(net930),
    .B(_04143_));
 sg13g2_nor4_1 _21793_ (.A(_04136_),
    .B(net86),
    .C(_04142_),
    .D(_04144_),
    .Y(_04145_));
 sg13g2_buf_1 _21794_ (.A(_04145_),
    .X(_04146_));
 sg13g2_buf_1 _21795_ (.A(_04146_),
    .X(_04147_));
 sg13g2_a22oi_1 _21796_ (.Y(_04148_),
    .B1(net32),
    .B2(net809),
    .A2(net86),
    .A1(_11524_));
 sg13g2_o21ai_1 _21797_ (.B1(_04148_),
    .Y(_00982_),
    .A1(net65),
    .A2(_04132_));
 sg13g2_buf_1 _21798_ (.A(_11674_),
    .X(_04149_));
 sg13g2_nand2_2 _21799_ (.Y(_04150_),
    .A(_04099_),
    .B(_04118_));
 sg13g2_nor2_1 _21800_ (.A(_03663_),
    .B(_03668_),
    .Y(_04151_));
 sg13g2_xnor2_1 _21801_ (.Y(_04152_),
    .A(_03672_),
    .B(_04151_));
 sg13g2_xnor2_1 _21802_ (.Y(_04153_),
    .A(_03568_),
    .B(_04151_));
 sg13g2_nor2_1 _21803_ (.A(_03620_),
    .B(_03635_),
    .Y(_04154_));
 sg13g2_a21o_1 _21804_ (.A2(_03602_),
    .A1(_11429_),
    .B1(_11584_),
    .X(_04155_));
 sg13g2_o21ai_1 _21805_ (.B1(_04155_),
    .Y(_04156_),
    .A1(_03633_),
    .A2(_04154_));
 sg13g2_buf_1 _21806_ (.A(_04156_),
    .X(_04157_));
 sg13g2_nand2_1 _21807_ (.Y(_04158_),
    .A(_03596_),
    .B(_03598_));
 sg13g2_xor2_1 _21808_ (.B(_04158_),
    .A(_04157_),
    .X(_04159_));
 sg13g2_a21oi_1 _21809_ (.A1(_09997_),
    .A2(_04159_),
    .Y(_04160_),
    .B1(_04125_));
 sg13g2_buf_1 _21810_ (.A(_04160_),
    .X(_04161_));
 sg13g2_nor2_2 _21811_ (.A(_08373_),
    .B(_03684_),
    .Y(_04162_));
 sg13g2_o21ai_1 _21812_ (.B1(_04162_),
    .Y(_04163_),
    .A1(net229),
    .A2(_11643_));
 sg13g2_buf_1 _21813_ (.A(_04163_),
    .X(_04164_));
 sg13g2_nor2_1 _21814_ (.A(_03591_),
    .B(_04056_),
    .Y(_04165_));
 sg13g2_nor2_1 _21815_ (.A(_11642_),
    .B(_03612_),
    .Y(_04166_));
 sg13g2_buf_1 _21816_ (.A(_04166_),
    .X(_04167_));
 sg13g2_a21oi_1 _21817_ (.A1(_03478_),
    .A2(net137),
    .Y(_04168_),
    .B1(net127));
 sg13g2_nand2b_1 _21818_ (.Y(_04169_),
    .B(_04168_),
    .A_N(_04165_));
 sg13g2_nor2_1 _21819_ (.A(_03684_),
    .B(_04034_),
    .Y(_04170_));
 sg13g2_o21ai_1 _21820_ (.B1(net1135),
    .Y(_04171_),
    .A1(_04169_),
    .A2(_04170_));
 sg13g2_nor2_1 _21821_ (.A(_03684_),
    .B(net138),
    .Y(_04172_));
 sg13g2_o21ai_1 _21822_ (.B1(net1046),
    .Y(_04173_),
    .A1(_04169_),
    .A2(_04172_));
 sg13g2_nand3_1 _21823_ (.B(_04171_),
    .C(_04173_),
    .A(_04164_),
    .Y(_04174_));
 sg13g2_o21ai_1 _21824_ (.B1(_04174_),
    .Y(_04175_),
    .A1(_03492_),
    .A2(net139));
 sg13g2_inv_1 _21825_ (.Y(_04176_),
    .A(_03520_));
 sg13g2_nor2_1 _21826_ (.A(_11640_),
    .B(net191),
    .Y(_04177_));
 sg13g2_buf_1 _21827_ (.A(_04177_),
    .X(_04178_));
 sg13g2_nor2_1 _21828_ (.A(_04034_),
    .B(net217),
    .Y(_04179_));
 sg13g2_buf_1 _21829_ (.A(_04179_),
    .X(_04180_));
 sg13g2_o21ai_1 _21830_ (.B1(_04089_),
    .Y(_04181_),
    .A1(net218),
    .A2(net138));
 sg13g2_a221oi_1 _21831_ (.B2(net193),
    .C1(_04181_),
    .B1(net135),
    .A1(net216),
    .Y(_04182_),
    .A2(net136));
 sg13g2_nor3_1 _21832_ (.A(net190),
    .B(_03612_),
    .C(_04070_),
    .Y(_04183_));
 sg13g2_or2_1 _21833_ (.X(_04184_),
    .B(_04034_),
    .A(_03612_));
 sg13g2_buf_1 _21834_ (.A(_04184_),
    .X(_04185_));
 sg13g2_nor2_1 _21835_ (.A(net219),
    .B(_04185_),
    .Y(_04186_));
 sg13g2_nor2_1 _21836_ (.A(net195),
    .B(_04074_),
    .Y(_04187_));
 sg13g2_nor3_1 _21837_ (.A(_04183_),
    .B(_04186_),
    .C(_04187_),
    .Y(_04188_));
 sg13g2_nand2_1 _21838_ (.Y(_04189_),
    .A(net221),
    .B(_11523_));
 sg13g2_o21ai_1 _21839_ (.B1(_04189_),
    .Y(_04190_),
    .A1(_11524_),
    .A2(_03474_));
 sg13g2_buf_1 _21840_ (.A(_04190_),
    .X(_04191_));
 sg13g2_buf_1 _21841_ (.A(_04191_),
    .X(_04192_));
 sg13g2_nor2_1 _21842_ (.A(_11642_),
    .B(net217),
    .Y(_04193_));
 sg13g2_buf_1 _21843_ (.A(_04193_),
    .X(_04194_));
 sg13g2_o21ai_1 _21844_ (.B1(_04061_),
    .Y(_04195_),
    .A1(_03542_),
    .A2(_04059_));
 sg13g2_a221oi_1 _21845_ (.B2(net141),
    .C1(_04195_),
    .B1(net134),
    .A1(net126),
    .Y(_04196_),
    .A2(_04080_));
 sg13g2_nand3_1 _21846_ (.B(_04188_),
    .C(_04196_),
    .A(_04182_),
    .Y(_04197_));
 sg13g2_nand2_1 _21847_ (.Y(_04198_),
    .A(net163),
    .B(net111));
 sg13g2_nand3_1 _21848_ (.B(_04197_),
    .C(_04198_),
    .A(net1118),
    .Y(_04199_));
 sg13g2_or2_1 _21849_ (.X(_04200_),
    .B(net192),
    .A(_11892_));
 sg13g2_buf_1 _21850_ (.A(_04200_),
    .X(_04201_));
 sg13g2_inv_1 _21851_ (.Y(_04202_),
    .A(_10019_));
 sg13g2_nand2b_1 _21852_ (.Y(_04203_),
    .B(net1125),
    .A_N(_03663_));
 sg13g2_nand2_1 _21853_ (.Y(_04204_),
    .A(net1117),
    .B(_03663_));
 sg13g2_nand3_1 _21854_ (.B(_04203_),
    .C(_04204_),
    .A(_04202_),
    .Y(_04205_));
 sg13g2_a22oi_1 _21855_ (.Y(_04206_),
    .B1(_04201_),
    .B2(_04205_),
    .A2(_11735_),
    .A1(_09156_));
 sg13g2_nand4_1 _21856_ (.B(_04175_),
    .C(_04199_),
    .A(_04161_),
    .Y(_04207_),
    .D(_04206_));
 sg13g2_a21oi_1 _21857_ (.A1(net877),
    .A2(_04153_),
    .Y(_04208_),
    .B1(_04207_));
 sg13g2_o21ai_1 _21858_ (.B1(_04208_),
    .Y(_04209_),
    .A1(_04150_),
    .A2(_04152_));
 sg13g2_o21ai_1 _21859_ (.B1(_04209_),
    .Y(_04210_),
    .A1(net157),
    .A2(\cpu.ex.c_mult[11] ));
 sg13g2_buf_1 _21860_ (.A(_08768_),
    .X(_04211_));
 sg13g2_nand2_2 _21861_ (.Y(_04212_),
    .A(net943),
    .B(_08976_));
 sg13g2_nor2_1 _21862_ (.A(net948),
    .B(_04212_),
    .Y(_04213_));
 sg13g2_buf_2 _21863_ (.A(_04213_),
    .X(_04214_));
 sg13g2_nand3_1 _21864_ (.B(_08806_),
    .C(_04214_),
    .A(net1127),
    .Y(_04215_));
 sg13g2_or2_1 _21865_ (.X(_04216_),
    .B(_04215_),
    .A(net980));
 sg13g2_or2_1 _21866_ (.X(_04217_),
    .B(_04216_),
    .A(_08779_));
 sg13g2_buf_1 _21867_ (.A(_04217_),
    .X(_04218_));
 sg13g2_nor2_1 _21868_ (.A(_08759_),
    .B(_04218_),
    .Y(_04219_));
 sg13g2_nand3_1 _21869_ (.B(_08791_),
    .C(_04219_),
    .A(_08738_),
    .Y(_04220_));
 sg13g2_xnor2_1 _21870_ (.Y(_04221_),
    .A(_00290_),
    .B(_04220_));
 sg13g2_inv_1 _21871_ (.Y(_04222_),
    .A(_04221_));
 sg13g2_buf_1 _21872_ (.A(net86),
    .X(_04223_));
 sg13g2_a22oi_1 _21873_ (.Y(_04224_),
    .B1(_04222_),
    .B2(net64),
    .A2(_04147_),
    .A1(_08746_));
 sg13g2_o21ai_1 _21874_ (.B1(_04224_),
    .Y(_00983_),
    .A1(net65),
    .A2(_04210_));
 sg13g2_buf_1 _21875_ (.A(_04120_),
    .X(_04225_));
 sg13g2_nand2_1 _21876_ (.Y(_04226_),
    .A(_10532_),
    .B(_03667_));
 sg13g2_nand2b_1 _21877_ (.Y(_04227_),
    .B(_04226_),
    .A_N(_03674_));
 sg13g2_buf_1 _21878_ (.A(_04227_),
    .X(_04228_));
 sg13g2_nand2_1 _21879_ (.Y(_04229_),
    .A(net174),
    .B(net163));
 sg13g2_o21ai_1 _21880_ (.B1(_04201_),
    .Y(_04230_),
    .A1(_04229_),
    .A2(_03663_));
 sg13g2_nand2b_1 _21881_ (.Y(_04231_),
    .B(_04230_),
    .A_N(_04228_));
 sg13g2_nand2_1 _21882_ (.Y(_04232_),
    .A(_03663_),
    .B(_04228_));
 sg13g2_nand2_1 _21883_ (.Y(_04233_),
    .A(net172),
    .B(_03657_));
 sg13g2_nand2_1 _21884_ (.Y(_04234_),
    .A(net160),
    .B(_03660_));
 sg13g2_nand2_1 _21885_ (.Y(_04235_),
    .A(_04233_),
    .B(_04234_));
 sg13g2_nor2_2 _21886_ (.A(_11638_),
    .B(net163),
    .Y(_04236_));
 sg13g2_nor3_1 _21887_ (.A(_04236_),
    .B(_03663_),
    .C(_04228_),
    .Y(_04237_));
 sg13g2_and2_1 _21888_ (.A(_04201_),
    .B(_04228_),
    .X(_04238_));
 sg13g2_a22oi_1 _21889_ (.Y(_04239_),
    .B1(_04238_),
    .B2(_03672_),
    .A2(_04237_),
    .A1(_04235_));
 sg13g2_nand3_1 _21890_ (.B(_04232_),
    .C(_04239_),
    .A(_04231_),
    .Y(_04240_));
 sg13g2_xor2_1 _21891_ (.B(_04228_),
    .A(_03573_),
    .X(_04241_));
 sg13g2_a221oi_1 _21892_ (.B2(net164),
    .C1(net111),
    .B1(net137),
    .A1(net131),
    .Y(_04242_),
    .A2(net134));
 sg13g2_o21ai_1 _21893_ (.B1(net164),
    .Y(_04243_),
    .A1(_03608_),
    .A2(_11642_));
 sg13g2_a21oi_1 _21894_ (.A1(_04242_),
    .A2(_04243_),
    .Y(_04244_),
    .B1(_08373_));
 sg13g2_nor2b_1 _21895_ (.A(_04242_),
    .B_N(net1046),
    .Y(_04245_));
 sg13g2_nand2_1 _21896_ (.Y(_04246_),
    .A(_03592_),
    .B(net99));
 sg13g2_o21ai_1 _21897_ (.B1(_04246_),
    .Y(_04247_),
    .A1(_04244_),
    .A2(_04245_));
 sg13g2_nor2_1 _21898_ (.A(net194),
    .B(_04053_),
    .Y(_04248_));
 sg13g2_nor2_1 _21899_ (.A(net163),
    .B(_04056_),
    .Y(_04249_));
 sg13g2_or2_1 _21900_ (.X(_04250_),
    .B(net191),
    .A(_04043_));
 sg13g2_buf_2 _21901_ (.A(_04250_),
    .X(_04251_));
 sg13g2_nor2_1 _21902_ (.A(net159),
    .B(_04251_),
    .Y(_04252_));
 sg13g2_nor2_1 _21903_ (.A(net158),
    .B(_04050_),
    .Y(_04253_));
 sg13g2_nor4_1 _21904_ (.A(_04248_),
    .B(_04249_),
    .C(_04252_),
    .D(_04253_),
    .Y(_04254_));
 sg13g2_nor2_1 _21905_ (.A(net191),
    .B(_04072_),
    .Y(_04255_));
 sg13g2_buf_1 _21906_ (.A(_04255_),
    .X(_04256_));
 sg13g2_nor2_1 _21907_ (.A(_03542_),
    .B(_04066_),
    .Y(_04257_));
 sg13g2_nand4_1 _21908_ (.B(_11700_),
    .C(net272),
    .A(net346),
    .Y(_04258_),
    .D(net277));
 sg13g2_buf_1 _21909_ (.A(_04258_),
    .X(_04259_));
 sg13g2_nor2_1 _21910_ (.A(net218),
    .B(net156),
    .Y(_04260_));
 sg13g2_or2_1 _21911_ (.X(_04261_),
    .B(_04260_),
    .A(_04257_));
 sg13g2_a221oi_1 _21912_ (.B2(net216),
    .C1(_04261_),
    .B1(net125),
    .A1(net193),
    .Y(_04262_),
    .A2(net140));
 sg13g2_a22oi_1 _21913_ (.Y(_04263_),
    .B1(_04082_),
    .B2(_04192_),
    .A2(net136),
    .A1(net274));
 sg13g2_a21oi_1 _21914_ (.A1(net141),
    .A2(net137),
    .Y(_04264_),
    .B1(net127));
 sg13g2_nand4_1 _21915_ (.B(_04262_),
    .C(_04263_),
    .A(_04254_),
    .Y(_04265_),
    .D(_04264_));
 sg13g2_or2_1 _21916_ (.X(_04266_),
    .B(net139),
    .A(net192));
 sg13g2_nand3_1 _21917_ (.B(_04265_),
    .C(_04266_),
    .A(net1118),
    .Y(_04267_));
 sg13g2_o21ai_1 _21918_ (.B1(net1057),
    .Y(_04268_),
    .A1(_03487_),
    .A2(_03667_));
 sg13g2_nand2_1 _21919_ (.Y(_04269_),
    .A(net1043),
    .B(_03674_));
 sg13g2_nand3_1 _21920_ (.B(_04268_),
    .C(_04269_),
    .A(_04202_),
    .Y(_04270_));
 sg13g2_a22oi_1 _21921_ (.Y(_04271_),
    .B1(_04226_),
    .B2(_04270_),
    .A2(_11653_),
    .A1(net1058));
 sg13g2_nand4_1 _21922_ (.B(_04247_),
    .C(_04267_),
    .A(_04161_),
    .Y(_04272_),
    .D(_04271_));
 sg13g2_a221oi_1 _21923_ (.B2(net877),
    .C1(_04272_),
    .B1(_04241_),
    .A1(net589),
    .Y(_04273_),
    .A2(_04240_));
 sg13g2_buf_1 _21924_ (.A(_04125_),
    .X(_04274_));
 sg13g2_nand2b_1 _21925_ (.Y(_04275_),
    .B(net155),
    .A_N(_11909_));
 sg13g2_a221oi_1 _21926_ (.B2(_11900_),
    .C1(_04275_),
    .B1(_11908_),
    .A1(_11902_),
    .Y(_04276_),
    .A2(_11906_));
 sg13g2_nor3_1 _21927_ (.A(net65),
    .B(_04273_),
    .C(_04276_),
    .Y(_04277_));
 sg13g2_inv_1 _21928_ (.Y(_04278_),
    .A(_08746_));
 sg13g2_nor2_2 _21929_ (.A(net979),
    .B(_04220_),
    .Y(_04279_));
 sg13g2_xnor2_1 _21930_ (.Y(_04280_),
    .A(_00289_),
    .B(_04279_));
 sg13g2_a22oi_1 _21931_ (.Y(_04281_),
    .B1(_04280_),
    .B2(net64),
    .A2(net32),
    .A1(net719));
 sg13g2_nand2b_1 _21932_ (.Y(_00984_),
    .B(_04281_),
    .A_N(_04277_));
 sg13g2_o21ai_1 _21933_ (.B1(_03487_),
    .Y(_04282_),
    .A1(net129),
    .A2(_03573_));
 sg13g2_and2_1 _21934_ (.A(net129),
    .B(_03573_),
    .X(_04283_));
 sg13g2_nor2_1 _21935_ (.A(net175),
    .B(_03484_),
    .Y(_04284_));
 sg13g2_nor2_2 _21936_ (.A(net199),
    .B(_03591_),
    .Y(_04285_));
 sg13g2_nor2_1 _21937_ (.A(_04284_),
    .B(_04285_),
    .Y(_04286_));
 sg13g2_nor3_1 _21938_ (.A(_09121_),
    .B(_04283_),
    .C(_04286_),
    .Y(_04287_));
 sg13g2_xnor2_1 _21939_ (.Y(_04288_),
    .A(_03677_),
    .B(_04286_));
 sg13g2_nand2_1 _21940_ (.Y(_04289_),
    .A(_09119_),
    .B(_04286_));
 sg13g2_nor2_1 _21941_ (.A(_03493_),
    .B(_04289_),
    .Y(_04290_));
 sg13g2_nand2_1 _21942_ (.Y(_04291_),
    .A(_03579_),
    .B(net111));
 sg13g2_o21ai_1 _21943_ (.B1(net1135),
    .Y(_04292_),
    .A1(net196),
    .A2(net127));
 sg13g2_inv_1 _21944_ (.Y(_04293_),
    .A(_04292_));
 sg13g2_nand2_1 _21945_ (.Y(_04294_),
    .A(_10532_),
    .B(net129));
 sg13g2_a22oi_1 _21946_ (.Y(_04295_),
    .B1(net127),
    .B2(net131),
    .A2(net134),
    .A1(net196));
 sg13g2_nand2b_1 _21947_ (.Y(_04296_),
    .B(net1046),
    .A_N(_04295_));
 sg13g2_o21ai_1 _21948_ (.B1(_04296_),
    .Y(_04297_),
    .A1(_04294_),
    .A2(_04289_));
 sg13g2_a221oi_1 _21949_ (.B2(_04293_),
    .C1(_04297_),
    .B1(_04291_),
    .A1(_09156_),
    .Y(_04298_),
    .A2(_11645_));
 sg13g2_mux2_1 _21950_ (.A0(net1125),
    .A1(net1117),
    .S(_04285_),
    .X(_04299_));
 sg13g2_nand2_1 _21951_ (.Y(_04300_),
    .A(net169),
    .B(net128));
 sg13g2_o21ai_1 _21952_ (.B1(_04300_),
    .Y(_04301_),
    .A1(net1045),
    .A2(_04299_));
 sg13g2_nor2_1 _21953_ (.A(net194),
    .B(_04185_),
    .Y(_04302_));
 sg13g2_nor2_1 _21954_ (.A(net161),
    .B(_04259_),
    .Y(_04303_));
 sg13g2_nand2_1 _21955_ (.Y(_04304_),
    .A(_11290_),
    .B(net134));
 sg13g2_o21ai_1 _21956_ (.B1(_04304_),
    .Y(_04305_),
    .A1(net190),
    .A2(_04086_));
 sg13g2_nor2_2 _21957_ (.A(_11640_),
    .B(_04034_),
    .Y(_04306_));
 sg13g2_a22oi_1 _21958_ (.Y(_04307_),
    .B1(_04306_),
    .B2(net141),
    .A2(_04178_),
    .A1(net193));
 sg13g2_o21ai_1 _21959_ (.B1(_04307_),
    .Y(_04308_),
    .A1(net266),
    .A2(_04251_));
 sg13g2_nor4_1 _21960_ (.A(_04302_),
    .B(_04303_),
    .C(_04305_),
    .D(_04308_),
    .Y(_04309_));
 sg13g2_nor2_2 _21961_ (.A(_11640_),
    .B(_04039_),
    .Y(_04310_));
 sg13g2_a21oi_1 _21962_ (.A1(_04192_),
    .A2(_04310_),
    .Y(_04311_),
    .B1(_04054_));
 sg13g2_a21oi_1 _21963_ (.A1(_11313_),
    .A2(net137),
    .Y(_04312_),
    .B1(net127));
 sg13g2_nor3_1 _21964_ (.A(net159),
    .B(_03612_),
    .C(net191),
    .Y(_04313_));
 sg13g2_a21oi_1 _21965_ (.A1(net274),
    .A2(net125),
    .Y(_04314_),
    .B1(_04313_));
 sg13g2_nand4_1 _21966_ (.B(_04311_),
    .C(_04312_),
    .A(_04309_),
    .Y(_04315_),
    .D(_04314_));
 sg13g2_a21oi_1 _21967_ (.A1(_03667_),
    .A2(net111),
    .Y(_04316_),
    .B1(net1044));
 sg13g2_nand2_1 _21968_ (.Y(_04317_),
    .A(_04315_),
    .B(_04316_));
 sg13g2_nand4_1 _21969_ (.B(_04298_),
    .C(_04301_),
    .A(_04161_),
    .Y(_04318_),
    .D(_04317_));
 sg13g2_a21o_1 _21970_ (.A2(_04290_),
    .A1(_03573_),
    .B1(_04318_),
    .X(_04319_));
 sg13g2_a221oi_1 _21971_ (.B2(net589),
    .C1(_04319_),
    .B1(_04288_),
    .A1(_04282_),
    .Y(_04320_),
    .A2(_04287_));
 sg13g2_o21ai_1 _21972_ (.B1(_04136_),
    .Y(_04321_),
    .A1(net157),
    .A2(\cpu.ex.c_mult[13] ));
 sg13g2_nand2_1 _21973_ (.Y(_04322_),
    .A(net719),
    .B(_04279_));
 sg13g2_xor2_1 _21974_ (.B(_04322_),
    .A(_00196_),
    .X(_04323_));
 sg13g2_a22oi_1 _21975_ (.Y(_04324_),
    .B1(_04323_),
    .B2(net64),
    .A2(net32),
    .A1(net816));
 sg13g2_o21ai_1 _21976_ (.B1(_04324_),
    .Y(_00985_),
    .A1(_04320_),
    .A2(_04321_));
 sg13g2_nand2_1 _21977_ (.Y(_04325_),
    .A(net145),
    .B(net128));
 sg13g2_nand2b_1 _21978_ (.Y(_04326_),
    .B(_03589_),
    .A_N(_03681_));
 sg13g2_nand3_1 _21979_ (.B(_04283_),
    .C(_04326_),
    .A(_04325_),
    .Y(_04327_));
 sg13g2_nand2_1 _21980_ (.Y(_04328_),
    .A(_03494_),
    .B(_03573_));
 sg13g2_inv_1 _21981_ (.Y(_04329_),
    .A(_03589_));
 sg13g2_nor2_2 _21982_ (.A(_03681_),
    .B(_04329_),
    .Y(_04330_));
 sg13g2_a21o_1 _21983_ (.A2(_04326_),
    .A1(_03573_),
    .B1(net129),
    .X(_04331_));
 sg13g2_nor2_1 _21984_ (.A(net171),
    .B(_03486_),
    .Y(_04332_));
 sg13g2_o21ai_1 _21985_ (.B1(net877),
    .Y(_04333_),
    .A1(_11914_),
    .A2(net128));
 sg13g2_a221oi_1 _21986_ (.B2(_04332_),
    .C1(_04333_),
    .B1(_04331_),
    .A1(_04328_),
    .Y(_04334_),
    .A2(_04330_));
 sg13g2_nor2_1 _21987_ (.A(_03668_),
    .B(_04284_),
    .Y(_04335_));
 sg13g2_nor2_1 _21988_ (.A(net128),
    .B(_03667_),
    .Y(_04336_));
 sg13g2_a21o_1 _21989_ (.A2(_04335_),
    .A1(_03665_),
    .B1(_04336_),
    .X(_04337_));
 sg13g2_nor2_1 _21990_ (.A(net147),
    .B(_04284_),
    .Y(_04338_));
 sg13g2_a21oi_1 _21991_ (.A1(_11638_),
    .A2(net163),
    .Y(_04339_),
    .B1(_03667_));
 sg13g2_nand4_1 _21992_ (.B(_04234_),
    .C(_04338_),
    .A(_04233_),
    .Y(_04340_),
    .D(_04339_));
 sg13g2_and2_1 _21993_ (.A(net233),
    .B(net142),
    .X(_04341_));
 sg13g2_buf_1 _21994_ (.A(_04341_),
    .X(_04342_));
 sg13g2_nand4_1 _21995_ (.B(_04233_),
    .C(_04234_),
    .A(_04229_),
    .Y(_04343_),
    .D(_04342_));
 sg13g2_nand3_1 _21996_ (.B(_04236_),
    .C(_04338_),
    .A(net129),
    .Y(_04344_));
 sg13g2_nand2_1 _21997_ (.Y(_04345_),
    .A(_04342_),
    .B(_04338_));
 sg13g2_nand2_1 _21998_ (.Y(_04346_),
    .A(_04344_),
    .B(_04345_));
 sg13g2_a21oi_1 _21999_ (.A1(_04236_),
    .A2(_04342_),
    .Y(_04347_),
    .B1(_04346_));
 sg13g2_nand4_1 _22000_ (.B(_04340_),
    .C(_04343_),
    .A(net143),
    .Y(_04348_),
    .D(_04347_));
 sg13g2_nand3_1 _22001_ (.B(_04337_),
    .C(_04348_),
    .A(_04330_),
    .Y(_04349_));
 sg13g2_xnor2_1 _22002_ (.Y(_04350_),
    .A(net128),
    .B(_03674_));
 sg13g2_a21oi_1 _22003_ (.A1(_03674_),
    .A2(_04300_),
    .Y(_04351_),
    .B1(_04330_));
 sg13g2_nand2_1 _22004_ (.Y(_04352_),
    .A(_03665_),
    .B(_04335_));
 sg13g2_o21ai_1 _22005_ (.B1(net589),
    .Y(_04353_),
    .A1(_04226_),
    .A2(_04330_));
 sg13g2_a221oi_1 _22006_ (.B2(_04352_),
    .C1(_04353_),
    .B1(_04351_),
    .A1(net145),
    .Y(_04354_),
    .A2(_04350_));
 sg13g2_nand2_1 _22007_ (.Y(_04355_),
    .A(net1135),
    .B(_03473_));
 sg13g2_nor2_1 _22008_ (.A(net161),
    .B(_04053_),
    .Y(_04356_));
 sg13g2_nor2_1 _22009_ (.A(net195),
    .B(_04050_),
    .Y(_04357_));
 sg13g2_nor2_1 _22010_ (.A(_03558_),
    .B(_04066_),
    .Y(_04358_));
 sg13g2_nor3_1 _22011_ (.A(_04356_),
    .B(_04357_),
    .C(_04358_),
    .Y(_04359_));
 sg13g2_o21ai_1 _22012_ (.B1(_04359_),
    .Y(_04360_),
    .A1(net219),
    .A2(_04251_));
 sg13g2_nor3_1 _22013_ (.A(net266),
    .B(_03612_),
    .C(_04070_),
    .Y(_04361_));
 sg13g2_nor3_1 _22014_ (.A(net190),
    .B(_04039_),
    .C(_04043_),
    .Y(_04362_));
 sg13g2_nand2_1 _22015_ (.Y(_04363_),
    .A(net142),
    .B(net134));
 sg13g2_o21ai_1 _22016_ (.B1(_04363_),
    .Y(_04364_),
    .A1(net194),
    .A2(_04078_));
 sg13g2_nor4_1 _22017_ (.A(_04360_),
    .B(_04361_),
    .C(_04362_),
    .D(_04364_),
    .Y(_04365_));
 sg13g2_o21ai_1 _22018_ (.B1(net139),
    .Y(_04366_),
    .A1(net218),
    .A2(_04185_));
 sg13g2_nor2_1 _22019_ (.A(_04039_),
    .B(_04072_),
    .Y(_04367_));
 sg13g2_nand2_1 _22020_ (.Y(_04368_),
    .A(net233),
    .B(net137));
 sg13g2_o21ai_1 _22021_ (.B1(_04368_),
    .Y(_04369_),
    .A1(net160),
    .A2(net156));
 sg13g2_a221oi_1 _22022_ (.B2(net193),
    .C1(_04369_),
    .B1(net125),
    .A1(net126),
    .Y(_04370_),
    .A2(_04367_));
 sg13g2_nor2b_1 _22023_ (.A(_04366_),
    .B_N(_04370_),
    .Y(_04371_));
 sg13g2_a221oi_1 _22024_ (.B2(_04371_),
    .C1(net1044),
    .B1(_04365_),
    .A1(_03592_),
    .Y(_04372_),
    .A2(net99));
 sg13g2_inv_1 _22025_ (.Y(_04373_),
    .A(_09156_));
 sg13g2_nand3_1 _22026_ (.B(net164),
    .C(net99),
    .A(net1046),
    .Y(_04374_));
 sg13g2_o21ai_1 _22027_ (.B1(_04374_),
    .Y(_04375_),
    .A1(_04373_),
    .A2(_11011_));
 sg13g2_and3_1 _22028_ (.X(_04376_),
    .A(net1059),
    .B(_03575_),
    .C(_04330_));
 sg13g2_nor2_1 _22029_ (.A(_11925_),
    .B(_04150_),
    .Y(_04377_));
 sg13g2_o21ai_1 _22030_ (.B1(_04377_),
    .Y(_04378_),
    .A1(net130),
    .A2(_03674_));
 sg13g2_nand3b_1 _22031_ (.B(_03681_),
    .C(_04378_),
    .Y(_04379_),
    .A_N(net1043));
 sg13g2_o21ai_1 _22032_ (.B1(_04379_),
    .Y(_04380_),
    .A1(net1057),
    .A2(_04326_));
 sg13g2_a22oi_1 _22033_ (.Y(_04381_),
    .B1(_04380_),
    .B2(_04202_),
    .A2(_04378_),
    .A1(_04329_));
 sg13g2_nor4_1 _22034_ (.A(_04372_),
    .B(_04375_),
    .C(_04376_),
    .D(_04381_),
    .Y(_04382_));
 sg13g2_nand3_1 _22035_ (.B(_04355_),
    .C(_04382_),
    .A(_04161_),
    .Y(_04383_));
 sg13g2_a221oi_1 _22036_ (.B2(_04354_),
    .C1(_04383_),
    .B1(_04349_),
    .A1(_04327_),
    .Y(_04384_),
    .A2(_04334_));
 sg13g2_o21ai_1 _22037_ (.B1(_04136_),
    .Y(_04385_),
    .A1(net157),
    .A2(\cpu.ex.c_mult[14] ));
 sg13g2_nand3_1 _22038_ (.B(net816),
    .C(_04279_),
    .A(net719),
    .Y(_04386_));
 sg13g2_xor2_1 _22039_ (.B(_04386_),
    .A(_00195_),
    .X(_04387_));
 sg13g2_a22oi_1 _22040_ (.Y(_04388_),
    .B1(_04387_),
    .B2(net64),
    .A2(net32),
    .A1(net815));
 sg13g2_o21ai_1 _22041_ (.B1(_04388_),
    .Y(_00986_),
    .A1(_04384_),
    .A2(_04385_));
 sg13g2_or2_1 _22042_ (.X(_04389_),
    .B(_03685_),
    .A(_03587_));
 sg13g2_buf_2 _22043_ (.A(_04389_),
    .X(_04390_));
 sg13g2_nand2b_1 _22044_ (.Y(_04391_),
    .B(_03580_),
    .A_N(_04390_));
 sg13g2_nand2_1 _22045_ (.Y(_04392_),
    .A(_03480_),
    .B(_04390_));
 sg13g2_mux2_1 _22046_ (.A0(_04391_),
    .A1(_04392_),
    .S(_03576_),
    .X(_04393_));
 sg13g2_nor2_1 _22047_ (.A(_09121_),
    .B(_04393_),
    .Y(_04394_));
 sg13g2_mux2_1 _22048_ (.A0(net1057),
    .A1(net1043),
    .S(_03685_),
    .X(_04395_));
 sg13g2_nor2_1 _22049_ (.A(net1045),
    .B(_04395_),
    .Y(_04396_));
 sg13g2_nand2_1 _22050_ (.Y(_04397_),
    .A(net1058),
    .B(_11587_));
 sg13g2_o21ai_1 _22051_ (.B1(_04397_),
    .Y(_04398_),
    .A1(_03587_),
    .A2(_04396_));
 sg13g2_mux2_1 _22052_ (.A0(_03480_),
    .A1(_03580_),
    .S(_04390_),
    .X(_04399_));
 sg13g2_nand2_1 _22053_ (.Y(_04400_),
    .A(_03681_),
    .B(_04390_));
 sg13g2_o21ai_1 _22054_ (.B1(_04400_),
    .Y(_04401_),
    .A1(_03589_),
    .A2(_04390_));
 sg13g2_nand2_1 _22055_ (.Y(_04402_),
    .A(net589),
    .B(_04401_));
 sg13g2_o21ai_1 _22056_ (.B1(_04402_),
    .Y(_04403_),
    .A1(_09121_),
    .A2(_04399_));
 sg13g2_nor2_1 _22057_ (.A(_03681_),
    .B(_04390_),
    .Y(_04404_));
 sg13g2_and2_1 _22058_ (.A(_03589_),
    .B(_04390_),
    .X(_04405_));
 sg13g2_a22oi_1 _22059_ (.Y(_04406_),
    .B1(_04405_),
    .B2(_04285_),
    .A2(_04404_),
    .A1(_04284_));
 sg13g2_nor2_1 _22060_ (.A(net159),
    .B(_04086_),
    .Y(_04407_));
 sg13g2_nor2_1 _22061_ (.A(net265),
    .B(net190),
    .Y(_04408_));
 sg13g2_a21oi_1 _22062_ (.A1(net265),
    .A2(net274),
    .Y(_04409_),
    .B1(_04408_));
 sg13g2_nand2_1 _22063_ (.Y(_04410_),
    .A(_11735_),
    .B(_04046_));
 sg13g2_a21oi_1 _22064_ (.A1(net142),
    .A2(net137),
    .Y(_04411_),
    .B1(net127));
 sg13g2_o21ai_1 _22065_ (.B1(_04411_),
    .Y(_04412_),
    .A1(_04409_),
    .A2(_04410_));
 sg13g2_nand2b_1 _22066_ (.Y(_04413_),
    .B(_11313_),
    .A_N(net156));
 sg13g2_nand2_1 _22067_ (.Y(_04414_),
    .A(_04037_),
    .B(_04413_));
 sg13g2_nor4_1 _22068_ (.A(_04165_),
    .B(_04407_),
    .C(_04412_),
    .D(_04414_),
    .Y(_04415_));
 sg13g2_nor2_1 _22069_ (.A(net160),
    .B(_04053_),
    .Y(_04416_));
 sg13g2_a21oi_1 _22070_ (.A1(_11429_),
    .A2(net125),
    .Y(_04417_),
    .B1(_04416_));
 sg13g2_nor2b_1 _22071_ (.A(net138),
    .B_N(net192),
    .Y(_04418_));
 sg13g2_a221oi_1 _22072_ (.B2(net216),
    .C1(_04418_),
    .B1(_04310_),
    .A1(net193),
    .Y(_04419_),
    .A2(_04080_));
 sg13g2_a22oi_1 _22073_ (.Y(_04420_),
    .B1(_04044_),
    .B2(net126),
    .A2(net136),
    .A1(_11454_));
 sg13g2_nand4_1 _22074_ (.B(_04417_),
    .C(_04419_),
    .A(_04415_),
    .Y(_04421_),
    .D(_04420_));
 sg13g2_nand3_1 _22075_ (.B(_04291_),
    .C(_04421_),
    .A(net1118),
    .Y(_04422_));
 sg13g2_o21ai_1 _22076_ (.B1(_04422_),
    .Y(_04423_),
    .A1(_04150_),
    .A2(_04406_));
 sg13g2_nor4_1 _22077_ (.A(_04162_),
    .B(_04398_),
    .C(_04403_),
    .D(_04423_),
    .Y(_04424_));
 sg13g2_nand3_1 _22078_ (.B(_04300_),
    .C(_04405_),
    .A(net589),
    .Y(_04425_));
 sg13g2_nand3b_1 _22079_ (.B(_04404_),
    .C(net589),
    .Y(_04426_),
    .A_N(_04285_));
 sg13g2_mux2_1 _22080_ (.A0(_04425_),
    .A1(_04426_),
    .S(_03677_),
    .X(_04427_));
 sg13g2_nand3_1 _22081_ (.B(_04424_),
    .C(_04427_),
    .A(_04161_),
    .Y(_04428_));
 sg13g2_nand4_1 _22082_ (.B(_11979_),
    .C(_12000_),
    .A(net155),
    .Y(_04429_),
    .D(_12002_));
 sg13g2_o21ai_1 _22083_ (.B1(_04429_),
    .Y(_04430_),
    .A1(_04394_),
    .A2(_04428_));
 sg13g2_nand4_1 _22084_ (.B(net816),
    .C(net815),
    .A(net719),
    .Y(_04431_),
    .D(_04279_));
 sg13g2_xnor2_1 _22085_ (.Y(_04432_),
    .A(_11146_),
    .B(_04431_));
 sg13g2_a22oi_1 _22086_ (.Y(_04433_),
    .B1(_04432_),
    .B2(net64),
    .A2(net32),
    .A1(_08679_));
 sg13g2_o21ai_1 _22087_ (.B1(_04433_),
    .Y(_00987_),
    .A1(net65),
    .A2(_04430_));
 sg13g2_nand3_1 _22088_ (.B(net282),
    .C(_11677_),
    .A(_09284_),
    .Y(_04434_));
 sg13g2_and2_1 _22089_ (.A(_09013_),
    .B(net86),
    .X(_04435_));
 sg13g2_o21ai_1 _22090_ (.B1(net712),
    .Y(_04436_),
    .A1(_04146_),
    .A2(_04435_));
 sg13g2_nand3_1 _22091_ (.B(net809),
    .C(net86),
    .A(net822),
    .Y(_04437_));
 sg13g2_nor2_1 _22092_ (.A(_04176_),
    .B(net139),
    .Y(_04438_));
 sg13g2_nor2_1 _22093_ (.A(net219),
    .B(_04056_),
    .Y(_04439_));
 sg13g2_nand2_1 _22094_ (.Y(_04440_),
    .A(_03479_),
    .B(_04310_));
 sg13g2_a22oi_1 _22095_ (.Y(_04441_),
    .B1(_04082_),
    .B2(net130),
    .A2(_04036_),
    .A1(net141));
 sg13g2_a22oi_1 _22096_ (.Y(_04442_),
    .B1(_04367_),
    .B2(net196),
    .A2(_04080_),
    .A1(net142));
 sg13g2_a22oi_1 _22097_ (.Y(_04443_),
    .B1(net125),
    .B2(net233),
    .A2(net136),
    .A1(_11313_));
 sg13g2_nand4_1 _22098_ (.B(_04441_),
    .C(_04442_),
    .A(_04440_),
    .Y(_04444_),
    .D(_04443_));
 sg13g2_nor2_1 _22099_ (.A(net194),
    .B(net138),
    .Y(_04445_));
 sg13g2_o21ai_1 _22100_ (.B1(_04061_),
    .Y(_04446_),
    .A1(_03532_),
    .A2(_04059_));
 sg13g2_or4_1 _22101_ (.A(_04260_),
    .B(_04356_),
    .C(_04445_),
    .D(_04446_),
    .X(_04447_));
 sg13g2_nor3_1 _22102_ (.A(_04439_),
    .B(_04444_),
    .C(_04447_),
    .Y(_04448_));
 sg13g2_inv_1 _22103_ (.Y(_04449_),
    .A(_04448_));
 sg13g2_a21oi_1 _22104_ (.A1(_03503_),
    .A2(_04045_),
    .Y(_04450_),
    .B1(_11643_));
 sg13g2_o21ai_1 _22105_ (.B1(_04448_),
    .Y(_04451_),
    .A1(_03684_),
    .A2(_04450_));
 sg13g2_a22oi_1 _22106_ (.Y(_04452_),
    .B1(_04451_),
    .B2(net1135),
    .A2(_04449_),
    .A1(_09992_));
 sg13g2_nor2_1 _22107_ (.A(_09997_),
    .B(_10045_),
    .Y(_04453_));
 sg13g2_nand2_1 _22108_ (.Y(_04454_),
    .A(_04453_),
    .B(_04150_));
 sg13g2_buf_2 _22109_ (.A(_04454_),
    .X(_04455_));
 sg13g2_a21o_1 _22110_ (.A2(_04112_),
    .A1(net220),
    .B1(_03610_),
    .X(_04456_));
 sg13g2_nand2_1 _22111_ (.Y(_04457_),
    .A(net265),
    .B(net159));
 sg13g2_nand2_1 _22112_ (.Y(_04458_),
    .A(_03616_),
    .B(_04457_));
 sg13g2_xnor2_1 _22113_ (.Y(_04459_),
    .A(_04456_),
    .B(_04458_));
 sg13g2_or2_1 _22114_ (.X(_04460_),
    .B(_03504_),
    .A(_03502_));
 sg13g2_xor2_1 _22115_ (.B(_04458_),
    .A(_04460_),
    .X(_04461_));
 sg13g2_mux2_1 _22116_ (.A0(net1117),
    .A1(net1125),
    .S(_03616_),
    .X(_04462_));
 sg13g2_o21ai_1 _22117_ (.B1(_04457_),
    .Y(_04463_),
    .A1(_10020_),
    .A2(_04462_));
 sg13g2_nand2_1 _22118_ (.Y(_04464_),
    .A(net126),
    .B(_04095_));
 sg13g2_o21ai_1 _22119_ (.B1(_04464_),
    .Y(_04465_),
    .A1(_04107_),
    .A2(_04056_));
 sg13g2_a221oi_1 _22120_ (.B2(net1118),
    .C1(_04125_),
    .B1(_04465_),
    .A1(_09156_),
    .Y(_04466_),
    .A2(_11840_));
 sg13g2_nand2_1 _22121_ (.Y(_04467_),
    .A(_04463_),
    .B(_04466_));
 sg13g2_a221oi_1 _22122_ (.B2(net1059),
    .C1(_04467_),
    .B1(_04461_),
    .A1(_04455_),
    .Y(_04468_),
    .A2(_04459_));
 sg13g2_o21ai_1 _22123_ (.B1(_04468_),
    .Y(_04469_),
    .A1(_04438_),
    .A2(_04452_));
 sg13g2_o21ai_1 _22124_ (.B1(_04469_),
    .Y(_04470_),
    .A1(net157),
    .A2(\cpu.ex.c_mult[2] ));
 sg13g2_or2_1 _22125_ (.X(_04471_),
    .B(_04470_),
    .A(net65));
 sg13g2_nand4_1 _22126_ (.B(_04436_),
    .C(_04437_),
    .A(_04434_),
    .Y(_00988_),
    .D(_04471_));
 sg13g2_nor2_1 _22127_ (.A(_04303_),
    .B(_04416_),
    .Y(_04472_));
 sg13g2_a22oi_1 _22128_ (.Y(_04473_),
    .B1(_04082_),
    .B2(net131),
    .A2(net136),
    .A1(net233));
 sg13g2_nand2_1 _22129_ (.Y(_04474_),
    .A(_03537_),
    .B(_04193_));
 sg13g2_o21ai_1 _22130_ (.B1(_04474_),
    .Y(_04475_),
    .A1(_03591_),
    .A2(_04251_));
 sg13g2_a221oi_1 _22131_ (.B2(net142),
    .C1(_04475_),
    .B1(net125),
    .A1(_11194_),
    .Y(_04476_),
    .A2(_04310_));
 sg13g2_o21ai_1 _22132_ (.B1(_04061_),
    .Y(_04477_),
    .A1(_03529_),
    .A2(_04059_));
 sg13g2_a221oi_1 _22133_ (.B2(_11454_),
    .C1(_04477_),
    .B1(_04306_),
    .A1(_11313_),
    .Y(_04478_),
    .A2(_04035_));
 sg13g2_nand4_1 _22134_ (.B(_04473_),
    .C(_04476_),
    .A(_04472_),
    .Y(_04479_),
    .D(_04478_));
 sg13g2_nand2_1 _22135_ (.Y(_04480_),
    .A(_09992_),
    .B(_04479_));
 sg13g2_a21oi_1 _22136_ (.A1(_04086_),
    .A2(_04450_),
    .Y(_04481_),
    .B1(_03684_));
 sg13g2_o21ai_1 _22137_ (.B1(net1135),
    .Y(_04482_),
    .A1(_04479_),
    .A2(_04481_));
 sg13g2_nor2_1 _22138_ (.A(net274),
    .B(net139),
    .Y(_04483_));
 sg13g2_a21o_1 _22139_ (.A2(_04482_),
    .A1(_04480_),
    .B1(_04483_),
    .X(_04484_));
 sg13g2_mux2_1 _22140_ (.A0(net1043),
    .A1(net1057),
    .S(_03627_),
    .X(_04485_));
 sg13g2_nand2_1 _22141_ (.Y(_04486_),
    .A(_11731_),
    .B(net266));
 sg13g2_o21ai_1 _22142_ (.B1(_04486_),
    .Y(_04487_),
    .A1(net1045),
    .A2(_04485_));
 sg13g2_a21oi_1 _22143_ (.A1(net126),
    .A2(_04194_),
    .Y(_04488_),
    .B1(net111));
 sg13g2_o21ai_1 _22144_ (.B1(_04488_),
    .Y(_04489_),
    .A1(_04107_),
    .A2(_04059_));
 sg13g2_a21oi_1 _22145_ (.A1(_04093_),
    .A2(net99),
    .Y(_04490_),
    .B1(net1044));
 sg13g2_a221oi_1 _22146_ (.B2(_04490_),
    .C1(_04125_),
    .B1(_04489_),
    .A1(net1058),
    .Y(_04491_),
    .A2(_11892_));
 sg13g2_and3_1 _22147_ (.X(_04492_),
    .A(_04484_),
    .B(_04487_),
    .C(_04491_));
 sg13g2_nand2_1 _22148_ (.Y(_04493_),
    .A(_04457_),
    .B(_04456_));
 sg13g2_nand2_1 _22149_ (.Y(_04494_),
    .A(_03616_),
    .B(_04493_));
 sg13g2_nand2_1 _22150_ (.Y(_04495_),
    .A(_03627_),
    .B(_04486_));
 sg13g2_xnor2_1 _22151_ (.Y(_04496_),
    .A(_04494_),
    .B(_04495_));
 sg13g2_nor2_1 _22152_ (.A(_11714_),
    .B(net195),
    .Y(_04497_));
 sg13g2_nand2_1 _22153_ (.Y(_04498_),
    .A(_11714_),
    .B(net195));
 sg13g2_o21ai_1 _22154_ (.B1(_04498_),
    .Y(_04499_),
    .A1(_04460_),
    .A2(_04497_));
 sg13g2_xnor2_1 _22155_ (.Y(_04500_),
    .A(_04495_),
    .B(_04499_));
 sg13g2_a22oi_1 _22156_ (.Y(_04501_),
    .B1(_04500_),
    .B2(net877),
    .A2(_04496_),
    .A1(_04455_));
 sg13g2_a22oi_1 _22157_ (.Y(_04502_),
    .B1(_04492_),
    .B2(_04501_),
    .A2(_11744_),
    .A1(net155));
 sg13g2_a21oi_1 _22158_ (.A1(_04135_),
    .A2(_04212_),
    .Y(_04503_),
    .B1(_04146_));
 sg13g2_nor2_1 _22159_ (.A(net711),
    .B(_04212_),
    .Y(_04504_));
 sg13g2_o21ai_1 _22160_ (.B1(_04143_),
    .Y(_04505_),
    .A1(_00274_),
    .A2(_04434_));
 sg13g2_a21oi_1 _22161_ (.A1(net86),
    .A2(_04504_),
    .Y(_04506_),
    .B1(_04505_));
 sg13g2_o21ai_1 _22162_ (.B1(_04506_),
    .Y(_04507_),
    .A1(net948),
    .A2(_04503_));
 sg13g2_a21o_1 _22163_ (.A2(_04502_),
    .A1(_04136_),
    .B1(_04507_),
    .X(_00989_));
 sg13g2_nor2b_1 _22164_ (.A(_04214_),
    .B_N(net86),
    .Y(_04508_));
 sg13g2_o21ai_1 _22165_ (.B1(net1127),
    .Y(_04509_),
    .A1(_04146_),
    .A2(_04508_));
 sg13g2_nand3_1 _22166_ (.B(net86),
    .C(_04214_),
    .A(_08562_),
    .Y(_04510_));
 sg13g2_or4_1 _22167_ (.A(_09357_),
    .B(net282),
    .C(_09388_),
    .D(_04139_),
    .X(_04511_));
 sg13g2_nand2_1 _22168_ (.Y(_04512_),
    .A(_03532_),
    .B(net127));
 sg13g2_o21ai_1 _22169_ (.B1(_04039_),
    .Y(_04513_),
    .A1(_11640_),
    .A2(_11642_));
 sg13g2_nand2_1 _22170_ (.Y(_04514_),
    .A(_03490_),
    .B(_04177_));
 sg13g2_nor3_1 _22171_ (.A(_03558_),
    .B(_04034_),
    .C(net217),
    .Y(_04515_));
 sg13g2_a221oi_1 _22172_ (.B2(_11194_),
    .C1(_04515_),
    .B1(_04082_),
    .A1(net233),
    .Y(_04516_),
    .A2(_04035_));
 sg13g2_o21ai_1 _22173_ (.B1(_04061_),
    .Y(_04517_),
    .A1(net218),
    .A2(_04059_));
 sg13g2_a221oi_1 _22174_ (.B2(_11429_),
    .C1(_04517_),
    .B1(_04193_),
    .A1(_03478_),
    .Y(_04518_),
    .A2(_04080_));
 sg13g2_a221oi_1 _22175_ (.B2(_03484_),
    .C1(_04257_),
    .B1(_04255_),
    .A1(_03566_),
    .Y(_04519_),
    .A2(_04088_));
 sg13g2_nand4_1 _22176_ (.B(_04516_),
    .C(_04518_),
    .A(_04514_),
    .Y(_04520_),
    .D(_04519_));
 sg13g2_a21oi_1 _22177_ (.A1(_03472_),
    .A2(_04513_),
    .Y(_04521_),
    .B1(_04520_));
 sg13g2_nand2_1 _22178_ (.Y(_04522_),
    .A(_09991_),
    .B(_04520_));
 sg13g2_o21ai_1 _22179_ (.B1(_04522_),
    .Y(_04523_),
    .A1(_08373_),
    .A2(_04521_));
 sg13g2_inv_1 _22180_ (.Y(_04524_),
    .A(_03634_));
 sg13g2_nor2_1 _22181_ (.A(_10908_),
    .B(net219),
    .Y(_04525_));
 sg13g2_nor2_1 _22182_ (.A(_04524_),
    .B(_04525_),
    .Y(_04526_));
 sg13g2_nand2_1 _22183_ (.Y(_04527_),
    .A(_11731_),
    .B(net216));
 sg13g2_o21ai_1 _22184_ (.B1(_04527_),
    .Y(_04528_),
    .A1(_03514_),
    .A2(_04499_));
 sg13g2_xnor2_1 _22185_ (.Y(_04529_),
    .A(_04526_),
    .B(_04528_));
 sg13g2_nand2b_1 _22186_ (.Y(_04530_),
    .B(net134),
    .A_N(net195));
 sg13g2_nor2_1 _22187_ (.A(_11559_),
    .B(_04066_),
    .Y(_04531_));
 sg13g2_a21oi_1 _22188_ (.A1(_04191_),
    .A2(_04167_),
    .Y(_04532_),
    .B1(_04531_));
 sg13g2_nand3_1 _22189_ (.B(_04530_),
    .C(_04532_),
    .A(_04062_),
    .Y(_04533_));
 sg13g2_nand3b_1 _22190_ (.B(_04533_),
    .C(_10023_),
    .Y(_04534_),
    .A_N(_04438_));
 sg13g2_a21oi_1 _22191_ (.A1(_09156_),
    .A2(net171),
    .Y(_04535_),
    .B1(_04120_));
 sg13g2_mux2_1 _22192_ (.A0(net1125),
    .A1(net1117),
    .S(_04525_),
    .X(_04536_));
 sg13g2_o21ai_1 _22193_ (.B1(_03634_),
    .Y(_04537_),
    .A1(_10019_),
    .A2(_04536_));
 sg13g2_nand3_1 _22194_ (.B(_04535_),
    .C(_04537_),
    .A(_04534_),
    .Y(_04538_));
 sg13g2_a221oi_1 _22195_ (.B2(net1059),
    .C1(_04538_),
    .B1(_04529_),
    .A1(_04512_),
    .Y(_04539_),
    .A2(_04523_));
 sg13g2_nand2_1 _22196_ (.Y(_04540_),
    .A(_03627_),
    .B(_03620_));
 sg13g2_xnor2_1 _22197_ (.Y(_04541_),
    .A(_04540_),
    .B(_04526_));
 sg13g2_a21oi_1 _22198_ (.A1(_04453_),
    .A2(_04539_),
    .Y(_04542_),
    .B1(_04541_));
 sg13g2_o21ai_1 _22199_ (.B1(_11674_),
    .Y(_04543_),
    .A1(_04225_),
    .A2(_04539_));
 sg13g2_nor2_1 _22200_ (.A(_04542_),
    .B(_04543_),
    .Y(_04544_));
 sg13g2_a21oi_1 _22201_ (.A1(net155),
    .A2(_11760_),
    .Y(_04545_),
    .B1(_04544_));
 sg13g2_nand2_1 _22202_ (.Y(_04546_),
    .A(_04136_),
    .B(_04545_));
 sg13g2_nand4_1 _22203_ (.B(_04510_),
    .C(_04511_),
    .A(_04509_),
    .Y(_00990_),
    .D(_04546_));
 sg13g2_mux2_1 _22204_ (.A0(net1043),
    .A1(net1057),
    .S(_03622_),
    .X(_04547_));
 sg13g2_o21ai_1 _22205_ (.B1(_03606_),
    .Y(_04548_),
    .A1(net1045),
    .A2(_04547_));
 sg13g2_o21ai_1 _22206_ (.B1(net139),
    .Y(_04549_),
    .A1(_11528_),
    .A2(net138));
 sg13g2_nor2_1 _22207_ (.A(net158),
    .B(net156),
    .Y(_04550_));
 sg13g2_nor3_1 _22208_ (.A(_04057_),
    .B(_04549_),
    .C(_04550_),
    .Y(_04551_));
 sg13g2_o21ai_1 _22209_ (.B1(_04551_),
    .Y(_04552_),
    .A1(net159),
    .A2(_04059_));
 sg13g2_nor2_1 _22210_ (.A(net1044),
    .B(_04483_),
    .Y(_04553_));
 sg13g2_a221oi_1 _22211_ (.B2(_04553_),
    .C1(_04125_),
    .B1(_04552_),
    .A1(net1058),
    .Y(_04554_),
    .A2(net145));
 sg13g2_and2_1 _22212_ (.A(_03516_),
    .B(_03525_),
    .X(_04555_));
 sg13g2_nand2_1 _22213_ (.Y(_04556_),
    .A(_03622_),
    .B(_03606_));
 sg13g2_xnor2_1 _22214_ (.Y(_04557_),
    .A(_04555_),
    .B(_04556_));
 sg13g2_a22oi_1 _22215_ (.Y(_04558_),
    .B1(net135),
    .B2(net192),
    .A2(_04080_),
    .A1(net196));
 sg13g2_o21ai_1 _22216_ (.B1(_04413_),
    .Y(_04559_),
    .A1(net160),
    .A2(_04066_));
 sg13g2_a221oi_1 _22217_ (.B2(_03478_),
    .C1(_04559_),
    .B1(_04256_),
    .A1(net142),
    .Y(_04560_),
    .A2(net140));
 sg13g2_a221oi_1 _22218_ (.B2(_11454_),
    .C1(_04195_),
    .B1(net134),
    .A1(net130),
    .Y(_04561_),
    .A2(net136));
 sg13g2_nand3_1 _22219_ (.B(_04560_),
    .C(_04561_),
    .A(_04558_),
    .Y(_04562_));
 sg13g2_o21ai_1 _22220_ (.B1(_03472_),
    .Y(_04563_),
    .A1(_04082_),
    .A2(_04513_));
 sg13g2_nand4_1 _22221_ (.B(_04560_),
    .C(_04561_),
    .A(_04558_),
    .Y(_04564_),
    .D(_04563_));
 sg13g2_a22oi_1 _22222_ (.Y(_04565_),
    .B1(_04564_),
    .B2(net1135),
    .A2(_04562_),
    .A1(net1046));
 sg13g2_a21oi_1 _22223_ (.A1(net194),
    .A2(_04097_),
    .Y(_04566_),
    .B1(_04565_));
 sg13g2_a21oi_1 _22224_ (.A1(_09120_),
    .A2(_04557_),
    .Y(_04567_),
    .B1(_04566_));
 sg13g2_o21ai_1 _22225_ (.B1(_03634_),
    .Y(_04568_),
    .A1(_04525_),
    .A2(_04540_));
 sg13g2_xor2_1 _22226_ (.B(_04568_),
    .A(_04556_),
    .X(_04569_));
 sg13g2_nand2_1 _22227_ (.Y(_04570_),
    .A(_04455_),
    .B(_04569_));
 sg13g2_nand4_1 _22228_ (.B(_04554_),
    .C(_04567_),
    .A(_04548_),
    .Y(_04571_),
    .D(_04570_));
 sg13g2_o21ai_1 _22229_ (.B1(_04571_),
    .Y(_04572_),
    .A1(_04149_),
    .A2(\cpu.ex.c_mult[5] ));
 sg13g2_nand2_1 _22230_ (.Y(_04573_),
    .A(net1127),
    .B(_04214_));
 sg13g2_xor2_1 _22231_ (.B(_04573_),
    .A(_11401_),
    .X(_04574_));
 sg13g2_a22oi_1 _22232_ (.Y(_04575_),
    .B1(_04574_),
    .B2(net64),
    .A2(net32),
    .A1(_08806_));
 sg13g2_o21ai_1 _22233_ (.B1(_04575_),
    .Y(_00991_),
    .A1(net65),
    .A2(_04572_));
 sg13g2_nand2_1 _22234_ (.Y(_04576_),
    .A(_03595_),
    .B(_04095_));
 sg13g2_a22oi_1 _22235_ (.Y(_04577_),
    .B1(_04256_),
    .B2(net196),
    .A2(_04088_),
    .A1(net192));
 sg13g2_a22oi_1 _22236_ (.Y(_04578_),
    .B1(net135),
    .B2(_03491_),
    .A2(net140),
    .A1(net130));
 sg13g2_nand3_1 _22237_ (.B(_04577_),
    .C(_04578_),
    .A(_04264_),
    .Y(_04579_));
 sg13g2_nor2_1 _22238_ (.A(net161),
    .B(_04056_),
    .Y(_04580_));
 sg13g2_a21oi_1 _22239_ (.A1(_03479_),
    .A2(net136),
    .Y(_04581_),
    .B1(_04580_));
 sg13g2_nand2b_1 _22240_ (.Y(_04582_),
    .B(_04581_),
    .A_N(_04358_));
 sg13g2_nor2_1 _22241_ (.A(_04082_),
    .B(_04513_),
    .Y(_04583_));
 sg13g2_a21oi_1 _22242_ (.A1(_04251_),
    .A2(_04583_),
    .Y(_04584_),
    .B1(_03684_));
 sg13g2_nor3_1 _22243_ (.A(_04579_),
    .B(_04582_),
    .C(_04584_),
    .Y(_04585_));
 sg13g2_o21ai_1 _22244_ (.B1(net1046),
    .Y(_04586_),
    .A1(_04579_),
    .A2(_04582_));
 sg13g2_o21ai_1 _22245_ (.B1(_04586_),
    .Y(_04587_),
    .A1(_08373_),
    .A2(_04585_));
 sg13g2_inv_1 _22246_ (.Y(_04588_),
    .A(_03533_));
 sg13g2_a21oi_1 _22247_ (.A1(_04555_),
    .A2(_04588_),
    .Y(_04589_),
    .B1(_03538_));
 sg13g2_nand2_1 _22248_ (.Y(_04590_),
    .A(_03640_),
    .B(_03643_));
 sg13g2_xor2_1 _22249_ (.B(_04590_),
    .A(_04589_),
    .X(_04591_));
 sg13g2_nor2_1 _22250_ (.A(_04093_),
    .B(_04067_),
    .Y(_04592_));
 sg13g2_nand2_1 _22251_ (.Y(_04593_),
    .A(net216),
    .B(_04167_));
 sg13g2_o21ai_1 _22252_ (.B1(_04593_),
    .Y(_04594_),
    .A1(_11528_),
    .A2(net156));
 sg13g2_o21ai_1 _22253_ (.B1(net139),
    .Y(_04595_),
    .A1(_04106_),
    .A2(_04053_));
 sg13g2_or4_1 _22254_ (.A(_04439_),
    .B(_04592_),
    .C(_04594_),
    .D(_04595_),
    .X(_04596_));
 sg13g2_nand3_1 _22255_ (.B(_04512_),
    .C(_04596_),
    .A(net1118),
    .Y(_04597_));
 sg13g2_mux2_1 _22256_ (.A0(net1043),
    .A1(net1057),
    .S(_03640_),
    .X(_04598_));
 sg13g2_o21ai_1 _22257_ (.B1(_03643_),
    .Y(_04599_),
    .A1(net1045),
    .A2(_04598_));
 sg13g2_a21oi_1 _22258_ (.A1(net1058),
    .A2(_11954_),
    .Y(_04600_),
    .B1(_04125_));
 sg13g2_nand3_1 _22259_ (.B(_04599_),
    .C(_04600_),
    .A(_04597_),
    .Y(_04601_));
 sg13g2_a221oi_1 _22260_ (.B2(net877),
    .C1(_04601_),
    .B1(_04591_),
    .A1(_04576_),
    .Y(_04602_),
    .A2(_04587_));
 sg13g2_a21oi_1 _22261_ (.A1(_03622_),
    .A2(_04568_),
    .Y(_04603_),
    .B1(_03607_));
 sg13g2_xnor2_1 _22262_ (.Y(_04604_),
    .A(_04590_),
    .B(_04603_));
 sg13g2_nand2_1 _22263_ (.Y(_04605_),
    .A(_04455_),
    .B(_04604_));
 sg13g2_a22oi_1 _22264_ (.Y(_04606_),
    .B1(_04602_),
    .B2(_04605_),
    .A2(_11790_),
    .A1(_04274_));
 sg13g2_inv_1 _22265_ (.Y(_04607_),
    .A(_04606_));
 sg13g2_xnor2_1 _22266_ (.Y(_04608_),
    .A(_11407_),
    .B(_04215_));
 sg13g2_a22oi_1 _22267_ (.Y(_04609_),
    .B1(_04608_),
    .B2(_04223_),
    .A2(net32),
    .A1(\cpu.ex.pc[6] ));
 sg13g2_o21ai_1 _22268_ (.B1(_04609_),
    .Y(_00992_),
    .A1(net65),
    .A2(_04607_));
 sg13g2_nand2_1 _22269_ (.Y(_04610_),
    .A(net161),
    .B(net99));
 sg13g2_a22oi_1 _22270_ (.Y(_04611_),
    .B1(net135),
    .B2(net130),
    .A2(net140),
    .A1(net131));
 sg13g2_a221oi_1 _22271_ (.B2(net129),
    .C1(_04418_),
    .B1(_04088_),
    .A1(_03566_),
    .Y(_04612_),
    .A2(net134));
 sg13g2_nand3_1 _22272_ (.B(_04611_),
    .C(_04612_),
    .A(_04312_),
    .Y(_04613_));
 sg13g2_a21oi_1 _22273_ (.A1(net164),
    .A2(net136),
    .Y(_04614_),
    .B1(_04613_));
 sg13g2_a21oi_1 _22274_ (.A1(_08372_),
    .A2(_04613_),
    .Y(_04615_),
    .B1(net1046));
 sg13g2_o21ai_1 _22275_ (.B1(_04164_),
    .Y(_04616_),
    .A1(_04614_),
    .A2(_04615_));
 sg13g2_mux2_1 _22276_ (.A0(net1057),
    .A1(net1043),
    .S(_03642_),
    .X(_04617_));
 sg13g2_o21ai_1 _22277_ (.B1(_03596_),
    .Y(_04618_),
    .A1(net1045),
    .A2(_04617_));
 sg13g2_nor2_1 _22278_ (.A(net158),
    .B(_04185_),
    .Y(_04619_));
 sg13g2_nor2_1 _22279_ (.A(net266),
    .B(net138),
    .Y(_04620_));
 sg13g2_nor3_1 _22280_ (.A(_04063_),
    .B(_04619_),
    .C(_04620_),
    .Y(_04621_));
 sg13g2_nor2_1 _22281_ (.A(net159),
    .B(net156),
    .Y(_04622_));
 sg13g2_a21oi_1 _22282_ (.A1(net126),
    .A2(net135),
    .Y(_04623_),
    .B1(_04622_));
 sg13g2_nand3_1 _22283_ (.B(_04621_),
    .C(_04623_),
    .A(_04474_),
    .Y(_04624_));
 sg13g2_a21oi_1 _22284_ (.A1(net194),
    .A2(net99),
    .Y(_04625_),
    .B1(net1044));
 sg13g2_a221oi_1 _22285_ (.B2(_04625_),
    .C1(_04125_),
    .B1(_04624_),
    .A1(_09157_),
    .Y(_04626_),
    .A2(_10461_));
 sg13g2_nand2_1 _22286_ (.Y(_04627_),
    .A(_04618_),
    .B(_04626_));
 sg13g2_a221oi_1 _22287_ (.B2(_04616_),
    .C1(_04627_),
    .B1(_04610_),
    .A1(_04159_),
    .Y(_04628_),
    .A2(_04455_));
 sg13g2_a21o_1 _22288_ (.A2(_04589_),
    .A1(_03536_),
    .B1(_03530_),
    .X(_04629_));
 sg13g2_xor2_1 _22289_ (.B(_04158_),
    .A(_04629_),
    .X(_04630_));
 sg13g2_nand2_1 _22290_ (.Y(_04631_),
    .A(_03586_),
    .B(_04630_));
 sg13g2_nor2_1 _22291_ (.A(net157),
    .B(\cpu.ex.c_mult[7] ),
    .Y(_04632_));
 sg13g2_a21oi_1 _22292_ (.A1(_04628_),
    .A2(_04631_),
    .Y(_04633_),
    .B1(_04632_));
 sg13g2_inv_1 _22293_ (.Y(_04634_),
    .A(_04633_));
 sg13g2_xnor2_1 _22294_ (.Y(_04635_),
    .A(_11430_),
    .B(_04216_));
 sg13g2_a22oi_1 _22295_ (.Y(_04636_),
    .B1(_04635_),
    .B2(net64),
    .A2(net32),
    .A1(_08777_));
 sg13g2_o21ai_1 _22296_ (.B1(_04636_),
    .Y(_00993_),
    .A1(net65),
    .A2(_04634_));
 sg13g2_nor3_1 _22297_ (.A(_11454_),
    .B(_03547_),
    .C(_03549_),
    .Y(_04637_));
 sg13g2_or3_1 _22298_ (.A(_04637_),
    .B(_03535_),
    .C(_03540_),
    .X(_04638_));
 sg13g2_nor2_1 _22299_ (.A(_10753_),
    .B(net161),
    .Y(_04639_));
 sg13g2_nand2_1 _22300_ (.Y(_04640_),
    .A(_10753_),
    .B(net161));
 sg13g2_nand2b_1 _22301_ (.Y(_04641_),
    .B(_04640_),
    .A_N(_04639_));
 sg13g2_xnor2_1 _22302_ (.Y(_04642_),
    .A(_04638_),
    .B(_04641_));
 sg13g2_nand2_1 _22303_ (.Y(_04643_),
    .A(_03586_),
    .B(_04642_));
 sg13g2_a21oi_1 _22304_ (.A1(_09997_),
    .A2(_04159_),
    .Y(_04644_),
    .B1(net589));
 sg13g2_a22oi_1 _22305_ (.Y(_04645_),
    .B1(_04306_),
    .B2(_03492_),
    .A2(net135),
    .A1(net131));
 sg13g2_a21oi_1 _22306_ (.A1(net196),
    .A2(net140),
    .Y(_04646_),
    .B1(net111));
 sg13g2_a221oi_1 _22307_ (.B2(_03485_),
    .C1(_04249_),
    .B1(_04088_),
    .A1(_03569_),
    .Y(_04647_),
    .A2(net137));
 sg13g2_nand4_1 _22308_ (.B(_04645_),
    .C(_04646_),
    .A(_04164_),
    .Y(_04648_),
    .D(_04647_));
 sg13g2_a21oi_1 _22309_ (.A1(_04076_),
    .A2(_04096_),
    .Y(_04649_),
    .B1(_04099_));
 sg13g2_nor2_1 _22310_ (.A(_03529_),
    .B(_04056_),
    .Y(_04650_));
 sg13g2_nor2_1 _22311_ (.A(_03507_),
    .B(_04067_),
    .Y(_04651_));
 sg13g2_nand2_1 _22312_ (.Y(_04652_),
    .A(_04191_),
    .B(_04036_));
 sg13g2_o21ai_1 _22313_ (.B1(_04652_),
    .Y(_04653_),
    .A1(net190),
    .A2(_04078_));
 sg13g2_a21oi_1 _22314_ (.A1(net216),
    .A2(_04088_),
    .Y(_04654_),
    .B1(_04446_));
 sg13g2_o21ai_1 _22315_ (.B1(_04654_),
    .Y(_04655_),
    .A1(_03510_),
    .A2(_04053_));
 sg13g2_nor4_1 _22316_ (.A(_04650_),
    .B(_04651_),
    .C(_04653_),
    .D(_04655_),
    .Y(_04656_));
 sg13g2_nand2_1 _22317_ (.Y(_04657_),
    .A(net1118),
    .B(_04576_));
 sg13g2_mux2_1 _22318_ (.A0(_09262_),
    .A1(_10036_),
    .S(_04639_),
    .X(_04658_));
 sg13g2_o21ai_1 _22319_ (.B1(_04640_),
    .Y(_04659_),
    .A1(_10019_),
    .A2(_04658_));
 sg13g2_o21ai_1 _22320_ (.B1(_04659_),
    .Y(_04660_),
    .A1(_04656_),
    .A2(_04657_));
 sg13g2_a221oi_1 _22321_ (.B2(_04649_),
    .C1(_04660_),
    .B1(_04648_),
    .A1(net1058),
    .Y(_04661_),
    .A2(_11660_));
 sg13g2_and2_1 _22322_ (.A(_04644_),
    .B(_04661_),
    .X(_04662_));
 sg13g2_o21ai_1 _22323_ (.B1(net218),
    .Y(_04663_),
    .A1(net276),
    .A2(_04157_));
 sg13g2_nand2_1 _22324_ (.Y(_04664_),
    .A(net276),
    .B(_04157_));
 sg13g2_nand2_1 _22325_ (.Y(_04665_),
    .A(_04663_),
    .B(_04664_));
 sg13g2_xnor2_1 _22326_ (.Y(_04666_),
    .A(_04641_),
    .B(_04665_));
 sg13g2_a221oi_1 _22327_ (.B2(_04225_),
    .C1(net155),
    .B1(_04666_),
    .A1(_04643_),
    .Y(_04667_),
    .A2(_04662_));
 sg13g2_a21o_1 _22328_ (.A2(\cpu.ex.c_mult[8] ),
    .A1(_04274_),
    .B1(_04667_),
    .X(_04668_));
 sg13g2_inv_1 _22329_ (.Y(_04669_),
    .A(_04668_));
 sg13g2_xor2_1 _22330_ (.B(_04218_),
    .A(_11317_),
    .X(_04670_));
 sg13g2_a22oi_1 _22331_ (.Y(_04671_),
    .B1(_04670_),
    .B2(net64),
    .A2(_04146_),
    .A1(_08757_));
 sg13g2_o21ai_1 _22332_ (.B1(_04671_),
    .Y(_00994_),
    .A1(_04031_),
    .A2(_04669_));
 sg13g2_nor2_1 _22333_ (.A(net172),
    .B(net160),
    .Y(_04672_));
 sg13g2_nand2_1 _22334_ (.Y(_04673_),
    .A(net172),
    .B(net160));
 sg13g2_nand2b_1 _22335_ (.Y(_04674_),
    .B(_04673_),
    .A_N(_04672_));
 sg13g2_xor2_1 _22336_ (.B(_04674_),
    .A(_03660_),
    .X(_04675_));
 sg13g2_nand2_1 _22337_ (.Y(_04676_),
    .A(net201),
    .B(net161));
 sg13g2_nand3_1 _22338_ (.B(_03545_),
    .C(_03551_),
    .A(_04676_),
    .Y(_04677_));
 sg13g2_xnor2_1 _22339_ (.Y(_04678_),
    .A(_04677_),
    .B(_04674_));
 sg13g2_nand2_1 _22340_ (.Y(_04679_),
    .A(net877),
    .B(_04678_));
 sg13g2_o21ai_1 _22341_ (.B1(_04304_),
    .Y(_04680_),
    .A1(net128),
    .A2(net138));
 sg13g2_a221oi_1 _22342_ (.B2(net131),
    .C1(_04680_),
    .B1(_04088_),
    .A1(net164),
    .Y(_04681_),
    .A2(net135));
 sg13g2_a21oi_1 _22343_ (.A1(_04411_),
    .A2(_04681_),
    .Y(_04682_),
    .B1(_04099_));
 sg13g2_o21ai_1 _22344_ (.B1(_04164_),
    .Y(_04683_),
    .A1(_04185_),
    .A2(_04355_));
 sg13g2_o21ai_1 _22345_ (.B1(_04198_),
    .Y(_04684_),
    .A1(_04682_),
    .A2(_04683_));
 sg13g2_nand2_1 _22346_ (.Y(_04685_),
    .A(_10037_),
    .B(_04672_));
 sg13g2_o21ai_1 _22347_ (.B1(_09262_),
    .Y(_04686_),
    .A1(_11829_),
    .A2(net160));
 sg13g2_nand3_1 _22348_ (.B(_04685_),
    .C(_04686_),
    .A(_04202_),
    .Y(_04687_));
 sg13g2_nand2b_1 _22349_ (.Y(_04688_),
    .B(_04035_),
    .A_N(_03510_));
 sg13g2_o21ai_1 _22350_ (.B1(_04688_),
    .Y(_04689_),
    .A1(_03507_),
    .A2(net156));
 sg13g2_a221oi_1 _22351_ (.B2(net216),
    .C1(_04689_),
    .B1(_04180_),
    .A1(_04191_),
    .Y(_04690_),
    .A2(_04178_));
 sg13g2_nor2b_1 _22352_ (.A(_04477_),
    .B_N(_04690_),
    .Y(_04691_));
 sg13g2_nor2_1 _22353_ (.A(_04106_),
    .B(_04074_),
    .Y(_04692_));
 sg13g2_a221oi_1 _22354_ (.B2(_03537_),
    .C1(_04692_),
    .B1(_04306_),
    .A1(_11454_),
    .Y(_04693_),
    .A2(_04194_));
 sg13g2_a221oi_1 _22355_ (.B2(_04693_),
    .C1(net1044),
    .B1(_04691_),
    .A1(_04032_),
    .Y(_04694_),
    .A2(net99));
 sg13g2_a221oi_1 _22356_ (.B2(_04687_),
    .C1(_04694_),
    .B1(_04673_),
    .A1(_09157_),
    .Y(_04695_),
    .A2(_03503_));
 sg13g2_nand4_1 _22357_ (.B(_04679_),
    .C(_04684_),
    .A(_04644_),
    .Y(_04696_),
    .D(_04695_));
 sg13g2_o21ai_1 _22358_ (.B1(_04696_),
    .Y(_04697_),
    .A1(_04150_),
    .A2(_04675_));
 sg13g2_nor2_1 _22359_ (.A(net157),
    .B(\cpu.ex.c_mult[9] ),
    .Y(_04698_));
 sg13g2_a21oi_1 _22360_ (.A1(_04149_),
    .A2(_04697_),
    .Y(_04699_),
    .B1(_04698_));
 sg13g2_nand2_1 _22361_ (.Y(_04700_),
    .A(_04136_),
    .B(_04699_));
 sg13g2_xnor2_1 _22362_ (.Y(_04701_),
    .A(_11316_),
    .B(_04219_));
 sg13g2_a22oi_1 _22363_ (.Y(_04702_),
    .B1(_04701_),
    .B2(_04223_),
    .A2(_04147_),
    .A1(_08738_));
 sg13g2_nand2_1 _22364_ (.Y(_00995_),
    .A(_04700_),
    .B(_04702_));
 sg13g2_inv_1 _22365_ (.Y(_04703_),
    .A(_04236_));
 sg13g2_and2_1 _22366_ (.A(_04229_),
    .B(_04703_),
    .X(_04704_));
 sg13g2_xnor2_1 _22367_ (.Y(_04705_),
    .A(_04235_),
    .B(_04704_));
 sg13g2_nor2_1 _22368_ (.A(_11829_),
    .B(net141),
    .Y(_04706_));
 sg13g2_a21oi_1 _22369_ (.A1(_04677_),
    .A2(_03563_),
    .Y(_04707_),
    .B1(_04706_));
 sg13g2_xnor2_1 _22370_ (.Y(_04708_),
    .A(_04707_),
    .B(_04704_));
 sg13g2_a21oi_1 _22371_ (.A1(net131),
    .A2(_04306_),
    .Y(_04709_),
    .B1(net111));
 sg13g2_a22oi_1 _22372_ (.Y(_04710_),
    .B1(_04088_),
    .B2(_03473_),
    .A2(net137),
    .A1(net130));
 sg13g2_nand3_1 _22373_ (.B(_04709_),
    .C(_04710_),
    .A(_04363_),
    .Y(_04711_));
 sg13g2_nand2b_1 _22374_ (.Y(_04712_),
    .B(_04711_),
    .A_N(_04099_));
 sg13g2_o21ai_1 _22375_ (.B1(_04162_),
    .Y(_04713_),
    .A1(net140),
    .A2(net135));
 sg13g2_nand3_1 _22376_ (.B(_04712_),
    .C(_04713_),
    .A(_04164_),
    .Y(_04714_));
 sg13g2_nand2_1 _22377_ (.Y(_04715_),
    .A(_04266_),
    .B(_04714_));
 sg13g2_a22oi_1 _22378_ (.Y(_04716_),
    .B1(net125),
    .B2(net126),
    .A2(net140),
    .A1(net216));
 sg13g2_nor2_1 _22379_ (.A(_04445_),
    .B(_04580_),
    .Y(_04717_));
 sg13g2_nor2_1 _22380_ (.A(_03532_),
    .B(net156),
    .Y(_04718_));
 sg13g2_nand2_1 _22381_ (.Y(_04719_),
    .A(_11382_),
    .B(_04180_));
 sg13g2_o21ai_1 _22382_ (.B1(_04719_),
    .Y(_04720_),
    .A1(net159),
    .A2(_04078_));
 sg13g2_nor2_1 _22383_ (.A(net158),
    .B(_04251_),
    .Y(_04721_));
 sg13g2_nor4_1 _22384_ (.A(_04517_),
    .B(_04718_),
    .C(_04720_),
    .D(_04721_),
    .Y(_04722_));
 sg13g2_nand3_1 _22385_ (.B(_04717_),
    .C(_04722_),
    .A(_04716_),
    .Y(_04723_));
 sg13g2_a21oi_1 _22386_ (.A1(net160),
    .A2(net99),
    .Y(_04724_),
    .B1(_10024_));
 sg13g2_mux2_1 _22387_ (.A0(net1125),
    .A1(net1117),
    .S(_04236_),
    .X(_04725_));
 sg13g2_o21ai_1 _22388_ (.B1(_04229_),
    .Y(_04726_),
    .A1(net1045),
    .A2(_04725_));
 sg13g2_o21ai_1 _22389_ (.B1(_04726_),
    .Y(_04727_),
    .A1(_04373_),
    .A2(net265));
 sg13g2_a21oi_1 _22390_ (.A1(_04723_),
    .A2(_04724_),
    .Y(_04728_),
    .B1(_04727_));
 sg13g2_nand3_1 _22391_ (.B(_04715_),
    .C(_04728_),
    .A(_04161_),
    .Y(_04729_));
 sg13g2_a221oi_1 _22392_ (.B2(net877),
    .C1(_04729_),
    .B1(_04708_),
    .A1(net589),
    .Y(_04730_),
    .A2(_04705_));
 sg13g2_a21o_1 _22393_ (.A2(_11855_),
    .A1(net155),
    .B1(_04730_),
    .X(_04731_));
 sg13g2_buf_1 _22394_ (.A(_08791_),
    .X(_04732_));
 sg13g2_nand2_1 _22395_ (.Y(_04733_),
    .A(_08738_),
    .B(_04219_));
 sg13g2_xnor2_1 _22396_ (.Y(_04734_),
    .A(_11292_),
    .B(_04733_));
 sg13g2_a22oi_1 _22397_ (.Y(_04735_),
    .B1(_04734_),
    .B2(_04135_),
    .A2(_04146_),
    .A1(net978));
 sg13g2_o21ai_1 _22398_ (.B1(_04735_),
    .Y(_00996_),
    .A1(_04031_),
    .A2(_04731_));
 sg13g2_mux2_1 _22399_ (.A0(\cpu.dec.r_set_cc ),
    .A1(_10359_),
    .S(_03583_),
    .X(_00999_));
 sg13g2_buf_1 _22400_ (.A(_00256_),
    .X(_04736_));
 sg13g2_nor4_1 _22401_ (.A(net1112),
    .B(net1111),
    .C(_04736_),
    .D(_03421_),
    .Y(_04737_));
 sg13g2_buf_2 _22402_ (.A(_04737_),
    .X(_04738_));
 sg13g2_buf_1 _22403_ (.A(_04738_),
    .X(_04739_));
 sg13g2_mux2_1 _22404_ (.A0(_10772_),
    .A1(_03431_),
    .S(net588),
    .X(_01000_));
 sg13g2_mux2_1 _22405_ (.A0(_10664_),
    .A1(net878),
    .S(net588),
    .X(_01001_));
 sg13g2_mux2_1 _22406_ (.A0(_10500_),
    .A1(net601),
    .S(net588),
    .X(_01002_));
 sg13g2_mux2_1 _22407_ (.A0(_10545_),
    .A1(_03428_),
    .S(net588),
    .X(_01003_));
 sg13g2_mux2_1 _22408_ (.A0(_10599_),
    .A1(net525),
    .S(net588),
    .X(_01004_));
 sg13g2_mux2_1 _22409_ (.A0(_10449_),
    .A1(net743),
    .S(net588),
    .X(_01005_));
 sg13g2_mux2_1 _22410_ (.A0(_10825_),
    .A1(net434),
    .S(net588),
    .X(_01006_));
 sg13g2_mux2_1 _22411_ (.A0(_10918_),
    .A1(_03434_),
    .S(_04739_),
    .X(_01007_));
 sg13g2_mux2_1 _22412_ (.A0(_10894_),
    .A1(net474),
    .S(_04739_),
    .X(_01008_));
 sg13g2_mux2_1 _22413_ (.A0(_10859_),
    .A1(net521),
    .S(net588),
    .X(_01009_));
 sg13g2_mux2_1 _22414_ (.A0(_10992_),
    .A1(_02995_),
    .S(_04738_),
    .X(_01010_));
 sg13g2_buf_1 _22415_ (.A(net983),
    .X(_04740_));
 sg13g2_mux2_1 _22416_ (.A0(_11021_),
    .A1(_04740_),
    .S(_04738_),
    .X(_01011_));
 sg13g2_buf_1 _22417_ (.A(net887),
    .X(_04741_));
 sg13g2_mux2_1 _22418_ (.A0(_10727_),
    .A1(_04741_),
    .S(_04738_),
    .X(_01012_));
 sg13g2_mux2_1 _22419_ (.A0(_10706_),
    .A1(net879),
    .S(_04738_),
    .X(_01013_));
 sg13g2_buf_1 _22420_ (.A(net982),
    .X(_04742_));
 sg13g2_mux2_1 _22421_ (.A0(_10633_),
    .A1(_04742_),
    .S(_04738_),
    .X(_01014_));
 sg13g2_or2_1 _22422_ (.X(_04743_),
    .B(_03421_),
    .A(_10356_));
 sg13g2_buf_1 _22423_ (.A(_04743_),
    .X(_04744_));
 sg13g2_buf_1 _22424_ (.A(_04744_),
    .X(_04745_));
 sg13g2_nor2b_1 _22425_ (.A(_04736_),
    .B_N(net955),
    .Y(_04746_));
 sg13g2_nand2_1 _22426_ (.Y(_04747_),
    .A(net744),
    .B(_04746_));
 sg13g2_and2_1 _22427_ (.A(net955),
    .B(net1111),
    .X(_04748_));
 sg13g2_a21oi_1 _22428_ (.A1(_10354_),
    .A2(\cpu.ex.r_wb_swapsp ),
    .Y(_04749_),
    .B1(_04748_));
 sg13g2_or4_1 _22429_ (.A(net1112),
    .B(_04736_),
    .C(_03421_),
    .D(_04749_),
    .X(_04750_));
 sg13g2_buf_1 _22430_ (.A(_04750_),
    .X(_04751_));
 sg13g2_buf_1 _22431_ (.A(net517),
    .X(_04752_));
 sg13g2_nand2_1 _22432_ (.Y(_04753_),
    .A(\cpu.ex.r_stmp[0] ),
    .B(net471));
 sg13g2_o21ai_1 _22433_ (.B1(_04753_),
    .Y(_01015_),
    .A1(net518),
    .A2(_04747_));
 sg13g2_buf_1 _22434_ (.A(net587),
    .X(_04754_));
 sg13g2_mux2_1 _22435_ (.A0(net1107),
    .A1(_10633_),
    .S(net516),
    .X(_04755_));
 sg13g2_mux2_1 _22436_ (.A0(_04755_),
    .A1(\cpu.ex.r_stmp[10] ),
    .S(net471),
    .X(_01016_));
 sg13g2_buf_1 _22437_ (.A(net517),
    .X(_04756_));
 sg13g2_nor2_1 _22438_ (.A(_02962_),
    .B(net516),
    .Y(_04757_));
 sg13g2_a21oi_1 _22439_ (.A1(_10664_),
    .A2(net518),
    .Y(_04758_),
    .B1(_04757_));
 sg13g2_nand2_1 _22440_ (.Y(_04759_),
    .A(\cpu.ex.r_stmp[11] ),
    .B(net471));
 sg13g2_o21ai_1 _22441_ (.B1(_04759_),
    .Y(_01017_),
    .A1(net470),
    .A2(_04758_));
 sg13g2_nor2_1 _22442_ (.A(_03694_),
    .B(net516),
    .Y(_04760_));
 sg13g2_a21oi_1 _22443_ (.A1(_10500_),
    .A2(net518),
    .Y(_04761_),
    .B1(_04760_));
 sg13g2_nand2_1 _22444_ (.Y(_04762_),
    .A(\cpu.ex.r_stmp[12] ),
    .B(net471));
 sg13g2_o21ai_1 _22445_ (.B1(_04762_),
    .Y(_01018_),
    .A1(net470),
    .A2(_04761_));
 sg13g2_nor2_1 _22446_ (.A(_03697_),
    .B(net516),
    .Y(_04763_));
 sg13g2_a21oi_1 _22447_ (.A1(_10545_),
    .A2(net518),
    .Y(_04764_),
    .B1(_04763_));
 sg13g2_nand2_1 _22448_ (.Y(_04765_),
    .A(\cpu.ex.r_stmp[13] ),
    .B(net471));
 sg13g2_o21ai_1 _22449_ (.B1(_04765_),
    .Y(_01019_),
    .A1(net470),
    .A2(_04764_));
 sg13g2_nor2_1 _22450_ (.A(_03700_),
    .B(net516),
    .Y(_04766_));
 sg13g2_a21oi_1 _22451_ (.A1(_10599_),
    .A2(net518),
    .Y(_04767_),
    .B1(_04766_));
 sg13g2_nand2_1 _22452_ (.Y(_04768_),
    .A(\cpu.ex.r_stmp[14] ),
    .B(net471));
 sg13g2_o21ai_1 _22453_ (.B1(_04768_),
    .Y(_01020_),
    .A1(net470),
    .A2(_04767_));
 sg13g2_nor2_1 _22454_ (.A(net670),
    .B(net516),
    .Y(_04769_));
 sg13g2_a21oi_1 _22455_ (.A1(_10449_),
    .A2(net518),
    .Y(_04770_),
    .B1(_04769_));
 sg13g2_nand2_1 _22456_ (.Y(_04771_),
    .A(\cpu.ex.r_stmp[15] ),
    .B(net517));
 sg13g2_o21ai_1 _22457_ (.B1(_04771_),
    .Y(_01021_),
    .A1(net470),
    .A2(_04770_));
 sg13g2_nor2_1 _22458_ (.A(net620),
    .B(net587),
    .Y(_04772_));
 sg13g2_a21oi_1 _22459_ (.A1(_10772_),
    .A2(net518),
    .Y(_04773_),
    .B1(_04772_));
 sg13g2_nand2_1 _22460_ (.Y(_04774_),
    .A(\cpu.ex.r_stmp[1] ),
    .B(net517));
 sg13g2_o21ai_1 _22461_ (.B1(_04774_),
    .Y(_01022_),
    .A1(net470),
    .A2(_04773_));
 sg13g2_nor2_1 _22462_ (.A(_09349_),
    .B(net587),
    .Y(_04775_));
 sg13g2_a21oi_1 _22463_ (.A1(_10825_),
    .A2(net518),
    .Y(_04776_),
    .B1(_04775_));
 sg13g2_nand2_1 _22464_ (.Y(_04777_),
    .A(\cpu.ex.r_stmp[2] ),
    .B(net517));
 sg13g2_o21ai_1 _22465_ (.B1(_04777_),
    .Y(_01023_),
    .A1(net470),
    .A2(_04776_));
 sg13g2_nor2_1 _22466_ (.A(_12656_),
    .B(net587),
    .Y(_04778_));
 sg13g2_a21oi_1 _22467_ (.A1(_10918_),
    .A2(_04745_),
    .Y(_04779_),
    .B1(_04778_));
 sg13g2_nand2_1 _22468_ (.Y(_04780_),
    .A(\cpu.ex.r_stmp[3] ),
    .B(net517));
 sg13g2_o21ai_1 _22469_ (.B1(_04780_),
    .Y(_01024_),
    .A1(_04756_),
    .A2(_04779_));
 sg13g2_nor2_1 _22470_ (.A(net656),
    .B(net587),
    .Y(_04781_));
 sg13g2_a21oi_1 _22471_ (.A1(_10894_),
    .A2(_04745_),
    .Y(_04782_),
    .B1(_04781_));
 sg13g2_nand2_1 _22472_ (.Y(_04783_),
    .A(\cpu.ex.r_stmp[4] ),
    .B(_04751_));
 sg13g2_o21ai_1 _22473_ (.B1(_04783_),
    .Y(_01025_),
    .A1(_04756_),
    .A2(_04782_));
 sg13g2_nor2_1 _22474_ (.A(_11383_),
    .B(net587),
    .Y(_04784_));
 sg13g2_a21oi_1 _22475_ (.A1(_10859_),
    .A2(_04754_),
    .Y(_04785_),
    .B1(_04784_));
 sg13g2_nand2_1 _22476_ (.Y(_04786_),
    .A(\cpu.ex.r_stmp[5] ),
    .B(_04751_));
 sg13g2_o21ai_1 _22477_ (.B1(_04786_),
    .Y(_01026_),
    .A1(_04752_),
    .A2(_04785_));
 sg13g2_mux2_1 _22478_ (.A0(net984),
    .A1(_10992_),
    .S(net516),
    .X(_04787_));
 sg13g2_mux2_1 _22479_ (.A0(_04787_),
    .A1(\cpu.ex.r_stmp[6] ),
    .S(_04752_),
    .X(_01027_));
 sg13g2_mux2_1 _22480_ (.A0(net983),
    .A1(_11021_),
    .S(net587),
    .X(_04788_));
 sg13g2_nor2_1 _22481_ (.A(net517),
    .B(_04788_),
    .Y(_04789_));
 sg13g2_a21oi_1 _22482_ (.A1(_11444_),
    .A2(net470),
    .Y(_01028_),
    .B1(_04789_));
 sg13g2_mux2_1 _22483_ (.A0(net1056),
    .A1(_10727_),
    .S(_04754_),
    .X(_04790_));
 sg13g2_mux2_1 _22484_ (.A0(_04790_),
    .A1(\cpu.ex.r_stmp[8] ),
    .S(net471),
    .X(_01029_));
 sg13g2_nor2_1 _22485_ (.A(_02958_),
    .B(net587),
    .Y(_04791_));
 sg13g2_a21oi_1 _22486_ (.A1(_10706_),
    .A2(net516),
    .Y(_04792_),
    .B1(_04791_));
 sg13g2_nand2_1 _22487_ (.Y(_04793_),
    .A(\cpu.ex.r_stmp[9] ),
    .B(net517));
 sg13g2_o21ai_1 _22488_ (.B1(_04793_),
    .Y(_01030_),
    .A1(net471),
    .A2(_04792_));
 sg13g2_nand2_1 _22489_ (.Y(_04794_),
    .A(net196),
    .B(_04046_));
 sg13g2_o21ai_1 _22490_ (.B1(_04794_),
    .Y(_04795_),
    .A1(_03579_),
    .A2(net217));
 sg13g2_a21oi_1 _22491_ (.A1(_04045_),
    .A2(_04795_),
    .Y(_04796_),
    .B1(_04366_));
 sg13g2_a21oi_1 _22492_ (.A1(_03485_),
    .A2(_04367_),
    .Y(_04797_),
    .B1(_04248_));
 sg13g2_and4_1 _22493_ (.A(_04530_),
    .B(_04593_),
    .C(_04796_),
    .D(_04797_),
    .X(_04798_));
 sg13g2_a22oi_1 _22494_ (.Y(_04799_),
    .B1(_04082_),
    .B2(_03569_),
    .A2(_04310_),
    .A1(_03491_));
 sg13g2_o21ai_1 _22495_ (.B1(_04799_),
    .Y(_04800_),
    .A1(_04032_),
    .A2(_04078_));
 sg13g2_nand2_1 _22496_ (.Y(_04801_),
    .A(net141),
    .B(net125));
 sg13g2_o21ai_1 _22497_ (.B1(_04801_),
    .Y(_04802_),
    .A1(net163),
    .A2(_04251_));
 sg13g2_nor4_1 _22498_ (.A(_04651_),
    .B(_04718_),
    .C(_04800_),
    .D(_04802_),
    .Y(_04803_));
 sg13g2_a21oi_1 _22499_ (.A1(_04798_),
    .A2(_04803_),
    .Y(_04804_),
    .B1(_04099_));
 sg13g2_a21o_1 _22500_ (.A2(_04162_),
    .A1(_11643_),
    .B1(_04804_),
    .X(_04805_));
 sg13g2_o21ai_1 _22501_ (.B1(_04805_),
    .Y(_04806_),
    .A1(net126),
    .A2(_04062_));
 sg13g2_nor3_1 _22502_ (.A(_10037_),
    .B(_10984_),
    .C(net158),
    .Y(_04807_));
 sg13g2_nor4_1 _22503_ (.A(net1059),
    .B(_09263_),
    .C(_11660_),
    .D(_04455_),
    .Y(_04808_));
 sg13g2_o21ai_1 _22504_ (.B1(_04202_),
    .Y(_04809_),
    .A1(_04807_),
    .A2(_04808_));
 sg13g2_nor4_1 _22505_ (.A(net1059),
    .B(_09263_),
    .C(_10020_),
    .D(_04455_),
    .Y(_04810_));
 sg13g2_o21ai_1 _22506_ (.B1(net158),
    .Y(_04811_),
    .A1(_10984_),
    .A2(_04810_));
 sg13g2_a221oi_1 _22507_ (.B2(_04811_),
    .C1(net155),
    .B1(_04809_),
    .A1(net1058),
    .Y(_04812_),
    .A2(net201));
 sg13g2_and2_1 _22508_ (.A(_10368_),
    .B(net155),
    .X(_04813_));
 sg13g2_a22oi_1 _22509_ (.Y(_04814_),
    .B1(_04813_),
    .B2(_11668_),
    .A2(_04812_),
    .A1(_04806_));
 sg13g2_inv_1 _22510_ (.Y(_04815_),
    .A(_04814_));
 sg13g2_a21oi_1 _22511_ (.A1(_11678_),
    .A2(_11679_),
    .Y(_04816_),
    .B1(_11680_));
 sg13g2_buf_1 _22512_ (.A(_04816_),
    .X(_04817_));
 sg13g2_buf_1 _22513_ (.A(_04817_),
    .X(_04818_));
 sg13g2_nand2_1 _22514_ (.Y(_04819_),
    .A(_04025_),
    .B(_11688_));
 sg13g2_buf_1 _22515_ (.A(_04819_),
    .X(_04820_));
 sg13g2_nor2_1 _22516_ (.A(_04818_),
    .B(_04820_),
    .Y(_04821_));
 sg13g2_buf_1 _22517_ (.A(_04025_),
    .X(_04822_));
 sg13g2_a21oi_1 _22518_ (.A1(net215),
    .A2(net762),
    .Y(_04823_),
    .B1(net745));
 sg13g2_buf_1 _22519_ (.A(net101),
    .X(_04824_));
 sg13g2_nand2_1 _22520_ (.Y(_04825_),
    .A(net1053),
    .B(_11694_));
 sg13g2_buf_2 _22521_ (.A(_04825_),
    .X(_04826_));
 sg13g2_buf_1 _22522_ (.A(_04826_),
    .X(_04827_));
 sg13g2_buf_2 _22523_ (.A(net84),
    .X(_04828_));
 sg13g2_buf_1 _22524_ (.A(_04826_),
    .X(_04829_));
 sg13g2_buf_1 _22525_ (.A(net548),
    .X(_04830_));
 sg13g2_buf_1 _22526_ (.A(net469),
    .X(_04831_));
 sg13g2_mux2_1 _22527_ (.A0(\cpu.dcache.r_data[4][8] ),
    .A1(\cpu.dcache.r_data[6][8] ),
    .S(net551),
    .X(_04832_));
 sg13g2_a22oi_1 _22528_ (.Y(_04833_),
    .B1(_04832_),
    .B2(net806),
    .A2(_09625_),
    .A1(\cpu.dcache.r_data[5][8] ));
 sg13g2_nand2b_1 _22529_ (.Y(_04834_),
    .B(net785),
    .A_N(_04833_));
 sg13g2_buf_1 _22530_ (.A(net488),
    .X(_04835_));
 sg13g2_a22oi_1 _22531_ (.Y(_04836_),
    .B1(net545),
    .B2(\cpu.dcache.r_data[7][8] ),
    .A2(net432),
    .A1(\cpu.dcache.r_data[2][8] ));
 sg13g2_buf_1 _22532_ (.A(net530),
    .X(_04837_));
 sg13g2_a22oi_1 _22533_ (.Y(_04838_),
    .B1(net468),
    .B2(\cpu.dcache.r_data[3][8] ),
    .A2(net439),
    .A1(\cpu.dcache.r_data[1][8] ));
 sg13g2_and3_1 _22534_ (.X(_04839_),
    .A(_04834_),
    .B(_04836_),
    .C(_04838_));
 sg13g2_o21ai_1 _22535_ (.B1(_04839_),
    .Y(_04840_),
    .A1(_00312_),
    .A2(net433));
 sg13g2_a22oi_1 _22536_ (.Y(_04841_),
    .B1(net493),
    .B2(\cpu.dcache.r_data[4][24] ),
    .A2(net487),
    .A1(\cpu.dcache.r_data[3][24] ));
 sg13g2_nand2_1 _22537_ (.Y(_04842_),
    .A(\cpu.dcache.r_data[5][24] ),
    .B(_12782_));
 sg13g2_a22oi_1 _22538_ (.Y(_04843_),
    .B1(net485),
    .B2(\cpu.dcache.r_data[6][24] ),
    .A2(net438),
    .A1(\cpu.dcache.r_data[2][24] ));
 sg13g2_buf_1 _22539_ (.A(net489),
    .X(_04844_));
 sg13g2_nor2_1 _22540_ (.A(_00311_),
    .B(net469),
    .Y(_04845_));
 sg13g2_a221oi_1 _22541_ (.B2(\cpu.dcache.r_data[7][24] ),
    .C1(_04845_),
    .B1(net545),
    .A1(\cpu.dcache.r_data[1][24] ),
    .Y(_04846_),
    .A2(net431));
 sg13g2_nand4_1 _22542_ (.B(_04842_),
    .C(_04843_),
    .A(_04841_),
    .Y(_04847_),
    .D(_04846_));
 sg13g2_or3_1 _22543_ (.A(_04026_),
    .B(_08393_),
    .C(_08504_),
    .X(_04848_));
 sg13g2_buf_2 _22544_ (.A(_04848_),
    .X(_04849_));
 sg13g2_a221oi_1 _22545_ (.B2(_12152_),
    .C1(_04849_),
    .B1(_04847_),
    .A1(net682),
    .Y(_04850_),
    .A2(_04840_));
 sg13g2_nor3_1 _22546_ (.A(_04026_),
    .B(_08393_),
    .C(_08504_),
    .Y(_04851_));
 sg13g2_buf_1 _22547_ (.A(_04851_),
    .X(_04852_));
 sg13g2_mux2_1 _22548_ (.A0(\cpu.dcache.r_data[5][16] ),
    .A1(\cpu.dcache.r_data[7][16] ),
    .S(net551),
    .X(_04853_));
 sg13g2_a22oi_1 _22549_ (.Y(_04854_),
    .B1(_04853_),
    .B2(net619),
    .A2(_12447_),
    .A1(\cpu.dcache.r_data[6][16] ));
 sg13g2_nand2b_1 _22550_ (.Y(_04855_),
    .B(net785),
    .A_N(_04854_));
 sg13g2_a22oi_1 _22551_ (.Y(_04856_),
    .B1(_10235_),
    .B2(\cpu.dcache.r_data[4][16] ),
    .A2(_04844_),
    .A1(\cpu.dcache.r_data[1][16] ));
 sg13g2_a22oi_1 _22552_ (.Y(_04857_),
    .B1(_12459_),
    .B2(\cpu.dcache.r_data[2][16] ),
    .A2(_12570_),
    .A1(\cpu.dcache.r_data[3][16] ));
 sg13g2_nand3_1 _22553_ (.B(_04856_),
    .C(_04857_),
    .A(_04855_),
    .Y(_04858_));
 sg13g2_a21oi_2 _22554_ (.B1(_04858_),
    .Y(_04859_),
    .A2(net546),
    .A1(\cpu.dcache.r_data[0][16] ));
 sg13g2_o21ai_1 _22555_ (.B1(_12152_),
    .Y(_04860_),
    .A1(_10171_),
    .A2(_04859_));
 sg13g2_nor2_1 _22556_ (.A(_04852_),
    .B(_04860_),
    .Y(_04861_));
 sg13g2_nand2_1 _22557_ (.Y(_04862_),
    .A(_08502_),
    .B(net654));
 sg13g2_buf_2 _22558_ (.A(_04862_),
    .X(_04863_));
 sg13g2_o21ai_1 _22559_ (.B1(_04863_),
    .Y(_04864_),
    .A1(_04850_),
    .A2(_04861_));
 sg13g2_and2_1 _22560_ (.A(_08502_),
    .B(_04851_),
    .X(_04865_));
 sg13g2_buf_1 _22561_ (.A(_04865_),
    .X(_04866_));
 sg13g2_nand3_1 _22562_ (.B(_04866_),
    .C(_04859_),
    .A(net542),
    .Y(_04867_));
 sg13g2_buf_1 _22563_ (.A(net686),
    .X(_04868_));
 sg13g2_a22oi_1 _22564_ (.Y(_04869_),
    .B1(net603),
    .B2(\cpu.dcache.r_data[6][0] ),
    .A2(net604),
    .A1(\cpu.dcache.r_data[5][0] ));
 sg13g2_a22oi_1 _22565_ (.Y(_04870_),
    .B1(net488),
    .B2(\cpu.dcache.r_data[2][0] ),
    .A2(net530),
    .A1(\cpu.dcache.r_data[3][0] ));
 sg13g2_a22oi_1 _22566_ (.Y(_04871_),
    .B1(net621),
    .B2(\cpu.dcache.r_data[7][0] ),
    .A2(net544),
    .A1(\cpu.dcache.r_data[4][0] ));
 sg13g2_nand3_1 _22567_ (.B(_04870_),
    .C(_04871_),
    .A(_04869_),
    .Y(_04872_));
 sg13g2_nand2b_1 _22568_ (.Y(_04873_),
    .B(net586),
    .A_N(\cpu.dcache.r_data[0][0] ));
 sg13g2_o21ai_1 _22569_ (.B1(_04873_),
    .Y(_04874_),
    .A1(net586),
    .A2(_04872_));
 sg13g2_o21ai_1 _22570_ (.B1(net389),
    .Y(_04875_),
    .A1(\cpu.dcache.r_data[1][0] ),
    .A2(_04872_));
 sg13g2_o21ai_1 _22571_ (.B1(_04875_),
    .Y(_04876_),
    .A1(net389),
    .A2(_04874_));
 sg13g2_nand2_1 _22572_ (.Y(_04877_),
    .A(_12120_),
    .B(_04849_));
 sg13g2_o21ai_1 _22573_ (.B1(_04877_),
    .Y(_04878_),
    .A1(net618),
    .A2(_04863_));
 sg13g2_nand2b_1 _22574_ (.Y(_04879_),
    .B(_04878_),
    .A_N(_04876_));
 sg13g2_nand3_1 _22575_ (.B(_04867_),
    .C(_04879_),
    .A(_04864_),
    .Y(_04880_));
 sg13g2_nand2_2 _22576_ (.Y(_04881_),
    .A(net929),
    .B(net708));
 sg13g2_or2_1 _22577_ (.X(_04882_),
    .B(_04881_),
    .A(_10252_));
 sg13g2_buf_2 _22578_ (.A(_04882_),
    .X(_04883_));
 sg13g2_nor2_2 _22579_ (.A(net1042),
    .B(_04883_),
    .Y(_04884_));
 sg13g2_nor3_2 _22580_ (.A(net1042),
    .B(net1051),
    .C(_09831_),
    .Y(_04885_));
 sg13g2_inv_1 _22581_ (.Y(_04886_),
    .A(_09828_));
 sg13g2_buf_1 _22582_ (.A(_04886_),
    .X(_04887_));
 sg13g2_nand2_1 _22583_ (.Y(_04888_),
    .A(net922),
    .B(net872));
 sg13g2_nand2_1 _22584_ (.Y(_04889_),
    .A(net633),
    .B(_04888_));
 sg13g2_buf_1 _22585_ (.A(_00228_),
    .X(_04890_));
 sg13g2_nor2_1 _22586_ (.A(net681),
    .B(net1048),
    .Y(_04891_));
 sg13g2_nand2_1 _22587_ (.Y(_04892_),
    .A(net1120),
    .B(_04891_));
 sg13g2_o21ai_1 _22588_ (.B1(_04892_),
    .Y(_04893_),
    .A1(_09343_),
    .A2(_04890_));
 sg13g2_a21oi_1 _22589_ (.A1(_09527_),
    .A2(_09505_),
    .Y(_04894_),
    .B1(_09380_));
 sg13g2_a221oi_1 _22590_ (.B2(net1051),
    .C1(_04894_),
    .B1(_04893_),
    .A1(net806),
    .Y(_04895_),
    .A2(_04889_));
 sg13g2_nor3_1 _22591_ (.A(_04884_),
    .B(_04885_),
    .C(_04895_),
    .Y(_04896_));
 sg13g2_buf_2 _22592_ (.A(_04896_),
    .X(_04897_));
 sg13g2_and3_1 _22593_ (.X(_04898_),
    .A(_09322_),
    .B(_10116_),
    .C(_04890_));
 sg13g2_inv_1 _22594_ (.Y(_04899_),
    .A(\cpu.spi.r_ready ));
 sg13g2_nor3_1 _22595_ (.A(_10116_),
    .B(net437),
    .C(_04899_),
    .Y(_04900_));
 sg13g2_o21ai_1 _22596_ (.B1(net531),
    .Y(_04901_),
    .A1(_04898_),
    .A2(_04900_));
 sg13g2_nand2_1 _22597_ (.Y(_04902_),
    .A(net681),
    .B(net1051));
 sg13g2_buf_1 _22598_ (.A(_04902_),
    .X(_04903_));
 sg13g2_nor2_1 _22599_ (.A(net758),
    .B(_04903_),
    .Y(_04904_));
 sg13g2_buf_1 _22600_ (.A(_04904_),
    .X(_04905_));
 sg13g2_nor2_1 _22601_ (.A(_09353_),
    .B(_04881_),
    .Y(_04906_));
 sg13g2_buf_1 _22602_ (.A(_04906_),
    .X(_04907_));
 sg13g2_nand2_1 _22603_ (.Y(_04908_),
    .A(net899),
    .B(\cpu.spi.r_mode[2][0] ));
 sg13g2_o21ai_1 _22604_ (.B1(_04908_),
    .Y(_04909_),
    .A1(net899),
    .A2(_00224_));
 sg13g2_a22oi_1 _22605_ (.Y(_04910_),
    .B1(_04907_),
    .B2(_04909_),
    .A2(net430),
    .A1(\cpu.spi.r_timeout[0] ));
 sg13g2_inv_1 _22606_ (.Y(_04911_),
    .A(_00314_));
 sg13g2_buf_1 _22607_ (.A(_04884_),
    .X(_04912_));
 sg13g2_buf_1 _22608_ (.A(net1120),
    .X(_04913_));
 sg13g2_nor2_1 _22609_ (.A(_04913_),
    .B(_04883_),
    .Y(_04914_));
 sg13g2_buf_2 _22610_ (.A(_04914_),
    .X(_04915_));
 sg13g2_buf_1 _22611_ (.A(\cpu.spi.r_clk_count[2][0] ),
    .X(_04916_));
 sg13g2_a22oi_1 _22612_ (.Y(_04917_),
    .B1(_04915_),
    .B2(_04916_),
    .A2(net383),
    .A1(_04911_));
 sg13g2_nand3_1 _22613_ (.B(net1120),
    .C(net603),
    .A(net923),
    .Y(_04918_));
 sg13g2_buf_2 _22614_ (.A(_04918_),
    .X(_04919_));
 sg13g2_nor2_1 _22615_ (.A(_00313_),
    .B(_04919_),
    .Y(_04920_));
 sg13g2_a21oi_1 _22616_ (.A1(\cpu.spi.r_mode[1][0] ),
    .A2(_04885_),
    .Y(_04921_),
    .B1(_04920_));
 sg13g2_nand4_1 _22617_ (.B(_04910_),
    .C(_04917_),
    .A(_04901_),
    .Y(_04922_),
    .D(_04921_));
 sg13g2_a21oi_1 _22618_ (.A1(_09417_),
    .A2(_04897_),
    .Y(_04923_),
    .B1(_04922_));
 sg13g2_nor2_1 _22619_ (.A(net709),
    .B(_04923_),
    .Y(_04924_));
 sg13g2_nand2b_1 _22620_ (.Y(_04925_),
    .B(_10125_),
    .A_N(_09281_));
 sg13g2_buf_2 _22621_ (.A(_04925_),
    .X(_04926_));
 sg13g2_o21ai_1 _22622_ (.B1(net929),
    .Y(_04927_),
    .A1(net928),
    .A2(_09625_));
 sg13g2_buf_2 _22623_ (.A(_04927_),
    .X(_04928_));
 sg13g2_nor2_1 _22624_ (.A(_10252_),
    .B(_04881_),
    .Y(_04929_));
 sg13g2_buf_1 _22625_ (.A(_04929_),
    .X(_04930_));
 sg13g2_nor3_1 _22626_ (.A(net922),
    .B(net633),
    .C(_04903_),
    .Y(_04931_));
 sg13g2_buf_2 _22627_ (.A(_04931_),
    .X(_04932_));
 sg13g2_a22oi_1 _22628_ (.Y(_04933_),
    .B1(_04932_),
    .B2(\cpu.uart.r_x_invert ),
    .A2(_04930_),
    .A1(\cpu.uart.r_div_value[8] ));
 sg13g2_buf_1 _22629_ (.A(_04907_),
    .X(_04934_));
 sg13g2_nand2_1 _22630_ (.Y(_04935_),
    .A(_10173_),
    .B(_09351_));
 sg13g2_buf_2 _22631_ (.A(_04935_),
    .X(_04936_));
 sg13g2_nor3_1 _22632_ (.A(net1048),
    .B(net708),
    .C(_04936_),
    .Y(_04937_));
 sg13g2_buf_2 _22633_ (.A(_04937_),
    .X(_04938_));
 sg13g2_buf_1 _22634_ (.A(_04938_),
    .X(_04939_));
 sg13g2_a22oi_1 _22635_ (.Y(_04940_),
    .B1(net382),
    .B2(_09328_),
    .A2(net429),
    .A1(\cpu.uart.r_div_value[0] ));
 sg13g2_nand2_1 _22636_ (.Y(_04941_),
    .A(_04933_),
    .B(_04940_));
 sg13g2_a21oi_1 _22637_ (.A1(\cpu.uart.r_in[0] ),
    .A2(_04928_),
    .Y(_04942_),
    .B1(_04941_));
 sg13g2_nor2_1 _22638_ (.A(_04926_),
    .B(_04942_),
    .Y(_04943_));
 sg13g2_a22oi_1 _22639_ (.Y(_04944_),
    .B1(net494),
    .B2(\cpu.intr.r_timer_reload[0] ),
    .A2(net444),
    .A1(_10260_));
 sg13g2_a221oi_1 _22640_ (.B2(_10105_),
    .C1(net786),
    .B1(net435),
    .A1(\cpu.intr.r_timer_reload[16] ),
    .Y(_04945_),
    .A2(_10120_));
 sg13g2_a21oi_1 _22641_ (.A1(net786),
    .A2(_04944_),
    .Y(_04946_),
    .B1(_04945_));
 sg13g2_nor3_1 _22642_ (.A(net684),
    .B(_00285_),
    .C(_09831_),
    .Y(_04947_));
 sg13g2_nor2_1 _22643_ (.A(_10173_),
    .B(_09351_),
    .Y(_04948_));
 sg13g2_buf_1 _22644_ (.A(_04948_),
    .X(_04949_));
 sg13g2_and2_1 _22645_ (.A(net686),
    .B(_04949_),
    .X(_04950_));
 sg13g2_buf_1 _22646_ (.A(_04950_),
    .X(_04951_));
 sg13g2_buf_1 _22647_ (.A(_04951_),
    .X(_04952_));
 sg13g2_o21ai_1 _22648_ (.B1(net381),
    .Y(_04953_),
    .A1(_09328_),
    .A2(_09329_));
 sg13g2_buf_1 _22649_ (.A(\cpu.intr.r_clock_count[16] ),
    .X(_04954_));
 sg13g2_mux2_1 _22650_ (.A0(\cpu.intr.r_clock_cmp[0] ),
    .A1(\cpu.intr.r_clock_cmp[16] ),
    .S(net787),
    .X(_04955_));
 sg13g2_a22oi_1 _22651_ (.Y(_04956_),
    .B1(_04955_),
    .B2(net486),
    .A2(net443),
    .A1(_04954_));
 sg13g2_nand2_1 _22652_ (.Y(_04957_),
    .A(_04953_),
    .B(_04956_));
 sg13g2_nor3_1 _22653_ (.A(_04946_),
    .B(_04947_),
    .C(_04957_),
    .Y(_04958_));
 sg13g2_and2_1 _22654_ (.A(_10252_),
    .B(_04936_),
    .X(_04959_));
 sg13g2_buf_1 _22655_ (.A(_04959_),
    .X(_04960_));
 sg13g2_nor2_1 _22656_ (.A(net633),
    .B(_04960_),
    .Y(_04961_));
 sg13g2_nor2_1 _22657_ (.A(net922),
    .B(_04961_),
    .Y(_04962_));
 sg13g2_buf_1 _22658_ (.A(_04962_),
    .X(_04963_));
 sg13g2_o21ai_1 _22659_ (.B1(net264),
    .Y(_04964_),
    .A1(_09328_),
    .A2(_09329_));
 sg13g2_inv_1 _22660_ (.Y(_04965_),
    .A(_04964_));
 sg13g2_o21ai_1 _22661_ (.B1(\cpu.intr.r_enable[0] ),
    .Y(_04966_),
    .A1(net382),
    .A2(_04965_));
 sg13g2_a21oi_1 _22662_ (.A1(_04958_),
    .A2(_04966_),
    .Y(_04967_),
    .B1(net683));
 sg13g2_o21ai_1 _22663_ (.B1(net1120),
    .Y(_04968_),
    .A1(net1051),
    .A2(_10175_));
 sg13g2_nor2_1 _22664_ (.A(net1042),
    .B(net708),
    .Y(_04969_));
 sg13g2_nor2_1 _22665_ (.A(_11383_),
    .B(net758),
    .Y(_04970_));
 sg13g2_a21oi_1 _22666_ (.A1(_04968_),
    .A2(_04969_),
    .Y(_04971_),
    .B1(_04970_));
 sg13g2_o21ai_1 _22667_ (.B1(_04888_),
    .Y(_04972_),
    .A1(net758),
    .A2(_04887_));
 sg13g2_nand2_1 _22668_ (.Y(_04973_),
    .A(net929),
    .B(net1120));
 sg13g2_o21ai_1 _22669_ (.B1(_04888_),
    .Y(_04974_),
    .A1(_04973_),
    .A2(_04936_));
 sg13g2_a22oi_1 _22670_ (.Y(_04975_),
    .B1(net872),
    .B2(_04969_),
    .A2(_09343_),
    .A1(_10175_));
 sg13g2_nor2_1 _22671_ (.A(net933),
    .B(_04975_),
    .Y(_04976_));
 sg13g2_a221oi_1 _22672_ (.B2(_10123_),
    .C1(_04976_),
    .B1(_04974_),
    .A1(net681),
    .Y(_04977_),
    .A2(_04972_));
 sg13g2_o21ai_1 _22673_ (.B1(_04977_),
    .Y(_04978_),
    .A1(_10174_),
    .A2(_04971_));
 sg13g2_buf_2 _22674_ (.A(_04978_),
    .X(_04979_));
 sg13g2_nand3_1 _22675_ (.B(_09288_),
    .C(_04979_),
    .A(_09287_),
    .Y(_04980_));
 sg13g2_buf_2 _22676_ (.A(\cpu.gpio.r_spi_miso_src[0][0] ),
    .X(_04981_));
 sg13g2_nor3_1 _22677_ (.A(net933),
    .B(net872),
    .C(_09836_),
    .Y(_04982_));
 sg13g2_buf_1 _22678_ (.A(_04982_),
    .X(_04983_));
 sg13g2_buf_2 _22679_ (.A(\cpu.gpio.r_src_o[4][0] ),
    .X(_04984_));
 sg13g2_and2_1 _22680_ (.A(net872),
    .B(_04938_),
    .X(_04985_));
 sg13g2_buf_2 _22681_ (.A(_04985_),
    .X(_04986_));
 sg13g2_nor3_1 _22682_ (.A(net1120),
    .B(_04881_),
    .C(_04936_),
    .Y(_04987_));
 sg13g2_buf_1 _22683_ (.A(_04987_),
    .X(_04988_));
 sg13g2_buf_2 _22684_ (.A(\cpu.gpio.r_src_io[4][0] ),
    .X(_04989_));
 sg13g2_a22oi_1 _22685_ (.Y(_04990_),
    .B1(net428),
    .B2(_04989_),
    .A2(_04986_),
    .A1(_04984_));
 sg13g2_and2_1 _22686_ (.A(_11383_),
    .B(_04938_),
    .X(_04991_));
 sg13g2_buf_2 _22687_ (.A(_04991_),
    .X(_04992_));
 sg13g2_nand3_1 _22688_ (.B(net708),
    .C(_09382_),
    .A(net929),
    .Y(_04993_));
 sg13g2_buf_1 _22689_ (.A(_04993_),
    .X(_04994_));
 sg13g2_nor2_1 _22690_ (.A(net1042),
    .B(_04994_),
    .Y(_04995_));
 sg13g2_buf_1 _22691_ (.A(_04995_),
    .X(_04996_));
 sg13g2_a22oi_1 _22692_ (.Y(_04997_),
    .B1(net380),
    .B2(_09287_),
    .A2(_04992_),
    .A1(_09288_));
 sg13g2_buf_2 _22693_ (.A(\cpu.gpio.r_uart_rx_src[0] ),
    .X(_04998_));
 sg13g2_nand2_1 _22694_ (.Y(_04999_),
    .A(_04998_),
    .B(_04885_));
 sg13g2_buf_2 _22695_ (.A(\cpu.gpio.r_src_o[6][0] ),
    .X(_05000_));
 sg13g2_nand2_1 _22696_ (.Y(_05001_),
    .A(net1042),
    .B(_04932_));
 sg13g2_buf_1 _22697_ (.A(_05001_),
    .X(_05002_));
 sg13g2_inv_1 _22698_ (.Y(_05003_),
    .A(_05002_));
 sg13g2_nor3_1 _22699_ (.A(net1120),
    .B(_04881_),
    .C(_04903_),
    .Y(_05004_));
 sg13g2_buf_1 _22700_ (.A(_05004_),
    .X(_05005_));
 sg13g2_buf_2 _22701_ (.A(\cpu.gpio.r_src_io[6][0] ),
    .X(_05006_));
 sg13g2_a22oi_1 _22702_ (.Y(_05007_),
    .B1(net427),
    .B2(_05006_),
    .A2(_05003_),
    .A1(_05000_));
 sg13g2_nand4_1 _22703_ (.B(_04997_),
    .C(_04999_),
    .A(_04990_),
    .Y(_05008_),
    .D(_05007_));
 sg13g2_a21oi_1 _22704_ (.A1(_04981_),
    .A2(_04983_),
    .Y(_05009_),
    .B1(_05008_));
 sg13g2_nand2b_1 _22705_ (.Y(_05010_),
    .B(_09281_),
    .A_N(net984));
 sg13g2_buf_2 _22706_ (.A(_05010_),
    .X(_05011_));
 sg13g2_a21oi_1 _22707_ (.A1(_04980_),
    .A2(_05009_),
    .Y(_05012_),
    .B1(_05011_));
 sg13g2_nor4_1 _22708_ (.A(_04924_),
    .B(_04943_),
    .C(_04967_),
    .D(_05012_),
    .Y(_05013_));
 sg13g2_mux2_1 _22709_ (.A0(_04880_),
    .A1(_05013_),
    .S(net891),
    .X(_05014_));
 sg13g2_nor2_1 _22710_ (.A(net83),
    .B(_05014_),
    .Y(_05015_));
 sg13g2_a221oi_1 _22711_ (.B2(_03418_),
    .C1(_05015_),
    .B1(net63),
    .A1(net803),
    .Y(_05016_),
    .A2(_11686_));
 sg13g2_a221oi_1 _22712_ (.B2(net85),
    .C1(_05016_),
    .B1(_04823_),
    .A1(_04815_),
    .Y(_01031_),
    .A2(_04821_));
 sg13g2_nor2_1 _22713_ (.A(net762),
    .B(_04734_),
    .Y(_05017_));
 sg13g2_nand2_1 _22714_ (.Y(_05018_),
    .A(_09443_),
    .B(_11686_));
 sg13g2_buf_1 _22715_ (.A(_05018_),
    .X(_05019_));
 sg13g2_nor2_1 _22716_ (.A(net398),
    .B(_05019_),
    .Y(_05020_));
 sg13g2_buf_1 _22717_ (.A(_05019_),
    .X(_05021_));
 sg13g2_buf_1 _22718_ (.A(\cpu.spi.r_clk_count[2][7] ),
    .X(_05022_));
 sg13g2_nand2b_1 _22719_ (.Y(_05023_),
    .B(_04884_),
    .A_N(_00157_));
 sg13g2_o21ai_1 _22720_ (.B1(_05023_),
    .Y(_05024_),
    .A1(_00156_),
    .A2(_04919_));
 sg13g2_a221oi_1 _22721_ (.B2(\cpu.spi.r_timeout[7] ),
    .C1(_05024_),
    .B1(net430),
    .A1(_05022_),
    .Y(_05025_),
    .A2(_04915_));
 sg13g2_nand2b_1 _22722_ (.Y(_05026_),
    .B(_04897_),
    .A_N(_00222_));
 sg13g2_a21oi_1 _22723_ (.A1(_05025_),
    .A2(_05026_),
    .Y(_05027_),
    .B1(net709));
 sg13g2_a22oi_1 _22724_ (.Y(_05028_),
    .B1(_04928_),
    .B2(\cpu.uart.r_in[7] ),
    .A2(_04907_),
    .A1(\cpu.uart.r_div_value[7] ));
 sg13g2_a22oi_1 _22725_ (.Y(_05029_),
    .B1(net603),
    .B2(_10106_),
    .A2(net621),
    .A1(\cpu.intr.r_timer_reload[23] ));
 sg13g2_a221oi_1 _22726_ (.B2(\cpu.intr.r_clock_cmp[7] ),
    .C1(net923),
    .B1(net604),
    .A1(\cpu.intr.r_timer_reload[7] ),
    .Y(_05030_),
    .A2(net621));
 sg13g2_a21oi_1 _22727_ (.A1(net923),
    .A2(_05029_),
    .Y(_05031_),
    .B1(_05030_));
 sg13g2_nor2_1 _22728_ (.A(net923),
    .B(_09831_),
    .Y(_05032_));
 sg13g2_buf_2 _22729_ (.A(_05032_),
    .X(_05033_));
 sg13g2_nor2_1 _22730_ (.A(_09380_),
    .B(_12657_),
    .Y(_05034_));
 sg13g2_buf_2 _22731_ (.A(_05034_),
    .X(_05035_));
 sg13g2_a22oi_1 _22732_ (.Y(_05036_),
    .B1(_05035_),
    .B2(_10293_),
    .A2(_05033_),
    .A1(\cpu.intr.r_timer_count[7] ));
 sg13g2_buf_1 _22733_ (.A(\cpu.intr.r_clock_count[23] ),
    .X(_05037_));
 sg13g2_nor2_1 _22734_ (.A(net933),
    .B(_09836_),
    .Y(_05038_));
 sg13g2_a22oi_1 _22735_ (.Y(_05039_),
    .B1(_05038_),
    .B2(\cpu.intr.r_clock_cmp[23] ),
    .A2(_10254_),
    .A1(_05037_));
 sg13g2_nand2_1 _22736_ (.Y(_05040_),
    .A(_05036_),
    .B(_05039_));
 sg13g2_nor2_1 _22737_ (.A(_10125_),
    .B(_04963_),
    .Y(_05041_));
 sg13g2_o21ai_1 _22738_ (.B1(_05041_),
    .Y(_05042_),
    .A1(_05031_),
    .A2(_05040_));
 sg13g2_o21ai_1 _22739_ (.B1(_05042_),
    .Y(_05043_),
    .A1(_04926_),
    .A2(_05028_));
 sg13g2_a21oi_1 _22740_ (.A1(_09293_),
    .A2(_04951_),
    .Y(_05044_),
    .B1(_04932_));
 sg13g2_nand2b_1 _22741_ (.Y(_05045_),
    .B(_09294_),
    .A_N(_05044_));
 sg13g2_nor2_1 _22742_ (.A(net933),
    .B(_00162_),
    .Y(_05046_));
 sg13g2_nor2b_1 _22743_ (.A(net923),
    .B_N(net10),
    .Y(_05047_));
 sg13g2_o21ai_1 _22744_ (.B1(_12780_),
    .Y(_05048_),
    .A1(_05046_),
    .A2(_05047_));
 sg13g2_a22oi_1 _22745_ (.Y(_05049_),
    .B1(_05035_),
    .B2(\cpu.gpio.genblk1[7].srcs_o[0] ),
    .A2(_10254_),
    .A1(\cpu.gpio.genblk2[7].srcs_io[0] ));
 sg13g2_nand3_1 _22746_ (.B(_05048_),
    .C(_05049_),
    .A(_05045_),
    .Y(_05050_));
 sg13g2_inv_1 _22747_ (.Y(_05051_),
    .A(_00158_));
 sg13g2_a22oi_1 _22748_ (.Y(_05052_),
    .B1(_05005_),
    .B2(_05051_),
    .A2(_04884_),
    .A1(_09293_));
 sg13g2_buf_1 _22749_ (.A(\cpu.gpio.r_src_io[5][3] ),
    .X(_05053_));
 sg13g2_nand2_1 _22750_ (.Y(_05054_),
    .A(net872),
    .B(_04938_));
 sg13g2_nor2_1 _22751_ (.A(_00160_),
    .B(_05054_),
    .Y(_05055_));
 sg13g2_a221oi_1 _22752_ (.B2(_09290_),
    .C1(_05055_),
    .B1(_04992_),
    .A1(_05053_),
    .Y(_05056_),
    .A2(net428));
 sg13g2_nand3_1 _22753_ (.B(net1051),
    .C(net686),
    .A(net681),
    .Y(_05057_));
 sg13g2_buf_2 _22754_ (.A(_05057_),
    .X(_05058_));
 sg13g2_nand2b_1 _22755_ (.Y(_05059_),
    .B(_04951_),
    .A_N(_00161_));
 sg13g2_o21ai_1 _22756_ (.B1(_05059_),
    .Y(_05060_),
    .A1(_00159_),
    .A2(_05058_));
 sg13g2_a22oi_1 _22757_ (.Y(_05061_),
    .B1(_05060_),
    .B2(net1042),
    .A2(net380),
    .A1(_09289_));
 sg13g2_nand3_1 _22758_ (.B(_05056_),
    .C(_05061_),
    .A(_05052_),
    .Y(_05062_));
 sg13g2_a21oi_1 _22759_ (.A1(net977),
    .A2(_05050_),
    .Y(_05063_),
    .B1(_05062_));
 sg13g2_nand3_1 _22760_ (.B(_09290_),
    .C(_04979_),
    .A(_09289_),
    .Y(_05064_));
 sg13g2_a21oi_1 _22761_ (.A1(_05063_),
    .A2(_05064_),
    .Y(_05065_),
    .B1(_05011_));
 sg13g2_or3_1 _22762_ (.A(_05027_),
    .B(_05043_),
    .C(_05065_),
    .X(_05066_));
 sg13g2_inv_1 _22763_ (.Y(_05067_),
    .A(_04877_));
 sg13g2_a22oi_1 _22764_ (.Y(_05068_),
    .B1(net603),
    .B2(\cpu.dcache.r_data[6][7] ),
    .A2(net627),
    .A1(\cpu.dcache.r_data[3][7] ));
 sg13g2_a22oi_1 _22765_ (.Y(_05069_),
    .B1(net604),
    .B2(\cpu.dcache.r_data[5][7] ),
    .A2(net699),
    .A1(\cpu.dcache.r_data[7][7] ));
 sg13g2_a22oi_1 _22766_ (.Y(_05070_),
    .B1(net549),
    .B2(\cpu.dcache.r_data[2][7] ),
    .A2(net626),
    .A1(\cpu.dcache.r_data[4][7] ));
 sg13g2_nand3_1 _22767_ (.B(_05069_),
    .C(_05070_),
    .A(_05068_),
    .Y(_05071_));
 sg13g2_nand2_1 _22768_ (.Y(_05072_),
    .A(_00152_),
    .B(net686));
 sg13g2_o21ai_1 _22769_ (.B1(_05072_),
    .Y(_05073_),
    .A1(net686),
    .A2(_05071_));
 sg13g2_o21ai_1 _22770_ (.B1(_12330_),
    .Y(_05074_),
    .A1(\cpu.dcache.r_data[1][7] ),
    .A2(_05071_));
 sg13g2_o21ai_1 _22771_ (.B1(_05074_),
    .Y(_05075_),
    .A1(_12330_),
    .A2(_05073_));
 sg13g2_and2_1 _22772_ (.A(net708),
    .B(\cpu.dcache.r_data[6][31] ),
    .X(_05076_));
 sg13g2_a21oi_1 _22773_ (.A1(net758),
    .A2(\cpu.dcache.r_data[4][31] ),
    .Y(_05077_),
    .B1(_05076_));
 sg13g2_nand3_1 _22774_ (.B(net633),
    .C(\cpu.dcache.r_data[7][31] ),
    .A(net681),
    .Y(_05078_));
 sg13g2_o21ai_1 _22775_ (.B1(_05078_),
    .Y(_05079_),
    .A1(net681),
    .A2(_05077_));
 sg13g2_a22oi_1 _22776_ (.Y(_05080_),
    .B1(net549),
    .B2(\cpu.dcache.r_data[2][31] ),
    .A2(net547),
    .A1(\cpu.dcache.r_data[1][31] ));
 sg13g2_a22oi_1 _22777_ (.Y(_05081_),
    .B1(net604),
    .B2(\cpu.dcache.r_data[5][31] ),
    .A2(net627),
    .A1(\cpu.dcache.r_data[3][31] ));
 sg13g2_nand2_1 _22778_ (.Y(_05082_),
    .A(_05080_),
    .B(_05081_));
 sg13g2_a21oi_1 _22779_ (.A1(net922),
    .A2(_05079_),
    .Y(_05083_),
    .B1(_05082_));
 sg13g2_o21ai_1 _22780_ (.B1(_05083_),
    .Y(_05084_),
    .A1(_00154_),
    .A2(net548));
 sg13g2_a22oi_1 _22781_ (.Y(_05085_),
    .B1(net626),
    .B2(\cpu.dcache.r_data[4][23] ),
    .A2(net627),
    .A1(\cpu.dcache.r_data[3][23] ));
 sg13g2_nand2_1 _22782_ (.Y(_05086_),
    .A(\cpu.dcache.r_data[7][23] ),
    .B(net699));
 sg13g2_a22oi_1 _22783_ (.Y(_05087_),
    .B1(_02731_),
    .B2(\cpu.dcache.r_data[6][23] ),
    .A2(net549),
    .A1(\cpu.dcache.r_data[2][23] ));
 sg13g2_nor2_1 _22784_ (.A(_00153_),
    .B(_09623_),
    .Y(_05088_));
 sg13g2_a221oi_1 _22785_ (.B2(\cpu.dcache.r_data[5][23] ),
    .C1(_05088_),
    .B1(net702),
    .A1(\cpu.dcache.r_data[1][23] ),
    .Y(_05089_),
    .A2(_09697_));
 sg13g2_nand4_1 _22786_ (.B(_05086_),
    .C(_05087_),
    .A(_05085_),
    .Y(_05090_),
    .D(_05089_));
 sg13g2_nand2_1 _22787_ (.Y(_05091_),
    .A(_10115_),
    .B(_05090_));
 sg13g2_nor2_1 _22788_ (.A(net654),
    .B(_05091_),
    .Y(_05092_));
 sg13g2_a21oi_1 _22789_ (.A1(net654),
    .A2(_05084_),
    .Y(_05093_),
    .B1(_05092_));
 sg13g2_a22oi_1 _22790_ (.Y(_05094_),
    .B1(net549),
    .B2(\cpu.dcache.r_data[2][15] ),
    .A2(net547),
    .A1(\cpu.dcache.r_data[1][15] ));
 sg13g2_a22oi_1 _22791_ (.Y(_05095_),
    .B1(net626),
    .B2(\cpu.dcache.r_data[4][15] ),
    .A2(net627),
    .A1(\cpu.dcache.r_data[3][15] ));
 sg13g2_mux2_1 _22792_ (.A0(\cpu.dcache.r_data[5][15] ),
    .A1(\cpu.dcache.r_data[7][15] ),
    .S(net708),
    .X(_05096_));
 sg13g2_a22oi_1 _22793_ (.Y(_05097_),
    .B1(_05096_),
    .B2(net681),
    .A2(net928),
    .A1(\cpu.dcache.r_data[6][15] ));
 sg13g2_nand2b_1 _22794_ (.Y(_05098_),
    .B(net922),
    .A_N(_05097_));
 sg13g2_and4_1 _22795_ (.A(net548),
    .B(_05094_),
    .C(_05095_),
    .D(_05098_),
    .X(_05099_));
 sg13g2_a21oi_1 _22796_ (.A1(_00155_),
    .A2(net546),
    .Y(_05100_),
    .B1(_05099_));
 sg13g2_and2_1 _22797_ (.A(_09352_),
    .B(_05100_),
    .X(_05101_));
 sg13g2_o21ai_1 _22798_ (.B1(net654),
    .Y(_05102_),
    .A1(_08502_),
    .A2(_05101_));
 sg13g2_o21ai_1 _22799_ (.B1(_05102_),
    .Y(_05103_),
    .A1(_12120_),
    .A2(_05093_));
 sg13g2_a21oi_1 _22800_ (.A1(_05067_),
    .A2(_05075_),
    .Y(_05104_),
    .B1(_05103_));
 sg13g2_nand2_1 _22801_ (.Y(_05105_),
    .A(_04866_),
    .B(_05091_));
 sg13g2_a21oi_1 _22802_ (.A1(_09352_),
    .A2(_05075_),
    .Y(_05106_),
    .B1(_05105_));
 sg13g2_nor3_1 _22803_ (.A(_12117_),
    .B(_05104_),
    .C(_05106_),
    .Y(_05107_));
 sg13g2_a21oi_2 _22804_ (.B1(_05107_),
    .Y(_05108_),
    .A2(_05066_),
    .A1(_12117_));
 sg13g2_nand2_1 _22805_ (.Y(_05109_),
    .A(_08499_),
    .B(_05108_));
 sg13g2_inv_1 _22806_ (.Y(_05110_),
    .A(_05109_));
 sg13g2_buf_1 _22807_ (.A(_04866_),
    .X(_05111_));
 sg13g2_mux2_1 _22808_ (.A0(\cpu.dcache.r_data[5][26] ),
    .A1(\cpu.dcache.r_data[7][26] ),
    .S(net633),
    .X(_05112_));
 sg13g2_a22oi_1 _22809_ (.Y(_05113_),
    .B1(_05112_),
    .B2(net619),
    .A2(net689),
    .A1(\cpu.dcache.r_data[4][26] ));
 sg13g2_nand2b_1 _22810_ (.Y(_05114_),
    .B(net922),
    .A_N(_05113_));
 sg13g2_a22oi_1 _22811_ (.Y(_05115_),
    .B1(net488),
    .B2(\cpu.dcache.r_data[2][26] ),
    .A2(net530),
    .A1(\cpu.dcache.r_data[3][26] ));
 sg13g2_a22oi_1 _22812_ (.Y(_05116_),
    .B1(net603),
    .B2(\cpu.dcache.r_data[6][26] ),
    .A2(net489),
    .A1(\cpu.dcache.r_data[1][26] ));
 sg13g2_and3_1 _22813_ (.X(_05117_),
    .A(_05114_),
    .B(_05115_),
    .C(_05116_));
 sg13g2_o21ai_1 _22814_ (.B1(_05117_),
    .Y(_05118_),
    .A1(_00102_),
    .A2(net433));
 sg13g2_a22oi_1 _22815_ (.Y(_05119_),
    .B1(net544),
    .B2(\cpu.dcache.r_data[4][10] ),
    .A2(net468),
    .A1(\cpu.dcache.r_data[3][10] ));
 sg13g2_nand2_1 _22816_ (.Y(_05120_),
    .A(\cpu.dcache.r_data[5][10] ),
    .B(net529));
 sg13g2_a22oi_1 _22817_ (.Y(_05121_),
    .B1(net528),
    .B2(\cpu.dcache.r_data[6][10] ),
    .A2(net432),
    .A1(\cpu.dcache.r_data[2][10] ));
 sg13g2_nor2_1 _22818_ (.A(_00103_),
    .B(net548),
    .Y(_05122_));
 sg13g2_a221oi_1 _22819_ (.B2(\cpu.dcache.r_data[7][10] ),
    .C1(_05122_),
    .B1(net545),
    .A1(\cpu.dcache.r_data[1][10] ),
    .Y(_05123_),
    .A2(net489));
 sg13g2_nand4_1 _22820_ (.B(_05120_),
    .C(_05121_),
    .A(_05119_),
    .Y(_05124_),
    .D(_05123_));
 sg13g2_mux2_1 _22821_ (.A0(_05118_),
    .A1(_05124_),
    .S(net682),
    .X(_05125_));
 sg13g2_and2_1 _22822_ (.A(net1011),
    .B(_05041_),
    .X(_05126_));
 sg13g2_buf_2 _22823_ (.A(_05126_),
    .X(_05127_));
 sg13g2_nand2_2 _22824_ (.Y(_05128_),
    .A(net786),
    .B(_10176_));
 sg13g2_mux2_1 _22825_ (.A0(\cpu.intr.r_clock_cmp[10] ),
    .A1(\cpu.intr.r_timer_reload[10] ),
    .S(net437),
    .X(_05129_));
 sg13g2_a22oi_1 _22826_ (.Y(_05130_),
    .B1(_05129_),
    .B2(net475),
    .A2(net759),
    .A1(\cpu.intr.r_timer_count[10] ));
 sg13g2_buf_1 _22827_ (.A(_05038_),
    .X(_05131_));
 sg13g2_buf_1 _22828_ (.A(_05035_),
    .X(_05132_));
 sg13g2_buf_2 _22829_ (.A(\cpu.intr.r_clock_count[26] ),
    .X(_05133_));
 sg13g2_and2_1 _22830_ (.A(_05133_),
    .B(net399),
    .X(_05134_));
 sg13g2_a221oi_1 _22831_ (.B2(_10309_),
    .C1(_05134_),
    .B1(net467),
    .A1(\cpu.intr.r_clock_cmp[26] ),
    .Y(_05135_),
    .A2(net653));
 sg13g2_o21ai_1 _22832_ (.B1(_05135_),
    .Y(_05136_),
    .A1(_05128_),
    .A2(_05130_));
 sg13g2_buf_1 _22833_ (.A(_08499_),
    .X(_05137_));
 sg13g2_a221oi_1 _22834_ (.B2(_05136_),
    .C1(net976),
    .B1(_05127_),
    .A1(net514),
    .Y(_05138_),
    .A2(_05125_));
 sg13g2_nor3_1 _22835_ (.A(net84),
    .B(_05110_),
    .C(_05138_),
    .Y(_05139_));
 sg13g2_a21oi_1 _22836_ (.A1(net1107),
    .A2(net83),
    .Y(_05140_),
    .B1(_05139_));
 sg13g2_nor3_1 _22837_ (.A(net978),
    .B(net215),
    .C(_05019_),
    .Y(_05141_));
 sg13g2_a21o_1 _22838_ (.A2(_05140_),
    .A1(net98),
    .B1(_05141_),
    .X(_05142_));
 sg13g2_a221oi_1 _22839_ (.B2(_05020_),
    .C1(_05142_),
    .B1(_05017_),
    .A1(_04731_),
    .Y(_01032_),
    .A2(_04821_));
 sg13g2_buf_1 _22840_ (.A(_05019_),
    .X(_05143_));
 sg13g2_a22oi_1 _22841_ (.Y(_05144_),
    .B1(net603),
    .B2(\cpu.dcache.r_data[6][11] ),
    .A2(net549),
    .A1(\cpu.dcache.r_data[2][11] ));
 sg13g2_a22oi_1 _22842_ (.Y(_05145_),
    .B1(net604),
    .B2(\cpu.dcache.r_data[5][11] ),
    .A2(net621),
    .A1(\cpu.dcache.r_data[7][11] ));
 sg13g2_a22oi_1 _22843_ (.Y(_05146_),
    .B1(net626),
    .B2(\cpu.dcache.r_data[4][11] ),
    .A2(net627),
    .A1(\cpu.dcache.r_data[3][11] ));
 sg13g2_nand3_1 _22844_ (.B(_05145_),
    .C(_05146_),
    .A(_05144_),
    .Y(_05147_));
 sg13g2_nand2_1 _22845_ (.Y(_05148_),
    .A(_00113_),
    .B(net686));
 sg13g2_o21ai_1 _22846_ (.B1(_05148_),
    .Y(_05149_),
    .A1(net686),
    .A2(_05147_));
 sg13g2_o21ai_1 _22847_ (.B1(net431),
    .Y(_05150_),
    .A1(\cpu.dcache.r_data[1][11] ),
    .A2(_05147_));
 sg13g2_o21ai_1 _22848_ (.B1(_05150_),
    .Y(_05151_),
    .A1(net431),
    .A2(_05149_));
 sg13g2_a22oi_1 _22849_ (.Y(_05152_),
    .B1(net603),
    .B2(\cpu.dcache.r_data[6][27] ),
    .A2(net549),
    .A1(\cpu.dcache.r_data[2][27] ));
 sg13g2_a22oi_1 _22850_ (.Y(_05153_),
    .B1(net604),
    .B2(\cpu.dcache.r_data[5][27] ),
    .A2(net621),
    .A1(\cpu.dcache.r_data[7][27] ));
 sg13g2_a22oi_1 _22851_ (.Y(_05154_),
    .B1(net544),
    .B2(\cpu.dcache.r_data[4][27] ),
    .A2(net627),
    .A1(\cpu.dcache.r_data[3][27] ));
 sg13g2_nand3_1 _22852_ (.B(_05153_),
    .C(_05154_),
    .A(_05152_),
    .Y(_05155_));
 sg13g2_nand2_1 _22853_ (.Y(_05156_),
    .A(_00112_),
    .B(net586));
 sg13g2_o21ai_1 _22854_ (.B1(_05156_),
    .Y(_05157_),
    .A1(net586),
    .A2(_05155_));
 sg13g2_o21ai_1 _22855_ (.B1(net431),
    .Y(_05158_),
    .A1(\cpu.dcache.r_data[1][27] ),
    .A2(_05155_));
 sg13g2_o21ai_1 _22856_ (.B1(_05158_),
    .Y(_05159_),
    .A1(net389),
    .A2(_05157_));
 sg13g2_mux2_1 _22857_ (.A0(_05151_),
    .A1(_05159_),
    .S(net618),
    .X(_05160_));
 sg13g2_nor2_1 _22858_ (.A(net923),
    .B(_09836_),
    .Y(_05161_));
 sg13g2_buf_1 _22859_ (.A(_05161_),
    .X(_05162_));
 sg13g2_a22oi_1 _22860_ (.Y(_05163_),
    .B1(net652),
    .B2(\cpu.intr.r_clock_cmp[11] ),
    .A2(net467),
    .A1(_10314_));
 sg13g2_buf_2 _22861_ (.A(\cpu.intr.r_clock_count[27] ),
    .X(_05164_));
 sg13g2_a22oi_1 _22862_ (.Y(_05165_),
    .B1(net653),
    .B2(\cpu.intr.r_clock_cmp[27] ),
    .A2(net399),
    .A1(_05164_));
 sg13g2_a22oi_1 _22863_ (.Y(_05166_),
    .B1(net435),
    .B2(_10090_),
    .A2(net445),
    .A1(\cpu.intr.r_timer_reload[11] ));
 sg13g2_or2_1 _22864_ (.X(_05167_),
    .B(_05166_),
    .A(net618));
 sg13g2_nand3_1 _22865_ (.B(_05165_),
    .C(_05167_),
    .A(_05163_),
    .Y(_05168_));
 sg13g2_a221oi_1 _22866_ (.B2(_05127_),
    .C1(net976),
    .B1(_05168_),
    .A1(net514),
    .Y(_05169_),
    .A2(_05160_));
 sg13g2_nor3_1 _22867_ (.A(_04827_),
    .B(_05110_),
    .C(_05169_),
    .Y(_05170_));
 sg13g2_a21oi_1 _22868_ (.A1(_10680_),
    .A2(net63),
    .Y(_05171_),
    .B1(_05170_));
 sg13g2_mux2_1 _22869_ (.A0(_04221_),
    .A1(_04210_),
    .S(net762),
    .X(_05172_));
 sg13g2_buf_1 _22870_ (.A(net215),
    .X(_05173_));
 sg13g2_nor3_1 _22871_ (.A(_08746_),
    .B(net189),
    .C(net98),
    .Y(_05174_));
 sg13g2_a221oi_1 _22872_ (.B2(_05020_),
    .C1(_05174_),
    .B1(_05172_),
    .A1(net97),
    .Y(_01033_),
    .A2(_05171_));
 sg13g2_nand2_1 _22873_ (.Y(_05175_),
    .A(net655),
    .B(_04280_));
 sg13g2_a22oi_1 _22874_ (.Y(_05176_),
    .B1(net493),
    .B2(\cpu.dcache.r_data[4][28] ),
    .A2(net468),
    .A1(\cpu.dcache.r_data[3][28] ));
 sg13g2_nand2_1 _22875_ (.Y(_05177_),
    .A(\cpu.dcache.r_data[5][28] ),
    .B(net529));
 sg13g2_a22oi_1 _22876_ (.Y(_05178_),
    .B1(net528),
    .B2(\cpu.dcache.r_data[6][28] ),
    .A2(net432),
    .A1(\cpu.dcache.r_data[2][28] ));
 sg13g2_nor2_1 _22877_ (.A(_00123_),
    .B(net469),
    .Y(_05179_));
 sg13g2_a221oi_1 _22878_ (.B2(\cpu.dcache.r_data[7][28] ),
    .C1(_05179_),
    .B1(net545),
    .A1(\cpu.dcache.r_data[1][28] ),
    .Y(_05180_),
    .A2(net439));
 sg13g2_nand4_1 _22879_ (.B(_05177_),
    .C(_05178_),
    .A(_05176_),
    .Y(_05181_),
    .D(_05180_));
 sg13g2_buf_1 _22880_ (.A(_05181_),
    .X(_05182_));
 sg13g2_a22oi_1 _22881_ (.Y(_05183_),
    .B1(net488),
    .B2(\cpu.dcache.r_data[2][12] ),
    .A2(net489),
    .A1(\cpu.dcache.r_data[1][12] ));
 sg13g2_a22oi_1 _22882_ (.Y(_05184_),
    .B1(net544),
    .B2(\cpu.dcache.r_data[4][12] ),
    .A2(net530),
    .A1(\cpu.dcache.r_data[3][12] ));
 sg13g2_mux2_1 _22883_ (.A0(\cpu.dcache.r_data[5][12] ),
    .A1(\cpu.dcache.r_data[7][12] ),
    .S(net633),
    .X(_05185_));
 sg13g2_a22oi_1 _22884_ (.Y(_05186_),
    .B1(_05185_),
    .B2(net619),
    .A2(net759),
    .A1(\cpu.dcache.r_data[6][12] ));
 sg13g2_nand2b_1 _22885_ (.Y(_05187_),
    .B(net922),
    .A_N(_05186_));
 sg13g2_and4_1 _22886_ (.A(net469),
    .B(_05183_),
    .C(_05184_),
    .D(_05187_),
    .X(_05188_));
 sg13g2_a21oi_1 _22887_ (.A1(_00124_),
    .A2(net546),
    .Y(_05189_),
    .B1(_05188_));
 sg13g2_and2_1 _22888_ (.A(net786),
    .B(_05189_),
    .X(_05190_));
 sg13g2_a21oi_1 _22889_ (.A1(net684),
    .A2(_05182_),
    .Y(_05191_),
    .B1(_05190_));
 sg13g2_mux2_1 _22890_ (.A0(\cpu.intr.r_clock_cmp[12] ),
    .A1(\cpu.intr.r_timer_reload[12] ),
    .S(net496),
    .X(_05192_));
 sg13g2_a22oi_1 _22891_ (.Y(_05193_),
    .B1(_05192_),
    .B2(net531),
    .A2(net689),
    .A1(_10321_));
 sg13g2_buf_1 _22892_ (.A(\cpu.intr.r_clock_count[28] ),
    .X(_05194_));
 sg13g2_and2_1 _22893_ (.A(_05194_),
    .B(_10254_),
    .X(_05195_));
 sg13g2_a221oi_1 _22894_ (.B2(\cpu.intr.r_clock_cmp[28] ),
    .C1(_05195_),
    .B1(_05038_),
    .A1(\cpu.intr.r_timer_count[12] ),
    .Y(_05196_),
    .A2(_05033_));
 sg13g2_o21ai_1 _22895_ (.B1(_05196_),
    .Y(_05197_),
    .A1(_05128_),
    .A2(_05193_));
 sg13g2_a21oi_1 _22896_ (.A1(_05127_),
    .A2(_05197_),
    .Y(_05198_),
    .B1(_08499_));
 sg13g2_o21ai_1 _22897_ (.B1(_05198_),
    .Y(_05199_),
    .A1(_04863_),
    .A2(_05191_));
 sg13g2_a21oi_1 _22898_ (.A1(_05109_),
    .A2(_05199_),
    .Y(_05200_),
    .B1(_04826_));
 sg13g2_a21oi_1 _22899_ (.A1(net876),
    .A2(_04826_),
    .Y(_05201_),
    .B1(_05200_));
 sg13g2_nand3b_1 _22900_ (.B(net398),
    .C(net101),
    .Y(_05202_),
    .A_N(_08530_));
 sg13g2_o21ai_1 _22901_ (.B1(_05202_),
    .Y(_05203_),
    .A1(net101),
    .A2(_05201_));
 sg13g2_a21oi_1 _22902_ (.A1(_05020_),
    .A2(_05175_),
    .Y(_05204_),
    .B1(_05203_));
 sg13g2_nor4_1 _22903_ (.A(net655),
    .B(_04273_),
    .C(_04276_),
    .D(_05203_),
    .Y(_05205_));
 sg13g2_or2_1 _22904_ (.X(_01034_),
    .B(_05205_),
    .A(_05204_));
 sg13g2_o21ai_1 _22905_ (.B1(_05019_),
    .Y(_05206_),
    .A1(_11680_),
    .A2(_05108_));
 sg13g2_buf_1 _22906_ (.A(_05206_),
    .X(_05207_));
 sg13g2_buf_1 _22907_ (.A(\cpu.intr.r_clock_count[29] ),
    .X(_05208_));
 sg13g2_a22oi_1 _22908_ (.Y(_05209_),
    .B1(net467),
    .B2(_10327_),
    .A2(net399),
    .A1(_05208_));
 sg13g2_a22oi_1 _22909_ (.Y(_05210_),
    .B1(net653),
    .B2(\cpu.intr.r_clock_cmp[29] ),
    .A2(_05033_),
    .A1(\cpu.intr.r_timer_count[13] ));
 sg13g2_a22oi_1 _22910_ (.Y(_05211_),
    .B1(net486),
    .B2(\cpu.intr.r_clock_cmp[13] ),
    .A2(net445),
    .A1(\cpu.intr.r_timer_reload[13] ));
 sg13g2_or2_1 _22911_ (.X(_05212_),
    .B(_05211_),
    .A(net684));
 sg13g2_nand3_1 _22912_ (.B(_05210_),
    .C(_05212_),
    .A(_05209_),
    .Y(_05213_));
 sg13g2_nand2_1 _22913_ (.Y(_05214_),
    .A(\cpu.dcache.r_data[7][29] ),
    .B(net545));
 sg13g2_a22oi_1 _22914_ (.Y(_05215_),
    .B1(net529),
    .B2(\cpu.dcache.r_data[5][29] ),
    .A2(net468),
    .A1(\cpu.dcache.r_data[3][29] ));
 sg13g2_a22oi_1 _22915_ (.Y(_05216_),
    .B1(net528),
    .B2(\cpu.dcache.r_data[6][29] ),
    .A2(net544),
    .A1(\cpu.dcache.r_data[4][29] ));
 sg13g2_a22oi_1 _22916_ (.Y(_05217_),
    .B1(net432),
    .B2(\cpu.dcache.r_data[2][29] ),
    .A2(net439),
    .A1(\cpu.dcache.r_data[1][29] ));
 sg13g2_nand4_1 _22917_ (.B(_05215_),
    .C(_05216_),
    .A(_05214_),
    .Y(_05218_),
    .D(_05217_));
 sg13g2_nand2_1 _22918_ (.Y(_05219_),
    .A(_00130_),
    .B(net546));
 sg13g2_o21ai_1 _22919_ (.B1(_05219_),
    .Y(_05220_),
    .A1(net546),
    .A2(_05218_));
 sg13g2_nor2_1 _22920_ (.A(_00131_),
    .B(net469),
    .Y(_05221_));
 sg13g2_mux2_1 _22921_ (.A0(\cpu.dcache.r_data[5][13] ),
    .A1(\cpu.dcache.r_data[7][13] ),
    .S(net551),
    .X(_05222_));
 sg13g2_a22oi_1 _22922_ (.Y(_05223_),
    .B1(_05222_),
    .B2(net619),
    .A2(net689),
    .A1(\cpu.dcache.r_data[4][13] ));
 sg13g2_nor2_1 _22923_ (.A(net929),
    .B(_05223_),
    .Y(_05224_));
 sg13g2_a22oi_1 _22924_ (.Y(_05225_),
    .B1(net528),
    .B2(\cpu.dcache.r_data[6][13] ),
    .A2(net530),
    .A1(\cpu.dcache.r_data[3][13] ));
 sg13g2_a22oi_1 _22925_ (.Y(_05226_),
    .B1(net488),
    .B2(\cpu.dcache.r_data[2][13] ),
    .A2(net489),
    .A1(\cpu.dcache.r_data[1][13] ));
 sg13g2_nand2_1 _22926_ (.Y(_05227_),
    .A(_05225_),
    .B(_05226_));
 sg13g2_nor3_1 _22927_ (.A(_05221_),
    .B(_05224_),
    .C(_05227_),
    .Y(_05228_));
 sg13g2_or2_1 _22928_ (.X(_05229_),
    .B(_05228_),
    .A(_12151_));
 sg13g2_o21ai_1 _22929_ (.B1(_05229_),
    .Y(_05230_),
    .A1(net682),
    .A2(_05220_));
 sg13g2_a22oi_1 _22930_ (.Y(_05231_),
    .B1(_05230_),
    .B2(net514),
    .A2(_05213_),
    .A1(_05127_));
 sg13g2_nor2_1 _22931_ (.A(net976),
    .B(_05231_),
    .Y(_05232_));
 sg13g2_nor3_1 _22932_ (.A(net84),
    .B(_05207_),
    .C(_05232_),
    .Y(_05233_));
 sg13g2_a21o_1 _22933_ (.A2(net63),
    .A1(_03697_),
    .B1(_05233_),
    .X(_05234_));
 sg13g2_nor2_1 _22934_ (.A(net157),
    .B(\cpu.ex.c_mult[13] ),
    .Y(_05235_));
 sg13g2_or3_1 _22935_ (.A(net655),
    .B(_04320_),
    .C(_05235_),
    .X(_05236_));
 sg13g2_a21oi_1 _22936_ (.A1(net655),
    .A2(_04323_),
    .Y(_05237_),
    .B1(_04820_));
 sg13g2_nor3_1 _22937_ (.A(_08689_),
    .B(net189),
    .C(net98),
    .Y(_05238_));
 sg13g2_a221oi_1 _22938_ (.B2(_05237_),
    .C1(_05238_),
    .B1(_05236_),
    .A1(net97),
    .Y(_01035_),
    .A2(_05234_));
 sg13g2_buf_1 _22939_ (.A(_11689_),
    .X(_05239_));
 sg13g2_a22oi_1 _22940_ (.Y(_05240_),
    .B1(net652),
    .B2(\cpu.intr.r_clock_cmp[14] ),
    .A2(net467),
    .A1(_10333_));
 sg13g2_buf_1 _22941_ (.A(\cpu.intr.r_clock_count[30] ),
    .X(_05241_));
 sg13g2_a22oi_1 _22942_ (.Y(_05242_),
    .B1(net653),
    .B2(\cpu.intr.r_clock_cmp[30] ),
    .A2(net399),
    .A1(_05241_));
 sg13g2_a22oi_1 _22943_ (.Y(_05243_),
    .B1(net435),
    .B2(_10089_),
    .A2(net494),
    .A1(\cpu.intr.r_timer_reload[14] ));
 sg13g2_or2_1 _22944_ (.X(_05244_),
    .B(_05243_),
    .A(net684));
 sg13g2_nand3_1 _22945_ (.B(_05242_),
    .C(_05244_),
    .A(_05240_),
    .Y(_05245_));
 sg13g2_inv_1 _22946_ (.Y(_05246_),
    .A(_00142_));
 sg13g2_a22oi_1 _22947_ (.Y(_05247_),
    .B1(net488),
    .B2(\cpu.dcache.r_data[2][30] ),
    .A2(net489),
    .A1(\cpu.dcache.r_data[1][30] ));
 sg13g2_a22oi_1 _22948_ (.Y(_05248_),
    .B1(net544),
    .B2(\cpu.dcache.r_data[4][30] ),
    .A2(net530),
    .A1(\cpu.dcache.r_data[3][30] ));
 sg13g2_mux2_1 _22949_ (.A0(\cpu.dcache.r_data[5][30] ),
    .A1(\cpu.dcache.r_data[7][30] ),
    .S(net551),
    .X(_05249_));
 sg13g2_a22oi_1 _22950_ (.Y(_05250_),
    .B1(_05249_),
    .B2(net619),
    .A2(net759),
    .A1(\cpu.dcache.r_data[6][30] ));
 sg13g2_nand2b_1 _22951_ (.Y(_05251_),
    .B(net785),
    .A_N(_05250_));
 sg13g2_nand4_1 _22952_ (.B(_05247_),
    .C(_05248_),
    .A(net469),
    .Y(_05252_),
    .D(_05251_));
 sg13g2_o21ai_1 _22953_ (.B1(_05252_),
    .Y(_05253_),
    .A1(_05246_),
    .A2(net433));
 sg13g2_a22oi_1 _22954_ (.Y(_05254_),
    .B1(net493),
    .B2(\cpu.dcache.r_data[4][14] ),
    .A2(net468),
    .A1(\cpu.dcache.r_data[3][14] ));
 sg13g2_nand2_1 _22955_ (.Y(_05255_),
    .A(\cpu.dcache.r_data[7][14] ),
    .B(net545));
 sg13g2_a22oi_1 _22956_ (.Y(_05256_),
    .B1(net528),
    .B2(\cpu.dcache.r_data[6][14] ),
    .A2(net432),
    .A1(\cpu.dcache.r_data[2][14] ));
 sg13g2_nor2_1 _22957_ (.A(_00143_),
    .B(net469),
    .Y(_05257_));
 sg13g2_a221oi_1 _22958_ (.B2(\cpu.dcache.r_data[5][14] ),
    .C1(_05257_),
    .B1(net529),
    .A1(\cpu.dcache.r_data[1][14] ),
    .Y(_05258_),
    .A2(net439));
 sg13g2_nand4_1 _22959_ (.B(_05255_),
    .C(_05256_),
    .A(_05254_),
    .Y(_05259_),
    .D(_05258_));
 sg13g2_nand2_1 _22960_ (.Y(_05260_),
    .A(net786),
    .B(_05259_));
 sg13g2_o21ai_1 _22961_ (.B1(_05260_),
    .Y(_05261_),
    .A1(net682),
    .A2(_05253_));
 sg13g2_a22oi_1 _22962_ (.Y(_05262_),
    .B1(_05261_),
    .B2(_04866_),
    .A2(_05245_),
    .A1(_05127_));
 sg13g2_nor2_1 _22963_ (.A(net976),
    .B(_05262_),
    .Y(_05263_));
 sg13g2_nor3_1 _22964_ (.A(_04826_),
    .B(_05207_),
    .C(_05263_),
    .Y(_05264_));
 sg13g2_a21o_1 _22965_ (.A2(net84),
    .A1(_03700_),
    .B1(_05264_),
    .X(_05265_));
 sg13g2_o21ai_1 _22966_ (.B1(_11689_),
    .Y(_05266_),
    .A1(net815),
    .A2(_04822_));
 sg13g2_o21ai_1 _22967_ (.B1(_05266_),
    .Y(_05267_),
    .A1(net82),
    .A2(_05265_));
 sg13g2_o21ai_1 _22968_ (.B1(net762),
    .Y(_05268_),
    .A1(net157),
    .A2(\cpu.ex.c_mult[14] ));
 sg13g2_a21oi_1 _22969_ (.A1(net655),
    .A2(_04387_),
    .Y(_05269_),
    .B1(_04820_));
 sg13g2_o21ai_1 _22970_ (.B1(_05269_),
    .Y(_05270_),
    .A1(_04384_),
    .A2(_05268_));
 sg13g2_and2_1 _22971_ (.A(_05267_),
    .B(_05270_),
    .X(_01036_));
 sg13g2_nand2b_1 _22972_ (.Y(_05271_),
    .B(net655),
    .A_N(_04432_));
 sg13g2_a21oi_1 _22973_ (.A1(net684),
    .A2(_05084_),
    .Y(_05272_),
    .B1(_05101_));
 sg13g2_mux2_1 _22974_ (.A0(\cpu.intr.r_clock_cmp[15] ),
    .A1(\cpu.intr.r_timer_reload[15] ),
    .S(net496),
    .X(_05273_));
 sg13g2_a22oi_1 _22975_ (.Y(_05274_),
    .B1(_05273_),
    .B2(net531),
    .A2(net689),
    .A1(_10341_));
 sg13g2_buf_1 _22976_ (.A(\cpu.intr.r_clock_count[31] ),
    .X(_05275_));
 sg13g2_and2_1 _22977_ (.A(_05275_),
    .B(net443),
    .X(_05276_));
 sg13g2_a221oi_1 _22978_ (.B2(\cpu.intr.r_clock_cmp[31] ),
    .C1(_05276_),
    .B1(net653),
    .A1(\cpu.intr.r_timer_count[15] ),
    .Y(_05277_),
    .A2(_05033_));
 sg13g2_o21ai_1 _22979_ (.B1(_05277_),
    .Y(_05278_),
    .A1(_05128_),
    .A2(_05274_));
 sg13g2_nand2_1 _22980_ (.Y(_05279_),
    .A(_05127_),
    .B(_05278_));
 sg13g2_o21ai_1 _22981_ (.B1(_05279_),
    .Y(_05280_),
    .A1(_04863_),
    .A2(_05272_));
 sg13g2_a21oi_1 _22982_ (.A1(_11680_),
    .A2(_05280_),
    .Y(_05281_),
    .B1(_05207_));
 sg13g2_nor2_1 _22983_ (.A(_04826_),
    .B(_05281_),
    .Y(_05282_));
 sg13g2_a21oi_1 _22984_ (.A1(net926),
    .A2(net84),
    .Y(_05283_),
    .B1(_05282_));
 sg13g2_o21ai_1 _22985_ (.B1(net101),
    .Y(_05284_),
    .A1(_08679_),
    .A2(net215));
 sg13g2_o21ai_1 _22986_ (.B1(_05284_),
    .Y(_05285_),
    .A1(net101),
    .A2(_05283_));
 sg13g2_o21ai_1 _22987_ (.B1(_05285_),
    .Y(_05286_),
    .A1(_04820_),
    .A2(_05271_));
 sg13g2_a21oi_1 _22988_ (.A1(_04430_),
    .A2(_04821_),
    .Y(_01037_),
    .B1(_05286_));
 sg13g2_a22oi_1 _22989_ (.Y(_05287_),
    .B1(_10236_),
    .B2(\cpu.dcache.r_data[4][17] ),
    .A2(net487),
    .A1(\cpu.dcache.r_data[3][17] ));
 sg13g2_nand2_1 _22990_ (.Y(_05288_),
    .A(\cpu.dcache.r_data[7][17] ),
    .B(_10120_));
 sg13g2_a22oi_1 _22991_ (.Y(_05289_),
    .B1(net485),
    .B2(\cpu.dcache.r_data[6][17] ),
    .A2(net438),
    .A1(\cpu.dcache.r_data[2][17] ));
 sg13g2_nor2_1 _22992_ (.A(_00091_),
    .B(net433),
    .Y(_05290_));
 sg13g2_a221oi_1 _22993_ (.B2(\cpu.dcache.r_data[5][17] ),
    .C1(_05290_),
    .B1(_12782_),
    .A1(\cpu.dcache.r_data[1][17] ),
    .Y(_05291_),
    .A2(net431));
 sg13g2_nand4_1 _22994_ (.B(_05288_),
    .C(_05289_),
    .A(_05287_),
    .Y(_05292_),
    .D(_05291_));
 sg13g2_buf_1 _22995_ (.A(_05292_),
    .X(_05293_));
 sg13g2_and2_1 _22996_ (.A(\cpu.dcache.r_data[7][1] ),
    .B(net621),
    .X(_05294_));
 sg13g2_a221oi_1 _22997_ (.B2(\cpu.dcache.r_data[4][1] ),
    .C1(_05294_),
    .B1(net544),
    .A1(\cpu.dcache.r_data[3][1] ),
    .Y(_05295_),
    .A2(_04837_));
 sg13g2_a22oi_1 _22998_ (.Y(_05296_),
    .B1(_02732_),
    .B2(\cpu.dcache.r_data[6][1] ),
    .A2(net529),
    .A1(\cpu.dcache.r_data[5][1] ));
 sg13g2_a22oi_1 _22999_ (.Y(_05297_),
    .B1(_04835_),
    .B2(\cpu.dcache.r_data[2][1] ),
    .A2(net439),
    .A1(\cpu.dcache.r_data[1][1] ));
 sg13g2_nand4_1 _23000_ (.B(_05295_),
    .C(_05296_),
    .A(net433),
    .Y(_05298_),
    .D(_05297_));
 sg13g2_o21ai_1 _23001_ (.B1(_05298_),
    .Y(_05299_),
    .A1(\cpu.dcache.r_data[0][1] ),
    .A2(_04831_));
 sg13g2_nor2_1 _23002_ (.A(net618),
    .B(_05299_),
    .Y(_05300_));
 sg13g2_a21oi_1 _23003_ (.A1(net542),
    .A2(_05293_),
    .Y(_05301_),
    .B1(_05300_));
 sg13g2_nand2_1 _23004_ (.Y(_05302_),
    .A(\cpu.dcache.r_data[1][9] ),
    .B(net431));
 sg13g2_a22oi_1 _23005_ (.Y(_05303_),
    .B1(net485),
    .B2(\cpu.dcache.r_data[6][9] ),
    .A2(net545),
    .A1(\cpu.dcache.r_data[7][9] ));
 sg13g2_a22oi_1 _23006_ (.Y(_05304_),
    .B1(net438),
    .B2(\cpu.dcache.r_data[2][9] ),
    .A2(net493),
    .A1(\cpu.dcache.r_data[4][9] ));
 sg13g2_nor2_1 _23007_ (.A(_00093_),
    .B(net469),
    .Y(_05305_));
 sg13g2_a221oi_1 _23008_ (.B2(\cpu.dcache.r_data[5][9] ),
    .C1(_05305_),
    .B1(net529),
    .A1(\cpu.dcache.r_data[3][9] ),
    .Y(_05306_),
    .A2(net468));
 sg13g2_nand4_1 _23009_ (.B(_05303_),
    .C(_05304_),
    .A(_05302_),
    .Y(_05307_),
    .D(_05306_));
 sg13g2_nor2_1 _23010_ (.A(_12151_),
    .B(_04849_),
    .Y(_05308_));
 sg13g2_nand2_1 _23011_ (.Y(_05309_),
    .A(_05307_),
    .B(_05308_));
 sg13g2_o21ai_1 _23012_ (.B1(_05309_),
    .Y(_05310_),
    .A1(_04877_),
    .A2(_05299_));
 sg13g2_buf_1 _23013_ (.A(_12120_),
    .X(_05311_));
 sg13g2_mux2_1 _23014_ (.A0(\cpu.dcache.r_data[5][25] ),
    .A1(\cpu.dcache.r_data[7][25] ),
    .S(net551),
    .X(_05312_));
 sg13g2_a22oi_1 _23015_ (.Y(_05313_),
    .B1(_05312_),
    .B2(net619),
    .A2(net689),
    .A1(\cpu.dcache.r_data[4][25] ));
 sg13g2_nand2b_1 _23016_ (.Y(_05314_),
    .B(net785),
    .A_N(_05313_));
 sg13g2_a22oi_1 _23017_ (.Y(_05315_),
    .B1(net432),
    .B2(\cpu.dcache.r_data[2][25] ),
    .A2(net468),
    .A1(\cpu.dcache.r_data[3][25] ));
 sg13g2_a22oi_1 _23018_ (.Y(_05316_),
    .B1(net528),
    .B2(\cpu.dcache.r_data[6][25] ),
    .A2(net439),
    .A1(\cpu.dcache.r_data[1][25] ));
 sg13g2_and3_1 _23019_ (.X(_05317_),
    .A(_05314_),
    .B(_05315_),
    .C(_05316_));
 sg13g2_o21ai_1 _23020_ (.B1(_05317_),
    .Y(_05318_),
    .A1(_00092_),
    .A2(net433));
 sg13g2_nor2_1 _23021_ (.A(_10170_),
    .B(net654),
    .Y(_05319_));
 sg13g2_a22oi_1 _23022_ (.Y(_05320_),
    .B1(_05293_),
    .B2(_05319_),
    .A2(_05318_),
    .A1(net654));
 sg13g2_nor2_1 _23023_ (.A(net975),
    .B(_05320_),
    .Y(_05321_));
 sg13g2_nor3_1 _23024_ (.A(net514),
    .B(_05310_),
    .C(_05321_),
    .Y(_05322_));
 sg13g2_a21oi_1 _23025_ (.A1(_05111_),
    .A2(_05301_),
    .Y(_05323_),
    .B1(_05322_));
 sg13g2_mux2_1 _23026_ (.A0(_12049_),
    .A1(_12054_),
    .S(net899),
    .X(_05324_));
 sg13g2_a22oi_1 _23027_ (.Y(_05325_),
    .B1(net429),
    .B2(_05324_),
    .A2(net430),
    .A1(\cpu.spi.r_timeout[1] ));
 sg13g2_buf_1 _23028_ (.A(\cpu.spi.r_clk_count[2][1] ),
    .X(_05326_));
 sg13g2_nand2_1 _23029_ (.Y(_05327_),
    .A(_05326_),
    .B(_04915_));
 sg13g2_inv_1 _23030_ (.Y(_05328_),
    .A(_00095_));
 sg13g2_nor2_1 _23031_ (.A(_00094_),
    .B(_04919_),
    .Y(_05329_));
 sg13g2_a21oi_1 _23032_ (.A1(_05328_),
    .A2(net383),
    .Y(_05330_),
    .B1(_05329_));
 sg13g2_nand3_1 _23033_ (.B(_05327_),
    .C(_05330_),
    .A(_05325_),
    .Y(_05331_));
 sg13g2_a221oi_1 _23034_ (.B2(_09416_),
    .C1(_05331_),
    .B1(_04897_),
    .A1(_12050_),
    .Y(_05332_),
    .A2(_04885_));
 sg13g2_a22oi_1 _23035_ (.Y(_05333_),
    .B1(net382),
    .B2(_09329_),
    .A2(_04907_),
    .A1(\cpu.uart.r_div_value[1] ));
 sg13g2_a22oi_1 _23036_ (.Y(_05334_),
    .B1(_04932_),
    .B2(\cpu.uart.r_r_invert ),
    .A2(_04930_),
    .A1(\cpu.uart.r_div_value[9] ));
 sg13g2_nand2_1 _23037_ (.Y(_05335_),
    .A(_05333_),
    .B(_05334_));
 sg13g2_a21oi_1 _23038_ (.A1(\cpu.uart.r_in[1] ),
    .A2(_04928_),
    .Y(_05336_),
    .B1(_05335_));
 sg13g2_o21ai_1 _23039_ (.B1(net1011),
    .Y(_05337_),
    .A1(_04926_),
    .A2(_05336_));
 sg13g2_nand3_1 _23040_ (.B(_09302_),
    .C(_04979_),
    .A(_09301_),
    .Y(_05338_));
 sg13g2_nor2b_1 _23041_ (.A(_00100_),
    .B_N(_04983_),
    .Y(_05339_));
 sg13g2_a22oi_1 _23042_ (.Y(_05340_),
    .B1(net380),
    .B2(_09301_),
    .A2(_04992_),
    .A1(_09302_));
 sg13g2_inv_1 _23043_ (.Y(_05341_),
    .A(_00098_));
 sg13g2_buf_2 _23044_ (.A(\cpu.gpio.r_src_io[4][1] ),
    .X(_05342_));
 sg13g2_a22oi_1 _23045_ (.Y(_05343_),
    .B1(net428),
    .B2(_05342_),
    .A2(_04986_),
    .A1(_05341_));
 sg13g2_nand2_1 _23046_ (.Y(_05344_),
    .A(_05340_),
    .B(_05343_));
 sg13g2_nand2_1 _23047_ (.Y(_05345_),
    .A(_11383_),
    .B(_05033_));
 sg13g2_buf_2 _23048_ (.A(_05345_),
    .X(_05346_));
 sg13g2_nor2_1 _23049_ (.A(_00099_),
    .B(_05346_),
    .Y(_05347_));
 sg13g2_nand2b_1 _23050_ (.Y(_05348_),
    .B(net427),
    .A_N(_00096_));
 sg13g2_o21ai_1 _23051_ (.B1(_05348_),
    .Y(_05349_),
    .A1(_00097_),
    .A2(_05002_));
 sg13g2_nor4_1 _23052_ (.A(_05339_),
    .B(_05344_),
    .C(_05347_),
    .D(_05349_),
    .Y(_05350_));
 sg13g2_a21oi_1 _23053_ (.A1(_05338_),
    .A2(_05350_),
    .Y(_05351_),
    .B1(_05011_));
 sg13g2_a21o_1 _23054_ (.A2(net264),
    .A1(_09325_),
    .B1(net381),
    .X(_05352_));
 sg13g2_nand2_1 _23055_ (.Y(_05353_),
    .A(\cpu.intr.r_clock_cmp[1] ),
    .B(net652));
 sg13g2_a22oi_1 _23056_ (.Y(_05354_),
    .B1(net485),
    .B2(_10104_),
    .A2(net486),
    .A1(\cpu.intr.r_clock_cmp[17] ));
 sg13g2_nand2b_1 _23057_ (.Y(_05355_),
    .B(net662),
    .A_N(_05354_));
 sg13g2_nand2_1 _23058_ (.Y(_05356_),
    .A(net787),
    .B(\cpu.intr.r_timer_reload[17] ));
 sg13g2_nand2_1 _23059_ (.Y(_05357_),
    .A(net933),
    .B(\cpu.intr.r_timer_reload[1] ));
 sg13g2_a21oi_1 _23060_ (.A1(_05356_),
    .A2(_05357_),
    .Y(_05358_),
    .B1(_10178_));
 sg13g2_a221oi_1 _23061_ (.B2(_10261_),
    .C1(_05358_),
    .B1(_05035_),
    .A1(_09325_),
    .Y(_05359_),
    .A2(net382));
 sg13g2_buf_1 _23062_ (.A(\cpu.intr.r_clock_count[17] ),
    .X(_05360_));
 sg13g2_a22oi_1 _23063_ (.Y(_05361_),
    .B1(_05033_),
    .B2(_10092_),
    .A2(net443),
    .A1(_05360_));
 sg13g2_nand4_1 _23064_ (.B(_05355_),
    .C(_05359_),
    .A(_05353_),
    .Y(_05362_),
    .D(_05361_));
 sg13g2_a21oi_1 _23065_ (.A1(\cpu.intr.r_clock ),
    .A2(_05352_),
    .Y(_05363_),
    .B1(_05362_));
 sg13g2_nor2_1 _23066_ (.A(net683),
    .B(_05363_),
    .Y(_05364_));
 sg13g2_nor3_1 _23067_ (.A(_05337_),
    .B(_05351_),
    .C(_05364_),
    .Y(_05365_));
 sg13g2_o21ai_1 _23068_ (.B1(_05365_),
    .Y(_05366_),
    .A1(_09283_),
    .A2(_05332_));
 sg13g2_o21ai_1 _23069_ (.B1(_05366_),
    .Y(_05367_),
    .A1(net891),
    .A2(_05323_));
 sg13g2_nor2_1 _23070_ (.A(net83),
    .B(_05367_),
    .Y(_05368_));
 sg13g2_a21oi_1 _23071_ (.A1(_10246_),
    .A2(net63),
    .Y(_05369_),
    .B1(_05368_));
 sg13g2_nand2_1 _23072_ (.Y(_05370_),
    .A(_11524_),
    .B(_04817_));
 sg13g2_o21ai_1 _23073_ (.B1(_05370_),
    .Y(_05371_),
    .A1(_04817_),
    .A2(_04132_));
 sg13g2_mux2_1 _23074_ (.A0(net809),
    .A1(_05371_),
    .S(net215),
    .X(_05372_));
 sg13g2_nand2_1 _23075_ (.Y(_05373_),
    .A(net82),
    .B(_05372_));
 sg13g2_o21ai_1 _23076_ (.B1(_05373_),
    .Y(_01038_),
    .A1(net85),
    .A2(_05369_));
 sg13g2_a22oi_1 _23077_ (.Y(_05374_),
    .B1(_02732_),
    .B2(\cpu.dcache.r_data[6][18] ),
    .A2(net604),
    .A1(\cpu.dcache.r_data[5][18] ));
 sg13g2_nand2_1 _23078_ (.Y(_05375_),
    .A(\cpu.dcache.r_data[7][18] ),
    .B(net621));
 sg13g2_a22oi_1 _23079_ (.Y(_05376_),
    .B1(net488),
    .B2(\cpu.dcache.r_data[2][18] ),
    .A2(_10234_),
    .A1(\cpu.dcache.r_data[4][18] ));
 sg13g2_nor2_1 _23080_ (.A(_00101_),
    .B(net548),
    .Y(_05377_));
 sg13g2_a221oi_1 _23081_ (.B2(\cpu.dcache.r_data[3][18] ),
    .C1(_05377_),
    .B1(_12569_),
    .A1(\cpu.dcache.r_data[1][18] ),
    .Y(_05378_),
    .A2(net489));
 sg13g2_nand4_1 _23082_ (.B(_05375_),
    .C(_05376_),
    .A(_05374_),
    .Y(_05379_),
    .D(_05378_));
 sg13g2_buf_1 _23083_ (.A(_05379_),
    .X(_05380_));
 sg13g2_a22oi_1 _23084_ (.Y(_05381_),
    .B1(_05319_),
    .B2(_05380_),
    .A2(_05118_),
    .A1(net654));
 sg13g2_mux2_1 _23085_ (.A0(\cpu.dcache.r_data[4][2] ),
    .A1(\cpu.dcache.r_data[6][2] ),
    .S(net551),
    .X(_05382_));
 sg13g2_a22oi_1 _23086_ (.Y(_05383_),
    .B1(_05382_),
    .B2(net806),
    .A2(_09625_),
    .A1(\cpu.dcache.r_data[5][2] ));
 sg13g2_a22oi_1 _23087_ (.Y(_05384_),
    .B1(_12458_),
    .B2(\cpu.dcache.r_data[2][2] ),
    .A2(net627),
    .A1(\cpu.dcache.r_data[3][2] ));
 sg13g2_a22oi_1 _23088_ (.Y(_05385_),
    .B1(_10118_),
    .B2(\cpu.dcache.r_data[7][2] ),
    .A2(net547),
    .A1(\cpu.dcache.r_data[1][2] ));
 sg13g2_nand2_1 _23089_ (.Y(_05386_),
    .A(_05384_),
    .B(_05385_));
 sg13g2_a21oi_1 _23090_ (.A1(\cpu.dcache.r_data[0][2] ),
    .A2(_09769_),
    .Y(_05387_),
    .B1(_05386_));
 sg13g2_o21ai_1 _23091_ (.B1(_05387_),
    .Y(_05388_),
    .A1(_09495_),
    .A2(_05383_));
 sg13g2_a22oi_1 _23092_ (.Y(_05389_),
    .B1(_05388_),
    .B2(_05067_),
    .A2(_05308_),
    .A1(_05124_));
 sg13g2_o21ai_1 _23093_ (.B1(_05389_),
    .Y(_05390_),
    .A1(net975),
    .A2(_05381_));
 sg13g2_mux2_1 _23094_ (.A0(_05380_),
    .A1(_05388_),
    .S(net682),
    .X(_05391_));
 sg13g2_mux2_1 _23095_ (.A0(_05390_),
    .A1(_05391_),
    .S(_05111_),
    .X(_05392_));
 sg13g2_inv_1 _23096_ (.Y(_05393_),
    .A(_00105_));
 sg13g2_buf_1 _23097_ (.A(\cpu.spi.r_clk_count[2][2] ),
    .X(_05394_));
 sg13g2_nand2_1 _23098_ (.Y(_05395_),
    .A(net899),
    .B(_12035_));
 sg13g2_o21ai_1 _23099_ (.B1(_05395_),
    .Y(_05396_),
    .A1(net899),
    .A2(_00282_));
 sg13g2_a22oi_1 _23100_ (.Y(_05397_),
    .B1(_04907_),
    .B2(_05396_),
    .A2(net430),
    .A1(\cpu.spi.r_timeout[2] ));
 sg13g2_o21ai_1 _23101_ (.B1(_05397_),
    .Y(_05398_),
    .A1(_00104_),
    .A2(_04919_));
 sg13g2_a221oi_1 _23102_ (.B2(_05394_),
    .C1(_05398_),
    .B1(_04915_),
    .A1(_05393_),
    .Y(_05399_),
    .A2(net383));
 sg13g2_o21ai_1 _23103_ (.B1(_05399_),
    .Y(_05400_),
    .A1(_00283_),
    .A2(_05346_));
 sg13g2_a21oi_1 _23104_ (.A1(_09420_),
    .A2(_04897_),
    .Y(_05401_),
    .B1(_05400_));
 sg13g2_nand3_1 _23105_ (.B(_09308_),
    .C(_04979_),
    .A(_09307_),
    .Y(_05402_));
 sg13g2_nand2b_1 _23106_ (.Y(_05403_),
    .B(_04983_),
    .A_N(_00110_));
 sg13g2_buf_1 _23107_ (.A(\cpu.gpio.r_src_io[4][2] ),
    .X(_05404_));
 sg13g2_nand2b_1 _23108_ (.Y(_05405_),
    .B(net427),
    .A_N(_00106_));
 sg13g2_o21ai_1 _23109_ (.B1(_05405_),
    .Y(_05406_),
    .A1(_00107_),
    .A2(net343));
 sg13g2_a221oi_1 _23110_ (.B2(_09308_),
    .C1(_05406_),
    .B1(_04992_),
    .A1(_05404_),
    .Y(_05407_),
    .A2(net428));
 sg13g2_inv_1 _23111_ (.Y(_05408_),
    .A(_00108_));
 sg13g2_nor2_1 _23112_ (.A(_00109_),
    .B(_05346_),
    .Y(_05409_));
 sg13g2_a221oi_1 _23113_ (.B2(_09307_),
    .C1(_05409_),
    .B1(net380),
    .A1(_05408_),
    .Y(_05410_),
    .A2(_04986_));
 sg13g2_nand4_1 _23114_ (.B(_05403_),
    .C(_05407_),
    .A(_05402_),
    .Y(_05411_),
    .D(_05410_));
 sg13g2_nor2b_1 _23115_ (.A(_05011_),
    .B_N(_05411_),
    .Y(_05412_));
 sg13g2_a21o_1 _23116_ (.A2(net264),
    .A1(_09321_),
    .B1(_04939_),
    .X(_05413_));
 sg13g2_mux2_1 _23117_ (.A0(\cpu.intr.r_clock_cmp[2] ),
    .A1(\cpu.intr.r_clock_cmp[18] ),
    .S(net787),
    .X(_05414_));
 sg13g2_a22oi_1 _23118_ (.Y(_05415_),
    .B1(_05414_),
    .B2(net486),
    .A2(net381),
    .A1(_09321_));
 sg13g2_buf_2 _23119_ (.A(\cpu.intr.r_clock_count[18] ),
    .X(_05416_));
 sg13g2_mux2_1 _23120_ (.A0(\cpu.intr.r_timer_count[2] ),
    .A1(_10107_),
    .S(net787),
    .X(_05417_));
 sg13g2_a22oi_1 _23121_ (.Y(_05418_),
    .B1(_05417_),
    .B2(net435),
    .A2(net443),
    .A1(_05416_));
 sg13g2_a22oi_1 _23122_ (.Y(_05419_),
    .B1(net494),
    .B2(\cpu.intr.r_timer_reload[2] ),
    .A2(net444),
    .A1(_10265_));
 sg13g2_or2_1 _23123_ (.X(_05420_),
    .B(_05419_),
    .A(net662));
 sg13g2_nand3_1 _23124_ (.B(\cpu.intr.r_timer_reload[18] ),
    .C(net445),
    .A(net662),
    .Y(_05421_));
 sg13g2_nand4_1 _23125_ (.B(_05418_),
    .C(_05420_),
    .A(_05415_),
    .Y(_05422_),
    .D(_05421_));
 sg13g2_a21oi_1 _23126_ (.A1(\cpu.intr.r_enable[2] ),
    .A2(_05413_),
    .Y(_05423_),
    .B1(_05422_));
 sg13g2_nor2_1 _23127_ (.A(net683),
    .B(_05423_),
    .Y(_05424_));
 sg13g2_and2_1 _23128_ (.A(_10080_),
    .B(_04930_),
    .X(_05425_));
 sg13g2_a221oi_1 _23129_ (.B2(\cpu.uart.r_in[2] ),
    .C1(_05425_),
    .B1(_04928_),
    .A1(\cpu.uart.r_div_value[2] ),
    .Y(_05426_),
    .A2(net429));
 sg13g2_o21ai_1 _23130_ (.B1(net1011),
    .Y(_05427_),
    .A1(_04926_),
    .A2(_05426_));
 sg13g2_nor3_1 _23131_ (.A(_05412_),
    .B(_05424_),
    .C(_05427_),
    .Y(_05428_));
 sg13g2_o21ai_1 _23132_ (.B1(_05428_),
    .Y(_05429_),
    .A1(net709),
    .A2(_05401_));
 sg13g2_o21ai_1 _23133_ (.B1(_05429_),
    .Y(_05430_),
    .A1(net891),
    .A2(_05392_));
 sg13g2_nor2_1 _23134_ (.A(net63),
    .B(_05430_),
    .Y(_05431_));
 sg13g2_a21oi_1 _23135_ (.A1(net475),
    .A2(net63),
    .Y(_05432_),
    .B1(_05431_));
 sg13g2_o21ai_1 _23136_ (.B1(net215),
    .Y(_05433_),
    .A1(net809),
    .A2(_11682_));
 sg13g2_buf_1 _23137_ (.A(_04817_),
    .X(_05434_));
 sg13g2_nand3_1 _23138_ (.B(net809),
    .C(net651),
    .A(net822),
    .Y(_05435_));
 sg13g2_o21ai_1 _23139_ (.B1(_05435_),
    .Y(_05436_),
    .A1(net651),
    .A2(_04470_));
 sg13g2_a221oi_1 _23140_ (.B2(net189),
    .C1(net98),
    .B1(_05436_),
    .A1(net712),
    .Y(_05437_),
    .A2(_05433_));
 sg13g2_a21oi_1 _23141_ (.A1(_05143_),
    .A2(_05432_),
    .Y(_01039_),
    .B1(_05437_));
 sg13g2_nand2_1 _23142_ (.Y(_05438_),
    .A(net651),
    .B(_04214_));
 sg13g2_o21ai_1 _23143_ (.B1(_05438_),
    .Y(_05439_),
    .A1(net651),
    .A2(_04502_));
 sg13g2_a21oi_1 _23144_ (.A1(net651),
    .A2(_04212_),
    .Y(_05440_),
    .B1(net398));
 sg13g2_nor2_1 _23145_ (.A(net711),
    .B(_05440_),
    .Y(_05441_));
 sg13g2_a21oi_1 _23146_ (.A1(_05173_),
    .A2(_05439_),
    .Y(_05442_),
    .B1(_05441_));
 sg13g2_mux2_1 _23147_ (.A0(\cpu.dcache.r_data[5][3] ),
    .A1(\cpu.dcache.r_data[7][3] ),
    .S(net496),
    .X(_05443_));
 sg13g2_a22oi_1 _23148_ (.Y(_05444_),
    .B1(_05443_),
    .B2(_12557_),
    .A2(net759),
    .A1(\cpu.dcache.r_data[6][3] ));
 sg13g2_a22oi_1 _23149_ (.Y(_05445_),
    .B1(_12458_),
    .B2(\cpu.dcache.r_data[2][3] ),
    .A2(net439),
    .A1(\cpu.dcache.r_data[1][3] ));
 sg13g2_a22oi_1 _23150_ (.Y(_05446_),
    .B1(_10234_),
    .B2(\cpu.dcache.r_data[4][3] ),
    .A2(_12569_),
    .A1(\cpu.dcache.r_data[3][3] ));
 sg13g2_nand2_1 _23151_ (.Y(_05447_),
    .A(_05445_),
    .B(_05446_));
 sg13g2_a21oi_1 _23152_ (.A1(\cpu.dcache.r_data[0][3] ),
    .A2(_09769_),
    .Y(_05448_),
    .B1(_05447_));
 sg13g2_o21ai_1 _23153_ (.B1(_05448_),
    .Y(_05449_),
    .A1(_12062_),
    .A2(_05444_));
 sg13g2_mux2_1 _23154_ (.A0(\cpu.dcache.r_data[4][19] ),
    .A1(\cpu.dcache.r_data[6][19] ),
    .S(_09344_),
    .X(_05450_));
 sg13g2_a22oi_1 _23155_ (.Y(_05451_),
    .B1(_05450_),
    .B2(net806),
    .A2(_09625_),
    .A1(\cpu.dcache.r_data[5][19] ));
 sg13g2_nand2b_1 _23156_ (.Y(_05452_),
    .B(net785),
    .A_N(_05451_));
 sg13g2_a22oi_1 _23157_ (.Y(_05453_),
    .B1(net468),
    .B2(\cpu.dcache.r_data[3][19] ),
    .A2(net439),
    .A1(\cpu.dcache.r_data[1][19] ));
 sg13g2_a22oi_1 _23158_ (.Y(_05454_),
    .B1(_10119_),
    .B2(\cpu.dcache.r_data[7][19] ),
    .A2(_04835_),
    .A1(\cpu.dcache.r_data[2][19] ));
 sg13g2_and3_1 _23159_ (.X(_05455_),
    .A(_05452_),
    .B(_05453_),
    .C(_05454_));
 sg13g2_o21ai_1 _23160_ (.B1(_05455_),
    .Y(_05456_),
    .A1(_00111_),
    .A2(_04831_));
 sg13g2_nor2_1 _23161_ (.A(_10170_),
    .B(_12120_),
    .Y(_05457_));
 sg13g2_a221oi_1 _23162_ (.B2(_05457_),
    .C1(net654),
    .B1(_05456_),
    .A1(net975),
    .Y(_05458_),
    .A2(_05449_));
 sg13g2_a221oi_1 _23163_ (.B2(_12152_),
    .C1(_04849_),
    .B1(_05159_),
    .A1(net682),
    .Y(_05459_),
    .A2(_05151_));
 sg13g2_nor3_1 _23164_ (.A(_04866_),
    .B(_05458_),
    .C(_05459_),
    .Y(_05460_));
 sg13g2_nor2_1 _23165_ (.A(net682),
    .B(_05456_),
    .Y(_05461_));
 sg13g2_nor2_1 _23166_ (.A(net618),
    .B(_05449_),
    .Y(_05462_));
 sg13g2_nor3_1 _23167_ (.A(_04863_),
    .B(_05461_),
    .C(_05462_),
    .Y(_05463_));
 sg13g2_nor3_1 _23168_ (.A(net891),
    .B(_05460_),
    .C(_05463_),
    .Y(_05464_));
 sg13g2_buf_1 _23169_ (.A(\cpu.gpio.r_src_io[4][3] ),
    .X(_05465_));
 sg13g2_a22oi_1 _23170_ (.Y(_05466_),
    .B1(_04992_),
    .B2(_09297_),
    .A2(net428),
    .A1(_05465_));
 sg13g2_inv_1 _23171_ (.Y(_05467_),
    .A(_00118_));
 sg13g2_a22oi_1 _23172_ (.Y(_05468_),
    .B1(net380),
    .B2(_09296_),
    .A2(_04986_),
    .A1(_05467_));
 sg13g2_nand2_1 _23173_ (.Y(_05469_),
    .A(_05466_),
    .B(_05468_));
 sg13g2_nand2b_1 _23174_ (.Y(_05470_),
    .B(net427),
    .A_N(_00116_));
 sg13g2_o21ai_1 _23175_ (.B1(_05470_),
    .Y(_05471_),
    .A1(_00117_),
    .A2(net343));
 sg13g2_inv_1 _23176_ (.Y(_05472_),
    .A(_00119_));
 sg13g2_a22oi_1 _23177_ (.Y(_05473_),
    .B1(net467),
    .B2(\cpu.gpio.genblk1[3].srcs_o[0] ),
    .A2(_05131_),
    .A1(_05472_));
 sg13g2_nor2_1 _23178_ (.A(net872),
    .B(_05473_),
    .Y(_05474_));
 sg13g2_nor3_1 _23179_ (.A(_05469_),
    .B(_05471_),
    .C(_05474_),
    .Y(_05475_));
 sg13g2_nand3_1 _23180_ (.B(_09297_),
    .C(_04979_),
    .A(_09296_),
    .Y(_05476_));
 sg13g2_a21oi_1 _23181_ (.A1(_05475_),
    .A2(_05476_),
    .Y(_05477_),
    .B1(_05011_));
 sg13g2_inv_1 _23182_ (.Y(_05478_),
    .A(_00115_));
 sg13g2_buf_1 _23183_ (.A(\cpu.spi.r_clk_count[2][3] ),
    .X(_05479_));
 sg13g2_nand2_1 _23184_ (.Y(_05480_),
    .A(\cpu.spi.r_timeout[3] ),
    .B(net430));
 sg13g2_o21ai_1 _23185_ (.B1(_05480_),
    .Y(_05481_),
    .A1(_00114_),
    .A2(_04919_));
 sg13g2_a221oi_1 _23186_ (.B2(_05479_),
    .C1(_05481_),
    .B1(_04915_),
    .A1(_05478_),
    .Y(_05482_),
    .A2(net383));
 sg13g2_nand2_1 _23187_ (.Y(_05483_),
    .A(_09414_),
    .B(_04897_));
 sg13g2_a21oi_1 _23188_ (.A1(_05482_),
    .A2(_05483_),
    .Y(_05484_),
    .B1(net709));
 sg13g2_a22oi_1 _23189_ (.Y(_05485_),
    .B1(net435),
    .B2(_10108_),
    .A2(net445),
    .A1(\cpu.intr.r_timer_reload[19] ));
 sg13g2_inv_1 _23190_ (.Y(_05486_),
    .A(_05485_));
 sg13g2_a22oi_1 _23191_ (.Y(_05487_),
    .B1(_02734_),
    .B2(\cpu.intr.r_timer_count[3] ),
    .A2(_10121_),
    .A1(\cpu.intr.r_timer_reload[3] ));
 sg13g2_buf_2 _23192_ (.A(\cpu.intr.r_clock_count[19] ),
    .X(_05488_));
 sg13g2_nand2_1 _23193_ (.Y(_05489_),
    .A(net787),
    .B(\cpu.intr.r_clock_cmp[19] ));
 sg13g2_nand2_1 _23194_ (.Y(_05490_),
    .A(net933),
    .B(\cpu.intr.r_clock_cmp[3] ));
 sg13g2_a21oi_1 _23195_ (.A1(_05489_),
    .A2(_05490_),
    .Y(_05491_),
    .B1(_09836_));
 sg13g2_a221oi_1 _23196_ (.B2(_09326_),
    .C1(_05491_),
    .B1(net381),
    .A1(_05488_),
    .Y(_05492_),
    .A2(net443));
 sg13g2_o21ai_1 _23197_ (.B1(_05492_),
    .Y(_05493_),
    .A1(net684),
    .A2(_05487_));
 sg13g2_a221oi_1 _23198_ (.B2(net618),
    .C1(_05493_),
    .B1(_05486_),
    .A1(_10270_),
    .Y(_05494_),
    .A2(net467));
 sg13g2_a21oi_1 _23199_ (.A1(_09326_),
    .A2(net264),
    .Y(_05495_),
    .B1(_04939_));
 sg13g2_nand2b_1 _23200_ (.Y(_05496_),
    .B(\cpu.intr.r_enable[3] ),
    .A_N(_05495_));
 sg13g2_a21oi_1 _23201_ (.A1(_05494_),
    .A2(_05496_),
    .Y(_05497_),
    .B1(net683));
 sg13g2_and2_1 _23202_ (.A(\cpu.uart.r_div_value[11] ),
    .B(_04930_),
    .X(_05498_));
 sg13g2_a221oi_1 _23203_ (.B2(\cpu.uart.r_in[3] ),
    .C1(_05498_),
    .B1(_04928_),
    .A1(\cpu.uart.r_div_value[3] ),
    .Y(_05499_),
    .A2(net429));
 sg13g2_o21ai_1 _23204_ (.B1(net1011),
    .Y(_05500_),
    .A1(_04926_),
    .A2(_05499_));
 sg13g2_nor4_1 _23205_ (.A(_05477_),
    .B(_05484_),
    .C(_05497_),
    .D(_05500_),
    .Y(_05501_));
 sg13g2_nor3_1 _23206_ (.A(net84),
    .B(_05464_),
    .C(_05501_),
    .Y(_05502_));
 sg13g2_a21oi_1 _23207_ (.A1(_12558_),
    .A2(net83),
    .Y(_05503_),
    .B1(_05502_));
 sg13g2_nor2_1 _23208_ (.A(net82),
    .B(_05503_),
    .Y(_05504_));
 sg13g2_a21o_1 _23209_ (.A2(_05442_),
    .A1(net85),
    .B1(_05504_),
    .X(_01040_));
 sg13g2_o21ai_1 _23210_ (.B1(_04822_),
    .Y(_05505_),
    .A1(net762),
    .A2(_04214_));
 sg13g2_nand3_1 _23211_ (.B(_04817_),
    .C(_04214_),
    .A(net1127),
    .Y(_05506_));
 sg13g2_o21ai_1 _23212_ (.B1(_05506_),
    .Y(_05507_),
    .A1(net651),
    .A2(_04545_));
 sg13g2_a22oi_1 _23213_ (.Y(_05508_),
    .B1(_05507_),
    .B2(_05173_),
    .A2(_05505_),
    .A1(_08562_));
 sg13g2_a21oi_1 _23214_ (.A1(_12152_),
    .A2(_05182_),
    .Y(_05509_),
    .B1(_05190_));
 sg13g2_a22oi_1 _23215_ (.Y(_05510_),
    .B1(_02731_),
    .B2(\cpu.dcache.r_data[6][20] ),
    .A2(net530),
    .A1(\cpu.dcache.r_data[3][20] ));
 sg13g2_a22oi_1 _23216_ (.Y(_05511_),
    .B1(_12780_),
    .B2(\cpu.dcache.r_data[5][20] ),
    .A2(_10118_),
    .A1(\cpu.dcache.r_data[7][20] ));
 sg13g2_a22oi_1 _23217_ (.Y(_05512_),
    .B1(net549),
    .B2(\cpu.dcache.r_data[2][20] ),
    .A2(net626),
    .A1(\cpu.dcache.r_data[4][20] ));
 sg13g2_nand3_1 _23218_ (.B(_05511_),
    .C(_05512_),
    .A(_05510_),
    .Y(_05513_));
 sg13g2_nand2_1 _23219_ (.Y(_05514_),
    .A(_00122_),
    .B(net586));
 sg13g2_o21ai_1 _23220_ (.B1(_05514_),
    .Y(_05515_),
    .A1(net586),
    .A2(_05513_));
 sg13g2_o21ai_1 _23221_ (.B1(net389),
    .Y(_05516_),
    .A1(\cpu.dcache.r_data[1][20] ),
    .A2(_05513_));
 sg13g2_o21ai_1 _23222_ (.B1(_05516_),
    .Y(_05517_),
    .A1(net389),
    .A2(_05515_));
 sg13g2_nand2_1 _23223_ (.Y(_05518_),
    .A(_05319_),
    .B(_05517_));
 sg13g2_o21ai_1 _23224_ (.B1(_05518_),
    .Y(_05519_),
    .A1(_04849_),
    .A2(_05509_));
 sg13g2_a22oi_1 _23225_ (.Y(_05520_),
    .B1(net438),
    .B2(\cpu.dcache.r_data[2][4] ),
    .A2(net431),
    .A1(\cpu.dcache.r_data[1][4] ));
 sg13g2_a22oi_1 _23226_ (.Y(_05521_),
    .B1(net493),
    .B2(\cpu.dcache.r_data[4][4] ),
    .A2(net487),
    .A1(\cpu.dcache.r_data[3][4] ));
 sg13g2_mux2_1 _23227_ (.A0(\cpu.dcache.r_data[5][4] ),
    .A1(\cpu.dcache.r_data[7][4] ),
    .S(net551),
    .X(_05522_));
 sg13g2_a22oi_1 _23228_ (.Y(_05523_),
    .B1(_05522_),
    .B2(_10174_),
    .A2(net759),
    .A1(\cpu.dcache.r_data[6][4] ));
 sg13g2_nand2b_1 _23229_ (.Y(_05524_),
    .B(_10176_),
    .A_N(_05523_));
 sg13g2_and4_1 _23230_ (.A(net433),
    .B(_05520_),
    .C(_05521_),
    .D(_05524_),
    .X(_05525_));
 sg13g2_a21oi_1 _23231_ (.A1(_00121_),
    .A2(net546),
    .Y(_05526_),
    .B1(_05525_));
 sg13g2_and2_1 _23232_ (.A(_05067_),
    .B(_05526_),
    .X(_05527_));
 sg13g2_a21oi_1 _23233_ (.A1(_04877_),
    .A2(_05519_),
    .Y(_05528_),
    .B1(_05527_));
 sg13g2_mux2_1 _23234_ (.A0(_05526_),
    .A1(_05517_),
    .S(_10117_),
    .X(_05529_));
 sg13g2_nand2_1 _23235_ (.Y(_05530_),
    .A(_04866_),
    .B(_05529_));
 sg13g2_o21ai_1 _23236_ (.B1(_05530_),
    .Y(_05531_),
    .A1(net514),
    .A2(_05528_));
 sg13g2_nor2_1 _23237_ (.A(net891),
    .B(_05531_),
    .Y(_05532_));
 sg13g2_nand3_1 _23238_ (.B(_09304_),
    .C(_04979_),
    .A(_09303_),
    .Y(_05533_));
 sg13g2_buf_2 _23239_ (.A(\cpu.gpio.r_src_o[5][0] ),
    .X(_05534_));
 sg13g2_a22oi_1 _23240_ (.Y(_05535_),
    .B1(net652),
    .B2(net7),
    .A2(net443),
    .A1(\cpu.gpio.genblk2[4].srcs_io[0] ));
 sg13g2_inv_1 _23241_ (.Y(_05536_),
    .A(_05535_));
 sg13g2_nand3_1 _23242_ (.B(\cpu.gpio.genblk1[4].srcs_o[0] ),
    .C(_05035_),
    .A(net977),
    .Y(_05537_));
 sg13g2_and3_1 _23243_ (.X(_05538_),
    .A(_09292_),
    .B(net977),
    .C(net381));
 sg13g2_o21ai_1 _23244_ (.B1(\cpu.gpio.r_enable_io[4] ),
    .Y(_05539_),
    .A1(net383),
    .A2(_05538_));
 sg13g2_buf_2 _23245_ (.A(\cpu.gpio.r_spi_miso_src[1][0] ),
    .X(_05540_));
 sg13g2_buf_2 _23246_ (.A(\cpu.gpio.r_src_o[3][0] ),
    .X(_05541_));
 sg13g2_and3_1 _23247_ (.X(_05542_),
    .A(_12057_),
    .B(_05541_),
    .C(net381));
 sg13g2_a221oi_1 _23248_ (.B2(_09303_),
    .C1(_05542_),
    .B1(net380),
    .A1(_05540_),
    .Y(_05543_),
    .A2(_04983_));
 sg13g2_buf_2 _23249_ (.A(\cpu.gpio.r_src_io[5][0] ),
    .X(_05544_));
 sg13g2_buf_2 _23250_ (.A(\cpu.gpio.r_src_o[7][0] ),
    .X(_05545_));
 sg13g2_a22oi_1 _23251_ (.Y(_05546_),
    .B1(_05545_),
    .B2(net899),
    .A2(net977),
    .A1(_09292_));
 sg13g2_buf_2 _23252_ (.A(\cpu.gpio.r_src_io[7][0] ),
    .X(_05547_));
 sg13g2_nand2_1 _23253_ (.Y(_05548_),
    .A(_05547_),
    .B(net427));
 sg13g2_o21ai_1 _23254_ (.B1(_05548_),
    .Y(_05549_),
    .A1(_05058_),
    .A2(_05546_));
 sg13g2_a221oi_1 _23255_ (.B2(_09304_),
    .C1(_05549_),
    .B1(_04992_),
    .A1(_05544_),
    .Y(_05550_),
    .A2(_04988_));
 sg13g2_nand4_1 _23256_ (.B(_05539_),
    .C(_05543_),
    .A(_05537_),
    .Y(_05551_),
    .D(_05550_));
 sg13g2_a221oi_1 _23257_ (.B2(_04913_),
    .C1(_05551_),
    .B1(_05536_),
    .A1(_05534_),
    .Y(_05552_),
    .A2(_04986_));
 sg13g2_a21oi_1 _23258_ (.A1(_05533_),
    .A2(_05552_),
    .Y(_05553_),
    .B1(_05011_));
 sg13g2_mux2_1 _23259_ (.A0(\cpu.intr.r_clock_cmp[20] ),
    .A1(\cpu.intr.r_timer_reload[20] ),
    .S(_09345_),
    .X(_05554_));
 sg13g2_a22oi_1 _23260_ (.Y(_05555_),
    .B1(_05554_),
    .B2(net531),
    .A2(net759),
    .A1(_10109_));
 sg13g2_nor3_1 _23261_ (.A(net786),
    .B(net760),
    .C(_05555_),
    .Y(_05556_));
 sg13g2_a22oi_1 _23262_ (.Y(_05557_),
    .B1(net485),
    .B2(\cpu.intr.r_timer_count[4] ),
    .A2(net494),
    .A1(\cpu.intr.r_timer_reload[4] ));
 sg13g2_nor2_1 _23263_ (.A(net787),
    .B(_05557_),
    .Y(_05558_));
 sg13g2_buf_2 _23264_ (.A(\cpu.intr.r_clock_count[20] ),
    .X(_05559_));
 sg13g2_a221oi_1 _23265_ (.B2(_10277_),
    .C1(net264),
    .B1(_05035_),
    .A1(_05559_),
    .Y(_05560_),
    .A2(_10254_));
 sg13g2_a22oi_1 _23266_ (.Y(_05561_),
    .B1(net652),
    .B2(\cpu.intr.r_clock_cmp[4] ),
    .A2(_04938_),
    .A1(_09318_));
 sg13g2_nand2_1 _23267_ (.Y(_05562_),
    .A(_05560_),
    .B(_05561_));
 sg13g2_nor3_1 _23268_ (.A(_05556_),
    .B(_05558_),
    .C(_05562_),
    .Y(_05563_));
 sg13g2_nand2_2 _23269_ (.Y(_05564_),
    .A(net586),
    .B(net515));
 sg13g2_a221oi_1 _23270_ (.B2(_05564_),
    .C1(net683),
    .B1(_05563_),
    .A1(_09319_),
    .Y(_05565_),
    .A2(_04963_));
 sg13g2_nor2_1 _23271_ (.A(_11124_),
    .B(_11125_),
    .Y(_05566_));
 sg13g2_o21ai_1 _23272_ (.B1(_05566_),
    .Y(_05567_),
    .A1(net264),
    .A2(_05563_));
 sg13g2_and2_1 _23273_ (.A(_05565_),
    .B(_05567_),
    .X(_05568_));
 sg13g2_inv_1 _23274_ (.Y(_05569_),
    .A(_00126_));
 sg13g2_buf_1 _23275_ (.A(\cpu.spi.r_clk_count[2][4] ),
    .X(_05570_));
 sg13g2_nand2_1 _23276_ (.Y(_05571_),
    .A(\cpu.spi.r_timeout[4] ),
    .B(net430));
 sg13g2_o21ai_1 _23277_ (.B1(_05571_),
    .Y(_05572_),
    .A1(_00125_),
    .A2(_04919_));
 sg13g2_a221oi_1 _23278_ (.B2(_05570_),
    .C1(_05572_),
    .B1(_04915_),
    .A1(_05569_),
    .Y(_05573_),
    .A2(net383));
 sg13g2_nand2_1 _23279_ (.Y(_05574_),
    .A(_09422_),
    .B(_04897_));
 sg13g2_a21oi_1 _23280_ (.A1(_05573_),
    .A2(_05574_),
    .Y(_05575_),
    .B1(net709));
 sg13g2_a22oi_1 _23281_ (.Y(_05576_),
    .B1(_04928_),
    .B2(\cpu.uart.r_in[4] ),
    .A2(net429),
    .A1(\cpu.uart.r_div_value[4] ));
 sg13g2_o21ai_1 _23282_ (.B1(net1011),
    .Y(_05577_),
    .A1(_04926_),
    .A2(_05576_));
 sg13g2_nor4_1 _23283_ (.A(_05553_),
    .B(_05568_),
    .C(_05575_),
    .D(_05577_),
    .Y(_05578_));
 sg13g2_nor3_1 _23284_ (.A(net84),
    .B(_05532_),
    .C(_05578_),
    .Y(_05579_));
 sg13g2_a21oi_1 _23285_ (.A1(net524),
    .A2(net83),
    .Y(_05580_),
    .B1(_05579_));
 sg13g2_nor2_1 _23286_ (.A(net82),
    .B(_05580_),
    .Y(_05581_));
 sg13g2_a21o_1 _23287_ (.A2(_05508_),
    .A1(net85),
    .B1(_05581_),
    .X(_01041_));
 sg13g2_nand2_1 _23288_ (.Y(_05582_),
    .A(net651),
    .B(_04574_));
 sg13g2_o21ai_1 _23289_ (.B1(_05582_),
    .Y(_05583_),
    .A1(_05434_),
    .A2(_04572_));
 sg13g2_nor2_1 _23290_ (.A(net398),
    .B(_05583_),
    .Y(_05584_));
 sg13g2_o21ai_1 _23291_ (.B1(net82),
    .Y(_05585_),
    .A1(_08806_),
    .A2(net189));
 sg13g2_a22oi_1 _23292_ (.Y(_05586_),
    .B1(net493),
    .B2(\cpu.dcache.r_data[4][5] ),
    .A2(net487),
    .A1(\cpu.dcache.r_data[3][5] ));
 sg13g2_nand2_1 _23293_ (.Y(_05587_),
    .A(\cpu.dcache.r_data[7][5] ),
    .B(net494));
 sg13g2_a22oi_1 _23294_ (.Y(_05588_),
    .B1(net485),
    .B2(\cpu.dcache.r_data[6][5] ),
    .A2(net438),
    .A1(\cpu.dcache.r_data[2][5] ));
 sg13g2_nor2_1 _23295_ (.A(_00128_),
    .B(_04830_),
    .Y(_05589_));
 sg13g2_a221oi_1 _23296_ (.B2(\cpu.dcache.r_data[5][5] ),
    .C1(_05589_),
    .B1(net529),
    .A1(\cpu.dcache.r_data[1][5] ),
    .Y(_05590_),
    .A2(net431));
 sg13g2_nand4_1 _23297_ (.B(_05587_),
    .C(_05588_),
    .A(_05586_),
    .Y(_05591_),
    .D(_05590_));
 sg13g2_buf_1 _23298_ (.A(_05591_),
    .X(_05592_));
 sg13g2_nor2_1 _23299_ (.A(_00129_),
    .B(net433),
    .Y(_05593_));
 sg13g2_mux2_1 _23300_ (.A0(\cpu.dcache.r_data[5][21] ),
    .A1(\cpu.dcache.r_data[7][21] ),
    .S(_09344_),
    .X(_05594_));
 sg13g2_a22oi_1 _23301_ (.Y(_05595_),
    .B1(_05594_),
    .B2(net531),
    .A2(net689),
    .A1(\cpu.dcache.r_data[4][21] ));
 sg13g2_nor2_1 _23302_ (.A(net929),
    .B(_05595_),
    .Y(_05596_));
 sg13g2_a22oi_1 _23303_ (.Y(_05597_),
    .B1(_02733_),
    .B2(\cpu.dcache.r_data[6][21] ),
    .A2(net487),
    .A1(\cpu.dcache.r_data[3][21] ));
 sg13g2_a22oi_1 _23304_ (.Y(_05598_),
    .B1(net438),
    .B2(\cpu.dcache.r_data[2][21] ),
    .A2(_04844_),
    .A1(\cpu.dcache.r_data[1][21] ));
 sg13g2_nand2_1 _23305_ (.Y(_05599_),
    .A(_05597_),
    .B(_05598_));
 sg13g2_nor3_2 _23306_ (.A(_05593_),
    .B(_05596_),
    .C(_05599_),
    .Y(_05600_));
 sg13g2_nor2_1 _23307_ (.A(_10171_),
    .B(_05600_),
    .Y(_05601_));
 sg13g2_a21oi_1 _23308_ (.A1(net620),
    .A2(_05592_),
    .Y(_05602_),
    .B1(_05601_));
 sg13g2_nor2b_1 _23309_ (.A(_05600_),
    .B_N(_05457_),
    .Y(_05603_));
 sg13g2_a21oi_1 _23310_ (.A1(net975),
    .A2(_05592_),
    .Y(_05604_),
    .B1(_05603_));
 sg13g2_o21ai_1 _23311_ (.B1(_05229_),
    .Y(_05605_),
    .A1(_12120_),
    .A2(_05220_));
 sg13g2_nor2_1 _23312_ (.A(_04849_),
    .B(_05605_),
    .Y(_05606_));
 sg13g2_a21oi_1 _23313_ (.A1(_04849_),
    .A2(_05604_),
    .Y(_05607_),
    .B1(_05606_));
 sg13g2_nand2_1 _23314_ (.Y(_05608_),
    .A(_04863_),
    .B(_05607_));
 sg13g2_o21ai_1 _23315_ (.B1(_05608_),
    .Y(_05609_),
    .A1(_04863_),
    .A2(_05602_));
 sg13g2_buf_1 _23316_ (.A(\cpu.spi.r_clk_count[2][5] ),
    .X(_05610_));
 sg13g2_nand2b_1 _23317_ (.Y(_05611_),
    .B(net383),
    .A_N(_00133_));
 sg13g2_o21ai_1 _23318_ (.B1(_05611_),
    .Y(_05612_),
    .A1(_00132_),
    .A2(_04919_));
 sg13g2_a221oi_1 _23319_ (.B2(\cpu.spi.r_timeout[5] ),
    .C1(_05612_),
    .B1(net430),
    .A1(_05610_),
    .Y(_05613_),
    .A2(_04915_));
 sg13g2_nand2_1 _23320_ (.Y(_05614_),
    .A(_09421_),
    .B(_04897_));
 sg13g2_a21oi_1 _23321_ (.A1(_05613_),
    .A2(_05614_),
    .Y(_05615_),
    .B1(net709));
 sg13g2_a22oi_1 _23322_ (.Y(_05616_),
    .B1(_04928_),
    .B2(\cpu.uart.r_in[5] ),
    .A2(net429),
    .A1(\cpu.uart.r_div_value[5] ));
 sg13g2_nor2_1 _23323_ (.A(_04926_),
    .B(_05616_),
    .Y(_05617_));
 sg13g2_a21o_1 _23324_ (.A2(net264),
    .A1(_09323_),
    .B1(net381),
    .X(_05618_));
 sg13g2_a22oi_1 _23325_ (.Y(_05619_),
    .B1(net486),
    .B2(\cpu.intr.r_clock_cmp[5] ),
    .A2(net444),
    .A1(_10283_));
 sg13g2_mux2_1 _23326_ (.A0(\cpu.intr.r_timer_count[5] ),
    .A1(\cpu.intr.r_timer_count[21] ),
    .S(net923),
    .X(_05620_));
 sg13g2_mux2_1 _23327_ (.A0(\cpu.intr.r_timer_reload[5] ),
    .A1(\cpu.intr.r_timer_reload[21] ),
    .S(net923),
    .X(_05621_));
 sg13g2_a22oi_1 _23328_ (.Y(_05622_),
    .B1(_05621_),
    .B2(net494),
    .A2(_05620_),
    .A1(net485));
 sg13g2_buf_1 _23329_ (.A(\cpu.intr.r_clock_count[21] ),
    .X(_05623_));
 sg13g2_a22oi_1 _23330_ (.Y(_05624_),
    .B1(_04938_),
    .B2(_09323_),
    .A2(net443),
    .A1(_05623_));
 sg13g2_and2_1 _23331_ (.A(_05622_),
    .B(_05624_),
    .X(_05625_));
 sg13g2_o21ai_1 _23332_ (.B1(_05625_),
    .Y(_05626_),
    .A1(net662),
    .A2(_05619_));
 sg13g2_a221oi_1 _23333_ (.B2(_09322_),
    .C1(_05626_),
    .B1(_05618_),
    .A1(\cpu.intr.r_clock_cmp[21] ),
    .Y(_05627_),
    .A2(_05131_));
 sg13g2_nor2_1 _23334_ (.A(net683),
    .B(_05627_),
    .Y(_05628_));
 sg13g2_nand3_1 _23335_ (.B(_09310_),
    .C(_04979_),
    .A(_09309_),
    .Y(_05629_));
 sg13g2_a22oi_1 _23336_ (.Y(_05630_),
    .B1(net652),
    .B2(net8),
    .A2(_10255_),
    .A1(\cpu.gpio.genblk2[5].srcs_io[0] ));
 sg13g2_a22oi_1 _23337_ (.Y(_05631_),
    .B1(_05035_),
    .B2(\cpu.gpio.genblk1[5].srcs_o[0] ),
    .A2(_04932_),
    .A1(_09313_));
 sg13g2_a21oi_1 _23338_ (.A1(_05630_),
    .A2(_05631_),
    .Y(_05632_),
    .B1(net872));
 sg13g2_nor2b_1 _23339_ (.A(_00138_),
    .B_N(_04983_),
    .Y(_05633_));
 sg13g2_a22oi_1 _23340_ (.Y(_05634_),
    .B1(_04992_),
    .B2(_09310_),
    .A2(_04912_),
    .A1(_09312_));
 sg13g2_nand3_1 _23341_ (.B(_09313_),
    .C(net977),
    .A(_09312_),
    .Y(_05635_));
 sg13g2_o21ai_1 _23342_ (.B1(_05635_),
    .Y(_05636_),
    .A1(_11383_),
    .A2(_00137_));
 sg13g2_a22oi_1 _23343_ (.Y(_05637_),
    .B1(_05636_),
    .B2(_04952_),
    .A2(net380),
    .A1(_09309_));
 sg13g2_inv_1 _23344_ (.Y(_05638_),
    .A(_00136_));
 sg13g2_buf_2 _23345_ (.A(\cpu.gpio.r_src_io[5][1] ),
    .X(_05639_));
 sg13g2_nand2b_1 _23346_ (.Y(_05640_),
    .B(net427),
    .A_N(_00134_));
 sg13g2_o21ai_1 _23347_ (.B1(_05640_),
    .Y(_05641_),
    .A1(_00135_),
    .A2(net343));
 sg13g2_a221oi_1 _23348_ (.B2(_05639_),
    .C1(_05641_),
    .B1(net428),
    .A1(_05638_),
    .Y(_05642_),
    .A2(_04986_));
 sg13g2_nand3_1 _23349_ (.B(_05637_),
    .C(_05642_),
    .A(_05634_),
    .Y(_05643_));
 sg13g2_nor3_1 _23350_ (.A(_05632_),
    .B(_05633_),
    .C(_05643_),
    .Y(_05644_));
 sg13g2_a21oi_1 _23351_ (.A1(_05629_),
    .A2(_05644_),
    .Y(_05645_),
    .B1(_05011_));
 sg13g2_nor4_1 _23352_ (.A(_05615_),
    .B(_05617_),
    .C(_05628_),
    .D(_05645_),
    .Y(_05646_));
 sg13g2_nand2_1 _23353_ (.Y(_05647_),
    .A(_02925_),
    .B(_05646_));
 sg13g2_o21ai_1 _23354_ (.B1(_05647_),
    .Y(_05648_),
    .A1(net891),
    .A2(_05609_));
 sg13g2_nand2_1 _23355_ (.Y(_05649_),
    .A(net659),
    .B(net83));
 sg13g2_o21ai_1 _23356_ (.B1(_05649_),
    .Y(_05650_),
    .A1(net63),
    .A2(_05648_));
 sg13g2_nand2_1 _23357_ (.Y(_05651_),
    .A(net97),
    .B(_05650_));
 sg13g2_o21ai_1 _23358_ (.B1(_05651_),
    .Y(_01042_),
    .A1(_05584_),
    .A2(_05585_));
 sg13g2_nand2_1 _23359_ (.Y(_05652_),
    .A(net762),
    .B(_04606_));
 sg13g2_a21oi_1 _23360_ (.A1(_05434_),
    .A2(_04608_),
    .Y(_05653_),
    .B1(net398));
 sg13g2_a22oi_1 _23361_ (.Y(_05654_),
    .B1(_05652_),
    .B2(_05653_),
    .A2(_11540_),
    .A1(net980));
 sg13g2_buf_1 _23362_ (.A(\cpu.intr.r_clock_count[22] ),
    .X(_05655_));
 sg13g2_mux2_1 _23363_ (.A0(\cpu.intr.r_clock_cmp[6] ),
    .A1(\cpu.intr.r_timer_reload[6] ),
    .S(net496),
    .X(_05656_));
 sg13g2_a221oi_1 _23364_ (.B2(net531),
    .C1(net662),
    .B1(_05656_),
    .A1(\cpu.intr.r_timer_count[6] ),
    .Y(_05657_),
    .A2(net759));
 sg13g2_mux2_1 _23365_ (.A0(\cpu.intr.r_clock_cmp[22] ),
    .A1(\cpu.intr.r_timer_reload[22] ),
    .S(_09345_),
    .X(_05658_));
 sg13g2_a221oi_1 _23366_ (.B2(net531),
    .C1(net786),
    .B1(_05658_),
    .A1(\cpu.intr.r_timer_count[22] ),
    .Y(_05659_),
    .A2(_12447_));
 sg13g2_nor3_1 _23367_ (.A(net760),
    .B(_05657_),
    .C(_05659_),
    .Y(_05660_));
 sg13g2_a221oi_1 _23368_ (.B2(_10289_),
    .C1(_05660_),
    .B1(net467),
    .A1(_05655_),
    .Y(_05661_),
    .A2(_10256_));
 sg13g2_nor3_1 _23369_ (.A(net683),
    .B(net264),
    .C(_05661_),
    .Y(_05662_));
 sg13g2_nand3_1 _23370_ (.B(_09299_),
    .C(_04979_),
    .A(_09298_),
    .Y(_05663_));
 sg13g2_nand2_1 _23371_ (.Y(_05664_),
    .A(\cpu.gpio.genblk1[6].srcs_o[0] ),
    .B(_05132_));
 sg13g2_a22oi_1 _23372_ (.Y(_05665_),
    .B1(_05162_),
    .B2(net9),
    .A2(_10255_),
    .A1(\cpu.gpio.genblk2[6].srcs_io[0] ));
 sg13g2_a21oi_1 _23373_ (.A1(_09314_),
    .A2(_04952_),
    .Y(_05666_),
    .B1(_04932_));
 sg13g2_nand2b_1 _23374_ (.Y(_05667_),
    .B(_09315_),
    .A_N(_05666_));
 sg13g2_nand3_1 _23375_ (.B(_05665_),
    .C(_05667_),
    .A(_05664_),
    .Y(_05668_));
 sg13g2_nand2b_1 _23376_ (.Y(_05669_),
    .B(_04983_),
    .A_N(_00150_));
 sg13g2_a22oi_1 _23377_ (.Y(_05670_),
    .B1(_04992_),
    .B2(_09299_),
    .A2(_04912_),
    .A1(_09314_));
 sg13g2_buf_1 _23378_ (.A(\cpu.gpio.r_src_io[5][2] ),
    .X(_05671_));
 sg13g2_inv_1 _23379_ (.Y(_05672_),
    .A(_00146_));
 sg13g2_a22oi_1 _23380_ (.Y(_05673_),
    .B1(net427),
    .B2(_05672_),
    .A2(net428),
    .A1(_05671_));
 sg13g2_nand2b_1 _23381_ (.Y(_05674_),
    .B(_04932_),
    .A_N(_00147_));
 sg13g2_o21ai_1 _23382_ (.B1(_05674_),
    .Y(_05675_),
    .A1(_00149_),
    .A2(_05564_));
 sg13g2_nor2_1 _23383_ (.A(_00148_),
    .B(_05054_),
    .Y(_05676_));
 sg13g2_a221oi_1 _23384_ (.B2(_12057_),
    .C1(_05676_),
    .B1(_05675_),
    .A1(_09298_),
    .Y(_05677_),
    .A2(net380));
 sg13g2_nand4_1 _23385_ (.B(_05670_),
    .C(_05673_),
    .A(_05669_),
    .Y(_05678_),
    .D(_05677_));
 sg13g2_a21oi_1 _23386_ (.A1(net977),
    .A2(_05668_),
    .Y(_05679_),
    .B1(_05678_));
 sg13g2_a21oi_1 _23387_ (.A1(_05663_),
    .A2(_05679_),
    .Y(_05680_),
    .B1(_05011_));
 sg13g2_a22oi_1 _23388_ (.Y(_05681_),
    .B1(_04928_),
    .B2(\cpu.uart.r_in[6] ),
    .A2(net429),
    .A1(\cpu.uart.r_div_value[6] ));
 sg13g2_o21ai_1 _23389_ (.B1(net1011),
    .Y(_05682_),
    .A1(_04926_),
    .A2(_05681_));
 sg13g2_buf_1 _23390_ (.A(\cpu.spi.r_clk_count[2][6] ),
    .X(_05683_));
 sg13g2_nand2b_1 _23391_ (.Y(_05684_),
    .B(net383),
    .A_N(_00145_));
 sg13g2_o21ai_1 _23392_ (.B1(_05684_),
    .Y(_05685_),
    .A1(_00144_),
    .A2(_04919_));
 sg13g2_a221oi_1 _23393_ (.B2(\cpu.spi.r_timeout[6] ),
    .C1(_05685_),
    .B1(net430),
    .A1(_05683_),
    .Y(_05686_),
    .A2(_04915_));
 sg13g2_nand2_1 _23394_ (.Y(_05687_),
    .A(_09415_),
    .B(_04897_));
 sg13g2_a21oi_1 _23395_ (.A1(_05686_),
    .A2(_05687_),
    .Y(_05688_),
    .B1(net709));
 sg13g2_nor4_1 _23396_ (.A(_05662_),
    .B(_05680_),
    .C(_05682_),
    .D(_05688_),
    .Y(_05689_));
 sg13g2_a22oi_1 _23397_ (.Y(_05690_),
    .B1(_10235_),
    .B2(\cpu.dcache.r_data[4][22] ),
    .A2(_04837_),
    .A1(\cpu.dcache.r_data[3][22] ));
 sg13g2_nand2_1 _23398_ (.Y(_05691_),
    .A(\cpu.dcache.r_data[7][22] ),
    .B(_10119_));
 sg13g2_a22oi_1 _23399_ (.Y(_05692_),
    .B1(net528),
    .B2(\cpu.dcache.r_data[6][22] ),
    .A2(net432),
    .A1(\cpu.dcache.r_data[2][22] ));
 sg13g2_nor2_1 _23400_ (.A(_00141_),
    .B(_04830_),
    .Y(_05693_));
 sg13g2_a221oi_1 _23401_ (.B2(\cpu.dcache.r_data[5][22] ),
    .C1(_05693_),
    .B1(net529),
    .A1(\cpu.dcache.r_data[1][22] ),
    .Y(_05694_),
    .A2(_12331_));
 sg13g2_nand4_1 _23402_ (.B(_05691_),
    .C(_05692_),
    .A(_05690_),
    .Y(_05695_),
    .D(_05694_));
 sg13g2_nand2_1 _23403_ (.Y(_05696_),
    .A(_10117_),
    .B(_05695_));
 sg13g2_mux2_1 _23404_ (.A0(_05253_),
    .A1(_05696_),
    .S(_04849_),
    .X(_05697_));
 sg13g2_nand2b_1 _23405_ (.Y(_05698_),
    .B(_05260_),
    .A_N(_08502_));
 sg13g2_a22oi_1 _23406_ (.Y(_05699_),
    .B1(net494),
    .B2(\cpu.dcache.r_data[7][6] ),
    .A2(net487),
    .A1(\cpu.dcache.r_data[3][6] ));
 sg13g2_a22oi_1 _23407_ (.Y(_05700_),
    .B1(net432),
    .B2(\cpu.dcache.r_data[2][6] ),
    .A2(net493),
    .A1(\cpu.dcache.r_data[4][6] ));
 sg13g2_a22oi_1 _23408_ (.Y(_05701_),
    .B1(_02733_),
    .B2(\cpu.dcache.r_data[6][6] ),
    .A2(_12781_),
    .A1(\cpu.dcache.r_data[5][6] ));
 sg13g2_nand3_1 _23409_ (.B(_05700_),
    .C(_05701_),
    .A(_05699_),
    .Y(_05702_));
 sg13g2_nand2_1 _23410_ (.Y(_05703_),
    .A(_00140_),
    .B(_04868_));
 sg13g2_o21ai_1 _23411_ (.B1(_05703_),
    .Y(_05704_),
    .A1(_04868_),
    .A2(_05702_));
 sg13g2_o21ai_1 _23412_ (.B1(_12332_),
    .Y(_05705_),
    .A1(\cpu.dcache.r_data[1][6] ),
    .A2(_05702_));
 sg13g2_o21ai_1 _23413_ (.B1(_05705_),
    .Y(_05706_),
    .A1(_12332_),
    .A2(_05704_));
 sg13g2_a22oi_1 _23414_ (.Y(_05707_),
    .B1(_05706_),
    .B2(_05067_),
    .A2(_05698_),
    .A1(_04852_));
 sg13g2_o21ai_1 _23415_ (.B1(_05707_),
    .Y(_05708_),
    .A1(net975),
    .A2(_05697_));
 sg13g2_nand2_1 _23416_ (.Y(_05709_),
    .A(net620),
    .B(_05706_));
 sg13g2_nand3_1 _23417_ (.B(_05696_),
    .C(_05709_),
    .A(net514),
    .Y(_05710_));
 sg13g2_a21oi_1 _23418_ (.A1(_05708_),
    .A2(_05710_),
    .Y(_05711_),
    .B1(net891));
 sg13g2_nor3_1 _23419_ (.A(net83),
    .B(_05689_),
    .C(_05711_),
    .Y(_05712_));
 sg13g2_a21o_1 _23420_ (.A2(net63),
    .A1(net984),
    .B1(_05712_),
    .X(_05713_));
 sg13g2_mux2_1 _23421_ (.A0(_05654_),
    .A1(_05713_),
    .S(net97),
    .X(_01043_));
 sg13g2_o21ai_1 _23422_ (.B1(net82),
    .Y(_05714_),
    .A1(_08777_),
    .A2(net189));
 sg13g2_nand2_1 _23423_ (.Y(_05715_),
    .A(_02953_),
    .B(net84));
 sg13g2_o21ai_1 _23424_ (.B1(_05715_),
    .Y(_05716_),
    .A1(net83),
    .A2(_05108_));
 sg13g2_nand2_1 _23425_ (.Y(_05717_),
    .A(net98),
    .B(_05716_));
 sg13g2_nand2_1 _23426_ (.Y(_05718_),
    .A(_11682_),
    .B(_04633_));
 sg13g2_a21oi_1 _23427_ (.A1(net655),
    .A2(_04635_),
    .Y(_05719_),
    .B1(_04820_));
 sg13g2_a22oi_1 _23428_ (.Y(_01044_),
    .B1(_05718_),
    .B2(_05719_),
    .A2(_05717_),
    .A1(_05714_));
 sg13g2_a21o_1 _23429_ (.A2(_04670_),
    .A1(net651),
    .B1(_11540_),
    .X(_05720_));
 sg13g2_a21oi_1 _23430_ (.A1(net762),
    .A2(_04668_),
    .Y(_05721_),
    .B1(_05720_));
 sg13g2_o21ai_1 _23431_ (.B1(net82),
    .Y(_05722_),
    .A1(_08757_),
    .A2(net189));
 sg13g2_nand2b_1 _23432_ (.Y(_05723_),
    .B(_04828_),
    .A_N(_09279_));
 sg13g2_a22oi_1 _23433_ (.Y(_05724_),
    .B1(net652),
    .B2(\cpu.intr.r_clock_cmp[8] ),
    .A2(net467),
    .A1(_10297_));
 sg13g2_buf_1 _23434_ (.A(\cpu.intr.r_clock_count[24] ),
    .X(_05725_));
 sg13g2_a22oi_1 _23435_ (.Y(_05726_),
    .B1(net653),
    .B2(\cpu.intr.r_clock_cmp[24] ),
    .A2(net399),
    .A1(_05725_));
 sg13g2_a22oi_1 _23436_ (.Y(_05727_),
    .B1(net435),
    .B2(_10091_),
    .A2(net445),
    .A1(\cpu.intr.r_timer_reload[8] ));
 sg13g2_or2_1 _23437_ (.X(_05728_),
    .B(_05727_),
    .A(net618));
 sg13g2_nand3_1 _23438_ (.B(_05726_),
    .C(_05728_),
    .A(_05724_),
    .Y(_05729_));
 sg13g2_mux2_1 _23439_ (.A0(_04840_),
    .A1(_04847_),
    .S(_10245_),
    .X(_05730_));
 sg13g2_a22oi_1 _23440_ (.Y(_05731_),
    .B1(_05730_),
    .B2(net514),
    .A2(_05729_),
    .A1(_05127_));
 sg13g2_nor2_1 _23441_ (.A(net976),
    .B(_05731_),
    .Y(_05732_));
 sg13g2_or3_1 _23442_ (.A(_04829_),
    .B(_05207_),
    .C(_05732_),
    .X(_05733_));
 sg13g2_nand3_1 _23443_ (.B(_05723_),
    .C(_05733_),
    .A(net98),
    .Y(_05734_));
 sg13g2_o21ai_1 _23444_ (.B1(_05734_),
    .Y(_01045_),
    .A1(_05721_),
    .A2(_05722_));
 sg13g2_nand2b_1 _23445_ (.Y(_05735_),
    .B(_04818_),
    .A_N(_04701_));
 sg13g2_o21ai_1 _23446_ (.B1(_05735_),
    .Y(_05736_),
    .A1(net655),
    .A2(_04699_));
 sg13g2_mux2_1 _23447_ (.A0(\cpu.intr.r_clock_cmp[9] ),
    .A1(\cpu.intr.r_timer_reload[9] ),
    .S(net437),
    .X(_05737_));
 sg13g2_a22oi_1 _23448_ (.Y(_05738_),
    .B1(_05737_),
    .B2(net475),
    .A2(net689),
    .A1(_10304_));
 sg13g2_buf_2 _23449_ (.A(\cpu.intr.r_clock_count[25] ),
    .X(_05739_));
 sg13g2_and2_1 _23450_ (.A(_05739_),
    .B(net399),
    .X(_05740_));
 sg13g2_a221oi_1 _23451_ (.B2(\cpu.intr.r_clock_cmp[25] ),
    .C1(_05740_),
    .B1(net653),
    .A1(\cpu.intr.r_timer_count[9] ),
    .Y(_05741_),
    .A2(_05033_));
 sg13g2_o21ai_1 _23452_ (.B1(_05741_),
    .Y(_05742_),
    .A1(_05128_),
    .A2(_05738_));
 sg13g2_mux2_1 _23453_ (.A0(_05307_),
    .A1(_05318_),
    .S(_10245_),
    .X(_05743_));
 sg13g2_a22oi_1 _23454_ (.Y(_05744_),
    .B1(_05743_),
    .B2(net514),
    .A2(_05742_),
    .A1(_05127_));
 sg13g2_nor2_1 _23455_ (.A(net976),
    .B(_05744_),
    .Y(_05745_));
 sg13g2_nor3_1 _23456_ (.A(_04827_),
    .B(_05207_),
    .C(_05745_),
    .Y(_05746_));
 sg13g2_a21oi_1 _23457_ (.A1(_02958_),
    .A2(_04829_),
    .Y(_05747_),
    .B1(_05746_));
 sg13g2_inv_1 _23458_ (.Y(_05748_),
    .A(_08738_));
 sg13g2_nor3_1 _23459_ (.A(net974),
    .B(net215),
    .C(_05021_),
    .Y(_05749_));
 sg13g2_a21oi_1 _23460_ (.A1(_05021_),
    .A2(_05747_),
    .Y(_05750_),
    .B1(_05749_));
 sg13g2_o21ai_1 _23461_ (.B1(_05750_),
    .Y(_01046_),
    .A1(_04820_),
    .A2(_05736_));
 sg13g2_nand2b_1 _23462_ (.Y(_05751_),
    .B(\cpu.dec.r_rd[0] ),
    .A_N(_03373_));
 sg13g2_a21oi_1 _23463_ (.A1(net189),
    .A2(_05751_),
    .Y(_05752_),
    .B1(net98));
 sg13g2_a21o_1 _23464_ (.A2(net97),
    .A1(_10350_),
    .B1(_05752_),
    .X(_01047_));
 sg13g2_nand2b_1 _23465_ (.Y(_05753_),
    .B(\cpu.dec.r_rd[1] ),
    .A_N(_03373_));
 sg13g2_a21oi_1 _23466_ (.A1(net189),
    .A2(_05753_),
    .Y(_05754_),
    .B1(net98));
 sg13g2_a21o_1 _23467_ (.A2(net97),
    .A1(_10349_),
    .B1(_05754_),
    .X(_01048_));
 sg13g2_nor3_1 _23468_ (.A(_03373_),
    .B(_09388_),
    .C(net398),
    .Y(_05755_));
 sg13g2_nand3_1 _23469_ (.B(_05239_),
    .C(_05755_),
    .A(\cpu.dec.r_rd[2] ),
    .Y(_05756_));
 sg13g2_o21ai_1 _23470_ (.B1(_05756_),
    .Y(_01049_),
    .A1(_10354_),
    .A2(net85));
 sg13g2_inv_1 _23471_ (.Y(_05757_),
    .A(net1112));
 sg13g2_nand3_1 _23472_ (.B(_05239_),
    .C(_05755_),
    .A(\cpu.dec.r_rd[3] ),
    .Y(_05758_));
 sg13g2_o21ai_1 _23473_ (.B1(_05758_),
    .Y(_01050_),
    .A1(_05757_),
    .A2(_04824_));
 sg13g2_mux2_1 _23474_ (.A0(\cpu.dec.r_swapsp ),
    .A1(\cpu.ex.r_wb_swapsp ),
    .S(_05143_),
    .X(_01051_));
 sg13g2_and2_1 _23475_ (.A(_10399_),
    .B(_10979_),
    .X(_05759_));
 sg13g2_a21o_1 _23476_ (.A2(_10389_),
    .A1(net880),
    .B1(_05759_),
    .X(_05760_));
 sg13g2_mux2_1 _23477_ (.A0(_12141_),
    .A1(_05760_),
    .S(net85),
    .X(_01052_));
 sg13g2_buf_1 _23478_ (.A(net976),
    .X(_05761_));
 sg13g2_nor2b_1 _23479_ (.A(_10644_),
    .B_N(_10646_),
    .Y(_05762_));
 sg13g2_nor2_2 _23480_ (.A(_10833_),
    .B(_10834_),
    .Y(_05763_));
 sg13g2_nand2_1 _23481_ (.Y(_05764_),
    .A(net871),
    .B(_05763_));
 sg13g2_o21ai_1 _23482_ (.B1(_05764_),
    .Y(_05765_),
    .A1(net871),
    .A2(_05762_));
 sg13g2_mux2_1 _23483_ (.A0(_10312_),
    .A1(_05765_),
    .S(net85),
    .X(_01053_));
 sg13g2_nand2_2 _23484_ (.Y(_05766_),
    .A(_10914_),
    .B(_10934_));
 sg13g2_a21oi_1 _23485_ (.A1(_10679_),
    .A2(_10681_),
    .Y(_05767_),
    .B1(net976));
 sg13g2_a21oi_1 _23486_ (.A1(net871),
    .A2(_05766_),
    .Y(_05768_),
    .B1(_05767_));
 sg13g2_nand2_1 _23487_ (.Y(_05769_),
    .A(_10319_),
    .B(net97));
 sg13g2_o21ai_1 _23488_ (.B1(_05769_),
    .Y(_01054_),
    .A1(net97),
    .A2(_05768_));
 sg13g2_nor2_2 _23489_ (.A(_10901_),
    .B(_10902_),
    .Y(_05770_));
 sg13g2_a21oi_1 _23490_ (.A1(_10523_),
    .A2(_10524_),
    .Y(_05771_),
    .B1(_05137_));
 sg13g2_a21o_1 _23491_ (.A2(_05770_),
    .A1(_05761_),
    .B1(_05771_),
    .X(_05772_));
 sg13g2_mux2_1 _23492_ (.A0(_10324_),
    .A1(_05772_),
    .S(net85),
    .X(_01055_));
 sg13g2_nand2_1 _23493_ (.Y(_05773_),
    .A(net871),
    .B(_10872_));
 sg13g2_o21ai_1 _23494_ (.B1(_05773_),
    .Y(_05774_),
    .A1(_05761_),
    .A2(_10562_));
 sg13g2_mux2_1 _23495_ (.A0(_10326_),
    .A1(_05774_),
    .S(_04824_),
    .X(_01056_));
 sg13g2_a21o_1 _23496_ (.A2(net541),
    .A1(_02950_),
    .B1(_11005_),
    .X(_05775_));
 sg13g2_mux2_1 _23497_ (.A0(_05775_),
    .A1(_10612_),
    .S(_11680_),
    .X(_05776_));
 sg13g2_buf_2 _23498_ (.A(net101),
    .X(_05777_));
 sg13g2_mux2_1 _23499_ (.A0(_10339_),
    .A1(_05776_),
    .S(net81),
    .X(_01057_));
 sg13g2_and2_1 _23500_ (.A(net540),
    .B(_11033_),
    .X(_05778_));
 sg13g2_a21o_1 _23501_ (.A2(net541),
    .A1(_02953_),
    .B1(_05778_),
    .X(_05779_));
 sg13g2_nand2_1 _23502_ (.Y(_05780_),
    .A(net871),
    .B(_05779_));
 sg13g2_o21ai_1 _23503_ (.B1(_05780_),
    .Y(_05781_),
    .A1(net871),
    .A2(_10455_));
 sg13g2_mux2_1 _23504_ (.A0(_10344_),
    .A1(_05781_),
    .S(_05777_),
    .X(_01058_));
 sg13g2_nand2_1 _23505_ (.Y(_05782_),
    .A(_10391_),
    .B(_10793_));
 sg13g2_nor2_1 _23506_ (.A(_10788_),
    .B(_10792_),
    .Y(_05783_));
 sg13g2_o21ai_1 _23507_ (.B1(net540),
    .Y(_05784_),
    .A1(_05783_),
    .A2(_10786_));
 sg13g2_nand2_2 _23508_ (.Y(_05785_),
    .A(_05782_),
    .B(_05784_));
 sg13g2_mux2_1 _23509_ (.A0(net918),
    .A1(_05785_),
    .S(net81),
    .X(_01059_));
 sg13g2_mux2_1 _23510_ (.A0(net917),
    .A1(_05763_),
    .S(net81),
    .X(_01060_));
 sg13g2_mux2_1 _23511_ (.A0(net1033),
    .A1(_05766_),
    .S(net81),
    .X(_01061_));
 sg13g2_mux2_1 _23512_ (.A0(net1032),
    .A1(_05770_),
    .S(net81),
    .X(_01062_));
 sg13g2_mux2_1 _23513_ (.A0(net916),
    .A1(_10872_),
    .S(net81),
    .X(_01063_));
 sg13g2_mux2_1 _23514_ (.A0(net1031),
    .A1(_05775_),
    .S(net81),
    .X(_01064_));
 sg13g2_mux2_1 _23515_ (.A0(net1034),
    .A1(_05779_),
    .S(net81),
    .X(_01065_));
 sg13g2_nor2b_1 _23516_ (.A(_10745_),
    .B_N(_10746_),
    .Y(_05786_));
 sg13g2_nand2_1 _23517_ (.Y(_05787_),
    .A(_05137_),
    .B(_05760_));
 sg13g2_o21ai_1 _23518_ (.B1(_05787_),
    .Y(_05788_),
    .A1(net871),
    .A2(_05786_));
 sg13g2_mux2_1 _23519_ (.A0(_10302_),
    .A1(_05788_),
    .S(_05777_),
    .X(_01066_));
 sg13g2_mux2_1 _23520_ (.A0(_10718_),
    .A1(_05785_),
    .S(net871),
    .X(_05789_));
 sg13g2_mux2_1 _23521_ (.A0(_10307_),
    .A1(_05789_),
    .S(net82),
    .X(_01067_));
 sg13g2_buf_1 _23522_ (.A(net282),
    .X(_05790_));
 sg13g2_nand2_1 _23523_ (.Y(_05791_),
    .A(_08456_),
    .B(_08489_));
 sg13g2_buf_2 _23524_ (.A(_05791_),
    .X(_05792_));
 sg13g2_nor2_1 _23525_ (.A(_08530_),
    .B(_05792_),
    .Y(_05793_));
 sg13g2_a21oi_1 _23526_ (.A1(_03694_),
    .A2(_05792_),
    .Y(_05794_),
    .B1(_05793_));
 sg13g2_nor3_1 _23527_ (.A(_10962_),
    .B(_10805_),
    .C(_10937_),
    .Y(_05795_));
 sg13g2_and2_1 _23528_ (.A(_10797_),
    .B(_05795_),
    .X(_05796_));
 sg13g2_buf_1 _23529_ (.A(_05796_),
    .X(_05797_));
 sg13g2_nand2b_1 _23530_ (.Y(_05798_),
    .B(\cpu.dec.do_inv_mmu ),
    .A_N(_05797_));
 sg13g2_buf_2 _23531_ (.A(_05798_),
    .X(_05799_));
 sg13g2_nor4_2 _23532_ (.A(_08388_),
    .B(_04736_),
    .C(_10356_),
    .Y(_05800_),
    .D(_03448_));
 sg13g2_and2_1 _23533_ (.A(_05799_),
    .B(_05800_),
    .X(_05801_));
 sg13g2_buf_1 _23534_ (.A(_05801_),
    .X(_05802_));
 sg13g2_buf_1 _23535_ (.A(_00288_),
    .X(_05803_));
 sg13g2_nand2b_1 _23536_ (.Y(_05804_),
    .B(net1052),
    .A_N(net1083));
 sg13g2_o21ai_1 _23537_ (.B1(_05804_),
    .Y(_05805_),
    .A1(net880),
    .A2(net687));
 sg13g2_nand3_1 _23538_ (.B(_05802_),
    .C(_05805_),
    .A(net282),
    .Y(_05806_));
 sg13g2_o21ai_1 _23539_ (.B1(_05806_),
    .Y(_05807_),
    .A1(net214),
    .A2(_05794_));
 sg13g2_nand2b_1 _23540_ (.Y(_05808_),
    .B(net282),
    .A_N(_05802_));
 sg13g2_nand2_1 _23541_ (.Y(_05809_),
    .A(_09444_),
    .B(_05808_));
 sg13g2_inv_2 _23542_ (.Y(_05810_),
    .A(_10483_));
 sg13g2_a22oi_1 _23543_ (.Y(_01070_),
    .B1(_05809_),
    .B2(_05810_),
    .A2(_05807_),
    .A1(_12004_));
 sg13g2_nor2_1 _23544_ (.A(_08689_),
    .B(_05792_),
    .Y(_05811_));
 sg13g2_a21oi_1 _23545_ (.A1(net875),
    .A2(_05792_),
    .Y(_05812_),
    .B1(_05811_));
 sg13g2_nor2_1 _23546_ (.A(_05810_),
    .B(_11224_),
    .Y(_05813_));
 sg13g2_buf_1 _23547_ (.A(_05813_),
    .X(_05814_));
 sg13g2_buf_1 _23548_ (.A(_10483_),
    .X(_05815_));
 sg13g2_nor2_1 _23549_ (.A(net973),
    .B(net1024),
    .Y(_05816_));
 sg13g2_buf_2 _23550_ (.A(_05816_),
    .X(_05817_));
 sg13g2_o21ai_1 _23551_ (.B1(net880),
    .Y(_05818_),
    .A1(_05814_),
    .A2(_05817_));
 sg13g2_o21ai_1 _23552_ (.B1(_05818_),
    .Y(_05819_),
    .A1(net880),
    .A2(net791));
 sg13g2_nand3_1 _23553_ (.B(_05802_),
    .C(_05819_),
    .A(net214),
    .Y(_05820_));
 sg13g2_o21ai_1 _23554_ (.B1(_05820_),
    .Y(_05821_),
    .A1(net214),
    .A2(_05812_));
 sg13g2_a22oi_1 _23555_ (.Y(_01071_),
    .B1(_05821_),
    .B2(net685),
    .A2(_05809_),
    .A1(_11224_));
 sg13g2_inv_1 _23556_ (.Y(_05822_),
    .A(net1109));
 sg13g2_buf_1 _23557_ (.A(_05822_),
    .X(_05823_));
 sg13g2_nor2_1 _23558_ (.A(net815),
    .B(_05792_),
    .Y(_05824_));
 sg13g2_a21oi_1 _23559_ (.A1(net740),
    .A2(_05792_),
    .Y(_05825_),
    .B1(_05824_));
 sg13g2_nand2_1 _23560_ (.Y(_05826_),
    .A(net973),
    .B(net1024));
 sg13g2_buf_2 _23561_ (.A(_05826_),
    .X(_05827_));
 sg13g2_nor2_2 _23562_ (.A(net870),
    .B(_05827_),
    .Y(_05828_));
 sg13g2_buf_1 _23563_ (.A(net1109),
    .X(_05829_));
 sg13g2_nor2_1 _23564_ (.A(net972),
    .B(_05814_),
    .Y(_05830_));
 sg13g2_o21ai_1 _23565_ (.B1(net880),
    .Y(_05831_),
    .A1(_05828_),
    .A2(_05830_));
 sg13g2_o21ai_1 _23566_ (.B1(_05831_),
    .Y(_05832_),
    .A1(net880),
    .A2(net622));
 sg13g2_nand3_1 _23567_ (.B(_05802_),
    .C(_05832_),
    .A(net282),
    .Y(_05833_));
 sg13g2_o21ai_1 _23568_ (.B1(_05833_),
    .Y(_05834_),
    .A1(net214),
    .A2(_05825_));
 sg13g2_buf_2 _23569_ (.A(net803),
    .X(_05835_));
 sg13g2_a22oi_1 _23570_ (.Y(_01072_),
    .B1(_05834_),
    .B2(_05835_),
    .A2(_05809_),
    .A1(_05823_));
 sg13g2_buf_1 _23571_ (.A(_10415_),
    .X(_05836_));
 sg13g2_inv_2 _23572_ (.Y(_05837_),
    .A(net971));
 sg13g2_nor2_1 _23573_ (.A(net941),
    .B(_05792_),
    .Y(_05838_));
 sg13g2_a21oi_1 _23574_ (.A1(_11147_),
    .A2(_05792_),
    .Y(_05839_),
    .B1(_05838_));
 sg13g2_xnor2_1 _23575_ (.Y(_05840_),
    .A(net971),
    .B(_05828_));
 sg13g2_nand2_1 _23576_ (.Y(_05841_),
    .A(net880),
    .B(_05840_));
 sg13g2_o21ai_1 _23577_ (.B1(_05841_),
    .Y(_05842_),
    .A1(net880),
    .A2(net926));
 sg13g2_nand3_1 _23578_ (.B(_05802_),
    .C(_05842_),
    .A(net282),
    .Y(_05843_));
 sg13g2_o21ai_1 _23579_ (.B1(_05843_),
    .Y(_05844_),
    .A1(net214),
    .A2(_05839_));
 sg13g2_a22oi_1 _23580_ (.Y(_01073_),
    .B1(_05844_),
    .B2(_05835_),
    .A2(_05809_),
    .A1(_05837_));
 sg13g2_buf_2 _23581_ (.A(_00188_),
    .X(_05845_));
 sg13g2_buf_1 _23582_ (.A(_10819_),
    .X(_05846_));
 sg13g2_nor2_1 _23583_ (.A(_05846_),
    .B(net971),
    .Y(_05847_));
 sg13g2_nand2_1 _23584_ (.Y(_05848_),
    .A(_05845_),
    .B(_05847_));
 sg13g2_nand2_1 _23585_ (.Y(_05849_),
    .A(net1052),
    .B(_05800_));
 sg13g2_nor2_1 _23586_ (.A(_10930_),
    .B(_05849_),
    .Y(_05850_));
 sg13g2_nand2_2 _23587_ (.Y(_05851_),
    .A(_05817_),
    .B(_05850_));
 sg13g2_nor2_1 _23588_ (.A(_05848_),
    .B(_05851_),
    .Y(_05852_));
 sg13g2_buf_1 _23589_ (.A(_05852_),
    .X(_05853_));
 sg13g2_buf_1 _23590_ (.A(_05853_),
    .X(_05854_));
 sg13g2_mux2_1 _23591_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][0] ),
    .A1(net474),
    .S(net342),
    .X(_01141_));
 sg13g2_mux2_1 _23592_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][10] ),
    .A1(_03429_),
    .S(net342),
    .X(_01142_));
 sg13g2_mux2_1 _23593_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][11] ),
    .A1(_03430_),
    .S(net342),
    .X(_01143_));
 sg13g2_mux2_1 _23594_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][1] ),
    .A1(net521),
    .S(_05854_),
    .X(_01144_));
 sg13g2_buf_1 _23595_ (.A(net889),
    .X(_05855_));
 sg13g2_mux2_1 _23596_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][2] ),
    .A1(net738),
    .S(net342),
    .X(_01145_));
 sg13g2_mux2_1 _23597_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][3] ),
    .A1(_04740_),
    .S(net342),
    .X(_01146_));
 sg13g2_mux2_1 _23598_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][4] ),
    .A1(net739),
    .S(net342),
    .X(_01147_));
 sg13g2_mux2_1 _23599_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][5] ),
    .A1(net879),
    .S(net342),
    .X(_01148_));
 sg13g2_mux2_1 _23600_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][6] ),
    .A1(_04742_),
    .S(net342),
    .X(_01149_));
 sg13g2_mux2_1 _23601_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][7] ),
    .A1(net878),
    .S(_05854_),
    .X(_01150_));
 sg13g2_mux2_1 _23602_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][8] ),
    .A1(_03427_),
    .S(_05853_),
    .X(_01151_));
 sg13g2_mux2_1 _23603_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][9] ),
    .A1(_03428_),
    .S(_05853_),
    .X(_01152_));
 sg13g2_buf_1 _23604_ (.A(_05850_),
    .X(_05856_));
 sg13g2_nor2_1 _23605_ (.A(_10483_),
    .B(_11224_),
    .Y(_05857_));
 sg13g2_buf_2 _23606_ (.A(_05857_),
    .X(_05858_));
 sg13g2_nand2_1 _23607_ (.Y(_05859_),
    .A(net870),
    .B(_05858_));
 sg13g2_buf_2 _23608_ (.A(_05859_),
    .X(_05860_));
 sg13g2_nand2_2 _23609_ (.Y(_05861_),
    .A(net1016),
    .B(net971));
 sg13g2_nor2_2 _23610_ (.A(_05860_),
    .B(_05861_),
    .Y(_05862_));
 sg13g2_and2_1 _23611_ (.A(net466),
    .B(_05862_),
    .X(_05863_));
 sg13g2_buf_1 _23612_ (.A(_05863_),
    .X(_05864_));
 sg13g2_buf_1 _23613_ (.A(_05864_),
    .X(_05865_));
 sg13g2_mux2_1 _23614_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][0] ),
    .A1(_03436_),
    .S(_05865_),
    .X(_01153_));
 sg13g2_buf_1 _23615_ (.A(net622),
    .X(_05866_));
 sg13g2_mux2_1 _23616_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][10] ),
    .A1(_05866_),
    .S(net341),
    .X(_01154_));
 sg13g2_mux2_1 _23617_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][11] ),
    .A1(_03430_),
    .S(net341),
    .X(_01155_));
 sg13g2_mux2_1 _23618_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][1] ),
    .A1(net521),
    .S(_05865_),
    .X(_01156_));
 sg13g2_mux2_1 _23619_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][2] ),
    .A1(net738),
    .S(net341),
    .X(_01157_));
 sg13g2_mux2_1 _23620_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][3] ),
    .A1(net874),
    .S(net341),
    .X(_01158_));
 sg13g2_mux2_1 _23621_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][4] ),
    .A1(net739),
    .S(net341),
    .X(_01159_));
 sg13g2_mux2_1 _23622_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][5] ),
    .A1(_03446_),
    .S(net341),
    .X(_01160_));
 sg13g2_mux2_1 _23623_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][6] ),
    .A1(net873),
    .S(net341),
    .X(_01161_));
 sg13g2_mux2_1 _23624_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][7] ),
    .A1(net878),
    .S(net341),
    .X(_01162_));
 sg13g2_buf_1 _23625_ (.A(net687),
    .X(_05867_));
 sg13g2_mux2_1 _23626_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][8] ),
    .A1(net585),
    .S(_05864_),
    .X(_01163_));
 sg13g2_buf_1 _23627_ (.A(net791),
    .X(_05868_));
 sg13g2_mux2_1 _23628_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][9] ),
    .A1(net649),
    .S(_05864_),
    .X(_01164_));
 sg13g2_nand2_1 _23629_ (.Y(_05869_),
    .A(net1016),
    .B(net973));
 sg13g2_nor4_1 _23630_ (.A(_11224_),
    .B(net1109),
    .C(_05837_),
    .D(_05869_),
    .Y(_05870_));
 sg13g2_buf_2 _23631_ (.A(_05870_),
    .X(_05871_));
 sg13g2_and2_1 _23632_ (.A(net466),
    .B(_05871_),
    .X(_05872_));
 sg13g2_buf_1 _23633_ (.A(_05872_),
    .X(_05873_));
 sg13g2_buf_1 _23634_ (.A(_05873_),
    .X(_05874_));
 sg13g2_mux2_1 _23635_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][0] ),
    .A1(_03436_),
    .S(_05874_),
    .X(_01165_));
 sg13g2_mux2_1 _23636_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][10] ),
    .A1(_05866_),
    .S(net340),
    .X(_01166_));
 sg13g2_buf_1 _23637_ (.A(net926),
    .X(_05875_));
 sg13g2_mux2_1 _23638_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][11] ),
    .A1(net737),
    .S(net340),
    .X(_01167_));
 sg13g2_mux2_1 _23639_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][1] ),
    .A1(net521),
    .S(_05874_),
    .X(_01168_));
 sg13g2_mux2_1 _23640_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][2] ),
    .A1(net738),
    .S(net340),
    .X(_01169_));
 sg13g2_mux2_1 _23641_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][3] ),
    .A1(net874),
    .S(net340),
    .X(_01170_));
 sg13g2_mux2_1 _23642_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][4] ),
    .A1(net739),
    .S(net340),
    .X(_01171_));
 sg13g2_mux2_1 _23643_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][5] ),
    .A1(_03446_),
    .S(net340),
    .X(_01172_));
 sg13g2_mux2_1 _23644_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][6] ),
    .A1(net873),
    .S(net340),
    .X(_01173_));
 sg13g2_mux2_1 _23645_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][7] ),
    .A1(net878),
    .S(net340),
    .X(_01174_));
 sg13g2_mux2_1 _23646_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][8] ),
    .A1(net585),
    .S(_05873_),
    .X(_01175_));
 sg13g2_mux2_1 _23647_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][9] ),
    .A1(net649),
    .S(_05873_),
    .X(_01176_));
 sg13g2_buf_1 _23648_ (.A(_03435_),
    .X(_05876_));
 sg13g2_nor2_1 _23649_ (.A(net970),
    .B(_05837_),
    .Y(_05877_));
 sg13g2_nand2b_1 _23650_ (.Y(_05878_),
    .B(_05877_),
    .A_N(_05845_));
 sg13g2_buf_1 _23651_ (.A(_05878_),
    .X(_05879_));
 sg13g2_nor2_1 _23652_ (.A(_05851_),
    .B(_05879_),
    .Y(_05880_));
 sg13g2_buf_1 _23653_ (.A(_05880_),
    .X(_05881_));
 sg13g2_buf_1 _23654_ (.A(_05881_),
    .X(_05882_));
 sg13g2_mux2_1 _23655_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][0] ),
    .A1(net465),
    .S(_05882_),
    .X(_01177_));
 sg13g2_mux2_1 _23656_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][10] ),
    .A1(net513),
    .S(net339),
    .X(_01178_));
 sg13g2_mux2_1 _23657_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][11] ),
    .A1(_05875_),
    .S(net339),
    .X(_01179_));
 sg13g2_mux2_1 _23658_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][1] ),
    .A1(net521),
    .S(net339),
    .X(_01180_));
 sg13g2_mux2_1 _23659_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][2] ),
    .A1(net738),
    .S(net339),
    .X(_01181_));
 sg13g2_mux2_1 _23660_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][3] ),
    .A1(net874),
    .S(net339),
    .X(_01182_));
 sg13g2_mux2_1 _23661_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][4] ),
    .A1(net739),
    .S(net339),
    .X(_01183_));
 sg13g2_buf_1 _23662_ (.A(_02973_),
    .X(_05883_));
 sg13g2_mux2_1 _23663_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][5] ),
    .A1(net869),
    .S(net339),
    .X(_01184_));
 sg13g2_mux2_1 _23664_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][6] ),
    .A1(net873),
    .S(net339),
    .X(_01185_));
 sg13g2_mux2_1 _23665_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][7] ),
    .A1(_03455_),
    .S(_05882_),
    .X(_01186_));
 sg13g2_mux2_1 _23666_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][8] ),
    .A1(net585),
    .S(_05881_),
    .X(_01187_));
 sg13g2_mux2_1 _23667_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][9] ),
    .A1(net649),
    .S(_05881_),
    .X(_01188_));
 sg13g2_nor2_2 _23668_ (.A(_05810_),
    .B(net1024),
    .Y(_05884_));
 sg13g2_nand2_1 _23669_ (.Y(_05885_),
    .A(_05884_),
    .B(_05850_));
 sg13g2_buf_2 _23670_ (.A(_05885_),
    .X(_05886_));
 sg13g2_nor2_1 _23671_ (.A(_05879_),
    .B(_05886_),
    .Y(_05887_));
 sg13g2_buf_1 _23672_ (.A(_05887_),
    .X(_05888_));
 sg13g2_buf_1 _23673_ (.A(_05888_),
    .X(_05889_));
 sg13g2_mux2_1 _23674_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][0] ),
    .A1(net465),
    .S(_05889_),
    .X(_01189_));
 sg13g2_mux2_1 _23675_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][10] ),
    .A1(net513),
    .S(net263),
    .X(_01190_));
 sg13g2_mux2_1 _23676_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][11] ),
    .A1(_05875_),
    .S(net263),
    .X(_01191_));
 sg13g2_mux2_1 _23677_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][1] ),
    .A1(net521),
    .S(net263),
    .X(_01192_));
 sg13g2_mux2_1 _23678_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][2] ),
    .A1(net738),
    .S(net263),
    .X(_01193_));
 sg13g2_mux2_1 _23679_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][3] ),
    .A1(net874),
    .S(net263),
    .X(_01194_));
 sg13g2_mux2_1 _23680_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][4] ),
    .A1(net739),
    .S(net263),
    .X(_01195_));
 sg13g2_mux2_1 _23681_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][5] ),
    .A1(net869),
    .S(net263),
    .X(_01196_));
 sg13g2_mux2_1 _23682_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][6] ),
    .A1(net873),
    .S(net263),
    .X(_01197_));
 sg13g2_mux2_1 _23683_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][7] ),
    .A1(_03455_),
    .S(_05889_),
    .X(_01198_));
 sg13g2_mux2_1 _23684_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][8] ),
    .A1(net585),
    .S(_05888_),
    .X(_01199_));
 sg13g2_mux2_1 _23685_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][9] ),
    .A1(net649),
    .S(_05888_),
    .X(_01200_));
 sg13g2_nand2_1 _23686_ (.Y(_05890_),
    .A(_05858_),
    .B(_05856_));
 sg13g2_nor2_1 _23687_ (.A(_05879_),
    .B(_05890_),
    .Y(_05891_));
 sg13g2_buf_1 _23688_ (.A(_05891_),
    .X(_05892_));
 sg13g2_buf_1 _23689_ (.A(_05892_),
    .X(_05893_));
 sg13g2_mux2_1 _23690_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][0] ),
    .A1(net465),
    .S(net262),
    .X(_01201_));
 sg13g2_mux2_1 _23691_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][10] ),
    .A1(net513),
    .S(net262),
    .X(_01202_));
 sg13g2_mux2_1 _23692_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][11] ),
    .A1(net737),
    .S(net262),
    .X(_01203_));
 sg13g2_mux2_1 _23693_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][1] ),
    .A1(_03465_),
    .S(_05893_),
    .X(_01204_));
 sg13g2_mux2_1 _23694_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][2] ),
    .A1(_05855_),
    .S(net262),
    .X(_01205_));
 sg13g2_mux2_1 _23695_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][3] ),
    .A1(net874),
    .S(net262),
    .X(_01206_));
 sg13g2_mux2_1 _23696_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][4] ),
    .A1(net739),
    .S(net262),
    .X(_01207_));
 sg13g2_mux2_1 _23697_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][5] ),
    .A1(net869),
    .S(net262),
    .X(_01208_));
 sg13g2_mux2_1 _23698_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][6] ),
    .A1(net873),
    .S(net262),
    .X(_01209_));
 sg13g2_buf_1 _23699_ (.A(net981),
    .X(_05894_));
 sg13g2_mux2_1 _23700_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][7] ),
    .A1(net868),
    .S(_05893_),
    .X(_01210_));
 sg13g2_mux2_1 _23701_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][8] ),
    .A1(_05867_),
    .S(_05892_),
    .X(_01211_));
 sg13g2_mux2_1 _23702_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][9] ),
    .A1(_05868_),
    .S(_05892_),
    .X(_01212_));
 sg13g2_or2_1 _23703_ (.X(_05895_),
    .B(_05849_),
    .A(_10930_));
 sg13g2_buf_2 _23704_ (.A(_05895_),
    .X(_05896_));
 sg13g2_nor3_1 _23705_ (.A(_05827_),
    .B(_05896_),
    .C(_05879_),
    .Y(_05897_));
 sg13g2_buf_1 _23706_ (.A(_05897_),
    .X(_05898_));
 sg13g2_buf_1 _23707_ (.A(_05898_),
    .X(_05899_));
 sg13g2_mux2_1 _23708_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][0] ),
    .A1(_05876_),
    .S(net338),
    .X(_01213_));
 sg13g2_mux2_1 _23709_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][10] ),
    .A1(net513),
    .S(net338),
    .X(_01214_));
 sg13g2_mux2_1 _23710_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][11] ),
    .A1(net737),
    .S(net338),
    .X(_01215_));
 sg13g2_mux2_1 _23711_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][1] ),
    .A1(_03465_),
    .S(_05899_),
    .X(_01216_));
 sg13g2_mux2_1 _23712_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][2] ),
    .A1(_05855_),
    .S(net338),
    .X(_01217_));
 sg13g2_mux2_1 _23713_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][3] ),
    .A1(net874),
    .S(net338),
    .X(_01218_));
 sg13g2_mux2_1 _23714_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][4] ),
    .A1(net739),
    .S(net338),
    .X(_01219_));
 sg13g2_mux2_1 _23715_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][5] ),
    .A1(_05883_),
    .S(net338),
    .X(_01220_));
 sg13g2_mux2_1 _23716_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][6] ),
    .A1(net873),
    .S(net338),
    .X(_01221_));
 sg13g2_mux2_1 _23717_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][7] ),
    .A1(_05894_),
    .S(_05899_),
    .X(_01222_));
 sg13g2_mux2_1 _23718_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][8] ),
    .A1(_05867_),
    .S(_05898_),
    .X(_01223_));
 sg13g2_mux2_1 _23719_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][9] ),
    .A1(_05868_),
    .S(_05898_),
    .X(_01224_));
 sg13g2_nand2_1 _23720_ (.Y(_05900_),
    .A(_10819_),
    .B(_05837_));
 sg13g2_buf_2 _23721_ (.A(_05900_),
    .X(_05901_));
 sg13g2_nand2_2 _23722_ (.Y(_05902_),
    .A(net870),
    .B(_05817_));
 sg13g2_nor3_1 _23723_ (.A(_05896_),
    .B(_05901_),
    .C(_05902_),
    .Y(_05903_));
 sg13g2_buf_1 _23724_ (.A(_05903_),
    .X(_05904_));
 sg13g2_buf_1 _23725_ (.A(_05904_),
    .X(_05905_));
 sg13g2_mux2_1 _23726_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][0] ),
    .A1(net465),
    .S(net337),
    .X(_01225_));
 sg13g2_mux2_1 _23727_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][10] ),
    .A1(net513),
    .S(net337),
    .X(_01226_));
 sg13g2_mux2_1 _23728_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][11] ),
    .A1(net737),
    .S(net337),
    .X(_01227_));
 sg13g2_buf_1 _23729_ (.A(net602),
    .X(_05906_));
 sg13g2_mux2_1 _23730_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][1] ),
    .A1(net512),
    .S(net337),
    .X(_01228_));
 sg13g2_mux2_1 _23731_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][2] ),
    .A1(net738),
    .S(_05905_),
    .X(_01229_));
 sg13g2_mux2_1 _23732_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][3] ),
    .A1(net874),
    .S(net337),
    .X(_01230_));
 sg13g2_mux2_1 _23733_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][4] ),
    .A1(_04741_),
    .S(net337),
    .X(_01231_));
 sg13g2_mux2_1 _23734_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][5] ),
    .A1(net869),
    .S(net337),
    .X(_01232_));
 sg13g2_mux2_1 _23735_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][6] ),
    .A1(net873),
    .S(net337),
    .X(_01233_));
 sg13g2_mux2_1 _23736_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][7] ),
    .A1(net868),
    .S(_05905_),
    .X(_01234_));
 sg13g2_mux2_1 _23737_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][8] ),
    .A1(net585),
    .S(_05904_),
    .X(_01235_));
 sg13g2_mux2_1 _23738_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][9] ),
    .A1(net649),
    .S(_05904_),
    .X(_01236_));
 sg13g2_nor3_1 _23739_ (.A(net972),
    .B(_05886_),
    .C(_05901_),
    .Y(_05907_));
 sg13g2_buf_1 _23740_ (.A(_05907_),
    .X(_05908_));
 sg13g2_buf_1 _23741_ (.A(_05908_),
    .X(_05909_));
 sg13g2_mux2_1 _23742_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][0] ),
    .A1(net465),
    .S(net261),
    .X(_01237_));
 sg13g2_mux2_1 _23743_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][10] ),
    .A1(net513),
    .S(net261),
    .X(_01238_));
 sg13g2_mux2_1 _23744_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][11] ),
    .A1(net737),
    .S(net261),
    .X(_01239_));
 sg13g2_mux2_1 _23745_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][1] ),
    .A1(_05906_),
    .S(net261),
    .X(_01240_));
 sg13g2_mux2_1 _23746_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][2] ),
    .A1(net738),
    .S(net261),
    .X(_01241_));
 sg13g2_mux2_1 _23747_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][3] ),
    .A1(net874),
    .S(net261),
    .X(_01242_));
 sg13g2_mux2_1 _23748_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][4] ),
    .A1(net739),
    .S(net261),
    .X(_01243_));
 sg13g2_mux2_1 _23749_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][5] ),
    .A1(net869),
    .S(_05909_),
    .X(_01244_));
 sg13g2_mux2_1 _23750_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][6] ),
    .A1(net873),
    .S(net261),
    .X(_01245_));
 sg13g2_mux2_1 _23751_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][7] ),
    .A1(net868),
    .S(_05909_),
    .X(_01246_));
 sg13g2_mux2_1 _23752_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][8] ),
    .A1(net585),
    .S(_05908_),
    .X(_01247_));
 sg13g2_mux2_1 _23753_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][9] ),
    .A1(net649),
    .S(_05908_),
    .X(_01248_));
 sg13g2_nor2_2 _23754_ (.A(_05860_),
    .B(_05901_),
    .Y(_05910_));
 sg13g2_and2_1 _23755_ (.A(net466),
    .B(_05910_),
    .X(_05911_));
 sg13g2_buf_1 _23756_ (.A(_05911_),
    .X(_05912_));
 sg13g2_buf_1 _23757_ (.A(_05912_),
    .X(_05913_));
 sg13g2_mux2_1 _23758_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][0] ),
    .A1(net465),
    .S(net336),
    .X(_01249_));
 sg13g2_mux2_1 _23759_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][10] ),
    .A1(net513),
    .S(net336),
    .X(_01250_));
 sg13g2_mux2_1 _23760_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][11] ),
    .A1(net737),
    .S(net336),
    .X(_01251_));
 sg13g2_mux2_1 _23761_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][1] ),
    .A1(net512),
    .S(net336),
    .X(_01252_));
 sg13g2_mux2_1 _23762_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][2] ),
    .A1(net738),
    .S(_05913_),
    .X(_01253_));
 sg13g2_buf_1 _23763_ (.A(net983),
    .X(_05914_));
 sg13g2_mux2_1 _23764_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][3] ),
    .A1(_05914_),
    .S(net336),
    .X(_01254_));
 sg13g2_buf_1 _23765_ (.A(_09279_),
    .X(_05915_));
 sg13g2_mux2_1 _23766_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][4] ),
    .A1(_05915_),
    .S(net336),
    .X(_01255_));
 sg13g2_mux2_1 _23767_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][5] ),
    .A1(net869),
    .S(net336),
    .X(_01256_));
 sg13g2_buf_1 _23768_ (.A(net1107),
    .X(_05916_));
 sg13g2_mux2_1 _23769_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][6] ),
    .A1(_05916_),
    .S(net336),
    .X(_01257_));
 sg13g2_mux2_1 _23770_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][7] ),
    .A1(net868),
    .S(_05913_),
    .X(_01258_));
 sg13g2_mux2_1 _23771_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][8] ),
    .A1(net585),
    .S(_05912_),
    .X(_01259_));
 sg13g2_mux2_1 _23772_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][9] ),
    .A1(net649),
    .S(_05912_),
    .X(_01260_));
 sg13g2_nor3_1 _23773_ (.A(net972),
    .B(_05827_),
    .C(_05901_),
    .Y(_05917_));
 sg13g2_buf_2 _23774_ (.A(_05917_),
    .X(_05918_));
 sg13g2_and2_1 _23775_ (.A(net466),
    .B(_05918_),
    .X(_05919_));
 sg13g2_buf_1 _23776_ (.A(_05919_),
    .X(_05920_));
 sg13g2_buf_1 _23777_ (.A(_05920_),
    .X(_05921_));
 sg13g2_mux2_1 _23778_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][0] ),
    .A1(net465),
    .S(net335),
    .X(_01261_));
 sg13g2_mux2_1 _23779_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][10] ),
    .A1(net513),
    .S(net335),
    .X(_01262_));
 sg13g2_mux2_1 _23780_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][11] ),
    .A1(net737),
    .S(net335),
    .X(_01263_));
 sg13g2_mux2_1 _23781_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][1] ),
    .A1(net512),
    .S(net335),
    .X(_01264_));
 sg13g2_buf_1 _23782_ (.A(_02950_),
    .X(_05922_));
 sg13g2_mux2_1 _23783_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][2] ),
    .A1(_05922_),
    .S(_05921_),
    .X(_01265_));
 sg13g2_mux2_1 _23784_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][3] ),
    .A1(net867),
    .S(net335),
    .X(_01266_));
 sg13g2_mux2_1 _23785_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][4] ),
    .A1(net866),
    .S(net335),
    .X(_01267_));
 sg13g2_mux2_1 _23786_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][5] ),
    .A1(net869),
    .S(net335),
    .X(_01268_));
 sg13g2_mux2_1 _23787_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][6] ),
    .A1(net969),
    .S(net335),
    .X(_01269_));
 sg13g2_mux2_1 _23788_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][7] ),
    .A1(net868),
    .S(_05921_),
    .X(_01270_));
 sg13g2_mux2_1 _23789_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][8] ),
    .A1(net585),
    .S(_05920_),
    .X(_01271_));
 sg13g2_mux2_1 _23790_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][9] ),
    .A1(net649),
    .S(_05920_),
    .X(_01272_));
 sg13g2_nor2_1 _23791_ (.A(_05848_),
    .B(_05886_),
    .Y(_05923_));
 sg13g2_buf_1 _23792_ (.A(_05923_),
    .X(_05924_));
 sg13g2_buf_1 _23793_ (.A(_05924_),
    .X(_05925_));
 sg13g2_mux2_1 _23794_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][0] ),
    .A1(_05876_),
    .S(net260),
    .X(_01273_));
 sg13g2_buf_1 _23795_ (.A(net622),
    .X(_05926_));
 sg13g2_mux2_1 _23796_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][10] ),
    .A1(_05926_),
    .S(net260),
    .X(_01274_));
 sg13g2_mux2_1 _23797_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][11] ),
    .A1(net737),
    .S(_05925_),
    .X(_01275_));
 sg13g2_mux2_1 _23798_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][1] ),
    .A1(_05906_),
    .S(net260),
    .X(_01276_));
 sg13g2_mux2_1 _23799_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][2] ),
    .A1(_05922_),
    .S(net260),
    .X(_01277_));
 sg13g2_mux2_1 _23800_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][3] ),
    .A1(_05914_),
    .S(net260),
    .X(_01278_));
 sg13g2_mux2_1 _23801_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][4] ),
    .A1(_05915_),
    .S(net260),
    .X(_01279_));
 sg13g2_mux2_1 _23802_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][5] ),
    .A1(_05883_),
    .S(net260),
    .X(_01280_));
 sg13g2_mux2_1 _23803_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][6] ),
    .A1(_05916_),
    .S(_05925_),
    .X(_01281_));
 sg13g2_mux2_1 _23804_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][7] ),
    .A1(_05894_),
    .S(net260),
    .X(_01282_));
 sg13g2_buf_1 _23805_ (.A(net687),
    .X(_05927_));
 sg13g2_mux2_1 _23806_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][8] ),
    .A1(_05927_),
    .S(_05924_),
    .X(_01283_));
 sg13g2_buf_1 _23807_ (.A(net791),
    .X(_05928_));
 sg13g2_mux2_1 _23808_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][9] ),
    .A1(_05928_),
    .S(_05924_),
    .X(_01284_));
 sg13g2_or2_1 _23809_ (.X(_05929_),
    .B(_05901_),
    .A(_05845_));
 sg13g2_buf_1 _23810_ (.A(_05929_),
    .X(_05930_));
 sg13g2_nor2_1 _23811_ (.A(_05851_),
    .B(_05930_),
    .Y(_05931_));
 sg13g2_buf_1 _23812_ (.A(_05931_),
    .X(_05932_));
 sg13g2_buf_1 _23813_ (.A(_05932_),
    .X(_05933_));
 sg13g2_mux2_1 _23814_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][0] ),
    .A1(net465),
    .S(net334),
    .X(_01285_));
 sg13g2_mux2_1 _23815_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][10] ),
    .A1(net511),
    .S(net334),
    .X(_01286_));
 sg13g2_buf_1 _23816_ (.A(_09632_),
    .X(_05934_));
 sg13g2_mux2_1 _23817_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][11] ),
    .A1(net736),
    .S(_05933_),
    .X(_01287_));
 sg13g2_mux2_1 _23818_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][1] ),
    .A1(net512),
    .S(net334),
    .X(_01288_));
 sg13g2_mux2_1 _23819_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][2] ),
    .A1(net865),
    .S(net334),
    .X(_01289_));
 sg13g2_mux2_1 _23820_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][3] ),
    .A1(net867),
    .S(net334),
    .X(_01290_));
 sg13g2_mux2_1 _23821_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][4] ),
    .A1(net866),
    .S(net334),
    .X(_01291_));
 sg13g2_mux2_1 _23822_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][5] ),
    .A1(net869),
    .S(_05933_),
    .X(_01292_));
 sg13g2_mux2_1 _23823_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][6] ),
    .A1(net969),
    .S(net334),
    .X(_01293_));
 sg13g2_mux2_1 _23824_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][7] ),
    .A1(net868),
    .S(net334),
    .X(_01294_));
 sg13g2_mux2_1 _23825_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][8] ),
    .A1(net584),
    .S(_05932_),
    .X(_01295_));
 sg13g2_mux2_1 _23826_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][9] ),
    .A1(net648),
    .S(_05932_),
    .X(_01296_));
 sg13g2_buf_1 _23827_ (.A(_03435_),
    .X(_05935_));
 sg13g2_nor2_1 _23828_ (.A(_05886_),
    .B(_05930_),
    .Y(_05936_));
 sg13g2_buf_1 _23829_ (.A(_05936_),
    .X(_05937_));
 sg13g2_buf_1 _23830_ (.A(_05937_),
    .X(_05938_));
 sg13g2_mux2_1 _23831_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][0] ),
    .A1(_05935_),
    .S(_05938_),
    .X(_01297_));
 sg13g2_mux2_1 _23832_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][10] ),
    .A1(net511),
    .S(net259),
    .X(_01298_));
 sg13g2_mux2_1 _23833_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][11] ),
    .A1(_05934_),
    .S(net259),
    .X(_01299_));
 sg13g2_mux2_1 _23834_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][1] ),
    .A1(net512),
    .S(net259),
    .X(_01300_));
 sg13g2_mux2_1 _23835_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][2] ),
    .A1(net865),
    .S(_05938_),
    .X(_01301_));
 sg13g2_mux2_1 _23836_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][3] ),
    .A1(net867),
    .S(net259),
    .X(_01302_));
 sg13g2_mux2_1 _23837_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][4] ),
    .A1(net866),
    .S(net259),
    .X(_01303_));
 sg13g2_buf_1 _23838_ (.A(_02973_),
    .X(_05939_));
 sg13g2_mux2_1 _23839_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][5] ),
    .A1(net864),
    .S(net259),
    .X(_01304_));
 sg13g2_mux2_1 _23840_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][6] ),
    .A1(net969),
    .S(net259),
    .X(_01305_));
 sg13g2_mux2_1 _23841_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][7] ),
    .A1(net868),
    .S(net259),
    .X(_01306_));
 sg13g2_mux2_1 _23842_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][8] ),
    .A1(net584),
    .S(_05937_),
    .X(_01307_));
 sg13g2_mux2_1 _23843_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][9] ),
    .A1(_05928_),
    .S(_05937_),
    .X(_01308_));
 sg13g2_nor2_1 _23844_ (.A(_05890_),
    .B(_05930_),
    .Y(_05940_));
 sg13g2_buf_1 _23845_ (.A(_05940_),
    .X(_05941_));
 sg13g2_buf_1 _23846_ (.A(_05941_),
    .X(_05942_));
 sg13g2_mux2_1 _23847_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][0] ),
    .A1(net464),
    .S(_05942_),
    .X(_01309_));
 sg13g2_mux2_1 _23848_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][10] ),
    .A1(net511),
    .S(net258),
    .X(_01310_));
 sg13g2_mux2_1 _23849_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][11] ),
    .A1(_05934_),
    .S(net258),
    .X(_01311_));
 sg13g2_mux2_1 _23850_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][1] ),
    .A1(net512),
    .S(net258),
    .X(_01312_));
 sg13g2_mux2_1 _23851_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][2] ),
    .A1(net865),
    .S(_05942_),
    .X(_01313_));
 sg13g2_mux2_1 _23852_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][3] ),
    .A1(net867),
    .S(net258),
    .X(_01314_));
 sg13g2_mux2_1 _23853_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][4] ),
    .A1(net866),
    .S(net258),
    .X(_01315_));
 sg13g2_mux2_1 _23854_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][5] ),
    .A1(net864),
    .S(net258),
    .X(_01316_));
 sg13g2_mux2_1 _23855_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][6] ),
    .A1(net969),
    .S(net258),
    .X(_01317_));
 sg13g2_mux2_1 _23856_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][7] ),
    .A1(net868),
    .S(net258),
    .X(_01318_));
 sg13g2_mux2_1 _23857_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][8] ),
    .A1(net584),
    .S(_05941_),
    .X(_01319_));
 sg13g2_mux2_1 _23858_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][9] ),
    .A1(net648),
    .S(_05941_),
    .X(_01320_));
 sg13g2_nor3_1 _23859_ (.A(_05827_),
    .B(_05896_),
    .C(_05930_),
    .Y(_05943_));
 sg13g2_buf_1 _23860_ (.A(_05943_),
    .X(_05944_));
 sg13g2_buf_1 _23861_ (.A(_05944_),
    .X(_05945_));
 sg13g2_mux2_1 _23862_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][0] ),
    .A1(net464),
    .S(_05945_),
    .X(_01321_));
 sg13g2_mux2_1 _23863_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][10] ),
    .A1(net511),
    .S(net333),
    .X(_01322_));
 sg13g2_mux2_1 _23864_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][11] ),
    .A1(net736),
    .S(net333),
    .X(_01323_));
 sg13g2_mux2_1 _23865_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][1] ),
    .A1(net512),
    .S(net333),
    .X(_01324_));
 sg13g2_mux2_1 _23866_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][2] ),
    .A1(net865),
    .S(_05945_),
    .X(_01325_));
 sg13g2_mux2_1 _23867_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][3] ),
    .A1(net867),
    .S(net333),
    .X(_01326_));
 sg13g2_mux2_1 _23868_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][4] ),
    .A1(net866),
    .S(net333),
    .X(_01327_));
 sg13g2_mux2_1 _23869_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][5] ),
    .A1(net864),
    .S(net333),
    .X(_01328_));
 sg13g2_mux2_1 _23870_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][6] ),
    .A1(net969),
    .S(net333),
    .X(_01329_));
 sg13g2_buf_1 _23871_ (.A(_10680_),
    .X(_05946_));
 sg13g2_mux2_1 _23872_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][7] ),
    .A1(net968),
    .S(net333),
    .X(_01330_));
 sg13g2_mux2_1 _23873_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][8] ),
    .A1(net584),
    .S(_05944_),
    .X(_01331_));
 sg13g2_mux2_1 _23874_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][9] ),
    .A1(net648),
    .S(_05944_),
    .X(_01332_));
 sg13g2_nand2_1 _23875_ (.Y(_05947_),
    .A(_10819_),
    .B(net971));
 sg13g2_buf_2 _23876_ (.A(_05947_),
    .X(_05948_));
 sg13g2_nor3_1 _23877_ (.A(_05896_),
    .B(_05902_),
    .C(_05948_),
    .Y(_05949_));
 sg13g2_buf_1 _23878_ (.A(_05949_),
    .X(_05950_));
 sg13g2_buf_1 _23879_ (.A(_05950_),
    .X(_05951_));
 sg13g2_mux2_1 _23880_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][0] ),
    .A1(net464),
    .S(net332),
    .X(_01333_));
 sg13g2_mux2_1 _23881_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][10] ),
    .A1(net511),
    .S(net332),
    .X(_01334_));
 sg13g2_mux2_1 _23882_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][11] ),
    .A1(net736),
    .S(net332),
    .X(_01335_));
 sg13g2_mux2_1 _23883_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][1] ),
    .A1(net512),
    .S(_05951_),
    .X(_01336_));
 sg13g2_mux2_1 _23884_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][2] ),
    .A1(net865),
    .S(net332),
    .X(_01337_));
 sg13g2_mux2_1 _23885_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][3] ),
    .A1(net867),
    .S(net332),
    .X(_01338_));
 sg13g2_mux2_1 _23886_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][4] ),
    .A1(net866),
    .S(net332),
    .X(_01339_));
 sg13g2_mux2_1 _23887_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][5] ),
    .A1(net864),
    .S(net332),
    .X(_01340_));
 sg13g2_mux2_1 _23888_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][6] ),
    .A1(net969),
    .S(net332),
    .X(_01341_));
 sg13g2_mux2_1 _23889_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][7] ),
    .A1(net968),
    .S(_05951_),
    .X(_01342_));
 sg13g2_mux2_1 _23890_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][8] ),
    .A1(net584),
    .S(_05950_),
    .X(_01343_));
 sg13g2_mux2_1 _23891_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][9] ),
    .A1(net648),
    .S(_05950_),
    .X(_01344_));
 sg13g2_nor3_1 _23892_ (.A(net972),
    .B(_05886_),
    .C(_05948_),
    .Y(_05952_));
 sg13g2_buf_1 _23893_ (.A(_05952_),
    .X(_05953_));
 sg13g2_buf_1 _23894_ (.A(_05953_),
    .X(_05954_));
 sg13g2_mux2_1 _23895_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][0] ),
    .A1(net464),
    .S(net257),
    .X(_01345_));
 sg13g2_mux2_1 _23896_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][10] ),
    .A1(net511),
    .S(net257),
    .X(_01346_));
 sg13g2_mux2_1 _23897_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][11] ),
    .A1(net736),
    .S(net257),
    .X(_01347_));
 sg13g2_buf_1 _23898_ (.A(_02965_),
    .X(_05955_));
 sg13g2_mux2_1 _23899_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][1] ),
    .A1(net583),
    .S(_05954_),
    .X(_01348_));
 sg13g2_mux2_1 _23900_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][2] ),
    .A1(net865),
    .S(net257),
    .X(_01349_));
 sg13g2_mux2_1 _23901_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][3] ),
    .A1(net867),
    .S(net257),
    .X(_01350_));
 sg13g2_mux2_1 _23902_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][4] ),
    .A1(net866),
    .S(net257),
    .X(_01351_));
 sg13g2_mux2_1 _23903_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][5] ),
    .A1(net864),
    .S(net257),
    .X(_01352_));
 sg13g2_mux2_1 _23904_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][6] ),
    .A1(net969),
    .S(net257),
    .X(_01353_));
 sg13g2_mux2_1 _23905_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][7] ),
    .A1(net968),
    .S(_05954_),
    .X(_01354_));
 sg13g2_mux2_1 _23906_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][8] ),
    .A1(net584),
    .S(_05953_),
    .X(_01355_));
 sg13g2_mux2_1 _23907_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][9] ),
    .A1(net648),
    .S(_05953_),
    .X(_01356_));
 sg13g2_nor2_2 _23908_ (.A(_05860_),
    .B(_05948_),
    .Y(_05956_));
 sg13g2_and2_1 _23909_ (.A(net466),
    .B(_05956_),
    .X(_05957_));
 sg13g2_buf_1 _23910_ (.A(_05957_),
    .X(_05958_));
 sg13g2_buf_1 _23911_ (.A(_05958_),
    .X(_05959_));
 sg13g2_mux2_1 _23912_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][0] ),
    .A1(net464),
    .S(net331),
    .X(_01357_));
 sg13g2_mux2_1 _23913_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][10] ),
    .A1(net511),
    .S(net331),
    .X(_01358_));
 sg13g2_mux2_1 _23914_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][11] ),
    .A1(net736),
    .S(net331),
    .X(_01359_));
 sg13g2_mux2_1 _23915_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][1] ),
    .A1(net583),
    .S(_05959_),
    .X(_01360_));
 sg13g2_mux2_1 _23916_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][2] ),
    .A1(net865),
    .S(net331),
    .X(_01361_));
 sg13g2_mux2_1 _23917_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][3] ),
    .A1(net867),
    .S(net331),
    .X(_01362_));
 sg13g2_mux2_1 _23918_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][4] ),
    .A1(net866),
    .S(net331),
    .X(_01363_));
 sg13g2_mux2_1 _23919_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][5] ),
    .A1(net864),
    .S(net331),
    .X(_01364_));
 sg13g2_mux2_1 _23920_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][6] ),
    .A1(net969),
    .S(net331),
    .X(_01365_));
 sg13g2_mux2_1 _23921_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][7] ),
    .A1(net968),
    .S(_05959_),
    .X(_01366_));
 sg13g2_mux2_1 _23922_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][8] ),
    .A1(net584),
    .S(_05958_),
    .X(_01367_));
 sg13g2_mux2_1 _23923_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][9] ),
    .A1(net648),
    .S(_05958_),
    .X(_01368_));
 sg13g2_nor3_1 _23924_ (.A(_05829_),
    .B(_05827_),
    .C(_05948_),
    .Y(_05960_));
 sg13g2_buf_2 _23925_ (.A(_05960_),
    .X(_05961_));
 sg13g2_and2_1 _23926_ (.A(net466),
    .B(_05961_),
    .X(_05962_));
 sg13g2_buf_1 _23927_ (.A(_05962_),
    .X(_05963_));
 sg13g2_buf_1 _23928_ (.A(_05963_),
    .X(_05964_));
 sg13g2_mux2_1 _23929_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][0] ),
    .A1(net464),
    .S(net330),
    .X(_01369_));
 sg13g2_mux2_1 _23930_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][10] ),
    .A1(net511),
    .S(net330),
    .X(_01370_));
 sg13g2_mux2_1 _23931_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][11] ),
    .A1(net736),
    .S(net330),
    .X(_01371_));
 sg13g2_mux2_1 _23932_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][1] ),
    .A1(net583),
    .S(_05964_),
    .X(_01372_));
 sg13g2_mux2_1 _23933_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][2] ),
    .A1(net865),
    .S(net330),
    .X(_01373_));
 sg13g2_buf_1 _23934_ (.A(net983),
    .X(_05965_));
 sg13g2_mux2_1 _23935_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][3] ),
    .A1(net863),
    .S(net330),
    .X(_01374_));
 sg13g2_buf_1 _23936_ (.A(net1056),
    .X(_05966_));
 sg13g2_mux2_1 _23937_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][4] ),
    .A1(net862),
    .S(net330),
    .X(_01375_));
 sg13g2_mux2_1 _23938_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][5] ),
    .A1(net864),
    .S(net330),
    .X(_01376_));
 sg13g2_buf_1 _23939_ (.A(_10645_),
    .X(_05967_));
 sg13g2_mux2_1 _23940_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][6] ),
    .A1(net967),
    .S(net330),
    .X(_01377_));
 sg13g2_mux2_1 _23941_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][7] ),
    .A1(net968),
    .S(_05964_),
    .X(_01378_));
 sg13g2_mux2_1 _23942_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][8] ),
    .A1(net584),
    .S(_05963_),
    .X(_01379_));
 sg13g2_mux2_1 _23943_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][9] ),
    .A1(net648),
    .S(_05963_),
    .X(_01380_));
 sg13g2_or2_1 _23944_ (.X(_05968_),
    .B(_05948_),
    .A(_05845_));
 sg13g2_buf_1 _23945_ (.A(_05968_),
    .X(_05969_));
 sg13g2_nor2_1 _23946_ (.A(_05851_),
    .B(_05969_),
    .Y(_05970_));
 sg13g2_buf_1 _23947_ (.A(_05970_),
    .X(_05971_));
 sg13g2_buf_1 _23948_ (.A(_05971_),
    .X(_05972_));
 sg13g2_mux2_1 _23949_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][0] ),
    .A1(net464),
    .S(net329),
    .X(_01381_));
 sg13g2_mux2_1 _23950_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][10] ),
    .A1(_05926_),
    .S(net329),
    .X(_01382_));
 sg13g2_mux2_1 _23951_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][11] ),
    .A1(net736),
    .S(net329),
    .X(_01383_));
 sg13g2_mux2_1 _23952_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][1] ),
    .A1(net583),
    .S(net329),
    .X(_01384_));
 sg13g2_buf_1 _23953_ (.A(net984),
    .X(_05973_));
 sg13g2_mux2_1 _23954_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][2] ),
    .A1(net861),
    .S(_05972_),
    .X(_01385_));
 sg13g2_mux2_1 _23955_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][3] ),
    .A1(net863),
    .S(net329),
    .X(_01386_));
 sg13g2_mux2_1 _23956_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][4] ),
    .A1(net862),
    .S(net329),
    .X(_01387_));
 sg13g2_mux2_1 _23957_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][5] ),
    .A1(_05939_),
    .S(net329),
    .X(_01388_));
 sg13g2_mux2_1 _23958_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][6] ),
    .A1(net967),
    .S(net329),
    .X(_01389_));
 sg13g2_mux2_1 _23959_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][7] ),
    .A1(net968),
    .S(_05972_),
    .X(_01390_));
 sg13g2_mux2_1 _23960_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][8] ),
    .A1(_05927_),
    .S(_05971_),
    .X(_01391_));
 sg13g2_mux2_1 _23961_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][9] ),
    .A1(net648),
    .S(_05971_),
    .X(_01392_));
 sg13g2_nor2_1 _23962_ (.A(_05886_),
    .B(_05969_),
    .Y(_05974_));
 sg13g2_buf_1 _23963_ (.A(_05974_),
    .X(_05975_));
 sg13g2_buf_1 _23964_ (.A(_05975_),
    .X(_05976_));
 sg13g2_mux2_1 _23965_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][0] ),
    .A1(net464),
    .S(net256),
    .X(_01393_));
 sg13g2_buf_1 _23966_ (.A(_09541_),
    .X(_05977_));
 sg13g2_mux2_1 _23967_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][10] ),
    .A1(net510),
    .S(net256),
    .X(_01394_));
 sg13g2_mux2_1 _23968_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][11] ),
    .A1(net736),
    .S(net256),
    .X(_01395_));
 sg13g2_mux2_1 _23969_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][1] ),
    .A1(net583),
    .S(net256),
    .X(_01396_));
 sg13g2_mux2_1 _23970_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][2] ),
    .A1(net861),
    .S(_05976_),
    .X(_01397_));
 sg13g2_mux2_1 _23971_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][3] ),
    .A1(net863),
    .S(net256),
    .X(_01398_));
 sg13g2_mux2_1 _23972_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][4] ),
    .A1(net862),
    .S(net256),
    .X(_01399_));
 sg13g2_mux2_1 _23973_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][5] ),
    .A1(net864),
    .S(net256),
    .X(_01400_));
 sg13g2_mux2_1 _23974_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][6] ),
    .A1(net967),
    .S(net256),
    .X(_01401_));
 sg13g2_mux2_1 _23975_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][7] ),
    .A1(_05946_),
    .S(_05976_),
    .X(_01402_));
 sg13g2_buf_1 _23976_ (.A(_09682_),
    .X(_05978_));
 sg13g2_mux2_1 _23977_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][8] ),
    .A1(net582),
    .S(_05975_),
    .X(_01403_));
 sg13g2_buf_1 _23978_ (.A(net791),
    .X(_05979_));
 sg13g2_mux2_1 _23979_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][9] ),
    .A1(net647),
    .S(_05975_),
    .X(_01404_));
 sg13g2_nor2_1 _23980_ (.A(_05848_),
    .B(_05890_),
    .Y(_05980_));
 sg13g2_buf_1 _23981_ (.A(_05980_),
    .X(_05981_));
 sg13g2_buf_1 _23982_ (.A(_05981_),
    .X(_05982_));
 sg13g2_mux2_1 _23983_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][0] ),
    .A1(_05935_),
    .S(net255),
    .X(_01405_));
 sg13g2_mux2_1 _23984_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][10] ),
    .A1(net510),
    .S(net255),
    .X(_01406_));
 sg13g2_buf_1 _23985_ (.A(_09632_),
    .X(_05983_));
 sg13g2_mux2_1 _23986_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][11] ),
    .A1(net735),
    .S(net255),
    .X(_01407_));
 sg13g2_mux2_1 _23987_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][1] ),
    .A1(_05955_),
    .S(net255),
    .X(_01408_));
 sg13g2_mux2_1 _23988_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][2] ),
    .A1(net861),
    .S(net255),
    .X(_01409_));
 sg13g2_mux2_1 _23989_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][3] ),
    .A1(net863),
    .S(net255),
    .X(_01410_));
 sg13g2_mux2_1 _23990_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][4] ),
    .A1(net862),
    .S(net255),
    .X(_01411_));
 sg13g2_mux2_1 _23991_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][5] ),
    .A1(_05939_),
    .S(net255),
    .X(_01412_));
 sg13g2_mux2_1 _23992_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][6] ),
    .A1(net967),
    .S(_05982_),
    .X(_01413_));
 sg13g2_mux2_1 _23993_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][7] ),
    .A1(_05946_),
    .S(_05982_),
    .X(_01414_));
 sg13g2_mux2_1 _23994_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][8] ),
    .A1(_05978_),
    .S(_05981_),
    .X(_01415_));
 sg13g2_mux2_1 _23995_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][9] ),
    .A1(net647),
    .S(_05981_),
    .X(_01416_));
 sg13g2_nor2_1 _23996_ (.A(_05890_),
    .B(_05969_),
    .Y(_05984_));
 sg13g2_buf_1 _23997_ (.A(_05984_),
    .X(_05985_));
 sg13g2_buf_1 _23998_ (.A(_05985_),
    .X(_05986_));
 sg13g2_mux2_1 _23999_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][0] ),
    .A1(net473),
    .S(net254),
    .X(_01417_));
 sg13g2_mux2_1 _24000_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][10] ),
    .A1(net510),
    .S(net254),
    .X(_01418_));
 sg13g2_mux2_1 _24001_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][11] ),
    .A1(net735),
    .S(_05986_),
    .X(_01419_));
 sg13g2_mux2_1 _24002_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][1] ),
    .A1(net583),
    .S(net254),
    .X(_01420_));
 sg13g2_mux2_1 _24003_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][2] ),
    .A1(net861),
    .S(_05986_),
    .X(_01421_));
 sg13g2_mux2_1 _24004_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][3] ),
    .A1(net863),
    .S(net254),
    .X(_01422_));
 sg13g2_mux2_1 _24005_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][4] ),
    .A1(net862),
    .S(net254),
    .X(_01423_));
 sg13g2_buf_1 _24006_ (.A(_02973_),
    .X(_05987_));
 sg13g2_mux2_1 _24007_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][5] ),
    .A1(net860),
    .S(net254),
    .X(_01424_));
 sg13g2_mux2_1 _24008_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][6] ),
    .A1(_05967_),
    .S(net254),
    .X(_01425_));
 sg13g2_mux2_1 _24009_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][7] ),
    .A1(net968),
    .S(net254),
    .X(_01426_));
 sg13g2_mux2_1 _24010_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][8] ),
    .A1(net582),
    .S(_05985_),
    .X(_01427_));
 sg13g2_mux2_1 _24011_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][9] ),
    .A1(net647),
    .S(_05985_),
    .X(_01428_));
 sg13g2_nor3_1 _24012_ (.A(_05827_),
    .B(_05896_),
    .C(_05969_),
    .Y(_05988_));
 sg13g2_buf_1 _24013_ (.A(_05988_),
    .X(_05989_));
 sg13g2_buf_1 _24014_ (.A(_05989_),
    .X(_05990_));
 sg13g2_mux2_1 _24015_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][0] ),
    .A1(net473),
    .S(_05990_),
    .X(_01429_));
 sg13g2_mux2_1 _24016_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][10] ),
    .A1(net510),
    .S(net328),
    .X(_01430_));
 sg13g2_mux2_1 _24017_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][11] ),
    .A1(net735),
    .S(net328),
    .X(_01431_));
 sg13g2_mux2_1 _24018_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][1] ),
    .A1(net583),
    .S(net328),
    .X(_01432_));
 sg13g2_mux2_1 _24019_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][2] ),
    .A1(net861),
    .S(_05990_),
    .X(_01433_));
 sg13g2_mux2_1 _24020_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][3] ),
    .A1(_05965_),
    .S(net328),
    .X(_01434_));
 sg13g2_mux2_1 _24021_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][4] ),
    .A1(net862),
    .S(net328),
    .X(_01435_));
 sg13g2_mux2_1 _24022_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][5] ),
    .A1(net860),
    .S(net328),
    .X(_01436_));
 sg13g2_mux2_1 _24023_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][6] ),
    .A1(net967),
    .S(net328),
    .X(_01437_));
 sg13g2_mux2_1 _24024_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][7] ),
    .A1(net968),
    .S(net328),
    .X(_01438_));
 sg13g2_mux2_1 _24025_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][8] ),
    .A1(net582),
    .S(_05989_),
    .X(_01439_));
 sg13g2_mux2_1 _24026_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][9] ),
    .A1(net647),
    .S(_05989_),
    .X(_01440_));
 sg13g2_nor3_1 _24027_ (.A(_05827_),
    .B(_05848_),
    .C(_05896_),
    .Y(_05991_));
 sg13g2_buf_1 _24028_ (.A(_05991_),
    .X(_05992_));
 sg13g2_buf_1 _24029_ (.A(_05992_),
    .X(_05993_));
 sg13g2_mux2_1 _24030_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][0] ),
    .A1(net473),
    .S(net327),
    .X(_01441_));
 sg13g2_mux2_1 _24031_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][10] ),
    .A1(net510),
    .S(net327),
    .X(_01442_));
 sg13g2_mux2_1 _24032_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][11] ),
    .A1(net735),
    .S(_05993_),
    .X(_01443_));
 sg13g2_mux2_1 _24033_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][1] ),
    .A1(net583),
    .S(net327),
    .X(_01444_));
 sg13g2_mux2_1 _24034_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][2] ),
    .A1(net861),
    .S(net327),
    .X(_01445_));
 sg13g2_mux2_1 _24035_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][3] ),
    .A1(net863),
    .S(net327),
    .X(_01446_));
 sg13g2_mux2_1 _24036_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][4] ),
    .A1(_05966_),
    .S(net327),
    .X(_01447_));
 sg13g2_mux2_1 _24037_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][5] ),
    .A1(net860),
    .S(net327),
    .X(_01448_));
 sg13g2_mux2_1 _24038_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][6] ),
    .A1(net967),
    .S(_05993_),
    .X(_01449_));
 sg13g2_mux2_1 _24039_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][7] ),
    .A1(net981),
    .S(net327),
    .X(_01450_));
 sg13g2_mux2_1 _24040_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][8] ),
    .A1(_05978_),
    .S(_05992_),
    .X(_01451_));
 sg13g2_mux2_1 _24041_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][9] ),
    .A1(_05979_),
    .S(_05992_),
    .X(_01452_));
 sg13g2_nand2_1 _24042_ (.Y(_05994_),
    .A(net1109),
    .B(_05837_));
 sg13g2_nor3_1 _24043_ (.A(net970),
    .B(_05851_),
    .C(_05994_),
    .Y(_05995_));
 sg13g2_buf_1 _24044_ (.A(_05995_),
    .X(_05996_));
 sg13g2_buf_1 _24045_ (.A(_05996_),
    .X(_05997_));
 sg13g2_mux2_1 _24046_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][0] ),
    .A1(net473),
    .S(net326),
    .X(_01453_));
 sg13g2_mux2_1 _24047_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][10] ),
    .A1(net510),
    .S(_05997_),
    .X(_01454_));
 sg13g2_mux2_1 _24048_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][11] ),
    .A1(net735),
    .S(net326),
    .X(_01455_));
 sg13g2_mux2_1 _24049_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][1] ),
    .A1(_05955_),
    .S(net326),
    .X(_01456_));
 sg13g2_mux2_1 _24050_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][2] ),
    .A1(net861),
    .S(net326),
    .X(_01457_));
 sg13g2_mux2_1 _24051_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][3] ),
    .A1(net863),
    .S(net326),
    .X(_01458_));
 sg13g2_mux2_1 _24052_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][4] ),
    .A1(net862),
    .S(net326),
    .X(_01459_));
 sg13g2_mux2_1 _24053_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][5] ),
    .A1(net860),
    .S(net326),
    .X(_01460_));
 sg13g2_mux2_1 _24054_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][6] ),
    .A1(net967),
    .S(_05997_),
    .X(_01461_));
 sg13g2_mux2_1 _24055_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][7] ),
    .A1(net981),
    .S(net326),
    .X(_01462_));
 sg13g2_mux2_1 _24056_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][8] ),
    .A1(net582),
    .S(_05996_),
    .X(_01463_));
 sg13g2_mux2_1 _24057_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][9] ),
    .A1(net647),
    .S(_05996_),
    .X(_01464_));
 sg13g2_nor3_1 _24058_ (.A(net1024),
    .B(_05869_),
    .C(_05994_),
    .Y(_05998_));
 sg13g2_buf_2 _24059_ (.A(_05998_),
    .X(_05999_));
 sg13g2_and2_1 _24060_ (.A(net466),
    .B(_05999_),
    .X(_06000_));
 sg13g2_buf_1 _24061_ (.A(_06000_),
    .X(_06001_));
 sg13g2_buf_1 _24062_ (.A(_06001_),
    .X(_06002_));
 sg13g2_mux2_1 _24063_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][0] ),
    .A1(net473),
    .S(net325),
    .X(_01465_));
 sg13g2_mux2_1 _24064_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][10] ),
    .A1(net510),
    .S(net325),
    .X(_01466_));
 sg13g2_mux2_1 _24065_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][11] ),
    .A1(net735),
    .S(net325),
    .X(_01467_));
 sg13g2_mux2_1 _24066_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][1] ),
    .A1(net602),
    .S(net325),
    .X(_01468_));
 sg13g2_mux2_1 _24067_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][2] ),
    .A1(net861),
    .S(_06002_),
    .X(_01469_));
 sg13g2_mux2_1 _24068_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][3] ),
    .A1(net863),
    .S(net325),
    .X(_01470_));
 sg13g2_mux2_1 _24069_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][4] ),
    .A1(_05966_),
    .S(net325),
    .X(_01471_));
 sg13g2_mux2_1 _24070_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][5] ),
    .A1(net860),
    .S(net325),
    .X(_01472_));
 sg13g2_mux2_1 _24071_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][6] ),
    .A1(net967),
    .S(_06002_),
    .X(_01473_));
 sg13g2_mux2_1 _24072_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][7] ),
    .A1(net981),
    .S(net325),
    .X(_01474_));
 sg13g2_mux2_1 _24073_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][8] ),
    .A1(net582),
    .S(_06001_),
    .X(_01475_));
 sg13g2_mux2_1 _24074_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][9] ),
    .A1(net647),
    .S(_06001_),
    .X(_01476_));
 sg13g2_nor2_1 _24075_ (.A(_05822_),
    .B(net971),
    .Y(_06003_));
 sg13g2_nand2_1 _24076_ (.Y(_06004_),
    .A(net1024),
    .B(_06003_));
 sg13g2_nor3_2 _24077_ (.A(net970),
    .B(net973),
    .C(_06004_),
    .Y(_06005_));
 sg13g2_and2_1 _24078_ (.A(_05856_),
    .B(_06005_),
    .X(_06006_));
 sg13g2_buf_1 _24079_ (.A(_06006_),
    .X(_06007_));
 sg13g2_buf_1 _24080_ (.A(_06007_),
    .X(_06008_));
 sg13g2_mux2_1 _24081_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][0] ),
    .A1(net473),
    .S(net324),
    .X(_01477_));
 sg13g2_mux2_1 _24082_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][10] ),
    .A1(_05977_),
    .S(_06008_),
    .X(_01478_));
 sg13g2_mux2_1 _24083_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][11] ),
    .A1(net735),
    .S(net324),
    .X(_01479_));
 sg13g2_mux2_1 _24084_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][1] ),
    .A1(net602),
    .S(net324),
    .X(_01480_));
 sg13g2_mux2_1 _24085_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][2] ),
    .A1(_05973_),
    .S(net324),
    .X(_01481_));
 sg13g2_mux2_1 _24086_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][3] ),
    .A1(_05965_),
    .S(net324),
    .X(_01482_));
 sg13g2_mux2_1 _24087_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][4] ),
    .A1(net862),
    .S(net324),
    .X(_01483_));
 sg13g2_mux2_1 _24088_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][5] ),
    .A1(net860),
    .S(net324),
    .X(_01484_));
 sg13g2_mux2_1 _24089_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][6] ),
    .A1(_05967_),
    .S(_06008_),
    .X(_01485_));
 sg13g2_mux2_1 _24090_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][7] ),
    .A1(net981),
    .S(net324),
    .X(_01486_));
 sg13g2_mux2_1 _24091_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][8] ),
    .A1(net582),
    .S(_06007_),
    .X(_01487_));
 sg13g2_mux2_1 _24092_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][9] ),
    .A1(net647),
    .S(_06007_),
    .X(_01488_));
 sg13g2_nor2_1 _24093_ (.A(_05869_),
    .B(_06004_),
    .Y(_06009_));
 sg13g2_buf_2 _24094_ (.A(_06009_),
    .X(_06010_));
 sg13g2_and2_1 _24095_ (.A(net466),
    .B(_06010_),
    .X(_06011_));
 sg13g2_buf_1 _24096_ (.A(_06011_),
    .X(_06012_));
 sg13g2_buf_1 _24097_ (.A(_06012_),
    .X(_06013_));
 sg13g2_mux2_1 _24098_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][0] ),
    .A1(_03463_),
    .S(net323),
    .X(_01489_));
 sg13g2_mux2_1 _24099_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][10] ),
    .A1(_05977_),
    .S(net323),
    .X(_01490_));
 sg13g2_mux2_1 _24100_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][11] ),
    .A1(net735),
    .S(net323),
    .X(_01491_));
 sg13g2_mux2_1 _24101_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][1] ),
    .A1(net602),
    .S(net323),
    .X(_01492_));
 sg13g2_mux2_1 _24102_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][2] ),
    .A1(_05973_),
    .S(net323),
    .X(_01493_));
 sg13g2_mux2_1 _24103_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][3] ),
    .A1(net888),
    .S(net323),
    .X(_01494_));
 sg13g2_mux2_1 _24104_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][4] ),
    .A1(net887),
    .S(net323),
    .X(_01495_));
 sg13g2_mux2_1 _24105_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][5] ),
    .A1(net860),
    .S(_06013_),
    .X(_01496_));
 sg13g2_mux2_1 _24106_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][6] ),
    .A1(net982),
    .S(_06013_),
    .X(_01497_));
 sg13g2_mux2_1 _24107_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][7] ),
    .A1(net981),
    .S(net323),
    .X(_01498_));
 sg13g2_mux2_1 _24108_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][8] ),
    .A1(net582),
    .S(_06012_),
    .X(_01499_));
 sg13g2_mux2_1 _24109_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][9] ),
    .A1(net647),
    .S(_06012_),
    .X(_01500_));
 sg13g2_nor3_1 _24110_ (.A(_05896_),
    .B(_05861_),
    .C(_05902_),
    .Y(_06014_));
 sg13g2_buf_1 _24111_ (.A(_06014_),
    .X(_06015_));
 sg13g2_buf_1 _24112_ (.A(_06015_),
    .X(_06016_));
 sg13g2_mux2_1 _24113_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][0] ),
    .A1(net473),
    .S(net322),
    .X(_01501_));
 sg13g2_mux2_1 _24114_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][10] ),
    .A1(net510),
    .S(net322),
    .X(_01502_));
 sg13g2_mux2_1 _24115_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][11] ),
    .A1(_05983_),
    .S(net322),
    .X(_01503_));
 sg13g2_mux2_1 _24116_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][1] ),
    .A1(_02966_),
    .S(_06016_),
    .X(_01504_));
 sg13g2_mux2_1 _24117_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][2] ),
    .A1(net889),
    .S(net322),
    .X(_01505_));
 sg13g2_mux2_1 _24118_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][3] ),
    .A1(net888),
    .S(net322),
    .X(_01506_));
 sg13g2_mux2_1 _24119_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][4] ),
    .A1(net887),
    .S(net322),
    .X(_01507_));
 sg13g2_mux2_1 _24120_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][5] ),
    .A1(net860),
    .S(net322),
    .X(_01508_));
 sg13g2_mux2_1 _24121_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][6] ),
    .A1(net982),
    .S(net322),
    .X(_01509_));
 sg13g2_mux2_1 _24122_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][7] ),
    .A1(_02976_),
    .S(_06016_),
    .X(_01510_));
 sg13g2_mux2_1 _24123_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][8] ),
    .A1(net582),
    .S(_06015_),
    .X(_01511_));
 sg13g2_mux2_1 _24124_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][9] ),
    .A1(_05979_),
    .S(_06015_),
    .X(_01512_));
 sg13g2_nor3_1 _24125_ (.A(_05829_),
    .B(_05861_),
    .C(_05886_),
    .Y(_06017_));
 sg13g2_buf_1 _24126_ (.A(_06017_),
    .X(_06018_));
 sg13g2_buf_1 _24127_ (.A(_06018_),
    .X(_06019_));
 sg13g2_mux2_1 _24128_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][0] ),
    .A1(net473),
    .S(net253),
    .X(_01513_));
 sg13g2_mux2_1 _24129_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][10] ),
    .A1(_09541_),
    .S(net253),
    .X(_01514_));
 sg13g2_mux2_1 _24130_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][11] ),
    .A1(_05983_),
    .S(net253),
    .X(_01515_));
 sg13g2_mux2_1 _24131_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][1] ),
    .A1(_02966_),
    .S(net253),
    .X(_01516_));
 sg13g2_mux2_1 _24132_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][2] ),
    .A1(_02951_),
    .S(_06019_),
    .X(_01517_));
 sg13g2_mux2_1 _24133_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][3] ),
    .A1(net888),
    .S(net253),
    .X(_01518_));
 sg13g2_mux2_1 _24134_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][4] ),
    .A1(_02956_),
    .S(net253),
    .X(_01519_));
 sg13g2_mux2_1 _24135_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][5] ),
    .A1(_05987_),
    .S(_06019_),
    .X(_01520_));
 sg13g2_mux2_1 _24136_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][6] ),
    .A1(_02960_),
    .S(net253),
    .X(_01521_));
 sg13g2_mux2_1 _24137_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][7] ),
    .A1(_02976_),
    .S(net253),
    .X(_01522_));
 sg13g2_mux2_1 _24138_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][8] ),
    .A1(_09682_),
    .S(_06018_),
    .X(_01523_));
 sg13g2_mux2_1 _24139_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][9] ),
    .A1(_09680_),
    .S(_06018_),
    .X(_01524_));
 sg13g2_and2_1 _24140_ (.A(_05845_),
    .B(_05847_),
    .X(_06020_));
 sg13g2_buf_1 _24141_ (.A(_06020_),
    .X(_06021_));
 sg13g2_and3_1 _24142_ (.X(_06022_),
    .A(net1052),
    .B(_10930_),
    .C(_05800_));
 sg13g2_buf_1 _24143_ (.A(_06022_),
    .X(_06023_));
 sg13g2_and2_1 _24144_ (.A(_05817_),
    .B(_06023_),
    .X(_06024_));
 sg13g2_buf_1 _24145_ (.A(_06024_),
    .X(_06025_));
 sg13g2_nand2_1 _24146_ (.Y(_06026_),
    .A(_06021_),
    .B(_06025_));
 sg13g2_buf_1 _24147_ (.A(_06026_),
    .X(_06027_));
 sg13g2_buf_1 _24148_ (.A(net321),
    .X(_06028_));
 sg13g2_nand2_1 _24149_ (.Y(_06029_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][0] ),
    .B(net321));
 sg13g2_o21ai_1 _24150_ (.B1(_06029_),
    .Y(_01525_),
    .A1(net592),
    .A2(net252));
 sg13g2_nand2_1 _24151_ (.Y(_06030_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][10] ),
    .B(net321));
 sg13g2_o21ai_1 _24152_ (.B1(_06030_),
    .Y(_01526_),
    .A1(net657),
    .A2(net252));
 sg13g2_nand2_1 _24153_ (.Y(_06031_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][11] ),
    .B(net321));
 sg13g2_o21ai_1 _24154_ (.B1(_06031_),
    .Y(_01527_),
    .A1(net593),
    .A2(net252));
 sg13g2_nand2_1 _24155_ (.Y(_06032_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][1] ),
    .B(net321));
 sg13g2_o21ai_1 _24156_ (.B1(_06032_),
    .Y(_01528_),
    .A1(net756),
    .A2(net252));
 sg13g2_mux2_1 _24157_ (.A0(net755),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][2] ),
    .S(net252),
    .X(_01529_));
 sg13g2_mux2_1 _24158_ (.A0(net754),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][3] ),
    .S(net252),
    .X(_01530_));
 sg13g2_mux2_1 _24159_ (.A0(net753),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][4] ),
    .S(net252),
    .X(_01531_));
 sg13g2_buf_1 _24160_ (.A(_05987_),
    .X(_06033_));
 sg13g2_mux2_1 _24161_ (.A0(_06033_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][5] ),
    .S(net321),
    .X(_01532_));
 sg13g2_mux2_1 _24162_ (.A0(net886),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][6] ),
    .S(_06027_),
    .X(_01533_));
 sg13g2_nand2_1 _24163_ (.Y(_06034_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][7] ),
    .B(net321));
 sg13g2_o21ai_1 _24164_ (.B1(_06034_),
    .Y(_01534_),
    .A1(net752),
    .A2(net252));
 sg13g2_nand2_1 _24165_ (.Y(_06035_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][8] ),
    .B(net321));
 sg13g2_o21ai_1 _24166_ (.B1(_06035_),
    .Y(_01535_),
    .A1(net742),
    .A2(_06028_));
 sg13g2_nand2_1 _24167_ (.Y(_06036_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][9] ),
    .B(_06027_));
 sg13g2_o21ai_1 _24168_ (.B1(_06036_),
    .Y(_01536_),
    .A1(net741),
    .A2(_06028_));
 sg13g2_buf_1 _24169_ (.A(_06023_),
    .X(_06037_));
 sg13g2_nand2_1 _24170_ (.Y(_06038_),
    .A(_05862_),
    .B(_06037_));
 sg13g2_buf_1 _24171_ (.A(_06038_),
    .X(_06039_));
 sg13g2_buf_1 _24172_ (.A(net379),
    .X(_06040_));
 sg13g2_nand2_1 _24173_ (.Y(_06041_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][0] ),
    .B(net379));
 sg13g2_o21ai_1 _24174_ (.B1(_06041_),
    .Y(_01537_),
    .A1(_03708_),
    .A2(net320));
 sg13g2_nand2_1 _24175_ (.Y(_06042_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][10] ),
    .B(net379));
 sg13g2_o21ai_1 _24176_ (.B1(_06042_),
    .Y(_01538_),
    .A1(net657),
    .A2(net320));
 sg13g2_nand2_1 _24177_ (.Y(_06043_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][11] ),
    .B(net379));
 sg13g2_o21ai_1 _24178_ (.B1(_06043_),
    .Y(_01539_),
    .A1(_03703_),
    .A2(net320));
 sg13g2_nand2_1 _24179_ (.Y(_06044_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][1] ),
    .B(net379));
 sg13g2_o21ai_1 _24180_ (.B1(_06044_),
    .Y(_01540_),
    .A1(net756),
    .A2(net320));
 sg13g2_mux2_1 _24181_ (.A0(net755),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][2] ),
    .S(net320),
    .X(_01541_));
 sg13g2_mux2_1 _24182_ (.A0(net754),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][3] ),
    .S(net320),
    .X(_01542_));
 sg13g2_mux2_1 _24183_ (.A0(net753),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][4] ),
    .S(net320),
    .X(_01543_));
 sg13g2_mux2_1 _24184_ (.A0(net734),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][5] ),
    .S(net379),
    .X(_01544_));
 sg13g2_mux2_1 _24185_ (.A0(net886),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][6] ),
    .S(net379),
    .X(_01545_));
 sg13g2_nand2_1 _24186_ (.Y(_06045_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][7] ),
    .B(net379));
 sg13g2_o21ai_1 _24187_ (.B1(_06045_),
    .Y(_01546_),
    .A1(net752),
    .A2(net320));
 sg13g2_nand2_1 _24188_ (.Y(_06046_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][8] ),
    .B(_06039_));
 sg13g2_o21ai_1 _24189_ (.B1(_06046_),
    .Y(_01547_),
    .A1(_03695_),
    .A2(_06040_));
 sg13g2_nand2_1 _24190_ (.Y(_06047_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][9] ),
    .B(_06039_));
 sg13g2_o21ai_1 _24191_ (.B1(_06047_),
    .Y(_01548_),
    .A1(_03698_),
    .A2(_06040_));
 sg13g2_nand2_1 _24192_ (.Y(_06048_),
    .A(_05871_),
    .B(net463));
 sg13g2_buf_1 _24193_ (.A(_06048_),
    .X(_06049_));
 sg13g2_buf_1 _24194_ (.A(net378),
    .X(_06050_));
 sg13g2_nand2_1 _24195_ (.Y(_06051_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][0] ),
    .B(net378));
 sg13g2_o21ai_1 _24196_ (.B1(_06051_),
    .Y(_01549_),
    .A1(_03708_),
    .A2(_06050_));
 sg13g2_nand2_1 _24197_ (.Y(_06052_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][10] ),
    .B(net378));
 sg13g2_o21ai_1 _24198_ (.B1(_06052_),
    .Y(_01550_),
    .A1(net657),
    .A2(net319));
 sg13g2_nand2_1 _24199_ (.Y(_06053_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][11] ),
    .B(net378));
 sg13g2_o21ai_1 _24200_ (.B1(_06053_),
    .Y(_01551_),
    .A1(_03703_),
    .A2(net319));
 sg13g2_nand2_1 _24201_ (.Y(_06054_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][1] ),
    .B(net378));
 sg13g2_o21ai_1 _24202_ (.B1(_06054_),
    .Y(_01552_),
    .A1(net756),
    .A2(_06050_));
 sg13g2_mux2_1 _24203_ (.A0(_02952_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][2] ),
    .S(net319),
    .X(_01553_));
 sg13g2_mux2_1 _24204_ (.A0(net754),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][3] ),
    .S(net319),
    .X(_01554_));
 sg13g2_mux2_1 _24205_ (.A0(net753),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][4] ),
    .S(net319),
    .X(_01555_));
 sg13g2_mux2_1 _24206_ (.A0(net734),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][5] ),
    .S(net378),
    .X(_01556_));
 sg13g2_mux2_1 _24207_ (.A0(net886),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][6] ),
    .S(net378),
    .X(_01557_));
 sg13g2_nand2_1 _24208_ (.Y(_06055_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][7] ),
    .B(net378));
 sg13g2_o21ai_1 _24209_ (.B1(_06055_),
    .Y(_01558_),
    .A1(net752),
    .A2(net319));
 sg13g2_nand2_1 _24210_ (.Y(_06056_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][8] ),
    .B(_06049_));
 sg13g2_o21ai_1 _24211_ (.B1(_06056_),
    .Y(_01559_),
    .A1(_03695_),
    .A2(net319));
 sg13g2_nand2_1 _24212_ (.Y(_06057_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][9] ),
    .B(_06049_));
 sg13g2_o21ai_1 _24213_ (.B1(_06057_),
    .Y(_01560_),
    .A1(_03698_),
    .A2(net319));
 sg13g2_nor2_1 _24214_ (.A(_05845_),
    .B(_05861_),
    .Y(_06058_));
 sg13g2_nand2_1 _24215_ (.Y(_06059_),
    .A(_06058_),
    .B(_06025_));
 sg13g2_buf_1 _24216_ (.A(_06059_),
    .X(_06060_));
 sg13g2_buf_1 _24217_ (.A(net318),
    .X(_06061_));
 sg13g2_nand2_1 _24218_ (.Y(_06062_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][0] ),
    .B(net318));
 sg13g2_o21ai_1 _24219_ (.B1(_06062_),
    .Y(_01561_),
    .A1(net592),
    .A2(net251));
 sg13g2_nand2_1 _24220_ (.Y(_06063_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][10] ),
    .B(net318));
 sg13g2_o21ai_1 _24221_ (.B1(_06063_),
    .Y(_01562_),
    .A1(net657),
    .A2(_06061_));
 sg13g2_nand2_1 _24222_ (.Y(_06064_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][11] ),
    .B(net318));
 sg13g2_o21ai_1 _24223_ (.B1(_06064_),
    .Y(_01563_),
    .A1(net593),
    .A2(net251));
 sg13g2_nand2_1 _24224_ (.Y(_06065_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][1] ),
    .B(net318));
 sg13g2_o21ai_1 _24225_ (.B1(_06065_),
    .Y(_01564_),
    .A1(net756),
    .A2(net251));
 sg13g2_mux2_1 _24226_ (.A0(net755),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][2] ),
    .S(net251),
    .X(_01565_));
 sg13g2_mux2_1 _24227_ (.A0(net754),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][3] ),
    .S(net251),
    .X(_01566_));
 sg13g2_mux2_1 _24228_ (.A0(net753),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][4] ),
    .S(net251),
    .X(_01567_));
 sg13g2_mux2_1 _24229_ (.A0(net734),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][5] ),
    .S(net318),
    .X(_01568_));
 sg13g2_mux2_1 _24230_ (.A0(net886),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][6] ),
    .S(_06060_),
    .X(_01569_));
 sg13g2_nand2_1 _24231_ (.Y(_06066_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][7] ),
    .B(net318));
 sg13g2_o21ai_1 _24232_ (.B1(_06066_),
    .Y(_01570_),
    .A1(net752),
    .A2(net251));
 sg13g2_nand2_1 _24233_ (.Y(_06067_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][8] ),
    .B(_06060_));
 sg13g2_o21ai_1 _24234_ (.B1(_06067_),
    .Y(_01571_),
    .A1(net742),
    .A2(_06061_));
 sg13g2_nand2_1 _24235_ (.Y(_06068_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][9] ),
    .B(net318));
 sg13g2_o21ai_1 _24236_ (.B1(_06068_),
    .Y(_01572_),
    .A1(net741),
    .A2(net251));
 sg13g2_and2_1 _24237_ (.A(_05884_),
    .B(_06023_),
    .X(_06069_));
 sg13g2_buf_2 _24238_ (.A(_06069_),
    .X(_06070_));
 sg13g2_nand2_1 _24239_ (.Y(_06071_),
    .A(_06058_),
    .B(_06070_));
 sg13g2_buf_1 _24240_ (.A(_06071_),
    .X(_06072_));
 sg13g2_buf_1 _24241_ (.A(_06072_),
    .X(_06073_));
 sg13g2_nand2_1 _24242_ (.Y(_06074_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][0] ),
    .B(net317));
 sg13g2_o21ai_1 _24243_ (.B1(_06074_),
    .Y(_01573_),
    .A1(net592),
    .A2(net250));
 sg13g2_nand2_1 _24244_ (.Y(_06075_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][10] ),
    .B(net317));
 sg13g2_o21ai_1 _24245_ (.B1(_06075_),
    .Y(_01574_),
    .A1(net657),
    .A2(_06073_));
 sg13g2_nand2_1 _24246_ (.Y(_06076_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][11] ),
    .B(net317));
 sg13g2_o21ai_1 _24247_ (.B1(_06076_),
    .Y(_01575_),
    .A1(net593),
    .A2(net250));
 sg13g2_nand2_1 _24248_ (.Y(_06077_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][1] ),
    .B(net317));
 sg13g2_o21ai_1 _24249_ (.B1(_06077_),
    .Y(_01576_),
    .A1(net756),
    .A2(net250));
 sg13g2_mux2_1 _24250_ (.A0(net755),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][2] ),
    .S(net250),
    .X(_01577_));
 sg13g2_mux2_1 _24251_ (.A0(net754),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][3] ),
    .S(net250),
    .X(_01578_));
 sg13g2_mux2_1 _24252_ (.A0(net753),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][4] ),
    .S(net250),
    .X(_01579_));
 sg13g2_mux2_1 _24253_ (.A0(net734),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][5] ),
    .S(net317),
    .X(_01580_));
 sg13g2_mux2_1 _24254_ (.A0(net886),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][6] ),
    .S(net317),
    .X(_01581_));
 sg13g2_nand2_1 _24255_ (.Y(_06078_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][7] ),
    .B(net317));
 sg13g2_o21ai_1 _24256_ (.B1(_06078_),
    .Y(_01582_),
    .A1(net752),
    .A2(net250));
 sg13g2_nand2_1 _24257_ (.Y(_06079_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][8] ),
    .B(_06072_));
 sg13g2_o21ai_1 _24258_ (.B1(_06079_),
    .Y(_01583_),
    .A1(net742),
    .A2(_06073_));
 sg13g2_nand2_1 _24259_ (.Y(_06080_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][9] ),
    .B(net317));
 sg13g2_o21ai_1 _24260_ (.B1(_06080_),
    .Y(_01584_),
    .A1(net741),
    .A2(net250));
 sg13g2_nand3_1 _24261_ (.B(_06058_),
    .C(net463),
    .A(_05858_),
    .Y(_06081_));
 sg13g2_buf_1 _24262_ (.A(_06081_),
    .X(_06082_));
 sg13g2_buf_1 _24263_ (.A(_06082_),
    .X(_06083_));
 sg13g2_nand2_1 _24264_ (.Y(_06084_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][0] ),
    .B(net377));
 sg13g2_o21ai_1 _24265_ (.B1(_06084_),
    .Y(_01585_),
    .A1(net592),
    .A2(net316));
 sg13g2_nand2_1 _24266_ (.Y(_06085_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][10] ),
    .B(net377));
 sg13g2_o21ai_1 _24267_ (.B1(_06085_),
    .Y(_01586_),
    .A1(net657),
    .A2(_06083_));
 sg13g2_nand2_1 _24268_ (.Y(_06086_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][11] ),
    .B(net377));
 sg13g2_o21ai_1 _24269_ (.B1(_06086_),
    .Y(_01587_),
    .A1(net593),
    .A2(net316));
 sg13g2_nand2_1 _24270_ (.Y(_06087_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][1] ),
    .B(net377));
 sg13g2_o21ai_1 _24271_ (.B1(_06087_),
    .Y(_01588_),
    .A1(net756),
    .A2(net316));
 sg13g2_mux2_1 _24272_ (.A0(net755),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][2] ),
    .S(net316),
    .X(_01589_));
 sg13g2_mux2_1 _24273_ (.A0(net754),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][3] ),
    .S(net316),
    .X(_01590_));
 sg13g2_mux2_1 _24274_ (.A0(net753),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][4] ),
    .S(net316),
    .X(_01591_));
 sg13g2_mux2_1 _24275_ (.A0(net734),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][5] ),
    .S(net377),
    .X(_01592_));
 sg13g2_mux2_1 _24276_ (.A0(net886),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][6] ),
    .S(net377),
    .X(_01593_));
 sg13g2_nand2_1 _24277_ (.Y(_06088_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][7] ),
    .B(net377));
 sg13g2_o21ai_1 _24278_ (.B1(_06088_),
    .Y(_01594_),
    .A1(net752),
    .A2(net316));
 sg13g2_nand2_1 _24279_ (.Y(_06089_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][8] ),
    .B(_06082_));
 sg13g2_o21ai_1 _24280_ (.B1(_06089_),
    .Y(_01595_),
    .A1(net742),
    .A2(_06083_));
 sg13g2_nand2_1 _24281_ (.Y(_06090_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][9] ),
    .B(net377));
 sg13g2_o21ai_1 _24282_ (.B1(_06090_),
    .Y(_01596_),
    .A1(net741),
    .A2(net316));
 sg13g2_buf_1 _24283_ (.A(_06023_),
    .X(_06091_));
 sg13g2_nand3_1 _24284_ (.B(_06058_),
    .C(net462),
    .A(_05814_),
    .Y(_06092_));
 sg13g2_buf_1 _24285_ (.A(_06092_),
    .X(_06093_));
 sg13g2_buf_1 _24286_ (.A(net376),
    .X(_06094_));
 sg13g2_nand2_1 _24287_ (.Y(_06095_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][0] ),
    .B(net376));
 sg13g2_o21ai_1 _24288_ (.B1(_06095_),
    .Y(_01597_),
    .A1(net592),
    .A2(net315));
 sg13g2_nand2_1 _24289_ (.Y(_06096_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][10] ),
    .B(net376));
 sg13g2_o21ai_1 _24290_ (.B1(_06096_),
    .Y(_01598_),
    .A1(net657),
    .A2(net315));
 sg13g2_nand2_1 _24291_ (.Y(_06097_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][11] ),
    .B(net376));
 sg13g2_o21ai_1 _24292_ (.B1(_06097_),
    .Y(_01599_),
    .A1(net593),
    .A2(net315));
 sg13g2_buf_1 _24293_ (.A(net890),
    .X(_06098_));
 sg13g2_nand2_1 _24294_ (.Y(_06099_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][1] ),
    .B(net376));
 sg13g2_o21ai_1 _24295_ (.B1(_06099_),
    .Y(_01600_),
    .A1(_06098_),
    .A2(net315));
 sg13g2_buf_1 _24296_ (.A(net889),
    .X(_06100_));
 sg13g2_mux2_1 _24297_ (.A0(_06100_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][2] ),
    .S(net315),
    .X(_01601_));
 sg13g2_buf_1 _24298_ (.A(net888),
    .X(_06101_));
 sg13g2_mux2_1 _24299_ (.A0(_06101_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][3] ),
    .S(net315),
    .X(_01602_));
 sg13g2_buf_1 _24300_ (.A(net887),
    .X(_06102_));
 sg13g2_mux2_1 _24301_ (.A0(_06102_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][4] ),
    .S(net315),
    .X(_01603_));
 sg13g2_mux2_1 _24302_ (.A0(_06033_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][5] ),
    .S(net376),
    .X(_01604_));
 sg13g2_buf_1 _24303_ (.A(net982),
    .X(_06103_));
 sg13g2_mux2_1 _24304_ (.A0(_06103_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][6] ),
    .S(_06093_),
    .X(_01605_));
 sg13g2_buf_1 _24305_ (.A(net885),
    .X(_06104_));
 sg13g2_nand2_1 _24306_ (.Y(_06105_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][7] ),
    .B(net376));
 sg13g2_o21ai_1 _24307_ (.B1(_06105_),
    .Y(_01606_),
    .A1(_06104_),
    .A2(net315));
 sg13g2_nand2_1 _24308_ (.Y(_06106_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][8] ),
    .B(_06093_));
 sg13g2_o21ai_1 _24309_ (.B1(_06106_),
    .Y(_01607_),
    .A1(net742),
    .A2(_06094_));
 sg13g2_nand2_1 _24310_ (.Y(_06107_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][9] ),
    .B(net376));
 sg13g2_o21ai_1 _24311_ (.B1(_06107_),
    .Y(_01608_),
    .A1(net741),
    .A2(_06094_));
 sg13g2_nand2_1 _24312_ (.Y(_06108_),
    .A(_11224_),
    .B(_05822_));
 sg13g2_nor2_1 _24313_ (.A(net973),
    .B(_06108_),
    .Y(_06109_));
 sg13g2_nand4_1 _24314_ (.B(_05837_),
    .C(_06109_),
    .A(net970),
    .Y(_06110_),
    .D(_06091_));
 sg13g2_buf_1 _24315_ (.A(_06110_),
    .X(_06111_));
 sg13g2_buf_1 _24316_ (.A(net375),
    .X(_06112_));
 sg13g2_nand2_1 _24317_ (.Y(_06113_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][0] ),
    .B(net375));
 sg13g2_o21ai_1 _24318_ (.B1(_06113_),
    .Y(_01609_),
    .A1(net592),
    .A2(net314));
 sg13g2_nand2_1 _24319_ (.Y(_06114_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][10] ),
    .B(net375));
 sg13g2_o21ai_1 _24320_ (.B1(_06114_),
    .Y(_01610_),
    .A1(net657),
    .A2(net314));
 sg13g2_nand2_1 _24321_ (.Y(_06115_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][11] ),
    .B(net375));
 sg13g2_o21ai_1 _24322_ (.B1(_06115_),
    .Y(_01611_),
    .A1(net593),
    .A2(_06112_));
 sg13g2_nand2_1 _24323_ (.Y(_06116_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][1] ),
    .B(net375));
 sg13g2_o21ai_1 _24324_ (.B1(_06116_),
    .Y(_01612_),
    .A1(net733),
    .A2(net314));
 sg13g2_mux2_1 _24325_ (.A0(net732),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][2] ),
    .S(net314),
    .X(_01613_));
 sg13g2_mux2_1 _24326_ (.A0(net731),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][3] ),
    .S(net314),
    .X(_01614_));
 sg13g2_mux2_1 _24327_ (.A0(net730),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][4] ),
    .S(net314),
    .X(_01615_));
 sg13g2_mux2_1 _24328_ (.A0(net734),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][5] ),
    .S(net375),
    .X(_01616_));
 sg13g2_mux2_1 _24329_ (.A0(net859),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][6] ),
    .S(net375),
    .X(_01617_));
 sg13g2_nand2_1 _24330_ (.Y(_06117_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][7] ),
    .B(net375));
 sg13g2_o21ai_1 _24331_ (.B1(_06117_),
    .Y(_01618_),
    .A1(net729),
    .A2(net314));
 sg13g2_nand2_1 _24332_ (.Y(_06118_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][8] ),
    .B(_06111_));
 sg13g2_o21ai_1 _24333_ (.B1(_06118_),
    .Y(_01619_),
    .A1(net742),
    .A2(_06112_));
 sg13g2_nand2_1 _24334_ (.Y(_06119_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][9] ),
    .B(_06111_));
 sg13g2_o21ai_1 _24335_ (.B1(_06119_),
    .Y(_01620_),
    .A1(net741),
    .A2(net314));
 sg13g2_buf_1 _24336_ (.A(net656),
    .X(_06120_));
 sg13g2_nand4_1 _24337_ (.B(net870),
    .C(_05837_),
    .A(net970),
    .Y(_06121_),
    .D(_06070_));
 sg13g2_buf_1 _24338_ (.A(_06121_),
    .X(_06122_));
 sg13g2_buf_1 _24339_ (.A(net313),
    .X(_06123_));
 sg13g2_nand2_1 _24340_ (.Y(_06124_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][0] ),
    .B(net313));
 sg13g2_o21ai_1 _24341_ (.B1(_06124_),
    .Y(_01621_),
    .A1(net581),
    .A2(net249));
 sg13g2_buf_1 _24342_ (.A(net740),
    .X(_06125_));
 sg13g2_nand2_1 _24343_ (.Y(_06126_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][10] ),
    .B(net313));
 sg13g2_o21ai_1 _24344_ (.B1(_06126_),
    .Y(_01622_),
    .A1(net646),
    .A2(net249));
 sg13g2_buf_1 _24345_ (.A(net670),
    .X(_06127_));
 sg13g2_nand2_1 _24346_ (.Y(_06128_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][11] ),
    .B(net313));
 sg13g2_o21ai_1 _24347_ (.B1(_06128_),
    .Y(_01623_),
    .A1(net580),
    .A2(_06123_));
 sg13g2_nand2_1 _24348_ (.Y(_06129_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][1] ),
    .B(_06122_));
 sg13g2_o21ai_1 _24349_ (.B1(_06129_),
    .Y(_01624_),
    .A1(net733),
    .A2(net249));
 sg13g2_mux2_1 _24350_ (.A0(net732),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][2] ),
    .S(net249),
    .X(_01625_));
 sg13g2_mux2_1 _24351_ (.A0(net731),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][3] ),
    .S(net249),
    .X(_01626_));
 sg13g2_mux2_1 _24352_ (.A0(net730),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][4] ),
    .S(net249),
    .X(_01627_));
 sg13g2_mux2_1 _24353_ (.A0(net734),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][5] ),
    .S(net313),
    .X(_01628_));
 sg13g2_mux2_1 _24354_ (.A0(net859),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][6] ),
    .S(net313),
    .X(_01629_));
 sg13g2_nand2_1 _24355_ (.Y(_06130_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][7] ),
    .B(net313));
 sg13g2_o21ai_1 _24356_ (.B1(_06130_),
    .Y(_01630_),
    .A1(net729),
    .A2(net249));
 sg13g2_buf_1 _24357_ (.A(net876),
    .X(_06131_));
 sg13g2_nand2_1 _24358_ (.Y(_06132_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][8] ),
    .B(net313));
 sg13g2_o21ai_1 _24359_ (.B1(_06132_),
    .Y(_01631_),
    .A1(net728),
    .A2(net249));
 sg13g2_buf_1 _24360_ (.A(net875),
    .X(_06133_));
 sg13g2_nand2_1 _24361_ (.Y(_06134_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][9] ),
    .B(_06122_));
 sg13g2_o21ai_1 _24362_ (.B1(_06134_),
    .Y(_01632_),
    .A1(net727),
    .A2(_06123_));
 sg13g2_nand2_1 _24363_ (.Y(_06135_),
    .A(_05910_),
    .B(net463));
 sg13g2_buf_1 _24364_ (.A(_06135_),
    .X(_06136_));
 sg13g2_buf_1 _24365_ (.A(net374),
    .X(_06137_));
 sg13g2_nand2_1 _24366_ (.Y(_06138_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][0] ),
    .B(net374));
 sg13g2_o21ai_1 _24367_ (.B1(_06138_),
    .Y(_01633_),
    .A1(net581),
    .A2(net312));
 sg13g2_nand2_1 _24368_ (.Y(_06139_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][10] ),
    .B(net374));
 sg13g2_o21ai_1 _24369_ (.B1(_06139_),
    .Y(_01634_),
    .A1(net646),
    .A2(net312));
 sg13g2_nand2_1 _24370_ (.Y(_06140_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][11] ),
    .B(net374));
 sg13g2_o21ai_1 _24371_ (.B1(_06140_),
    .Y(_01635_),
    .A1(net580),
    .A2(_06137_));
 sg13g2_nand2_1 _24372_ (.Y(_06141_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][1] ),
    .B(_06136_));
 sg13g2_o21ai_1 _24373_ (.B1(_06141_),
    .Y(_01636_),
    .A1(net733),
    .A2(net312));
 sg13g2_mux2_1 _24374_ (.A0(net732),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][2] ),
    .S(net312),
    .X(_01637_));
 sg13g2_mux2_1 _24375_ (.A0(net731),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][3] ),
    .S(net312),
    .X(_01638_));
 sg13g2_mux2_1 _24376_ (.A0(net730),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][4] ),
    .S(net312),
    .X(_01639_));
 sg13g2_mux2_1 _24377_ (.A0(net734),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][5] ),
    .S(net374),
    .X(_01640_));
 sg13g2_mux2_1 _24378_ (.A0(net859),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][6] ),
    .S(net374),
    .X(_01641_));
 sg13g2_nand2_1 _24379_ (.Y(_06142_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][7] ),
    .B(net374));
 sg13g2_o21ai_1 _24380_ (.B1(_06142_),
    .Y(_01642_),
    .A1(net729),
    .A2(net312));
 sg13g2_nand2_1 _24381_ (.Y(_06143_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][8] ),
    .B(net374));
 sg13g2_o21ai_1 _24382_ (.B1(_06143_),
    .Y(_01643_),
    .A1(net728),
    .A2(net312));
 sg13g2_nand2_1 _24383_ (.Y(_06144_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][9] ),
    .B(_06136_));
 sg13g2_o21ai_1 _24384_ (.B1(_06144_),
    .Y(_01644_),
    .A1(net727),
    .A2(_06137_));
 sg13g2_nand2_1 _24385_ (.Y(_06145_),
    .A(_05918_),
    .B(net463));
 sg13g2_buf_1 _24386_ (.A(_06145_),
    .X(_06146_));
 sg13g2_buf_1 _24387_ (.A(net373),
    .X(_06147_));
 sg13g2_nand2_1 _24388_ (.Y(_06148_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][0] ),
    .B(net373));
 sg13g2_o21ai_1 _24389_ (.B1(_06148_),
    .Y(_01645_),
    .A1(net581),
    .A2(net311));
 sg13g2_nand2_1 _24390_ (.Y(_06149_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][10] ),
    .B(net373));
 sg13g2_o21ai_1 _24391_ (.B1(_06149_),
    .Y(_01646_),
    .A1(net646),
    .A2(net311));
 sg13g2_nand2_1 _24392_ (.Y(_06150_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][11] ),
    .B(net373));
 sg13g2_o21ai_1 _24393_ (.B1(_06150_),
    .Y(_01647_),
    .A1(net580),
    .A2(_06147_));
 sg13g2_nand2_1 _24394_ (.Y(_06151_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][1] ),
    .B(_06146_));
 sg13g2_o21ai_1 _24395_ (.B1(_06151_),
    .Y(_01648_),
    .A1(net733),
    .A2(net311));
 sg13g2_mux2_1 _24396_ (.A0(net732),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][2] ),
    .S(net311),
    .X(_01649_));
 sg13g2_mux2_1 _24397_ (.A0(net731),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][3] ),
    .S(net311),
    .X(_01650_));
 sg13g2_mux2_1 _24398_ (.A0(net730),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][4] ),
    .S(net311),
    .X(_01651_));
 sg13g2_buf_1 _24399_ (.A(_02973_),
    .X(_06152_));
 sg13g2_mux2_1 _24400_ (.A0(_06152_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][5] ),
    .S(net373),
    .X(_01652_));
 sg13g2_mux2_1 _24401_ (.A0(net859),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][6] ),
    .S(net373),
    .X(_01653_));
 sg13g2_nand2_1 _24402_ (.Y(_06153_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][7] ),
    .B(net373));
 sg13g2_o21ai_1 _24403_ (.B1(_06153_),
    .Y(_01654_),
    .A1(net729),
    .A2(net311));
 sg13g2_nand2_1 _24404_ (.Y(_06154_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][8] ),
    .B(net373));
 sg13g2_o21ai_1 _24405_ (.B1(_06154_),
    .Y(_01655_),
    .A1(net728),
    .A2(net311));
 sg13g2_nand2_1 _24406_ (.Y(_06155_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][9] ),
    .B(_06146_));
 sg13g2_o21ai_1 _24407_ (.B1(_06155_),
    .Y(_01656_),
    .A1(net727),
    .A2(_06147_));
 sg13g2_nand2_1 _24408_ (.Y(_06156_),
    .A(_06021_),
    .B(_06070_));
 sg13g2_buf_1 _24409_ (.A(_06156_),
    .X(_06157_));
 sg13g2_buf_1 _24410_ (.A(_06157_),
    .X(_06158_));
 sg13g2_nand2_1 _24411_ (.Y(_06159_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][0] ),
    .B(net310));
 sg13g2_o21ai_1 _24412_ (.B1(_06159_),
    .Y(_01657_),
    .A1(net581),
    .A2(net248));
 sg13g2_nand2_1 _24413_ (.Y(_06160_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][10] ),
    .B(net310));
 sg13g2_o21ai_1 _24414_ (.B1(_06160_),
    .Y(_01658_),
    .A1(_06125_),
    .A2(_06158_));
 sg13g2_nand2_1 _24415_ (.Y(_06161_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][11] ),
    .B(net310));
 sg13g2_o21ai_1 _24416_ (.B1(_06161_),
    .Y(_01659_),
    .A1(net580),
    .A2(net248));
 sg13g2_nand2_1 _24417_ (.Y(_06162_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][1] ),
    .B(net310));
 sg13g2_o21ai_1 _24418_ (.B1(_06162_),
    .Y(_01660_),
    .A1(_06098_),
    .A2(net248));
 sg13g2_mux2_1 _24419_ (.A0(_06100_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][2] ),
    .S(net248),
    .X(_01661_));
 sg13g2_mux2_1 _24420_ (.A0(_06101_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][3] ),
    .S(net248),
    .X(_01662_));
 sg13g2_mux2_1 _24421_ (.A0(_06102_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][4] ),
    .S(net248),
    .X(_01663_));
 sg13g2_mux2_1 _24422_ (.A0(_06152_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][5] ),
    .S(net310),
    .X(_01664_));
 sg13g2_mux2_1 _24423_ (.A0(_06103_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][6] ),
    .S(_06157_),
    .X(_01665_));
 sg13g2_nand2_1 _24424_ (.Y(_06163_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][7] ),
    .B(net310));
 sg13g2_o21ai_1 _24425_ (.B1(_06163_),
    .Y(_01666_),
    .A1(_06104_),
    .A2(net248));
 sg13g2_nand2_1 _24426_ (.Y(_06164_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][8] ),
    .B(net310));
 sg13g2_o21ai_1 _24427_ (.B1(_06164_),
    .Y(_01667_),
    .A1(net728),
    .A2(_06158_));
 sg13g2_nand2_1 _24428_ (.Y(_06165_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][9] ),
    .B(net310));
 sg13g2_o21ai_1 _24429_ (.B1(_06165_),
    .Y(_01668_),
    .A1(_06133_),
    .A2(net248));
 sg13g2_nor2_1 _24430_ (.A(_05845_),
    .B(_05901_),
    .Y(_06166_));
 sg13g2_nand2_1 _24431_ (.Y(_06167_),
    .A(_06166_),
    .B(_06025_));
 sg13g2_buf_1 _24432_ (.A(_06167_),
    .X(_06168_));
 sg13g2_buf_1 _24433_ (.A(net309),
    .X(_06169_));
 sg13g2_nand2_1 _24434_ (.Y(_06170_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][0] ),
    .B(net309));
 sg13g2_o21ai_1 _24435_ (.B1(_06170_),
    .Y(_01669_),
    .A1(net581),
    .A2(net247));
 sg13g2_nand2_1 _24436_ (.Y(_06171_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][10] ),
    .B(net309));
 sg13g2_o21ai_1 _24437_ (.B1(_06171_),
    .Y(_01670_),
    .A1(net646),
    .A2(net247));
 sg13g2_nand2_1 _24438_ (.Y(_06172_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][11] ),
    .B(net309));
 sg13g2_o21ai_1 _24439_ (.B1(_06172_),
    .Y(_01671_),
    .A1(net580),
    .A2(_06169_));
 sg13g2_nand2_1 _24440_ (.Y(_06173_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][1] ),
    .B(net309));
 sg13g2_o21ai_1 _24441_ (.B1(_06173_),
    .Y(_01672_),
    .A1(net733),
    .A2(net247));
 sg13g2_mux2_1 _24442_ (.A0(net732),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][2] ),
    .S(net247),
    .X(_01673_));
 sg13g2_mux2_1 _24443_ (.A0(net731),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][3] ),
    .S(net247),
    .X(_01674_));
 sg13g2_mux2_1 _24444_ (.A0(net730),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][4] ),
    .S(net247),
    .X(_01675_));
 sg13g2_mux2_1 _24445_ (.A0(net858),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][5] ),
    .S(_06168_),
    .X(_01676_));
 sg13g2_mux2_1 _24446_ (.A0(net859),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][6] ),
    .S(_06168_),
    .X(_01677_));
 sg13g2_nand2_1 _24447_ (.Y(_06174_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][7] ),
    .B(net309));
 sg13g2_o21ai_1 _24448_ (.B1(_06174_),
    .Y(_01678_),
    .A1(net729),
    .A2(net247));
 sg13g2_nand2_1 _24449_ (.Y(_06175_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][8] ),
    .B(net309));
 sg13g2_o21ai_1 _24450_ (.B1(_06175_),
    .Y(_01679_),
    .A1(net728),
    .A2(net247));
 sg13g2_nand2_1 _24451_ (.Y(_06176_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][9] ),
    .B(net309));
 sg13g2_o21ai_1 _24452_ (.B1(_06176_),
    .Y(_01680_),
    .A1(net727),
    .A2(_06169_));
 sg13g2_nand2_1 _24453_ (.Y(_06177_),
    .A(_06166_),
    .B(_06070_));
 sg13g2_buf_1 _24454_ (.A(_06177_),
    .X(_06178_));
 sg13g2_buf_1 _24455_ (.A(net308),
    .X(_06179_));
 sg13g2_nand2_1 _24456_ (.Y(_06180_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][0] ),
    .B(net308));
 sg13g2_o21ai_1 _24457_ (.B1(_06180_),
    .Y(_01681_),
    .A1(net581),
    .A2(net246));
 sg13g2_nand2_1 _24458_ (.Y(_06181_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][10] ),
    .B(net308));
 sg13g2_o21ai_1 _24459_ (.B1(_06181_),
    .Y(_01682_),
    .A1(net646),
    .A2(net246));
 sg13g2_nand2_1 _24460_ (.Y(_06182_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][11] ),
    .B(net308));
 sg13g2_o21ai_1 _24461_ (.B1(_06182_),
    .Y(_01683_),
    .A1(net580),
    .A2(_06179_));
 sg13g2_nand2_1 _24462_ (.Y(_06183_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][1] ),
    .B(net308));
 sg13g2_o21ai_1 _24463_ (.B1(_06183_),
    .Y(_01684_),
    .A1(net733),
    .A2(net246));
 sg13g2_mux2_1 _24464_ (.A0(net732),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][2] ),
    .S(net246),
    .X(_01685_));
 sg13g2_mux2_1 _24465_ (.A0(net731),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][3] ),
    .S(net246),
    .X(_01686_));
 sg13g2_mux2_1 _24466_ (.A0(net730),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][4] ),
    .S(net246),
    .X(_01687_));
 sg13g2_mux2_1 _24467_ (.A0(net858),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][5] ),
    .S(_06178_),
    .X(_01688_));
 sg13g2_mux2_1 _24468_ (.A0(net859),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][6] ),
    .S(_06178_),
    .X(_01689_));
 sg13g2_nand2_1 _24469_ (.Y(_06184_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][7] ),
    .B(net308));
 sg13g2_o21ai_1 _24470_ (.B1(_06184_),
    .Y(_01690_),
    .A1(net729),
    .A2(net246));
 sg13g2_nand2_1 _24471_ (.Y(_06185_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][8] ),
    .B(net308));
 sg13g2_o21ai_1 _24472_ (.B1(_06185_),
    .Y(_01691_),
    .A1(net728),
    .A2(net246));
 sg13g2_nand2_1 _24473_ (.Y(_06186_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][9] ),
    .B(net308));
 sg13g2_o21ai_1 _24474_ (.B1(_06186_),
    .Y(_01692_),
    .A1(net727),
    .A2(_06179_));
 sg13g2_nand3_1 _24475_ (.B(_06166_),
    .C(net462),
    .A(_05858_),
    .Y(_06187_));
 sg13g2_buf_1 _24476_ (.A(_06187_),
    .X(_06188_));
 sg13g2_buf_1 _24477_ (.A(net372),
    .X(_06189_));
 sg13g2_nand2_1 _24478_ (.Y(_06190_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][0] ),
    .B(net372));
 sg13g2_o21ai_1 _24479_ (.B1(_06190_),
    .Y(_01693_),
    .A1(_06120_),
    .A2(net307));
 sg13g2_nand2_1 _24480_ (.Y(_06191_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][10] ),
    .B(net372));
 sg13g2_o21ai_1 _24481_ (.B1(_06191_),
    .Y(_01694_),
    .A1(_06125_),
    .A2(net307));
 sg13g2_nand2_1 _24482_ (.Y(_06192_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][11] ),
    .B(net372));
 sg13g2_o21ai_1 _24483_ (.B1(_06192_),
    .Y(_01695_),
    .A1(_06127_),
    .A2(_06189_));
 sg13g2_nand2_1 _24484_ (.Y(_06193_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][1] ),
    .B(net372));
 sg13g2_o21ai_1 _24485_ (.B1(_06193_),
    .Y(_01696_),
    .A1(net733),
    .A2(net307));
 sg13g2_mux2_1 _24486_ (.A0(net732),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][2] ),
    .S(net307),
    .X(_01697_));
 sg13g2_mux2_1 _24487_ (.A0(net731),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][3] ),
    .S(net307),
    .X(_01698_));
 sg13g2_mux2_1 _24488_ (.A0(net730),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][4] ),
    .S(net307),
    .X(_01699_));
 sg13g2_mux2_1 _24489_ (.A0(net858),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][5] ),
    .S(_06188_),
    .X(_01700_));
 sg13g2_mux2_1 _24490_ (.A0(net859),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][6] ),
    .S(_06188_),
    .X(_01701_));
 sg13g2_nand2_1 _24491_ (.Y(_06194_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][7] ),
    .B(net372));
 sg13g2_o21ai_1 _24492_ (.B1(_06194_),
    .Y(_01702_),
    .A1(net729),
    .A2(net307));
 sg13g2_nand2_1 _24493_ (.Y(_06195_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][8] ),
    .B(net372));
 sg13g2_o21ai_1 _24494_ (.B1(_06195_),
    .Y(_01703_),
    .A1(_06131_),
    .A2(net307));
 sg13g2_nand2_1 _24495_ (.Y(_06196_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][9] ),
    .B(net372));
 sg13g2_o21ai_1 _24496_ (.B1(_06196_),
    .Y(_01704_),
    .A1(net727),
    .A2(_06189_));
 sg13g2_nand3_1 _24497_ (.B(_06166_),
    .C(net462),
    .A(_05814_),
    .Y(_06197_));
 sg13g2_buf_1 _24498_ (.A(_06197_),
    .X(_06198_));
 sg13g2_buf_1 _24499_ (.A(net371),
    .X(_06199_));
 sg13g2_nand2_1 _24500_ (.Y(_06200_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][0] ),
    .B(net371));
 sg13g2_o21ai_1 _24501_ (.B1(_06200_),
    .Y(_01705_),
    .A1(_06120_),
    .A2(net306));
 sg13g2_nand2_1 _24502_ (.Y(_06201_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][10] ),
    .B(net371));
 sg13g2_o21ai_1 _24503_ (.B1(_06201_),
    .Y(_01706_),
    .A1(net646),
    .A2(net306));
 sg13g2_nand2_1 _24504_ (.Y(_06202_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][11] ),
    .B(net371));
 sg13g2_o21ai_1 _24505_ (.B1(_06202_),
    .Y(_01707_),
    .A1(_06127_),
    .A2(_06199_));
 sg13g2_nand2_1 _24506_ (.Y(_06203_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][1] ),
    .B(net371));
 sg13g2_o21ai_1 _24507_ (.B1(_06203_),
    .Y(_01708_),
    .A1(net733),
    .A2(net306));
 sg13g2_mux2_1 _24508_ (.A0(net732),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][2] ),
    .S(net306),
    .X(_01709_));
 sg13g2_mux2_1 _24509_ (.A0(net731),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][3] ),
    .S(net306),
    .X(_01710_));
 sg13g2_mux2_1 _24510_ (.A0(net730),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][4] ),
    .S(net306),
    .X(_01711_));
 sg13g2_mux2_1 _24511_ (.A0(net858),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][5] ),
    .S(_06198_),
    .X(_01712_));
 sg13g2_mux2_1 _24512_ (.A0(net859),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][6] ),
    .S(_06198_),
    .X(_01713_));
 sg13g2_nand2_1 _24513_ (.Y(_06204_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][7] ),
    .B(net371));
 sg13g2_o21ai_1 _24514_ (.B1(_06204_),
    .Y(_01714_),
    .A1(net729),
    .A2(net306));
 sg13g2_nand2_1 _24515_ (.Y(_06205_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][8] ),
    .B(net371));
 sg13g2_o21ai_1 _24516_ (.B1(_06205_),
    .Y(_01715_),
    .A1(_06131_),
    .A2(net306));
 sg13g2_nand2_1 _24517_ (.Y(_06206_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][9] ),
    .B(net371));
 sg13g2_o21ai_1 _24518_ (.B1(_06206_),
    .Y(_01716_),
    .A1(_06133_),
    .A2(_06199_));
 sg13g2_inv_1 _24519_ (.Y(_06207_),
    .A(_05948_));
 sg13g2_nand3_1 _24520_ (.B(_06207_),
    .C(_06091_),
    .A(_06109_),
    .Y(_06208_));
 sg13g2_buf_1 _24521_ (.A(_06208_),
    .X(_06209_));
 sg13g2_buf_1 _24522_ (.A(net370),
    .X(_06210_));
 sg13g2_nand2_1 _24523_ (.Y(_06211_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][0] ),
    .B(net370));
 sg13g2_o21ai_1 _24524_ (.B1(_06211_),
    .Y(_01717_),
    .A1(net581),
    .A2(net305));
 sg13g2_nand2_1 _24525_ (.Y(_06212_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][10] ),
    .B(net370));
 sg13g2_o21ai_1 _24526_ (.B1(_06212_),
    .Y(_01718_),
    .A1(net646),
    .A2(_06210_));
 sg13g2_nand2_1 _24527_ (.Y(_06213_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][11] ),
    .B(net370));
 sg13g2_o21ai_1 _24528_ (.B1(_06213_),
    .Y(_01719_),
    .A1(net580),
    .A2(_06210_));
 sg13g2_buf_1 _24529_ (.A(net890),
    .X(_06214_));
 sg13g2_nand2_1 _24530_ (.Y(_06215_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][1] ),
    .B(net370));
 sg13g2_o21ai_1 _24531_ (.B1(_06215_),
    .Y(_01720_),
    .A1(net726),
    .A2(net305));
 sg13g2_buf_1 _24532_ (.A(net889),
    .X(_06216_));
 sg13g2_mux2_1 _24533_ (.A0(net725),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][2] ),
    .S(net305),
    .X(_01721_));
 sg13g2_buf_1 _24534_ (.A(net888),
    .X(_06217_));
 sg13g2_mux2_1 _24535_ (.A0(net724),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][3] ),
    .S(net305),
    .X(_01722_));
 sg13g2_buf_1 _24536_ (.A(net887),
    .X(_06218_));
 sg13g2_mux2_1 _24537_ (.A0(net723),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][4] ),
    .S(net305),
    .X(_01723_));
 sg13g2_mux2_1 _24538_ (.A0(net858),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][5] ),
    .S(_06209_),
    .X(_01724_));
 sg13g2_buf_1 _24539_ (.A(net982),
    .X(_06219_));
 sg13g2_mux2_1 _24540_ (.A0(net857),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][6] ),
    .S(_06209_),
    .X(_01725_));
 sg13g2_buf_1 _24541_ (.A(net885),
    .X(_06220_));
 sg13g2_nand2_1 _24542_ (.Y(_06221_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][7] ),
    .B(net370));
 sg13g2_o21ai_1 _24543_ (.B1(_06221_),
    .Y(_01726_),
    .A1(net722),
    .A2(net305));
 sg13g2_nand2_1 _24544_ (.Y(_06222_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][8] ),
    .B(net370));
 sg13g2_o21ai_1 _24545_ (.B1(_06222_),
    .Y(_01727_),
    .A1(net728),
    .A2(net305));
 sg13g2_nand2_1 _24546_ (.Y(_06223_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][9] ),
    .B(net370));
 sg13g2_o21ai_1 _24547_ (.B1(_06223_),
    .Y(_01728_),
    .A1(net727),
    .A2(net305));
 sg13g2_nand3_1 _24548_ (.B(_06207_),
    .C(_06070_),
    .A(net870),
    .Y(_06224_));
 sg13g2_buf_1 _24549_ (.A(_06224_),
    .X(_06225_));
 sg13g2_buf_1 _24550_ (.A(net304),
    .X(_06226_));
 sg13g2_nand2_1 _24551_ (.Y(_06227_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][0] ),
    .B(net304));
 sg13g2_o21ai_1 _24552_ (.B1(_06227_),
    .Y(_01729_),
    .A1(net581),
    .A2(net245));
 sg13g2_nand2_1 _24553_ (.Y(_06228_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][10] ),
    .B(net304));
 sg13g2_o21ai_1 _24554_ (.B1(_06228_),
    .Y(_01730_),
    .A1(net646),
    .A2(_06226_));
 sg13g2_nand2_1 _24555_ (.Y(_06229_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][11] ),
    .B(net304));
 sg13g2_o21ai_1 _24556_ (.B1(_06229_),
    .Y(_01731_),
    .A1(net580),
    .A2(_06226_));
 sg13g2_nand2_1 _24557_ (.Y(_06230_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][1] ),
    .B(net304));
 sg13g2_o21ai_1 _24558_ (.B1(_06230_),
    .Y(_01732_),
    .A1(net726),
    .A2(net245));
 sg13g2_mux2_1 _24559_ (.A0(net725),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][2] ),
    .S(net245),
    .X(_01733_));
 sg13g2_mux2_1 _24560_ (.A0(net724),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][3] ),
    .S(net245),
    .X(_01734_));
 sg13g2_mux2_1 _24561_ (.A0(net723),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][4] ),
    .S(net245),
    .X(_01735_));
 sg13g2_mux2_1 _24562_ (.A0(net858),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][5] ),
    .S(_06225_),
    .X(_01736_));
 sg13g2_mux2_1 _24563_ (.A0(net857),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][6] ),
    .S(_06225_),
    .X(_01737_));
 sg13g2_nand2_1 _24564_ (.Y(_06231_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][7] ),
    .B(net304));
 sg13g2_o21ai_1 _24565_ (.B1(_06231_),
    .Y(_01738_),
    .A1(net722),
    .A2(net245));
 sg13g2_nand2_1 _24566_ (.Y(_06232_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][8] ),
    .B(net304));
 sg13g2_o21ai_1 _24567_ (.B1(_06232_),
    .Y(_01739_),
    .A1(net728),
    .A2(net245));
 sg13g2_nand2_1 _24568_ (.Y(_06233_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][9] ),
    .B(net304));
 sg13g2_o21ai_1 _24569_ (.B1(_06233_),
    .Y(_01740_),
    .A1(net727),
    .A2(net245));
 sg13g2_buf_1 _24570_ (.A(net656),
    .X(_06234_));
 sg13g2_nand2_1 _24571_ (.Y(_06235_),
    .A(_05956_),
    .B(net463));
 sg13g2_buf_1 _24572_ (.A(_06235_),
    .X(_06236_));
 sg13g2_buf_1 _24573_ (.A(net369),
    .X(_06237_));
 sg13g2_nand2_1 _24574_ (.Y(_06238_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][0] ),
    .B(net369));
 sg13g2_o21ai_1 _24575_ (.B1(_06238_),
    .Y(_01741_),
    .A1(net579),
    .A2(net303));
 sg13g2_buf_1 _24576_ (.A(net740),
    .X(_06239_));
 sg13g2_nand2_1 _24577_ (.Y(_06240_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][10] ),
    .B(net369));
 sg13g2_o21ai_1 _24578_ (.B1(_06240_),
    .Y(_01742_),
    .A1(net645),
    .A2(net303));
 sg13g2_buf_1 _24579_ (.A(net670),
    .X(_06241_));
 sg13g2_nand2_1 _24580_ (.Y(_06242_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][11] ),
    .B(net369));
 sg13g2_o21ai_1 _24581_ (.B1(_06242_),
    .Y(_01743_),
    .A1(net578),
    .A2(_06237_));
 sg13g2_nand2_1 _24582_ (.Y(_06243_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][1] ),
    .B(net369));
 sg13g2_o21ai_1 _24583_ (.B1(_06243_),
    .Y(_01744_),
    .A1(net726),
    .A2(net303));
 sg13g2_mux2_1 _24584_ (.A0(_06216_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][2] ),
    .S(net303),
    .X(_01745_));
 sg13g2_mux2_1 _24585_ (.A0(_06217_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][3] ),
    .S(net303),
    .X(_01746_));
 sg13g2_mux2_1 _24586_ (.A0(net723),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][4] ),
    .S(net303),
    .X(_01747_));
 sg13g2_mux2_1 _24587_ (.A0(net858),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][5] ),
    .S(_06236_),
    .X(_01748_));
 sg13g2_mux2_1 _24588_ (.A0(net857),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][6] ),
    .S(_06236_),
    .X(_01749_));
 sg13g2_nand2_1 _24589_ (.Y(_06244_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][7] ),
    .B(net369));
 sg13g2_o21ai_1 _24590_ (.B1(_06244_),
    .Y(_01750_),
    .A1(net722),
    .A2(net303));
 sg13g2_buf_1 _24591_ (.A(net876),
    .X(_06245_));
 sg13g2_nand2_1 _24592_ (.Y(_06246_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][8] ),
    .B(net369));
 sg13g2_o21ai_1 _24593_ (.B1(_06246_),
    .Y(_01751_),
    .A1(net721),
    .A2(net303));
 sg13g2_buf_1 _24594_ (.A(net875),
    .X(_06247_));
 sg13g2_nand2_1 _24595_ (.Y(_06248_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][9] ),
    .B(net369));
 sg13g2_o21ai_1 _24596_ (.B1(_06248_),
    .Y(_01752_),
    .A1(net720),
    .A2(_06237_));
 sg13g2_nand2_1 _24597_ (.Y(_06249_),
    .A(_05961_),
    .B(net463));
 sg13g2_buf_1 _24598_ (.A(_06249_),
    .X(_06250_));
 sg13g2_buf_1 _24599_ (.A(net368),
    .X(_06251_));
 sg13g2_nand2_1 _24600_ (.Y(_06252_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][0] ),
    .B(net368));
 sg13g2_o21ai_1 _24601_ (.B1(_06252_),
    .Y(_01753_),
    .A1(net579),
    .A2(net302));
 sg13g2_nand2_1 _24602_ (.Y(_06253_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][10] ),
    .B(net368));
 sg13g2_o21ai_1 _24603_ (.B1(_06253_),
    .Y(_01754_),
    .A1(net645),
    .A2(net302));
 sg13g2_nand2_1 _24604_ (.Y(_06254_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][11] ),
    .B(net368));
 sg13g2_o21ai_1 _24605_ (.B1(_06254_),
    .Y(_01755_),
    .A1(net578),
    .A2(_06251_));
 sg13g2_nand2_1 _24606_ (.Y(_06255_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][1] ),
    .B(net368));
 sg13g2_o21ai_1 _24607_ (.B1(_06255_),
    .Y(_01756_),
    .A1(net726),
    .A2(net302));
 sg13g2_mux2_1 _24608_ (.A0(_06216_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][2] ),
    .S(net302),
    .X(_01757_));
 sg13g2_mux2_1 _24609_ (.A0(_06217_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][3] ),
    .S(net302),
    .X(_01758_));
 sg13g2_mux2_1 _24610_ (.A0(_06218_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][4] ),
    .S(net302),
    .X(_01759_));
 sg13g2_mux2_1 _24611_ (.A0(net858),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][5] ),
    .S(_06250_),
    .X(_01760_));
 sg13g2_mux2_1 _24612_ (.A0(net857),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][6] ),
    .S(_06250_),
    .X(_01761_));
 sg13g2_nand2_1 _24613_ (.Y(_06256_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][7] ),
    .B(net368));
 sg13g2_o21ai_1 _24614_ (.B1(_06256_),
    .Y(_01762_),
    .A1(net722),
    .A2(net302));
 sg13g2_nand2_1 _24615_ (.Y(_06257_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][8] ),
    .B(net368));
 sg13g2_o21ai_1 _24616_ (.B1(_06257_),
    .Y(_01763_),
    .A1(net721),
    .A2(net302));
 sg13g2_nand2_1 _24617_ (.Y(_06258_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][9] ),
    .B(net368));
 sg13g2_o21ai_1 _24618_ (.B1(_06258_),
    .Y(_01764_),
    .A1(net720),
    .A2(_06251_));
 sg13g2_nor2_1 _24619_ (.A(_05845_),
    .B(_05948_),
    .Y(_06259_));
 sg13g2_nand2_1 _24620_ (.Y(_06260_),
    .A(_06259_),
    .B(_06025_));
 sg13g2_buf_1 _24621_ (.A(_06260_),
    .X(_06261_));
 sg13g2_buf_1 _24622_ (.A(net301),
    .X(_06262_));
 sg13g2_nand2_1 _24623_ (.Y(_06263_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][0] ),
    .B(net301));
 sg13g2_o21ai_1 _24624_ (.B1(_06263_),
    .Y(_01765_),
    .A1(net579),
    .A2(net244));
 sg13g2_nand2_1 _24625_ (.Y(_06264_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][10] ),
    .B(net301));
 sg13g2_o21ai_1 _24626_ (.B1(_06264_),
    .Y(_01766_),
    .A1(net645),
    .A2(net244));
 sg13g2_nand2_1 _24627_ (.Y(_06265_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][11] ),
    .B(net301));
 sg13g2_o21ai_1 _24628_ (.B1(_06265_),
    .Y(_01767_),
    .A1(net578),
    .A2(_06262_));
 sg13g2_nand2_1 _24629_ (.Y(_06266_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][1] ),
    .B(net301));
 sg13g2_o21ai_1 _24630_ (.B1(_06266_),
    .Y(_01768_),
    .A1(net726),
    .A2(net244));
 sg13g2_mux2_1 _24631_ (.A0(net725),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][2] ),
    .S(net244),
    .X(_01769_));
 sg13g2_mux2_1 _24632_ (.A0(net724),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][3] ),
    .S(net244),
    .X(_01770_));
 sg13g2_mux2_1 _24633_ (.A0(net723),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][4] ),
    .S(net244),
    .X(_01771_));
 sg13g2_buf_1 _24634_ (.A(_02973_),
    .X(_06267_));
 sg13g2_mux2_1 _24635_ (.A0(net856),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][5] ),
    .S(_06261_),
    .X(_01772_));
 sg13g2_mux2_1 _24636_ (.A0(net857),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][6] ),
    .S(_06261_),
    .X(_01773_));
 sg13g2_nand2_1 _24637_ (.Y(_06268_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][7] ),
    .B(net301));
 sg13g2_o21ai_1 _24638_ (.B1(_06268_),
    .Y(_01774_),
    .A1(net722),
    .A2(net244));
 sg13g2_nand2_1 _24639_ (.Y(_06269_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][8] ),
    .B(net301));
 sg13g2_o21ai_1 _24640_ (.B1(_06269_),
    .Y(_01775_),
    .A1(net721),
    .A2(_06262_));
 sg13g2_nand2_1 _24641_ (.Y(_06270_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][9] ),
    .B(net301));
 sg13g2_o21ai_1 _24642_ (.B1(_06270_),
    .Y(_01776_),
    .A1(net720),
    .A2(net244));
 sg13g2_nand2_1 _24643_ (.Y(_06271_),
    .A(_06259_),
    .B(_06070_));
 sg13g2_buf_1 _24644_ (.A(_06271_),
    .X(_06272_));
 sg13g2_buf_1 _24645_ (.A(net300),
    .X(_06273_));
 sg13g2_nand2_1 _24646_ (.Y(_06274_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][0] ),
    .B(net300));
 sg13g2_o21ai_1 _24647_ (.B1(_06274_),
    .Y(_01777_),
    .A1(net579),
    .A2(net243));
 sg13g2_nand2_1 _24648_ (.Y(_06275_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][10] ),
    .B(net300));
 sg13g2_o21ai_1 _24649_ (.B1(_06275_),
    .Y(_01778_),
    .A1(net645),
    .A2(net243));
 sg13g2_nand2_1 _24650_ (.Y(_06276_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][11] ),
    .B(net300));
 sg13g2_o21ai_1 _24651_ (.B1(_06276_),
    .Y(_01779_),
    .A1(net578),
    .A2(_06273_));
 sg13g2_nand2_1 _24652_ (.Y(_06277_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][1] ),
    .B(net300));
 sg13g2_o21ai_1 _24653_ (.B1(_06277_),
    .Y(_01780_),
    .A1(net726),
    .A2(net243));
 sg13g2_mux2_1 _24654_ (.A0(net725),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][2] ),
    .S(net243),
    .X(_01781_));
 sg13g2_mux2_1 _24655_ (.A0(net724),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][3] ),
    .S(net243),
    .X(_01782_));
 sg13g2_mux2_1 _24656_ (.A0(net723),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][4] ),
    .S(net243),
    .X(_01783_));
 sg13g2_mux2_1 _24657_ (.A0(net856),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][5] ),
    .S(_06272_),
    .X(_01784_));
 sg13g2_mux2_1 _24658_ (.A0(net857),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][6] ),
    .S(_06272_),
    .X(_01785_));
 sg13g2_nand2_1 _24659_ (.Y(_06278_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][7] ),
    .B(net300));
 sg13g2_o21ai_1 _24660_ (.B1(_06278_),
    .Y(_01786_),
    .A1(net722),
    .A2(net243));
 sg13g2_nand2_1 _24661_ (.Y(_06279_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][8] ),
    .B(net300));
 sg13g2_o21ai_1 _24662_ (.B1(_06279_),
    .Y(_01787_),
    .A1(net721),
    .A2(_06273_));
 sg13g2_nand2_1 _24663_ (.Y(_06280_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][9] ),
    .B(net300));
 sg13g2_o21ai_1 _24664_ (.B1(_06280_),
    .Y(_01788_),
    .A1(net720),
    .A2(net243));
 sg13g2_nand3_1 _24665_ (.B(_06021_),
    .C(net462),
    .A(_05858_),
    .Y(_06281_));
 sg13g2_buf_1 _24666_ (.A(_06281_),
    .X(_06282_));
 sg13g2_buf_1 _24667_ (.A(net367),
    .X(_06283_));
 sg13g2_nand2_1 _24668_ (.Y(_06284_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][0] ),
    .B(net367));
 sg13g2_o21ai_1 _24669_ (.B1(_06284_),
    .Y(_01789_),
    .A1(net579),
    .A2(net299));
 sg13g2_nand2_1 _24670_ (.Y(_06285_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][10] ),
    .B(net367));
 sg13g2_o21ai_1 _24671_ (.B1(_06285_),
    .Y(_01790_),
    .A1(_06239_),
    .A2(_06283_));
 sg13g2_nand2_1 _24672_ (.Y(_06286_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][11] ),
    .B(net367));
 sg13g2_o21ai_1 _24673_ (.B1(_06286_),
    .Y(_01791_),
    .A1(_06241_),
    .A2(net299));
 sg13g2_nand2_1 _24674_ (.Y(_06287_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][1] ),
    .B(net367));
 sg13g2_o21ai_1 _24675_ (.B1(_06287_),
    .Y(_01792_),
    .A1(_06214_),
    .A2(net299));
 sg13g2_mux2_1 _24676_ (.A0(net725),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][2] ),
    .S(net299),
    .X(_01793_));
 sg13g2_mux2_1 _24677_ (.A0(net724),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][3] ),
    .S(net299),
    .X(_01794_));
 sg13g2_mux2_1 _24678_ (.A0(net723),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][4] ),
    .S(net299),
    .X(_01795_));
 sg13g2_mux2_1 _24679_ (.A0(_06267_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][5] ),
    .S(_06282_),
    .X(_01796_));
 sg13g2_mux2_1 _24680_ (.A0(_06219_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][6] ),
    .S(_06282_),
    .X(_01797_));
 sg13g2_nand2_1 _24681_ (.Y(_06288_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][7] ),
    .B(net367));
 sg13g2_o21ai_1 _24682_ (.B1(_06288_),
    .Y(_01798_),
    .A1(_06220_),
    .A2(net299));
 sg13g2_nand2_1 _24683_ (.Y(_06289_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][8] ),
    .B(net367));
 sg13g2_o21ai_1 _24684_ (.B1(_06289_),
    .Y(_01799_),
    .A1(net721),
    .A2(_06283_));
 sg13g2_nand2_1 _24685_ (.Y(_06290_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][9] ),
    .B(net367));
 sg13g2_o21ai_1 _24686_ (.B1(_06290_),
    .Y(_01800_),
    .A1(net720),
    .A2(net299));
 sg13g2_nand3_1 _24687_ (.B(_06259_),
    .C(net462),
    .A(_05858_),
    .Y(_06291_));
 sg13g2_buf_1 _24688_ (.A(_06291_),
    .X(_06292_));
 sg13g2_buf_1 _24689_ (.A(net366),
    .X(_06293_));
 sg13g2_nand2_1 _24690_ (.Y(_06294_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][0] ),
    .B(net366));
 sg13g2_o21ai_1 _24691_ (.B1(_06294_),
    .Y(_01801_),
    .A1(net579),
    .A2(net298));
 sg13g2_nand2_1 _24692_ (.Y(_06295_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][10] ),
    .B(net366));
 sg13g2_o21ai_1 _24693_ (.B1(_06295_),
    .Y(_01802_),
    .A1(net645),
    .A2(net298));
 sg13g2_nand2_1 _24694_ (.Y(_06296_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][11] ),
    .B(net366));
 sg13g2_o21ai_1 _24695_ (.B1(_06296_),
    .Y(_01803_),
    .A1(net578),
    .A2(_06293_));
 sg13g2_nand2_1 _24696_ (.Y(_06297_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][1] ),
    .B(net366));
 sg13g2_o21ai_1 _24697_ (.B1(_06297_),
    .Y(_01804_),
    .A1(net726),
    .A2(net298));
 sg13g2_mux2_1 _24698_ (.A0(net725),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][2] ),
    .S(net298),
    .X(_01805_));
 sg13g2_mux2_1 _24699_ (.A0(net724),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][3] ),
    .S(net298),
    .X(_01806_));
 sg13g2_mux2_1 _24700_ (.A0(net723),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][4] ),
    .S(net298),
    .X(_01807_));
 sg13g2_mux2_1 _24701_ (.A0(net856),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][5] ),
    .S(_06292_),
    .X(_01808_));
 sg13g2_mux2_1 _24702_ (.A0(net857),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][6] ),
    .S(_06292_),
    .X(_01809_));
 sg13g2_nand2_1 _24703_ (.Y(_06298_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][7] ),
    .B(net366));
 sg13g2_o21ai_1 _24704_ (.B1(_06298_),
    .Y(_01810_),
    .A1(net722),
    .A2(net298));
 sg13g2_nand2_1 _24705_ (.Y(_06299_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][8] ),
    .B(net366));
 sg13g2_o21ai_1 _24706_ (.B1(_06299_),
    .Y(_01811_),
    .A1(net721),
    .A2(_06293_));
 sg13g2_nand2_1 _24707_ (.Y(_06300_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][9] ),
    .B(net366));
 sg13g2_o21ai_1 _24708_ (.B1(_06300_),
    .Y(_01812_),
    .A1(net720),
    .A2(net298));
 sg13g2_nand3_1 _24709_ (.B(_06259_),
    .C(net462),
    .A(_05814_),
    .Y(_06301_));
 sg13g2_buf_1 _24710_ (.A(_06301_),
    .X(_06302_));
 sg13g2_buf_1 _24711_ (.A(net365),
    .X(_06303_));
 sg13g2_nand2_1 _24712_ (.Y(_06304_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][0] ),
    .B(net365));
 sg13g2_o21ai_1 _24713_ (.B1(_06304_),
    .Y(_01813_),
    .A1(net579),
    .A2(net297));
 sg13g2_nand2_1 _24714_ (.Y(_06305_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][10] ),
    .B(net365));
 sg13g2_o21ai_1 _24715_ (.B1(_06305_),
    .Y(_01814_),
    .A1(net645),
    .A2(net297));
 sg13g2_nand2_1 _24716_ (.Y(_06306_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][11] ),
    .B(net365));
 sg13g2_o21ai_1 _24717_ (.B1(_06306_),
    .Y(_01815_),
    .A1(net578),
    .A2(_06303_));
 sg13g2_nand2_1 _24718_ (.Y(_06307_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][1] ),
    .B(net365));
 sg13g2_o21ai_1 _24719_ (.B1(_06307_),
    .Y(_01816_),
    .A1(net726),
    .A2(net297));
 sg13g2_mux2_1 _24720_ (.A0(net725),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][2] ),
    .S(net297),
    .X(_01817_));
 sg13g2_mux2_1 _24721_ (.A0(net724),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][3] ),
    .S(net297),
    .X(_01818_));
 sg13g2_mux2_1 _24722_ (.A0(net723),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][4] ),
    .S(net297),
    .X(_01819_));
 sg13g2_mux2_1 _24723_ (.A0(net856),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][5] ),
    .S(_06302_),
    .X(_01820_));
 sg13g2_mux2_1 _24724_ (.A0(net857),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][6] ),
    .S(_06302_),
    .X(_01821_));
 sg13g2_nand2_1 _24725_ (.Y(_06308_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][7] ),
    .B(net365));
 sg13g2_o21ai_1 _24726_ (.B1(_06308_),
    .Y(_01822_),
    .A1(net722),
    .A2(net297));
 sg13g2_nand2_1 _24727_ (.Y(_06309_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][8] ),
    .B(net365));
 sg13g2_o21ai_1 _24728_ (.B1(_06309_),
    .Y(_01823_),
    .A1(net721),
    .A2(_06303_));
 sg13g2_nand2_1 _24729_ (.Y(_06310_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][9] ),
    .B(net365));
 sg13g2_o21ai_1 _24730_ (.B1(_06310_),
    .Y(_01824_),
    .A1(net720),
    .A2(net297));
 sg13g2_nand3_1 _24731_ (.B(_06021_),
    .C(net462),
    .A(_05814_),
    .Y(_06311_));
 sg13g2_buf_1 _24732_ (.A(_06311_),
    .X(_06312_));
 sg13g2_buf_1 _24733_ (.A(net364),
    .X(_06313_));
 sg13g2_nand2_1 _24734_ (.Y(_06314_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][0] ),
    .B(net364));
 sg13g2_o21ai_1 _24735_ (.B1(_06314_),
    .Y(_01825_),
    .A1(net579),
    .A2(net296));
 sg13g2_nand2_1 _24736_ (.Y(_06315_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][10] ),
    .B(net364));
 sg13g2_o21ai_1 _24737_ (.B1(_06315_),
    .Y(_01826_),
    .A1(_06239_),
    .A2(_06313_));
 sg13g2_nand2_1 _24738_ (.Y(_06316_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][11] ),
    .B(net364));
 sg13g2_o21ai_1 _24739_ (.B1(_06316_),
    .Y(_01827_),
    .A1(_06241_),
    .A2(net296));
 sg13g2_nand2_1 _24740_ (.Y(_06317_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][1] ),
    .B(net364));
 sg13g2_o21ai_1 _24741_ (.B1(_06317_),
    .Y(_01828_),
    .A1(_06214_),
    .A2(net296));
 sg13g2_mux2_1 _24742_ (.A0(net725),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][2] ),
    .S(net296),
    .X(_01829_));
 sg13g2_mux2_1 _24743_ (.A0(net724),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][3] ),
    .S(net296),
    .X(_01830_));
 sg13g2_mux2_1 _24744_ (.A0(_06218_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][4] ),
    .S(net296),
    .X(_01831_));
 sg13g2_mux2_1 _24745_ (.A0(_06267_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][5] ),
    .S(_06312_),
    .X(_01832_));
 sg13g2_mux2_1 _24746_ (.A0(_06219_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][6] ),
    .S(_06312_),
    .X(_01833_));
 sg13g2_nand2_1 _24747_ (.Y(_06318_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][7] ),
    .B(net364));
 sg13g2_o21ai_1 _24748_ (.B1(_06318_),
    .Y(_01834_),
    .A1(_06220_),
    .A2(net296));
 sg13g2_nand2_1 _24749_ (.Y(_06319_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][8] ),
    .B(net364));
 sg13g2_o21ai_1 _24750_ (.B1(_06319_),
    .Y(_01835_),
    .A1(net721),
    .A2(_06313_));
 sg13g2_nand2_1 _24751_ (.Y(_06320_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][9] ),
    .B(net364));
 sg13g2_o21ai_1 _24752_ (.B1(_06320_),
    .Y(_01836_),
    .A1(net720),
    .A2(net296));
 sg13g2_nand3_1 _24753_ (.B(_06003_),
    .C(_06025_),
    .A(net1016),
    .Y(_06321_));
 sg13g2_buf_1 _24754_ (.A(_06321_),
    .X(_06322_));
 sg13g2_buf_1 _24755_ (.A(net295),
    .X(_06323_));
 sg13g2_nand2_1 _24756_ (.Y(_06324_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][0] ),
    .B(net295));
 sg13g2_o21ai_1 _24757_ (.B1(_06324_),
    .Y(_01837_),
    .A1(_06234_),
    .A2(net242));
 sg13g2_nand2_1 _24758_ (.Y(_06325_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][10] ),
    .B(net295));
 sg13g2_o21ai_1 _24759_ (.B1(_06325_),
    .Y(_01838_),
    .A1(net645),
    .A2(net242));
 sg13g2_nand2_1 _24760_ (.Y(_06326_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][11] ),
    .B(net295));
 sg13g2_o21ai_1 _24761_ (.B1(_06326_),
    .Y(_01839_),
    .A1(net578),
    .A2(net242));
 sg13g2_nand2_1 _24762_ (.Y(_06327_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][1] ),
    .B(net295));
 sg13g2_o21ai_1 _24763_ (.B1(_06327_),
    .Y(_01840_),
    .A1(net890),
    .A2(net242));
 sg13g2_mux2_1 _24764_ (.A0(net751),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][2] ),
    .S(net242),
    .X(_01841_));
 sg13g2_mux2_1 _24765_ (.A0(net750),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][3] ),
    .S(net242),
    .X(_01842_));
 sg13g2_mux2_1 _24766_ (.A0(net749),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][4] ),
    .S(net242),
    .X(_01843_));
 sg13g2_mux2_1 _24767_ (.A0(net856),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][5] ),
    .S(net295),
    .X(_01844_));
 sg13g2_mux2_1 _24768_ (.A0(net883),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][6] ),
    .S(net295),
    .X(_01845_));
 sg13g2_nand2_1 _24769_ (.Y(_06328_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][7] ),
    .B(net295));
 sg13g2_o21ai_1 _24770_ (.B1(_06328_),
    .Y(_01846_),
    .A1(net885),
    .A2(net242));
 sg13g2_nand2_1 _24771_ (.Y(_06329_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][8] ),
    .B(_06322_));
 sg13g2_o21ai_1 _24772_ (.B1(_06329_),
    .Y(_01847_),
    .A1(_06245_),
    .A2(_06323_));
 sg13g2_nand2_1 _24773_ (.Y(_06330_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][9] ),
    .B(_06322_));
 sg13g2_o21ai_1 _24774_ (.B1(_06330_),
    .Y(_01848_),
    .A1(_06247_),
    .A2(_06323_));
 sg13g2_nand2_1 _24775_ (.Y(_06331_),
    .A(_05999_),
    .B(net463));
 sg13g2_buf_1 _24776_ (.A(_06331_),
    .X(_06332_));
 sg13g2_buf_1 _24777_ (.A(net363),
    .X(_06333_));
 sg13g2_nand2_1 _24778_ (.Y(_06334_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][0] ),
    .B(net363));
 sg13g2_o21ai_1 _24779_ (.B1(_06334_),
    .Y(_01849_),
    .A1(_06234_),
    .A2(net294));
 sg13g2_nand2_1 _24780_ (.Y(_06335_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][10] ),
    .B(net363));
 sg13g2_o21ai_1 _24781_ (.B1(_06335_),
    .Y(_01850_),
    .A1(net645),
    .A2(net294));
 sg13g2_nand2_1 _24782_ (.Y(_06336_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][11] ),
    .B(net363));
 sg13g2_o21ai_1 _24783_ (.B1(_06336_),
    .Y(_01851_),
    .A1(net578),
    .A2(net294));
 sg13g2_nand2_1 _24784_ (.Y(_06337_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][1] ),
    .B(net363));
 sg13g2_o21ai_1 _24785_ (.B1(_06337_),
    .Y(_01852_),
    .A1(net890),
    .A2(_06333_));
 sg13g2_mux2_1 _24786_ (.A0(net751),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][2] ),
    .S(net294),
    .X(_01853_));
 sg13g2_mux2_1 _24787_ (.A0(net750),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][3] ),
    .S(net294),
    .X(_01854_));
 sg13g2_mux2_1 _24788_ (.A0(net749),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][4] ),
    .S(net294),
    .X(_01855_));
 sg13g2_mux2_1 _24789_ (.A0(net856),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][5] ),
    .S(net363),
    .X(_01856_));
 sg13g2_mux2_1 _24790_ (.A0(net883),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][6] ),
    .S(net363),
    .X(_01857_));
 sg13g2_nand2_1 _24791_ (.Y(_06338_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][7] ),
    .B(net363));
 sg13g2_o21ai_1 _24792_ (.B1(_06338_),
    .Y(_01858_),
    .A1(net885),
    .A2(net294));
 sg13g2_nand2_1 _24793_ (.Y(_06339_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][8] ),
    .B(_06332_));
 sg13g2_o21ai_1 _24794_ (.B1(_06339_),
    .Y(_01859_),
    .A1(_06245_),
    .A2(_06333_));
 sg13g2_nand2_1 _24795_ (.Y(_06340_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][9] ),
    .B(_06332_));
 sg13g2_o21ai_1 _24796_ (.B1(_06340_),
    .Y(_01860_),
    .A1(_06247_),
    .A2(net294));
 sg13g2_nand2_1 _24797_ (.Y(_06341_),
    .A(_06005_),
    .B(net463));
 sg13g2_buf_1 _24798_ (.A(_06341_),
    .X(_06342_));
 sg13g2_buf_1 _24799_ (.A(net362),
    .X(_06343_));
 sg13g2_nand2_1 _24800_ (.Y(_06344_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][0] ),
    .B(net362));
 sg13g2_o21ai_1 _24801_ (.B1(_06344_),
    .Y(_01861_),
    .A1(net656),
    .A2(net293));
 sg13g2_nand2_1 _24802_ (.Y(_06345_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][10] ),
    .B(net362));
 sg13g2_o21ai_1 _24803_ (.B1(_06345_),
    .Y(_01862_),
    .A1(net740),
    .A2(net293));
 sg13g2_nand2_1 _24804_ (.Y(_06346_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][11] ),
    .B(net362));
 sg13g2_o21ai_1 _24805_ (.B1(_06346_),
    .Y(_01863_),
    .A1(net670),
    .A2(net293));
 sg13g2_nand2_1 _24806_ (.Y(_06347_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][1] ),
    .B(net362));
 sg13g2_o21ai_1 _24807_ (.B1(_06347_),
    .Y(_01864_),
    .A1(net890),
    .A2(net293));
 sg13g2_mux2_1 _24808_ (.A0(net751),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][2] ),
    .S(net293),
    .X(_01865_));
 sg13g2_mux2_1 _24809_ (.A0(net750),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][3] ),
    .S(net293),
    .X(_01866_));
 sg13g2_mux2_1 _24810_ (.A0(net749),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][4] ),
    .S(net293),
    .X(_01867_));
 sg13g2_mux2_1 _24811_ (.A0(net856),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][5] ),
    .S(net362),
    .X(_01868_));
 sg13g2_mux2_1 _24812_ (.A0(net883),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][6] ),
    .S(net362),
    .X(_01869_));
 sg13g2_nand2_1 _24813_ (.Y(_06348_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][7] ),
    .B(net362));
 sg13g2_o21ai_1 _24814_ (.B1(_06348_),
    .Y(_01870_),
    .A1(_02962_),
    .A2(net293));
 sg13g2_nand2_1 _24815_ (.Y(_06349_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][8] ),
    .B(_06342_));
 sg13g2_o21ai_1 _24816_ (.B1(_06349_),
    .Y(_01871_),
    .A1(net876),
    .A2(_06343_));
 sg13g2_nand2_1 _24817_ (.Y(_06350_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][9] ),
    .B(_06342_));
 sg13g2_o21ai_1 _24818_ (.B1(_06350_),
    .Y(_01872_),
    .A1(net875),
    .A2(_06343_));
 sg13g2_nand2_1 _24819_ (.Y(_06351_),
    .A(_06010_),
    .B(_06037_));
 sg13g2_buf_1 _24820_ (.A(_06351_),
    .X(_06352_));
 sg13g2_buf_1 _24821_ (.A(net361),
    .X(_06353_));
 sg13g2_nand2_1 _24822_ (.Y(_06354_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][0] ),
    .B(net361));
 sg13g2_o21ai_1 _24823_ (.B1(_06354_),
    .Y(_01873_),
    .A1(net656),
    .A2(net292));
 sg13g2_nand2_1 _24824_ (.Y(_06355_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][10] ),
    .B(net361));
 sg13g2_o21ai_1 _24825_ (.B1(_06355_),
    .Y(_01874_),
    .A1(net740),
    .A2(net292));
 sg13g2_nand2_1 _24826_ (.Y(_06356_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][11] ),
    .B(net361));
 sg13g2_o21ai_1 _24827_ (.B1(_06356_),
    .Y(_01875_),
    .A1(net670),
    .A2(net292));
 sg13g2_nand2_1 _24828_ (.Y(_06357_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][1] ),
    .B(net361));
 sg13g2_o21ai_1 _24829_ (.B1(_06357_),
    .Y(_01876_),
    .A1(net890),
    .A2(net292));
 sg13g2_mux2_1 _24830_ (.A0(net751),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][2] ),
    .S(net292),
    .X(_01877_));
 sg13g2_mux2_1 _24831_ (.A0(net750),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][3] ),
    .S(net292),
    .X(_01878_));
 sg13g2_mux2_1 _24832_ (.A0(net749),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][4] ),
    .S(net292),
    .X(_01879_));
 sg13g2_mux2_1 _24833_ (.A0(net856),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][5] ),
    .S(net361),
    .X(_01880_));
 sg13g2_mux2_1 _24834_ (.A0(net883),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][6] ),
    .S(net361),
    .X(_01881_));
 sg13g2_nand2_1 _24835_ (.Y(_06358_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][7] ),
    .B(net361));
 sg13g2_o21ai_1 _24836_ (.B1(_06358_),
    .Y(_01882_),
    .A1(net885),
    .A2(net292));
 sg13g2_nand2_1 _24837_ (.Y(_06359_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][8] ),
    .B(_06352_));
 sg13g2_o21ai_1 _24838_ (.B1(_06359_),
    .Y(_01883_),
    .A1(net876),
    .A2(_06353_));
 sg13g2_nand2_1 _24839_ (.Y(_06360_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][9] ),
    .B(_06352_));
 sg13g2_o21ai_1 _24840_ (.B1(_06360_),
    .Y(_01884_),
    .A1(net875),
    .A2(_06353_));
 sg13g2_nand3_1 _24841_ (.B(_06109_),
    .C(net462),
    .A(_05877_),
    .Y(_06361_));
 sg13g2_buf_1 _24842_ (.A(_06361_),
    .X(_06362_));
 sg13g2_buf_1 _24843_ (.A(net360),
    .X(_06363_));
 sg13g2_nand2_1 _24844_ (.Y(_06364_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][0] ),
    .B(net360));
 sg13g2_o21ai_1 _24845_ (.B1(_06364_),
    .Y(_01885_),
    .A1(net656),
    .A2(net291));
 sg13g2_nand2_1 _24846_ (.Y(_06365_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][10] ),
    .B(net360));
 sg13g2_o21ai_1 _24847_ (.B1(_06365_),
    .Y(_01886_),
    .A1(net740),
    .A2(net291));
 sg13g2_nand2_1 _24848_ (.Y(_06366_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][11] ),
    .B(net360));
 sg13g2_o21ai_1 _24849_ (.B1(_06366_),
    .Y(_01887_),
    .A1(net670),
    .A2(net291));
 sg13g2_nand2_1 _24850_ (.Y(_06367_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][1] ),
    .B(net360));
 sg13g2_o21ai_1 _24851_ (.B1(_06367_),
    .Y(_01888_),
    .A1(net890),
    .A2(net291));
 sg13g2_mux2_1 _24852_ (.A0(net751),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][2] ),
    .S(net291),
    .X(_01889_));
 sg13g2_mux2_1 _24853_ (.A0(net750),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][3] ),
    .S(net291),
    .X(_01890_));
 sg13g2_mux2_1 _24854_ (.A0(net749),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][4] ),
    .S(net291),
    .X(_01891_));
 sg13g2_mux2_1 _24855_ (.A0(net884),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][5] ),
    .S(net360),
    .X(_01892_));
 sg13g2_mux2_1 _24856_ (.A0(net883),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][6] ),
    .S(net360),
    .X(_01893_));
 sg13g2_nand2_1 _24857_ (.Y(_06368_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][7] ),
    .B(net360));
 sg13g2_o21ai_1 _24858_ (.B1(_06368_),
    .Y(_01894_),
    .A1(net885),
    .A2(net291));
 sg13g2_nand2_1 _24859_ (.Y(_06369_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][8] ),
    .B(_06362_));
 sg13g2_o21ai_1 _24860_ (.B1(_06369_),
    .Y(_01895_),
    .A1(net876),
    .A2(_06363_));
 sg13g2_nand2_1 _24861_ (.Y(_06370_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][9] ),
    .B(_06362_));
 sg13g2_o21ai_1 _24862_ (.B1(_06370_),
    .Y(_01896_),
    .A1(net875),
    .A2(_06363_));
 sg13g2_nand3_1 _24863_ (.B(_05877_),
    .C(_06070_),
    .A(net870),
    .Y(_06371_));
 sg13g2_buf_1 _24864_ (.A(_06371_),
    .X(_06372_));
 sg13g2_buf_1 _24865_ (.A(net290),
    .X(_06373_));
 sg13g2_nand2_1 _24866_ (.Y(_06374_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][0] ),
    .B(net290));
 sg13g2_o21ai_1 _24867_ (.B1(_06374_),
    .Y(_01897_),
    .A1(_03707_),
    .A2(_06373_));
 sg13g2_nand2_1 _24868_ (.Y(_06375_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][10] ),
    .B(net290));
 sg13g2_o21ai_1 _24869_ (.B1(_06375_),
    .Y(_01898_),
    .A1(net740),
    .A2(net241));
 sg13g2_nand2_1 _24870_ (.Y(_06376_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][11] ),
    .B(net290));
 sg13g2_o21ai_1 _24871_ (.B1(_06376_),
    .Y(_01899_),
    .A1(net670),
    .A2(net241));
 sg13g2_nand2_1 _24872_ (.Y(_06377_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][1] ),
    .B(net290));
 sg13g2_o21ai_1 _24873_ (.B1(_06377_),
    .Y(_01900_),
    .A1(_02943_),
    .A2(net241));
 sg13g2_mux2_1 _24874_ (.A0(net751),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][2] ),
    .S(net241),
    .X(_01901_));
 sg13g2_mux2_1 _24875_ (.A0(net750),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][3] ),
    .S(net241),
    .X(_01902_));
 sg13g2_mux2_1 _24876_ (.A0(net749),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][4] ),
    .S(net241),
    .X(_01903_));
 sg13g2_mux2_1 _24877_ (.A0(net884),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][5] ),
    .S(net290),
    .X(_01904_));
 sg13g2_mux2_1 _24878_ (.A0(net883),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][6] ),
    .S(net290),
    .X(_01905_));
 sg13g2_nand2_1 _24879_ (.Y(_06378_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][7] ),
    .B(net290));
 sg13g2_o21ai_1 _24880_ (.B1(_06378_),
    .Y(_01906_),
    .A1(net885),
    .A2(net241));
 sg13g2_nand2_1 _24881_ (.Y(_06379_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][8] ),
    .B(_06372_));
 sg13g2_o21ai_1 _24882_ (.B1(_06379_),
    .Y(_01907_),
    .A1(net876),
    .A2(net241));
 sg13g2_nand2_1 _24883_ (.Y(_06380_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][9] ),
    .B(_06372_));
 sg13g2_o21ai_1 _24884_ (.B1(_06380_),
    .Y(_01908_),
    .A1(net875),
    .A2(_06373_));
 sg13g2_mux2_1 _24885_ (.A0(\cpu.genblk1.mmu.r_writeable_d[0] ),
    .A1(net434),
    .S(_05853_),
    .X(_01909_));
 sg13g2_buf_1 _24886_ (.A(net475),
    .X(_06381_));
 sg13g2_mux2_1 _24887_ (.A0(\cpu.genblk1.mmu.r_writeable_d[10] ),
    .A1(_06381_),
    .S(_05864_),
    .X(_01910_));
 sg13g2_mux2_1 _24888_ (.A0(\cpu.genblk1.mmu.r_writeable_d[11] ),
    .A1(net426),
    .S(_05873_),
    .X(_01911_));
 sg13g2_mux2_1 _24889_ (.A0(\cpu.genblk1.mmu.r_writeable_d[12] ),
    .A1(net426),
    .S(_05881_),
    .X(_01912_));
 sg13g2_mux2_1 _24890_ (.A0(\cpu.genblk1.mmu.r_writeable_d[13] ),
    .A1(net426),
    .S(_05888_),
    .X(_01913_));
 sg13g2_mux2_1 _24891_ (.A0(\cpu.genblk1.mmu.r_writeable_d[14] ),
    .A1(net426),
    .S(_05892_),
    .X(_01914_));
 sg13g2_mux2_1 _24892_ (.A0(\cpu.genblk1.mmu.r_writeable_d[15] ),
    .A1(_06381_),
    .S(_05898_),
    .X(_01915_));
 sg13g2_mux2_1 _24893_ (.A0(\cpu.genblk1.mmu.r_writeable_d[16] ),
    .A1(net426),
    .S(_05904_),
    .X(_01916_));
 sg13g2_mux2_1 _24894_ (.A0(\cpu.genblk1.mmu.r_writeable_d[17] ),
    .A1(net426),
    .S(_05908_),
    .X(_01917_));
 sg13g2_mux2_1 _24895_ (.A0(\cpu.genblk1.mmu.r_writeable_d[18] ),
    .A1(net426),
    .S(_05912_),
    .X(_01918_));
 sg13g2_mux2_1 _24896_ (.A0(\cpu.genblk1.mmu.r_writeable_d[19] ),
    .A1(net426),
    .S(_05920_),
    .X(_01919_));
 sg13g2_buf_1 _24897_ (.A(net475),
    .X(_06382_));
 sg13g2_mux2_1 _24898_ (.A0(\cpu.genblk1.mmu.r_writeable_d[1] ),
    .A1(_06382_),
    .S(_05924_),
    .X(_01920_));
 sg13g2_mux2_1 _24899_ (.A0(\cpu.genblk1.mmu.r_writeable_d[20] ),
    .A1(net425),
    .S(_05932_),
    .X(_01921_));
 sg13g2_mux2_1 _24900_ (.A0(\cpu.genblk1.mmu.r_writeable_d[21] ),
    .A1(net425),
    .S(_05937_),
    .X(_01922_));
 sg13g2_mux2_1 _24901_ (.A0(\cpu.genblk1.mmu.r_writeable_d[22] ),
    .A1(net425),
    .S(_05941_),
    .X(_01923_));
 sg13g2_mux2_1 _24902_ (.A0(\cpu.genblk1.mmu.r_writeable_d[23] ),
    .A1(_06382_),
    .S(_05944_),
    .X(_01924_));
 sg13g2_mux2_1 _24903_ (.A0(\cpu.genblk1.mmu.r_writeable_d[24] ),
    .A1(net425),
    .S(_05950_),
    .X(_01925_));
 sg13g2_mux2_1 _24904_ (.A0(\cpu.genblk1.mmu.r_writeable_d[25] ),
    .A1(net425),
    .S(_05953_),
    .X(_01926_));
 sg13g2_mux2_1 _24905_ (.A0(\cpu.genblk1.mmu.r_writeable_d[26] ),
    .A1(net425),
    .S(_05958_),
    .X(_01927_));
 sg13g2_mux2_1 _24906_ (.A0(\cpu.genblk1.mmu.r_writeable_d[27] ),
    .A1(net425),
    .S(_05963_),
    .X(_01928_));
 sg13g2_mux2_1 _24907_ (.A0(\cpu.genblk1.mmu.r_writeable_d[28] ),
    .A1(net425),
    .S(_05971_),
    .X(_01929_));
 sg13g2_buf_1 _24908_ (.A(_03432_),
    .X(_06383_));
 sg13g2_mux2_1 _24909_ (.A0(\cpu.genblk1.mmu.r_writeable_d[29] ),
    .A1(net424),
    .S(_05975_),
    .X(_01930_));
 sg13g2_mux2_1 _24910_ (.A0(\cpu.genblk1.mmu.r_writeable_d[2] ),
    .A1(_06383_),
    .S(_05981_),
    .X(_01931_));
 sg13g2_mux2_1 _24911_ (.A0(\cpu.genblk1.mmu.r_writeable_d[30] ),
    .A1(net424),
    .S(_05985_),
    .X(_01932_));
 sg13g2_mux2_1 _24912_ (.A0(\cpu.genblk1.mmu.r_writeable_d[31] ),
    .A1(net424),
    .S(_05989_),
    .X(_01933_));
 sg13g2_mux2_1 _24913_ (.A0(\cpu.genblk1.mmu.r_writeable_d[3] ),
    .A1(net424),
    .S(_05992_),
    .X(_01934_));
 sg13g2_mux2_1 _24914_ (.A0(\cpu.genblk1.mmu.r_writeable_d[4] ),
    .A1(net424),
    .S(_05996_),
    .X(_01935_));
 sg13g2_mux2_1 _24915_ (.A0(\cpu.genblk1.mmu.r_writeable_d[5] ),
    .A1(net424),
    .S(_06001_),
    .X(_01936_));
 sg13g2_mux2_1 _24916_ (.A0(\cpu.genblk1.mmu.r_writeable_d[6] ),
    .A1(net424),
    .S(_06007_),
    .X(_01937_));
 sg13g2_mux2_1 _24917_ (.A0(\cpu.genblk1.mmu.r_writeable_d[7] ),
    .A1(_06383_),
    .S(_06012_),
    .X(_01938_));
 sg13g2_mux2_1 _24918_ (.A0(\cpu.genblk1.mmu.r_writeable_d[8] ),
    .A1(net424),
    .S(_06015_),
    .X(_01939_));
 sg13g2_mux2_1 _24919_ (.A0(\cpu.genblk1.mmu.r_writeable_d[9] ),
    .A1(_03432_),
    .S(_06018_),
    .X(_01940_));
 sg13g2_nor2_1 _24920_ (.A(net984),
    .B(_09368_),
    .Y(_06384_));
 sg13g2_buf_2 _24921_ (.A(_06384_),
    .X(_06385_));
 sg13g2_nand3_1 _24922_ (.B(_09866_),
    .C(_06385_),
    .A(_09280_),
    .Y(_06386_));
 sg13g2_buf_1 _24923_ (.A(_06386_),
    .X(_06387_));
 sg13g2_nor2_1 _24924_ (.A(net931),
    .B(_06387_),
    .Y(_06388_));
 sg13g2_buf_2 _24925_ (.A(_06388_),
    .X(_06389_));
 sg13g2_nand3_1 _24926_ (.B(_10256_),
    .C(_06389_),
    .A(net977),
    .Y(_06390_));
 sg13g2_buf_1 _24927_ (.A(_06390_),
    .X(_06391_));
 sg13g2_mux2_1 _24928_ (.A0(net1032),
    .A1(\cpu.gpio.genblk2[4].srcs_io[0] ),
    .S(_06391_),
    .X(_01957_));
 sg13g2_mux2_1 _24929_ (.A0(net916),
    .A1(\cpu.gpio.genblk2[5].srcs_io[0] ),
    .S(_06391_),
    .X(_01958_));
 sg13g2_mux2_1 _24930_ (.A0(net1031),
    .A1(\cpu.gpio.genblk2[6].srcs_io[0] ),
    .S(_06391_),
    .X(_01959_));
 sg13g2_mux2_1 _24931_ (.A0(net1034),
    .A1(\cpu.gpio.genblk2[7].srcs_io[0] ),
    .S(_06391_),
    .X(_01960_));
 sg13g2_nand3_1 _24932_ (.B(_05132_),
    .C(_06389_),
    .A(net977),
    .Y(_06392_));
 sg13g2_buf_2 _24933_ (.A(_06392_),
    .X(_06393_));
 sg13g2_mux2_1 _24934_ (.A0(net1033),
    .A1(\cpu.gpio.genblk1[3].srcs_o[0] ),
    .S(_06393_),
    .X(_01961_));
 sg13g2_mux2_1 _24935_ (.A0(net1032),
    .A1(\cpu.gpio.genblk1[4].srcs_o[0] ),
    .S(_06393_),
    .X(_01962_));
 sg13g2_mux2_1 _24936_ (.A0(net916),
    .A1(\cpu.gpio.genblk1[5].srcs_o[0] ),
    .S(_06393_),
    .X(_01963_));
 sg13g2_mux2_1 _24937_ (.A0(net1031),
    .A1(\cpu.gpio.genblk1[6].srcs_o[0] ),
    .S(_06393_),
    .X(_01964_));
 sg13g2_mux2_1 _24938_ (.A0(net1034),
    .A1(\cpu.gpio.genblk1[7].srcs_o[0] ),
    .S(_06393_),
    .X(_01965_));
 sg13g2_nand2_1 _24939_ (.Y(_06394_),
    .A(_04983_),
    .B(_06389_));
 sg13g2_buf_4 _24940_ (.X(_06395_),
    .A(_06394_));
 sg13g2_mux2_1 _24941_ (.A0(net897),
    .A1(_04981_),
    .S(_06395_),
    .X(_01966_));
 sg13g2_buf_1 _24942_ (.A(\cpu.gpio.r_spi_miso_src[0][1] ),
    .X(_06396_));
 sg13g2_mux2_1 _24943_ (.A0(net918),
    .A1(_06396_),
    .S(_06395_),
    .X(_01967_));
 sg13g2_mux2_1 _24944_ (.A0(net917),
    .A1(\cpu.gpio.r_spi_miso_src[0][2] ),
    .S(_06395_),
    .X(_01968_));
 sg13g2_mux2_1 _24945_ (.A0(net1033),
    .A1(\cpu.gpio.r_spi_miso_src[0][3] ),
    .S(_06395_),
    .X(_01969_));
 sg13g2_mux2_1 _24946_ (.A0(net1032),
    .A1(_05540_),
    .S(_06395_),
    .X(_01970_));
 sg13g2_buf_1 _24947_ (.A(\cpu.gpio.r_spi_miso_src[1][1] ),
    .X(_06397_));
 sg13g2_mux2_1 _24948_ (.A0(net916),
    .A1(_06397_),
    .S(_06395_),
    .X(_01971_));
 sg13g2_mux2_1 _24949_ (.A0(net1031),
    .A1(\cpu.gpio.r_spi_miso_src[1][2] ),
    .S(_06395_),
    .X(_01972_));
 sg13g2_mux2_1 _24950_ (.A0(net1034),
    .A1(\cpu.gpio.r_spi_miso_src[1][3] ),
    .S(_06395_),
    .X(_01973_));
 sg13g2_nand2_1 _24951_ (.Y(_06398_),
    .A(net428),
    .B(_06389_));
 sg13g2_buf_4 _24952_ (.X(_06399_),
    .A(_06398_));
 sg13g2_mux2_1 _24953_ (.A0(net897),
    .A1(_04989_),
    .S(_06399_),
    .X(_01974_));
 sg13g2_mux2_1 _24954_ (.A0(net918),
    .A1(_05342_),
    .S(_06399_),
    .X(_01975_));
 sg13g2_mux2_1 _24955_ (.A0(net917),
    .A1(_05404_),
    .S(_06399_),
    .X(_01976_));
 sg13g2_mux2_1 _24956_ (.A0(net1033),
    .A1(_05465_),
    .S(_06399_),
    .X(_01977_));
 sg13g2_mux2_1 _24957_ (.A0(net1032),
    .A1(_05544_),
    .S(_06399_),
    .X(_01978_));
 sg13g2_mux2_1 _24958_ (.A0(net916),
    .A1(_05639_),
    .S(_06399_),
    .X(_01979_));
 sg13g2_mux2_1 _24959_ (.A0(net1031),
    .A1(_05671_),
    .S(_06399_),
    .X(_01980_));
 sg13g2_mux2_1 _24960_ (.A0(net1034),
    .A1(_05053_),
    .S(_06399_),
    .X(_01981_));
 sg13g2_nand2_1 _24961_ (.Y(_06400_),
    .A(net427),
    .B(_06389_));
 sg13g2_buf_4 _24962_ (.X(_06401_),
    .A(_06400_));
 sg13g2_mux2_1 _24963_ (.A0(net897),
    .A1(_05006_),
    .S(_06401_),
    .X(_01982_));
 sg13g2_buf_1 _24964_ (.A(\cpu.gpio.r_src_io[6][1] ),
    .X(_06402_));
 sg13g2_mux2_1 _24965_ (.A0(_10244_),
    .A1(_06402_),
    .S(_06401_),
    .X(_01983_));
 sg13g2_mux2_1 _24966_ (.A0(_10264_),
    .A1(\cpu.gpio.r_src_io[6][2] ),
    .S(_06401_),
    .X(_01984_));
 sg13g2_mux2_1 _24967_ (.A0(_10269_),
    .A1(\cpu.gpio.r_src_io[6][3] ),
    .S(_06401_),
    .X(_01985_));
 sg13g2_mux2_1 _24968_ (.A0(net1032),
    .A1(_05547_),
    .S(_06401_),
    .X(_01986_));
 sg13g2_buf_1 _24969_ (.A(\cpu.gpio.r_src_io[7][1] ),
    .X(_06403_));
 sg13g2_mux2_1 _24970_ (.A0(net916),
    .A1(_06403_),
    .S(_06401_),
    .X(_01987_));
 sg13g2_mux2_1 _24971_ (.A0(net1031),
    .A1(\cpu.gpio.r_src_io[7][2] ),
    .S(_06401_),
    .X(_01988_));
 sg13g2_mux2_1 _24972_ (.A0(net1034),
    .A1(\cpu.gpio.r_src_io[7][3] ),
    .S(_06401_),
    .X(_01989_));
 sg13g2_buf_1 _24973_ (.A(_06387_),
    .X(_06404_));
 sg13g2_nor4_2 _24974_ (.A(_11383_),
    .B(net931),
    .C(_05564_),
    .Y(_06405_),
    .D(net96));
 sg13g2_mux2_1 _24975_ (.A0(_05541_),
    .A1(net1002),
    .S(_06405_),
    .X(_01990_));
 sg13g2_buf_1 _24976_ (.A(\cpu.gpio.r_src_o[3][1] ),
    .X(_06406_));
 sg13g2_mux2_1 _24977_ (.A0(_06406_),
    .A1(net1001),
    .S(_06405_),
    .X(_01991_));
 sg13g2_mux2_1 _24978_ (.A0(\cpu.gpio.r_src_o[3][2] ),
    .A1(net1000),
    .S(_06405_),
    .X(_01992_));
 sg13g2_mux2_1 _24979_ (.A0(\cpu.gpio.r_src_o[3][3] ),
    .A1(net991),
    .S(_06405_),
    .X(_01993_));
 sg13g2_nand2_1 _24980_ (.Y(_06407_),
    .A(_04986_),
    .B(_06389_));
 sg13g2_buf_4 _24981_ (.X(_06408_),
    .A(_06407_));
 sg13g2_mux2_1 _24982_ (.A0(net897),
    .A1(_04984_),
    .S(_06408_),
    .X(_01994_));
 sg13g2_buf_1 _24983_ (.A(\cpu.gpio.r_src_o[4][1] ),
    .X(_06409_));
 sg13g2_mux2_1 _24984_ (.A0(_10244_),
    .A1(_06409_),
    .S(_06408_),
    .X(_01995_));
 sg13g2_mux2_1 _24985_ (.A0(net917),
    .A1(\cpu.gpio.r_src_o[4][2] ),
    .S(_06408_),
    .X(_01996_));
 sg13g2_mux2_1 _24986_ (.A0(_10269_),
    .A1(\cpu.gpio.r_src_o[4][3] ),
    .S(_06408_),
    .X(_01997_));
 sg13g2_mux2_1 _24987_ (.A0(_10275_),
    .A1(_05534_),
    .S(_06408_),
    .X(_01998_));
 sg13g2_buf_1 _24988_ (.A(\cpu.gpio.r_src_o[5][1] ),
    .X(_06410_));
 sg13g2_mux2_1 _24989_ (.A0(_10282_),
    .A1(_06410_),
    .S(_06408_),
    .X(_01999_));
 sg13g2_mux2_1 _24990_ (.A0(_10288_),
    .A1(\cpu.gpio.r_src_o[5][2] ),
    .S(_06408_),
    .X(_02000_));
 sg13g2_mux2_1 _24991_ (.A0(_10230_),
    .A1(\cpu.gpio.r_src_o[5][3] ),
    .S(_06408_),
    .X(_02001_));
 sg13g2_nand2_2 _24992_ (.Y(_06411_),
    .A(_05003_),
    .B(_06389_));
 sg13g2_mux2_1 _24993_ (.A0(_10275_),
    .A1(_05545_),
    .S(_06411_),
    .X(_02006_));
 sg13g2_buf_1 _24994_ (.A(\cpu.gpio.r_src_o[7][1] ),
    .X(_06412_));
 sg13g2_mux2_1 _24995_ (.A0(_10282_),
    .A1(_06412_),
    .S(_06411_),
    .X(_02007_));
 sg13g2_mux2_1 _24996_ (.A0(_10288_),
    .A1(\cpu.gpio.r_src_o[7][2] ),
    .S(_06411_),
    .X(_02008_));
 sg13g2_mux2_1 _24997_ (.A0(_10230_),
    .A1(\cpu.gpio.r_src_o[7][3] ),
    .S(_06411_),
    .X(_02009_));
 sg13g2_buf_1 _24998_ (.A(_02836_),
    .X(_06413_));
 sg13g2_and2_1 _24999_ (.A(_08601_),
    .B(_08673_),
    .X(_06414_));
 sg13g2_buf_4 _25000_ (.X(_06415_),
    .A(_06414_));
 sg13g2_buf_1 _25001_ (.A(_00253_),
    .X(_06416_));
 sg13g2_nor2_1 _25002_ (.A(\cpu.icache.r_offset[2] ),
    .B(_06416_),
    .Y(_06417_));
 sg13g2_buf_2 _25003_ (.A(_06417_),
    .X(_06418_));
 sg13g2_buf_1 _25004_ (.A(\cpu.icache.r_offset[1] ),
    .X(_06419_));
 sg13g2_buf_1 _25005_ (.A(\cpu.icache.r_offset[0] ),
    .X(_06420_));
 sg13g2_nor2b_1 _25006_ (.A(_06419_),
    .B_N(_06420_),
    .Y(_06421_));
 sg13g2_buf_1 _25007_ (.A(_06421_),
    .X(_06422_));
 sg13g2_and2_1 _25008_ (.A(_06418_),
    .B(_06422_),
    .X(_06423_));
 sg13g2_buf_2 _25009_ (.A(_06423_),
    .X(_06424_));
 sg13g2_nand2_2 _25010_ (.Y(_06425_),
    .A(_06415_),
    .B(_06424_));
 sg13g2_mux2_1 _25011_ (.A0(net855),
    .A1(\cpu.icache.r_data[0][0] ),
    .S(_06425_),
    .X(_02013_));
 sg13g2_buf_1 _25012_ (.A(_02870_),
    .X(_06426_));
 sg13g2_inv_1 _25013_ (.Y(_06427_),
    .A(_00254_));
 sg13g2_nand2_1 _25014_ (.Y(_06428_),
    .A(_06419_),
    .B(_06420_));
 sg13g2_buf_2 _25015_ (.A(_06428_),
    .X(_06429_));
 sg13g2_nor3_2 _25016_ (.A(_06416_),
    .B(_06427_),
    .C(_06429_),
    .Y(_06430_));
 sg13g2_nand2_2 _25017_ (.Y(_06431_),
    .A(_06415_),
    .B(_06430_));
 sg13g2_mux2_1 _25018_ (.A0(_06426_),
    .A1(\cpu.icache.r_data[0][10] ),
    .S(_06431_),
    .X(_02014_));
 sg13g2_buf_1 _25019_ (.A(_02874_),
    .X(_06432_));
 sg13g2_mux2_1 _25020_ (.A0(net853),
    .A1(\cpu.icache.r_data[0][11] ),
    .S(_06431_),
    .X(_02015_));
 sg13g2_nor2b_1 _25021_ (.A(_06420_),
    .B_N(_06419_),
    .Y(_06433_));
 sg13g2_buf_1 _25022_ (.A(_06433_),
    .X(_06434_));
 sg13g2_and2_1 _25023_ (.A(_06418_),
    .B(_06434_),
    .X(_06435_));
 sg13g2_buf_2 _25024_ (.A(_06435_),
    .X(_06436_));
 sg13g2_nand2_2 _25025_ (.Y(_06437_),
    .A(_06415_),
    .B(_06436_));
 sg13g2_mux2_1 _25026_ (.A0(net855),
    .A1(\cpu.icache.r_data[0][12] ),
    .S(_06437_),
    .X(_02016_));
 sg13g2_buf_1 _25027_ (.A(_02866_),
    .X(_06438_));
 sg13g2_mux2_1 _25028_ (.A0(net852),
    .A1(\cpu.icache.r_data[0][13] ),
    .S(_06437_),
    .X(_02017_));
 sg13g2_mux2_1 _25029_ (.A0(_06426_),
    .A1(\cpu.icache.r_data[0][14] ),
    .S(_06437_),
    .X(_02018_));
 sg13g2_mux2_1 _25030_ (.A0(net853),
    .A1(\cpu.icache.r_data[0][15] ),
    .S(_06437_),
    .X(_02019_));
 sg13g2_nor2_1 _25031_ (.A(_06416_),
    .B(_00254_),
    .Y(_06439_));
 sg13g2_buf_2 _25032_ (.A(_06439_),
    .X(_06440_));
 sg13g2_and2_1 _25033_ (.A(_06422_),
    .B(_06440_),
    .X(_06441_));
 sg13g2_buf_2 _25034_ (.A(_06441_),
    .X(_06442_));
 sg13g2_nand2_2 _25035_ (.Y(_06443_),
    .A(_06415_),
    .B(_06442_));
 sg13g2_mux2_1 _25036_ (.A0(net855),
    .A1(\cpu.icache.r_data[0][16] ),
    .S(_06443_),
    .X(_02020_));
 sg13g2_mux2_1 _25037_ (.A0(net852),
    .A1(\cpu.icache.r_data[0][17] ),
    .S(_06443_),
    .X(_02021_));
 sg13g2_mux2_1 _25038_ (.A0(net854),
    .A1(\cpu.icache.r_data[0][18] ),
    .S(_06443_),
    .X(_02022_));
 sg13g2_mux2_1 _25039_ (.A0(net853),
    .A1(\cpu.icache.r_data[0][19] ),
    .S(_06443_),
    .X(_02023_));
 sg13g2_mux2_1 _25040_ (.A0(net852),
    .A1(\cpu.icache.r_data[0][1] ),
    .S(_06425_),
    .X(_02024_));
 sg13g2_nor2_2 _25041_ (.A(_06419_),
    .B(_06420_),
    .Y(_06444_));
 sg13g2_and2_1 _25042_ (.A(_06440_),
    .B(_06444_),
    .X(_06445_));
 sg13g2_buf_2 _25043_ (.A(_06445_),
    .X(_06446_));
 sg13g2_nand2_2 _25044_ (.Y(_06447_),
    .A(_06415_),
    .B(_06446_));
 sg13g2_mux2_1 _25045_ (.A0(net855),
    .A1(\cpu.icache.r_data[0][20] ),
    .S(_06447_),
    .X(_02025_));
 sg13g2_mux2_1 _25046_ (.A0(net852),
    .A1(\cpu.icache.r_data[0][21] ),
    .S(_06447_),
    .X(_02026_));
 sg13g2_mux2_1 _25047_ (.A0(net854),
    .A1(\cpu.icache.r_data[0][22] ),
    .S(_06447_),
    .X(_02027_));
 sg13g2_mux2_1 _25048_ (.A0(net853),
    .A1(\cpu.icache.r_data[0][23] ),
    .S(_06447_),
    .X(_02028_));
 sg13g2_inv_1 _25049_ (.Y(_06448_),
    .A(\cpu.i_wstrobe_d ));
 sg13g2_nor3_2 _25050_ (.A(_00254_),
    .B(_06448_),
    .C(_06429_),
    .Y(_06449_));
 sg13g2_nand2_1 _25051_ (.Y(_06450_),
    .A(_06415_),
    .B(_06449_));
 sg13g2_buf_1 _25052_ (.A(_06450_),
    .X(_06451_));
 sg13g2_buf_1 _25053_ (.A(_06451_),
    .X(_06452_));
 sg13g2_mux2_1 _25054_ (.A0(net855),
    .A1(\cpu.icache.r_data[0][24] ),
    .S(net423),
    .X(_02029_));
 sg13g2_buf_1 _25055_ (.A(_06451_),
    .X(_06453_));
 sg13g2_mux2_1 _25056_ (.A0(_06438_),
    .A1(\cpu.icache.r_data[0][25] ),
    .S(net422),
    .X(_02030_));
 sg13g2_mux2_1 _25057_ (.A0(net854),
    .A1(\cpu.icache.r_data[0][26] ),
    .S(net422),
    .X(_02031_));
 sg13g2_mux2_1 _25058_ (.A0(_06432_),
    .A1(\cpu.icache.r_data[0][27] ),
    .S(net422),
    .X(_02032_));
 sg13g2_and2_1 _25059_ (.A(_06434_),
    .B(_06440_),
    .X(_06454_));
 sg13g2_buf_2 _25060_ (.A(_06454_),
    .X(_06455_));
 sg13g2_nand2_2 _25061_ (.Y(_06456_),
    .A(_06415_),
    .B(_06455_));
 sg13g2_mux2_1 _25062_ (.A0(_06413_),
    .A1(\cpu.icache.r_data[0][28] ),
    .S(_06456_),
    .X(_02033_));
 sg13g2_mux2_1 _25063_ (.A0(net852),
    .A1(\cpu.icache.r_data[0][29] ),
    .S(_06456_),
    .X(_02034_));
 sg13g2_mux2_1 _25064_ (.A0(net854),
    .A1(\cpu.icache.r_data[0][2] ),
    .S(_06425_),
    .X(_02035_));
 sg13g2_mux2_1 _25065_ (.A0(net854),
    .A1(\cpu.icache.r_data[0][30] ),
    .S(_06456_),
    .X(_02036_));
 sg13g2_mux2_1 _25066_ (.A0(_06432_),
    .A1(\cpu.icache.r_data[0][31] ),
    .S(_06456_),
    .X(_02037_));
 sg13g2_mux2_1 _25067_ (.A0(net853),
    .A1(\cpu.icache.r_data[0][3] ),
    .S(_06425_),
    .X(_02038_));
 sg13g2_and2_1 _25068_ (.A(_06418_),
    .B(_06444_),
    .X(_06457_));
 sg13g2_buf_2 _25069_ (.A(_06457_),
    .X(_06458_));
 sg13g2_nand2_2 _25070_ (.Y(_06459_),
    .A(_06415_),
    .B(_06458_));
 sg13g2_mux2_1 _25071_ (.A0(net855),
    .A1(\cpu.icache.r_data[0][4] ),
    .S(_06459_),
    .X(_02039_));
 sg13g2_mux2_1 _25072_ (.A0(net852),
    .A1(\cpu.icache.r_data[0][5] ),
    .S(_06459_),
    .X(_02040_));
 sg13g2_mux2_1 _25073_ (.A0(net854),
    .A1(\cpu.icache.r_data[0][6] ),
    .S(_06459_),
    .X(_02041_));
 sg13g2_mux2_1 _25074_ (.A0(net853),
    .A1(\cpu.icache.r_data[0][7] ),
    .S(_06459_),
    .X(_02042_));
 sg13g2_mux2_1 _25075_ (.A0(_06413_),
    .A1(\cpu.icache.r_data[0][8] ),
    .S(_06431_),
    .X(_02043_));
 sg13g2_mux2_1 _25076_ (.A0(_06438_),
    .A1(\cpu.icache.r_data[0][9] ),
    .S(_06431_),
    .X(_02044_));
 sg13g2_buf_1 _25077_ (.A(_02836_),
    .X(_06460_));
 sg13g2_nand2_1 _25078_ (.Y(_06461_),
    .A(_08562_),
    .B(_09061_));
 sg13g2_buf_4 _25079_ (.X(_06462_),
    .A(_06461_));
 sg13g2_nand2_2 _25080_ (.Y(_06463_),
    .A(_06418_),
    .B(_06422_));
 sg13g2_nor2_2 _25081_ (.A(_06462_),
    .B(_06463_),
    .Y(_06464_));
 sg13g2_mux2_1 _25082_ (.A0(\cpu.icache.r_data[1][0] ),
    .A1(net851),
    .S(_06464_),
    .X(_02045_));
 sg13g2_buf_1 _25083_ (.A(_02870_),
    .X(_06465_));
 sg13g2_or3_1 _25084_ (.A(_06416_),
    .B(_06427_),
    .C(_06429_),
    .X(_06466_));
 sg13g2_buf_2 _25085_ (.A(_06466_),
    .X(_06467_));
 sg13g2_nor2_2 _25086_ (.A(_06462_),
    .B(_06467_),
    .Y(_06468_));
 sg13g2_mux2_1 _25087_ (.A0(\cpu.icache.r_data[1][10] ),
    .A1(net850),
    .S(_06468_),
    .X(_02046_));
 sg13g2_buf_1 _25088_ (.A(_02874_),
    .X(_06469_));
 sg13g2_mux2_1 _25089_ (.A0(\cpu.icache.r_data[1][11] ),
    .A1(net849),
    .S(_06468_),
    .X(_02047_));
 sg13g2_buf_1 _25090_ (.A(_02836_),
    .X(_06470_));
 sg13g2_nand2_2 _25091_ (.Y(_06471_),
    .A(_06418_),
    .B(_06434_));
 sg13g2_nor2_2 _25092_ (.A(_06462_),
    .B(_06471_),
    .Y(_06472_));
 sg13g2_mux2_1 _25093_ (.A0(\cpu.icache.r_data[1][12] ),
    .A1(_06470_),
    .S(_06472_),
    .X(_02048_));
 sg13g2_buf_1 _25094_ (.A(_02866_),
    .X(_06473_));
 sg13g2_mux2_1 _25095_ (.A0(\cpu.icache.r_data[1][13] ),
    .A1(net847),
    .S(_06472_),
    .X(_02049_));
 sg13g2_buf_1 _25096_ (.A(_02870_),
    .X(_06474_));
 sg13g2_mux2_1 _25097_ (.A0(\cpu.icache.r_data[1][14] ),
    .A1(net846),
    .S(_06472_),
    .X(_02050_));
 sg13g2_buf_1 _25098_ (.A(_02874_),
    .X(_06475_));
 sg13g2_mux2_1 _25099_ (.A0(\cpu.icache.r_data[1][15] ),
    .A1(net845),
    .S(_06472_),
    .X(_02051_));
 sg13g2_nand2_2 _25100_ (.Y(_06476_),
    .A(_06422_),
    .B(_06440_));
 sg13g2_nor2_2 _25101_ (.A(_06462_),
    .B(_06476_),
    .Y(_06477_));
 sg13g2_mux2_1 _25102_ (.A0(\cpu.icache.r_data[1][16] ),
    .A1(net848),
    .S(_06477_),
    .X(_02052_));
 sg13g2_buf_1 _25103_ (.A(_02866_),
    .X(_06478_));
 sg13g2_mux2_1 _25104_ (.A0(\cpu.icache.r_data[1][17] ),
    .A1(net844),
    .S(_06477_),
    .X(_02053_));
 sg13g2_mux2_1 _25105_ (.A0(\cpu.icache.r_data[1][18] ),
    .A1(net846),
    .S(_06477_),
    .X(_02054_));
 sg13g2_mux2_1 _25106_ (.A0(\cpu.icache.r_data[1][19] ),
    .A1(net845),
    .S(_06477_),
    .X(_02055_));
 sg13g2_mux2_1 _25107_ (.A0(\cpu.icache.r_data[1][1] ),
    .A1(net844),
    .S(_06464_),
    .X(_02056_));
 sg13g2_nand2_2 _25108_ (.Y(_06479_),
    .A(_06440_),
    .B(_06444_));
 sg13g2_nor2_2 _25109_ (.A(_06462_),
    .B(_06479_),
    .Y(_06480_));
 sg13g2_mux2_1 _25110_ (.A0(\cpu.icache.r_data[1][20] ),
    .A1(net848),
    .S(_06480_),
    .X(_02057_));
 sg13g2_mux2_1 _25111_ (.A0(\cpu.icache.r_data[1][21] ),
    .A1(net844),
    .S(_06480_),
    .X(_02058_));
 sg13g2_mux2_1 _25112_ (.A0(\cpu.icache.r_data[1][22] ),
    .A1(net846),
    .S(_06480_),
    .X(_02059_));
 sg13g2_mux2_1 _25113_ (.A0(\cpu.icache.r_data[1][23] ),
    .A1(net845),
    .S(_06480_),
    .X(_02060_));
 sg13g2_nand4_1 _25114_ (.B(_06420_),
    .C(_06427_),
    .A(_06419_),
    .Y(_06481_),
    .D(\cpu.i_wstrobe_d ));
 sg13g2_buf_1 _25115_ (.A(_06481_),
    .X(_06482_));
 sg13g2_nor2_1 _25116_ (.A(_06462_),
    .B(_06482_),
    .Y(_06483_));
 sg13g2_buf_2 _25117_ (.A(_06483_),
    .X(_06484_));
 sg13g2_mux2_1 _25118_ (.A0(\cpu.icache.r_data[1][24] ),
    .A1(_06470_),
    .S(_06484_),
    .X(_02061_));
 sg13g2_mux2_1 _25119_ (.A0(\cpu.icache.r_data[1][25] ),
    .A1(net844),
    .S(_06484_),
    .X(_02062_));
 sg13g2_mux2_1 _25120_ (.A0(\cpu.icache.r_data[1][26] ),
    .A1(_06474_),
    .S(_06484_),
    .X(_02063_));
 sg13g2_mux2_1 _25121_ (.A0(\cpu.icache.r_data[1][27] ),
    .A1(net845),
    .S(_06484_),
    .X(_02064_));
 sg13g2_nand2_2 _25122_ (.Y(_06485_),
    .A(_06434_),
    .B(_06440_));
 sg13g2_nor2_2 _25123_ (.A(_06462_),
    .B(_06485_),
    .Y(_06486_));
 sg13g2_mux2_1 _25124_ (.A0(\cpu.icache.r_data[1][28] ),
    .A1(net848),
    .S(_06486_),
    .X(_02065_));
 sg13g2_mux2_1 _25125_ (.A0(\cpu.icache.r_data[1][29] ),
    .A1(net844),
    .S(_06486_),
    .X(_02066_));
 sg13g2_mux2_1 _25126_ (.A0(\cpu.icache.r_data[1][2] ),
    .A1(net846),
    .S(_06464_),
    .X(_02067_));
 sg13g2_mux2_1 _25127_ (.A0(\cpu.icache.r_data[1][30] ),
    .A1(net846),
    .S(_06486_),
    .X(_02068_));
 sg13g2_mux2_1 _25128_ (.A0(\cpu.icache.r_data[1][31] ),
    .A1(_06475_),
    .S(_06486_),
    .X(_02069_));
 sg13g2_mux2_1 _25129_ (.A0(\cpu.icache.r_data[1][3] ),
    .A1(net845),
    .S(_06464_),
    .X(_02070_));
 sg13g2_nand2_2 _25130_ (.Y(_06487_),
    .A(_06418_),
    .B(_06444_));
 sg13g2_nor2_2 _25131_ (.A(_06462_),
    .B(_06487_),
    .Y(_06488_));
 sg13g2_mux2_1 _25132_ (.A0(\cpu.icache.r_data[1][4] ),
    .A1(net848),
    .S(_06488_),
    .X(_02071_));
 sg13g2_mux2_1 _25133_ (.A0(\cpu.icache.r_data[1][5] ),
    .A1(_06478_),
    .S(_06488_),
    .X(_02072_));
 sg13g2_mux2_1 _25134_ (.A0(\cpu.icache.r_data[1][6] ),
    .A1(net846),
    .S(_06488_),
    .X(_02073_));
 sg13g2_mux2_1 _25135_ (.A0(\cpu.icache.r_data[1][7] ),
    .A1(net845),
    .S(_06488_),
    .X(_02074_));
 sg13g2_mux2_1 _25136_ (.A0(\cpu.icache.r_data[1][8] ),
    .A1(net848),
    .S(_06468_),
    .X(_02075_));
 sg13g2_mux2_1 _25137_ (.A0(\cpu.icache.r_data[1][9] ),
    .A1(net844),
    .S(_06468_),
    .X(_02076_));
 sg13g2_nand2_1 _25138_ (.Y(_06489_),
    .A(_08562_),
    .B(_08784_));
 sg13g2_buf_4 _25139_ (.X(_06490_),
    .A(_06489_));
 sg13g2_nor2_2 _25140_ (.A(_06490_),
    .B(_06463_),
    .Y(_06491_));
 sg13g2_mux2_1 _25141_ (.A0(\cpu.icache.r_data[2][0] ),
    .A1(net848),
    .S(_06491_),
    .X(_02077_));
 sg13g2_nor2_2 _25142_ (.A(_06490_),
    .B(_06467_),
    .Y(_06492_));
 sg13g2_mux2_1 _25143_ (.A0(\cpu.icache.r_data[2][10] ),
    .A1(net846),
    .S(_06492_),
    .X(_02078_));
 sg13g2_mux2_1 _25144_ (.A0(\cpu.icache.r_data[2][11] ),
    .A1(net845),
    .S(_06492_),
    .X(_02079_));
 sg13g2_nor2_2 _25145_ (.A(_06490_),
    .B(_06471_),
    .Y(_06493_));
 sg13g2_mux2_1 _25146_ (.A0(\cpu.icache.r_data[2][12] ),
    .A1(net848),
    .S(_06493_),
    .X(_02080_));
 sg13g2_mux2_1 _25147_ (.A0(\cpu.icache.r_data[2][13] ),
    .A1(_06478_),
    .S(_06493_),
    .X(_02081_));
 sg13g2_mux2_1 _25148_ (.A0(\cpu.icache.r_data[2][14] ),
    .A1(_06474_),
    .S(_06493_),
    .X(_02082_));
 sg13g2_mux2_1 _25149_ (.A0(\cpu.icache.r_data[2][15] ),
    .A1(_06475_),
    .S(_06493_),
    .X(_02083_));
 sg13g2_nor2_2 _25150_ (.A(_06490_),
    .B(_06476_),
    .Y(_06494_));
 sg13g2_mux2_1 _25151_ (.A0(\cpu.icache.r_data[2][16] ),
    .A1(net848),
    .S(_06494_),
    .X(_02084_));
 sg13g2_mux2_1 _25152_ (.A0(\cpu.icache.r_data[2][17] ),
    .A1(net844),
    .S(_06494_),
    .X(_02085_));
 sg13g2_mux2_1 _25153_ (.A0(\cpu.icache.r_data[2][18] ),
    .A1(net846),
    .S(_06494_),
    .X(_02086_));
 sg13g2_mux2_1 _25154_ (.A0(\cpu.icache.r_data[2][19] ),
    .A1(net845),
    .S(_06494_),
    .X(_02087_));
 sg13g2_mux2_1 _25155_ (.A0(\cpu.icache.r_data[2][1] ),
    .A1(net844),
    .S(_06491_),
    .X(_02088_));
 sg13g2_buf_1 _25156_ (.A(_02836_),
    .X(_06495_));
 sg13g2_nor2_2 _25157_ (.A(_06490_),
    .B(_06479_),
    .Y(_06496_));
 sg13g2_mux2_1 _25158_ (.A0(\cpu.icache.r_data[2][20] ),
    .A1(net843),
    .S(_06496_),
    .X(_02089_));
 sg13g2_buf_1 _25159_ (.A(_02866_),
    .X(_06497_));
 sg13g2_mux2_1 _25160_ (.A0(\cpu.icache.r_data[2][21] ),
    .A1(net842),
    .S(_06496_),
    .X(_02090_));
 sg13g2_buf_1 _25161_ (.A(_02870_),
    .X(_06498_));
 sg13g2_mux2_1 _25162_ (.A0(\cpu.icache.r_data[2][22] ),
    .A1(net841),
    .S(_06496_),
    .X(_02091_));
 sg13g2_buf_1 _25163_ (.A(_02874_),
    .X(_06499_));
 sg13g2_mux2_1 _25164_ (.A0(\cpu.icache.r_data[2][23] ),
    .A1(net840),
    .S(_06496_),
    .X(_02092_));
 sg13g2_nor2_1 _25165_ (.A(_06490_),
    .B(_06482_),
    .Y(_06500_));
 sg13g2_buf_2 _25166_ (.A(_06500_),
    .X(_06501_));
 sg13g2_mux2_1 _25167_ (.A0(\cpu.icache.r_data[2][24] ),
    .A1(net843),
    .S(_06501_),
    .X(_02093_));
 sg13g2_mux2_1 _25168_ (.A0(\cpu.icache.r_data[2][25] ),
    .A1(net842),
    .S(_06501_),
    .X(_02094_));
 sg13g2_mux2_1 _25169_ (.A0(\cpu.icache.r_data[2][26] ),
    .A1(net841),
    .S(_06501_),
    .X(_02095_));
 sg13g2_mux2_1 _25170_ (.A0(\cpu.icache.r_data[2][27] ),
    .A1(net840),
    .S(_06501_),
    .X(_02096_));
 sg13g2_nor2_2 _25171_ (.A(_06490_),
    .B(_06485_),
    .Y(_06502_));
 sg13g2_mux2_1 _25172_ (.A0(\cpu.icache.r_data[2][28] ),
    .A1(net843),
    .S(_06502_),
    .X(_02097_));
 sg13g2_mux2_1 _25173_ (.A0(\cpu.icache.r_data[2][29] ),
    .A1(net842),
    .S(_06502_),
    .X(_02098_));
 sg13g2_mux2_1 _25174_ (.A0(\cpu.icache.r_data[2][2] ),
    .A1(net841),
    .S(_06491_),
    .X(_02099_));
 sg13g2_mux2_1 _25175_ (.A0(\cpu.icache.r_data[2][30] ),
    .A1(net841),
    .S(_06502_),
    .X(_02100_));
 sg13g2_mux2_1 _25176_ (.A0(\cpu.icache.r_data[2][31] ),
    .A1(net840),
    .S(_06502_),
    .X(_02101_));
 sg13g2_mux2_1 _25177_ (.A0(\cpu.icache.r_data[2][3] ),
    .A1(_06499_),
    .S(_06491_),
    .X(_02102_));
 sg13g2_nor2_2 _25178_ (.A(_06490_),
    .B(_06487_),
    .Y(_06503_));
 sg13g2_mux2_1 _25179_ (.A0(\cpu.icache.r_data[2][4] ),
    .A1(net843),
    .S(_06503_),
    .X(_02103_));
 sg13g2_mux2_1 _25180_ (.A0(\cpu.icache.r_data[2][5] ),
    .A1(net842),
    .S(_06503_),
    .X(_02104_));
 sg13g2_mux2_1 _25181_ (.A0(\cpu.icache.r_data[2][6] ),
    .A1(net841),
    .S(_06503_),
    .X(_02105_));
 sg13g2_mux2_1 _25182_ (.A0(\cpu.icache.r_data[2][7] ),
    .A1(net840),
    .S(_06503_),
    .X(_02106_));
 sg13g2_mux2_1 _25183_ (.A0(\cpu.icache.r_data[2][8] ),
    .A1(_06495_),
    .S(_06492_),
    .X(_02107_));
 sg13g2_mux2_1 _25184_ (.A0(\cpu.icache.r_data[2][9] ),
    .A1(net842),
    .S(_06492_),
    .X(_02108_));
 sg13g2_nand2_2 _25185_ (.Y(_06504_),
    .A(net498),
    .B(_06424_));
 sg13g2_mux2_1 _25186_ (.A0(net855),
    .A1(\cpu.icache.r_data[3][0] ),
    .S(_06504_),
    .X(_02109_));
 sg13g2_and2_1 _25187_ (.A(_09000_),
    .B(_06430_),
    .X(_06505_));
 sg13g2_buf_1 _25188_ (.A(_06505_),
    .X(_06506_));
 sg13g2_mux2_1 _25189_ (.A0(\cpu.icache.r_data[3][10] ),
    .A1(_06498_),
    .S(_06506_),
    .X(_02110_));
 sg13g2_mux2_1 _25190_ (.A0(\cpu.icache.r_data[3][11] ),
    .A1(net840),
    .S(_06506_),
    .X(_02111_));
 sg13g2_nand2_2 _25191_ (.Y(_06507_),
    .A(net498),
    .B(_06436_));
 sg13g2_mux2_1 _25192_ (.A0(net855),
    .A1(\cpu.icache.r_data[3][12] ),
    .S(_06507_),
    .X(_02112_));
 sg13g2_mux2_1 _25193_ (.A0(net852),
    .A1(\cpu.icache.r_data[3][13] ),
    .S(_06507_),
    .X(_02113_));
 sg13g2_mux2_1 _25194_ (.A0(net854),
    .A1(\cpu.icache.r_data[3][14] ),
    .S(_06507_),
    .X(_02114_));
 sg13g2_mux2_1 _25195_ (.A0(net853),
    .A1(\cpu.icache.r_data[3][15] ),
    .S(_06507_),
    .X(_02115_));
 sg13g2_buf_1 _25196_ (.A(_02836_),
    .X(_06508_));
 sg13g2_nand2_2 _25197_ (.Y(_06509_),
    .A(net498),
    .B(_06442_));
 sg13g2_mux2_1 _25198_ (.A0(net839),
    .A1(\cpu.icache.r_data[3][16] ),
    .S(_06509_),
    .X(_02116_));
 sg13g2_mux2_1 _25199_ (.A0(net852),
    .A1(\cpu.icache.r_data[3][17] ),
    .S(_06509_),
    .X(_02117_));
 sg13g2_mux2_1 _25200_ (.A0(net854),
    .A1(\cpu.icache.r_data[3][18] ),
    .S(_06509_),
    .X(_02118_));
 sg13g2_mux2_1 _25201_ (.A0(net853),
    .A1(\cpu.icache.r_data[3][19] ),
    .S(_06509_),
    .X(_02119_));
 sg13g2_buf_1 _25202_ (.A(_02866_),
    .X(_06510_));
 sg13g2_mux2_1 _25203_ (.A0(net838),
    .A1(\cpu.icache.r_data[3][1] ),
    .S(_06504_),
    .X(_02120_));
 sg13g2_nand2_2 _25204_ (.Y(_06511_),
    .A(net498),
    .B(_06446_));
 sg13g2_mux2_1 _25205_ (.A0(net839),
    .A1(\cpu.icache.r_data[3][20] ),
    .S(_06511_),
    .X(_02121_));
 sg13g2_mux2_1 _25206_ (.A0(net838),
    .A1(\cpu.icache.r_data[3][21] ),
    .S(_06511_),
    .X(_02122_));
 sg13g2_buf_1 _25207_ (.A(_02870_),
    .X(_06512_));
 sg13g2_mux2_1 _25208_ (.A0(net837),
    .A1(\cpu.icache.r_data[3][22] ),
    .S(_06511_),
    .X(_02123_));
 sg13g2_buf_1 _25209_ (.A(_02874_),
    .X(_06513_));
 sg13g2_mux2_1 _25210_ (.A0(net836),
    .A1(\cpu.icache.r_data[3][23] ),
    .S(_06511_),
    .X(_02124_));
 sg13g2_nand2_1 _25211_ (.Y(_06514_),
    .A(_09000_),
    .B(_06449_));
 sg13g2_buf_1 _25212_ (.A(_06514_),
    .X(_06515_));
 sg13g2_buf_1 _25213_ (.A(_06515_),
    .X(_06516_));
 sg13g2_mux2_1 _25214_ (.A0(_06508_),
    .A1(\cpu.icache.r_data[3][24] ),
    .S(net289),
    .X(_02125_));
 sg13g2_buf_1 _25215_ (.A(_06515_),
    .X(_06517_));
 sg13g2_mux2_1 _25216_ (.A0(net838),
    .A1(\cpu.icache.r_data[3][25] ),
    .S(net288),
    .X(_02126_));
 sg13g2_mux2_1 _25217_ (.A0(_06512_),
    .A1(\cpu.icache.r_data[3][26] ),
    .S(net288),
    .X(_02127_));
 sg13g2_mux2_1 _25218_ (.A0(net836),
    .A1(\cpu.icache.r_data[3][27] ),
    .S(net288),
    .X(_02128_));
 sg13g2_nand2_2 _25219_ (.Y(_06518_),
    .A(net498),
    .B(_06455_));
 sg13g2_mux2_1 _25220_ (.A0(net839),
    .A1(\cpu.icache.r_data[3][28] ),
    .S(_06518_),
    .X(_02129_));
 sg13g2_mux2_1 _25221_ (.A0(net838),
    .A1(\cpu.icache.r_data[3][29] ),
    .S(_06518_),
    .X(_02130_));
 sg13g2_mux2_1 _25222_ (.A0(net837),
    .A1(\cpu.icache.r_data[3][2] ),
    .S(_06504_),
    .X(_02131_));
 sg13g2_mux2_1 _25223_ (.A0(net837),
    .A1(\cpu.icache.r_data[3][30] ),
    .S(_06518_),
    .X(_02132_));
 sg13g2_mux2_1 _25224_ (.A0(net836),
    .A1(\cpu.icache.r_data[3][31] ),
    .S(_06518_),
    .X(_02133_));
 sg13g2_mux2_1 _25225_ (.A0(_06513_),
    .A1(\cpu.icache.r_data[3][3] ),
    .S(_06504_),
    .X(_02134_));
 sg13g2_nand2_2 _25226_ (.Y(_06519_),
    .A(net498),
    .B(_06458_));
 sg13g2_mux2_1 _25227_ (.A0(net839),
    .A1(\cpu.icache.r_data[3][4] ),
    .S(_06519_),
    .X(_02135_));
 sg13g2_mux2_1 _25228_ (.A0(_06510_),
    .A1(\cpu.icache.r_data[3][5] ),
    .S(_06519_),
    .X(_02136_));
 sg13g2_mux2_1 _25229_ (.A0(net837),
    .A1(\cpu.icache.r_data[3][6] ),
    .S(_06519_),
    .X(_02137_));
 sg13g2_mux2_1 _25230_ (.A0(net836),
    .A1(\cpu.icache.r_data[3][7] ),
    .S(_06519_),
    .X(_02138_));
 sg13g2_mux2_1 _25231_ (.A0(\cpu.icache.r_data[3][8] ),
    .A1(_06495_),
    .S(_06506_),
    .X(_02139_));
 sg13g2_mux2_1 _25232_ (.A0(\cpu.icache.r_data[3][9] ),
    .A1(net842),
    .S(_06506_),
    .X(_02140_));
 sg13g2_nand2_2 _25233_ (.Y(_06520_),
    .A(net710),
    .B(_06424_));
 sg13g2_mux2_1 _25234_ (.A0(net839),
    .A1(\cpu.icache.r_data[4][0] ),
    .S(_06520_),
    .X(_02141_));
 sg13g2_and2_1 _25235_ (.A(net710),
    .B(_06430_),
    .X(_06521_));
 sg13g2_buf_1 _25236_ (.A(_06521_),
    .X(_06522_));
 sg13g2_mux2_1 _25237_ (.A0(\cpu.icache.r_data[4][10] ),
    .A1(net841),
    .S(_06522_),
    .X(_02142_));
 sg13g2_mux2_1 _25238_ (.A0(\cpu.icache.r_data[4][11] ),
    .A1(net840),
    .S(_06522_),
    .X(_02143_));
 sg13g2_nand2_2 _25239_ (.Y(_06523_),
    .A(net710),
    .B(_06436_));
 sg13g2_mux2_1 _25240_ (.A0(_06508_),
    .A1(\cpu.icache.r_data[4][12] ),
    .S(_06523_),
    .X(_02144_));
 sg13g2_mux2_1 _25241_ (.A0(net838),
    .A1(\cpu.icache.r_data[4][13] ),
    .S(_06523_),
    .X(_02145_));
 sg13g2_mux2_1 _25242_ (.A0(_06512_),
    .A1(\cpu.icache.r_data[4][14] ),
    .S(_06523_),
    .X(_02146_));
 sg13g2_mux2_1 _25243_ (.A0(net836),
    .A1(\cpu.icache.r_data[4][15] ),
    .S(_06523_),
    .X(_02147_));
 sg13g2_nand2_2 _25244_ (.Y(_06524_),
    .A(net710),
    .B(_06442_));
 sg13g2_mux2_1 _25245_ (.A0(net839),
    .A1(\cpu.icache.r_data[4][16] ),
    .S(_06524_),
    .X(_02148_));
 sg13g2_mux2_1 _25246_ (.A0(net838),
    .A1(\cpu.icache.r_data[4][17] ),
    .S(_06524_),
    .X(_02149_));
 sg13g2_mux2_1 _25247_ (.A0(net837),
    .A1(\cpu.icache.r_data[4][18] ),
    .S(_06524_),
    .X(_02150_));
 sg13g2_mux2_1 _25248_ (.A0(net836),
    .A1(\cpu.icache.r_data[4][19] ),
    .S(_06524_),
    .X(_02151_));
 sg13g2_mux2_1 _25249_ (.A0(net838),
    .A1(\cpu.icache.r_data[4][1] ),
    .S(_06520_),
    .X(_02152_));
 sg13g2_nand2_2 _25250_ (.Y(_06525_),
    .A(net710),
    .B(_06446_));
 sg13g2_mux2_1 _25251_ (.A0(net839),
    .A1(\cpu.icache.r_data[4][20] ),
    .S(_06525_),
    .X(_02153_));
 sg13g2_mux2_1 _25252_ (.A0(net838),
    .A1(\cpu.icache.r_data[4][21] ),
    .S(_06525_),
    .X(_02154_));
 sg13g2_mux2_1 _25253_ (.A0(net837),
    .A1(\cpu.icache.r_data[4][22] ),
    .S(_06525_),
    .X(_02155_));
 sg13g2_mux2_1 _25254_ (.A0(net836),
    .A1(\cpu.icache.r_data[4][23] ),
    .S(_06525_),
    .X(_02156_));
 sg13g2_and2_1 _25255_ (.A(_09007_),
    .B(_06449_),
    .X(_06526_));
 sg13g2_buf_2 _25256_ (.A(_06526_),
    .X(_06527_));
 sg13g2_mux2_1 _25257_ (.A0(\cpu.icache.r_data[4][24] ),
    .A1(net843),
    .S(_06527_),
    .X(_02157_));
 sg13g2_mux2_1 _25258_ (.A0(\cpu.icache.r_data[4][25] ),
    .A1(_06497_),
    .S(_06527_),
    .X(_02158_));
 sg13g2_mux2_1 _25259_ (.A0(\cpu.icache.r_data[4][26] ),
    .A1(net841),
    .S(_06527_),
    .X(_02159_));
 sg13g2_mux2_1 _25260_ (.A0(\cpu.icache.r_data[4][27] ),
    .A1(_06499_),
    .S(_06527_),
    .X(_02160_));
 sg13g2_nand2_2 _25261_ (.Y(_06528_),
    .A(net710),
    .B(_06455_));
 sg13g2_mux2_1 _25262_ (.A0(net839),
    .A1(\cpu.icache.r_data[4][28] ),
    .S(_06528_),
    .X(_02161_));
 sg13g2_mux2_1 _25263_ (.A0(_06510_),
    .A1(\cpu.icache.r_data[4][29] ),
    .S(_06528_),
    .X(_02162_));
 sg13g2_mux2_1 _25264_ (.A0(net837),
    .A1(\cpu.icache.r_data[4][2] ),
    .S(_06520_),
    .X(_02163_));
 sg13g2_mux2_1 _25265_ (.A0(net837),
    .A1(\cpu.icache.r_data[4][30] ),
    .S(_06528_),
    .X(_02164_));
 sg13g2_mux2_1 _25266_ (.A0(net836),
    .A1(\cpu.icache.r_data[4][31] ),
    .S(_06528_),
    .X(_02165_));
 sg13g2_mux2_1 _25267_ (.A0(_06513_),
    .A1(\cpu.icache.r_data[4][3] ),
    .S(_06520_),
    .X(_02166_));
 sg13g2_nand2_2 _25268_ (.Y(_06529_),
    .A(net710),
    .B(_06458_));
 sg13g2_mux2_1 _25269_ (.A0(_06460_),
    .A1(\cpu.icache.r_data[4][4] ),
    .S(_06529_),
    .X(_02167_));
 sg13g2_mux2_1 _25270_ (.A0(_06473_),
    .A1(\cpu.icache.r_data[4][5] ),
    .S(_06529_),
    .X(_02168_));
 sg13g2_mux2_1 _25271_ (.A0(net850),
    .A1(\cpu.icache.r_data[4][6] ),
    .S(_06529_),
    .X(_02169_));
 sg13g2_mux2_1 _25272_ (.A0(_06469_),
    .A1(\cpu.icache.r_data[4][7] ),
    .S(_06529_),
    .X(_02170_));
 sg13g2_mux2_1 _25273_ (.A0(\cpu.icache.r_data[4][8] ),
    .A1(net843),
    .S(_06522_),
    .X(_02171_));
 sg13g2_mux2_1 _25274_ (.A0(\cpu.icache.r_data[4][9] ),
    .A1(_06497_),
    .S(_06522_),
    .X(_02172_));
 sg13g2_nand2_2 _25275_ (.Y(_06530_),
    .A(net552),
    .B(_06424_));
 sg13g2_mux2_1 _25276_ (.A0(net851),
    .A1(\cpu.icache.r_data[5][0] ),
    .S(_06530_),
    .X(_02173_));
 sg13g2_nand2_2 _25277_ (.Y(_06531_),
    .A(net552),
    .B(_06430_));
 sg13g2_mux2_1 _25278_ (.A0(net850),
    .A1(\cpu.icache.r_data[5][10] ),
    .S(_06531_),
    .X(_02174_));
 sg13g2_mux2_1 _25279_ (.A0(net849),
    .A1(\cpu.icache.r_data[5][11] ),
    .S(_06531_),
    .X(_02175_));
 sg13g2_nand2_2 _25280_ (.Y(_06532_),
    .A(net552),
    .B(_06436_));
 sg13g2_mux2_1 _25281_ (.A0(net851),
    .A1(\cpu.icache.r_data[5][12] ),
    .S(_06532_),
    .X(_02176_));
 sg13g2_mux2_1 _25282_ (.A0(net847),
    .A1(\cpu.icache.r_data[5][13] ),
    .S(_06532_),
    .X(_02177_));
 sg13g2_mux2_1 _25283_ (.A0(_06465_),
    .A1(\cpu.icache.r_data[5][14] ),
    .S(_06532_),
    .X(_02178_));
 sg13g2_mux2_1 _25284_ (.A0(net849),
    .A1(\cpu.icache.r_data[5][15] ),
    .S(_06532_),
    .X(_02179_));
 sg13g2_nand2_2 _25285_ (.Y(_06533_),
    .A(net552),
    .B(_06442_));
 sg13g2_mux2_1 _25286_ (.A0(net851),
    .A1(\cpu.icache.r_data[5][16] ),
    .S(_06533_),
    .X(_02180_));
 sg13g2_mux2_1 _25287_ (.A0(net847),
    .A1(\cpu.icache.r_data[5][17] ),
    .S(_06533_),
    .X(_02181_));
 sg13g2_mux2_1 _25288_ (.A0(net850),
    .A1(\cpu.icache.r_data[5][18] ),
    .S(_06533_),
    .X(_02182_));
 sg13g2_mux2_1 _25289_ (.A0(net849),
    .A1(\cpu.icache.r_data[5][19] ),
    .S(_06533_),
    .X(_02183_));
 sg13g2_mux2_1 _25290_ (.A0(net847),
    .A1(\cpu.icache.r_data[5][1] ),
    .S(_06530_),
    .X(_02184_));
 sg13g2_nand2_2 _25291_ (.Y(_06534_),
    .A(net552),
    .B(_06446_));
 sg13g2_mux2_1 _25292_ (.A0(net851),
    .A1(\cpu.icache.r_data[5][20] ),
    .S(_06534_),
    .X(_02185_));
 sg13g2_mux2_1 _25293_ (.A0(net847),
    .A1(\cpu.icache.r_data[5][21] ),
    .S(_06534_),
    .X(_02186_));
 sg13g2_mux2_1 _25294_ (.A0(net850),
    .A1(\cpu.icache.r_data[5][22] ),
    .S(_06534_),
    .X(_02187_));
 sg13g2_mux2_1 _25295_ (.A0(net849),
    .A1(\cpu.icache.r_data[5][23] ),
    .S(_06534_),
    .X(_02188_));
 sg13g2_nand2_1 _25296_ (.Y(_06535_),
    .A(_08992_),
    .B(_06449_));
 sg13g2_buf_2 _25297_ (.A(_06535_),
    .X(_06536_));
 sg13g2_mux2_1 _25298_ (.A0(net851),
    .A1(\cpu.icache.r_data[5][24] ),
    .S(_06536_),
    .X(_02189_));
 sg13g2_mux2_1 _25299_ (.A0(net847),
    .A1(\cpu.icache.r_data[5][25] ),
    .S(_06536_),
    .X(_02190_));
 sg13g2_mux2_1 _25300_ (.A0(net850),
    .A1(\cpu.icache.r_data[5][26] ),
    .S(_06536_),
    .X(_02191_));
 sg13g2_mux2_1 _25301_ (.A0(net849),
    .A1(\cpu.icache.r_data[5][27] ),
    .S(_06536_),
    .X(_02192_));
 sg13g2_nand2_2 _25302_ (.Y(_06537_),
    .A(net552),
    .B(_06455_));
 sg13g2_mux2_1 _25303_ (.A0(net851),
    .A1(\cpu.icache.r_data[5][28] ),
    .S(_06537_),
    .X(_02193_));
 sg13g2_mux2_1 _25304_ (.A0(net847),
    .A1(\cpu.icache.r_data[5][29] ),
    .S(_06537_),
    .X(_02194_));
 sg13g2_mux2_1 _25305_ (.A0(net850),
    .A1(\cpu.icache.r_data[5][2] ),
    .S(_06530_),
    .X(_02195_));
 sg13g2_mux2_1 _25306_ (.A0(net850),
    .A1(\cpu.icache.r_data[5][30] ),
    .S(_06537_),
    .X(_02196_));
 sg13g2_mux2_1 _25307_ (.A0(net849),
    .A1(\cpu.icache.r_data[5][31] ),
    .S(_06537_),
    .X(_02197_));
 sg13g2_mux2_1 _25308_ (.A0(net849),
    .A1(\cpu.icache.r_data[5][3] ),
    .S(_06530_),
    .X(_02198_));
 sg13g2_nand2_2 _25309_ (.Y(_06538_),
    .A(net552),
    .B(_06458_));
 sg13g2_mux2_1 _25310_ (.A0(_06460_),
    .A1(\cpu.icache.r_data[5][4] ),
    .S(_06538_),
    .X(_02199_));
 sg13g2_mux2_1 _25311_ (.A0(_06473_),
    .A1(\cpu.icache.r_data[5][5] ),
    .S(_06538_),
    .X(_02200_));
 sg13g2_mux2_1 _25312_ (.A0(_06465_),
    .A1(\cpu.icache.r_data[5][6] ),
    .S(_06538_),
    .X(_02201_));
 sg13g2_mux2_1 _25313_ (.A0(_06469_),
    .A1(\cpu.icache.r_data[5][7] ),
    .S(_06538_),
    .X(_02202_));
 sg13g2_mux2_1 _25314_ (.A0(net851),
    .A1(\cpu.icache.r_data[5][8] ),
    .S(_06531_),
    .X(_02203_));
 sg13g2_mux2_1 _25315_ (.A0(net847),
    .A1(\cpu.icache.r_data[5][9] ),
    .S(_06531_),
    .X(_02204_));
 sg13g2_nand2_1 _25316_ (.Y(_06539_),
    .A(net808),
    .B(_08784_));
 sg13g2_buf_4 _25317_ (.X(_06540_),
    .A(_06539_));
 sg13g2_nor2_2 _25318_ (.A(_06540_),
    .B(_06463_),
    .Y(_06541_));
 sg13g2_mux2_1 _25319_ (.A0(\cpu.icache.r_data[6][0] ),
    .A1(net843),
    .S(_06541_),
    .X(_02205_));
 sg13g2_nor2_2 _25320_ (.A(_06540_),
    .B(_06467_),
    .Y(_06542_));
 sg13g2_mux2_1 _25321_ (.A0(\cpu.icache.r_data[6][10] ),
    .A1(net841),
    .S(_06542_),
    .X(_02206_));
 sg13g2_mux2_1 _25322_ (.A0(\cpu.icache.r_data[6][11] ),
    .A1(net840),
    .S(_06542_),
    .X(_02207_));
 sg13g2_nor2_2 _25323_ (.A(_06540_),
    .B(_06471_),
    .Y(_06543_));
 sg13g2_mux2_1 _25324_ (.A0(\cpu.icache.r_data[6][12] ),
    .A1(net843),
    .S(_06543_),
    .X(_02208_));
 sg13g2_mux2_1 _25325_ (.A0(\cpu.icache.r_data[6][13] ),
    .A1(net842),
    .S(_06543_),
    .X(_02209_));
 sg13g2_mux2_1 _25326_ (.A0(\cpu.icache.r_data[6][14] ),
    .A1(_06498_),
    .S(_06543_),
    .X(_02210_));
 sg13g2_mux2_1 _25327_ (.A0(\cpu.icache.r_data[6][15] ),
    .A1(net840),
    .S(_06543_),
    .X(_02211_));
 sg13g2_buf_1 _25328_ (.A(_02836_),
    .X(_06544_));
 sg13g2_nor2_2 _25329_ (.A(_06540_),
    .B(_06476_),
    .Y(_06545_));
 sg13g2_mux2_1 _25330_ (.A0(\cpu.icache.r_data[6][16] ),
    .A1(net835),
    .S(_06545_),
    .X(_02212_));
 sg13g2_mux2_1 _25331_ (.A0(\cpu.icache.r_data[6][17] ),
    .A1(net842),
    .S(_06545_),
    .X(_02213_));
 sg13g2_buf_1 _25332_ (.A(_02870_),
    .X(_06546_));
 sg13g2_mux2_1 _25333_ (.A0(\cpu.icache.r_data[6][18] ),
    .A1(net834),
    .S(_06545_),
    .X(_02214_));
 sg13g2_buf_1 _25334_ (.A(_02874_),
    .X(_06547_));
 sg13g2_mux2_1 _25335_ (.A0(\cpu.icache.r_data[6][19] ),
    .A1(net833),
    .S(_06545_),
    .X(_02215_));
 sg13g2_buf_1 _25336_ (.A(_02866_),
    .X(_06548_));
 sg13g2_mux2_1 _25337_ (.A0(\cpu.icache.r_data[6][1] ),
    .A1(net832),
    .S(_06541_),
    .X(_02216_));
 sg13g2_nor2_2 _25338_ (.A(_06540_),
    .B(_06479_),
    .Y(_06549_));
 sg13g2_mux2_1 _25339_ (.A0(\cpu.icache.r_data[6][20] ),
    .A1(net835),
    .S(_06549_),
    .X(_02217_));
 sg13g2_mux2_1 _25340_ (.A0(\cpu.icache.r_data[6][21] ),
    .A1(net832),
    .S(_06549_),
    .X(_02218_));
 sg13g2_mux2_1 _25341_ (.A0(\cpu.icache.r_data[6][22] ),
    .A1(net834),
    .S(_06549_),
    .X(_02219_));
 sg13g2_mux2_1 _25342_ (.A0(\cpu.icache.r_data[6][23] ),
    .A1(net833),
    .S(_06549_),
    .X(_02220_));
 sg13g2_nor2_1 _25343_ (.A(_06540_),
    .B(_06482_),
    .Y(_06550_));
 sg13g2_buf_2 _25344_ (.A(_06550_),
    .X(_06551_));
 sg13g2_mux2_1 _25345_ (.A0(\cpu.icache.r_data[6][24] ),
    .A1(net835),
    .S(_06551_),
    .X(_02221_));
 sg13g2_mux2_1 _25346_ (.A0(\cpu.icache.r_data[6][25] ),
    .A1(net832),
    .S(_06551_),
    .X(_02222_));
 sg13g2_mux2_1 _25347_ (.A0(\cpu.icache.r_data[6][26] ),
    .A1(net834),
    .S(_06551_),
    .X(_02223_));
 sg13g2_mux2_1 _25348_ (.A0(\cpu.icache.r_data[6][27] ),
    .A1(net833),
    .S(_06551_),
    .X(_02224_));
 sg13g2_nor2_2 _25349_ (.A(_06540_),
    .B(_06485_),
    .Y(_06552_));
 sg13g2_mux2_1 _25350_ (.A0(\cpu.icache.r_data[6][28] ),
    .A1(net835),
    .S(_06552_),
    .X(_02225_));
 sg13g2_mux2_1 _25351_ (.A0(\cpu.icache.r_data[6][29] ),
    .A1(net832),
    .S(_06552_),
    .X(_02226_));
 sg13g2_mux2_1 _25352_ (.A0(\cpu.icache.r_data[6][2] ),
    .A1(net834),
    .S(_06541_),
    .X(_02227_));
 sg13g2_mux2_1 _25353_ (.A0(\cpu.icache.r_data[6][30] ),
    .A1(net834),
    .S(_06552_),
    .X(_02228_));
 sg13g2_mux2_1 _25354_ (.A0(\cpu.icache.r_data[6][31] ),
    .A1(net833),
    .S(_06552_),
    .X(_02229_));
 sg13g2_mux2_1 _25355_ (.A0(\cpu.icache.r_data[6][3] ),
    .A1(net833),
    .S(_06541_),
    .X(_02230_));
 sg13g2_nor2_2 _25356_ (.A(_06540_),
    .B(_06487_),
    .Y(_06553_));
 sg13g2_mux2_1 _25357_ (.A0(\cpu.icache.r_data[6][4] ),
    .A1(net835),
    .S(_06553_),
    .X(_02231_));
 sg13g2_mux2_1 _25358_ (.A0(\cpu.icache.r_data[6][5] ),
    .A1(_06548_),
    .S(_06553_),
    .X(_02232_));
 sg13g2_mux2_1 _25359_ (.A0(\cpu.icache.r_data[6][6] ),
    .A1(net834),
    .S(_06553_),
    .X(_02233_));
 sg13g2_mux2_1 _25360_ (.A0(\cpu.icache.r_data[6][7] ),
    .A1(net833),
    .S(_06553_),
    .X(_02234_));
 sg13g2_mux2_1 _25361_ (.A0(\cpu.icache.r_data[6][8] ),
    .A1(_06544_),
    .S(_06542_),
    .X(_02235_));
 sg13g2_mux2_1 _25362_ (.A0(\cpu.icache.r_data[6][9] ),
    .A1(net832),
    .S(_06542_),
    .X(_02236_));
 sg13g2_nand2_1 _25363_ (.Y(_06554_),
    .A(net808),
    .B(net637));
 sg13g2_buf_4 _25364_ (.X(_06555_),
    .A(_06554_));
 sg13g2_nor2_2 _25365_ (.A(_06555_),
    .B(_06463_),
    .Y(_06556_));
 sg13g2_mux2_1 _25366_ (.A0(\cpu.icache.r_data[7][0] ),
    .A1(net835),
    .S(_06556_),
    .X(_02237_));
 sg13g2_nor2_2 _25367_ (.A(_06555_),
    .B(_06467_),
    .Y(_06557_));
 sg13g2_mux2_1 _25368_ (.A0(\cpu.icache.r_data[7][10] ),
    .A1(_06546_),
    .S(_06557_),
    .X(_02238_));
 sg13g2_mux2_1 _25369_ (.A0(\cpu.icache.r_data[7][11] ),
    .A1(_06547_),
    .S(_06557_),
    .X(_02239_));
 sg13g2_nor2_2 _25370_ (.A(_06555_),
    .B(_06471_),
    .Y(_06558_));
 sg13g2_mux2_1 _25371_ (.A0(\cpu.icache.r_data[7][12] ),
    .A1(_06544_),
    .S(_06558_),
    .X(_02240_));
 sg13g2_mux2_1 _25372_ (.A0(\cpu.icache.r_data[7][13] ),
    .A1(_06548_),
    .S(_06558_),
    .X(_02241_));
 sg13g2_mux2_1 _25373_ (.A0(\cpu.icache.r_data[7][14] ),
    .A1(_06546_),
    .S(_06558_),
    .X(_02242_));
 sg13g2_mux2_1 _25374_ (.A0(\cpu.icache.r_data[7][15] ),
    .A1(_06547_),
    .S(_06558_),
    .X(_02243_));
 sg13g2_nor2_2 _25375_ (.A(_06555_),
    .B(_06476_),
    .Y(_06559_));
 sg13g2_mux2_1 _25376_ (.A0(\cpu.icache.r_data[7][16] ),
    .A1(net835),
    .S(_06559_),
    .X(_02244_));
 sg13g2_mux2_1 _25377_ (.A0(\cpu.icache.r_data[7][17] ),
    .A1(net832),
    .S(_06559_),
    .X(_02245_));
 sg13g2_mux2_1 _25378_ (.A0(\cpu.icache.r_data[7][18] ),
    .A1(net834),
    .S(_06559_),
    .X(_02246_));
 sg13g2_mux2_1 _25379_ (.A0(\cpu.icache.r_data[7][19] ),
    .A1(net833),
    .S(_06559_),
    .X(_02247_));
 sg13g2_mux2_1 _25380_ (.A0(\cpu.icache.r_data[7][1] ),
    .A1(net832),
    .S(_06556_),
    .X(_02248_));
 sg13g2_nor2_2 _25381_ (.A(_06555_),
    .B(_06479_),
    .Y(_06560_));
 sg13g2_mux2_1 _25382_ (.A0(\cpu.icache.r_data[7][20] ),
    .A1(net835),
    .S(_06560_),
    .X(_02249_));
 sg13g2_mux2_1 _25383_ (.A0(\cpu.icache.r_data[7][21] ),
    .A1(net832),
    .S(_06560_),
    .X(_02250_));
 sg13g2_mux2_1 _25384_ (.A0(\cpu.icache.r_data[7][22] ),
    .A1(net834),
    .S(_06560_),
    .X(_02251_));
 sg13g2_mux2_1 _25385_ (.A0(\cpu.icache.r_data[7][23] ),
    .A1(net833),
    .S(_06560_),
    .X(_02252_));
 sg13g2_nor2_1 _25386_ (.A(_06555_),
    .B(_06482_),
    .Y(_06561_));
 sg13g2_buf_2 _25387_ (.A(_06561_),
    .X(_06562_));
 sg13g2_mux2_1 _25388_ (.A0(\cpu.icache.r_data[7][24] ),
    .A1(net1010),
    .S(_06562_),
    .X(_02253_));
 sg13g2_mux2_1 _25389_ (.A0(\cpu.icache.r_data[7][25] ),
    .A1(net1006),
    .S(_06562_),
    .X(_02254_));
 sg13g2_mux2_1 _25390_ (.A0(\cpu.icache.r_data[7][26] ),
    .A1(net1005),
    .S(_06562_),
    .X(_02255_));
 sg13g2_mux2_1 _25391_ (.A0(\cpu.icache.r_data[7][27] ),
    .A1(net1004),
    .S(_06562_),
    .X(_02256_));
 sg13g2_nor2_2 _25392_ (.A(_06555_),
    .B(_06485_),
    .Y(_06563_));
 sg13g2_mux2_1 _25393_ (.A0(\cpu.icache.r_data[7][28] ),
    .A1(net1010),
    .S(_06563_),
    .X(_02257_));
 sg13g2_mux2_1 _25394_ (.A0(\cpu.icache.r_data[7][29] ),
    .A1(net1006),
    .S(_06563_),
    .X(_02258_));
 sg13g2_mux2_1 _25395_ (.A0(\cpu.icache.r_data[7][2] ),
    .A1(net1005),
    .S(_06556_),
    .X(_02259_));
 sg13g2_mux2_1 _25396_ (.A0(\cpu.icache.r_data[7][30] ),
    .A1(_12223_),
    .S(_06563_),
    .X(_02260_));
 sg13g2_mux2_1 _25397_ (.A0(\cpu.icache.r_data[7][31] ),
    .A1(net1004),
    .S(_06563_),
    .X(_02261_));
 sg13g2_mux2_1 _25398_ (.A0(\cpu.icache.r_data[7][3] ),
    .A1(_12229_),
    .S(_06556_),
    .X(_02262_));
 sg13g2_nor2_2 _25399_ (.A(_06555_),
    .B(_06487_),
    .Y(_06564_));
 sg13g2_mux2_1 _25400_ (.A0(\cpu.icache.r_data[7][4] ),
    .A1(_12127_),
    .S(_06564_),
    .X(_02263_));
 sg13g2_mux2_1 _25401_ (.A0(\cpu.icache.r_data[7][5] ),
    .A1(_12218_),
    .S(_06564_),
    .X(_02264_));
 sg13g2_mux2_1 _25402_ (.A0(\cpu.icache.r_data[7][6] ),
    .A1(_12223_),
    .S(_06564_),
    .X(_02265_));
 sg13g2_mux2_1 _25403_ (.A0(\cpu.icache.r_data[7][7] ),
    .A1(_12229_),
    .S(_06564_),
    .X(_02266_));
 sg13g2_mux2_1 _25404_ (.A0(\cpu.icache.r_data[7][8] ),
    .A1(_12127_),
    .S(_06557_),
    .X(_02267_));
 sg13g2_mux2_1 _25405_ (.A0(\cpu.icache.r_data[7][9] ),
    .A1(_12218_),
    .S(_06557_),
    .X(_02268_));
 sg13g2_buf_1 _25406_ (.A(_06451_),
    .X(_06565_));
 sg13g2_nand2_1 _25407_ (.Y(_06566_),
    .A(\cpu.icache.r_tag[0][5] ),
    .B(net422));
 sg13g2_o21ai_1 _25408_ (.B1(_06566_),
    .Y(_02272_),
    .A1(net938),
    .A2(net421));
 sg13g2_nand2_1 _25409_ (.Y(_06567_),
    .A(\cpu.icache.r_tag[0][15] ),
    .B(net422));
 sg13g2_o21ai_1 _25410_ (.B1(_06567_),
    .Y(_02273_),
    .A1(net450),
    .A2(net421));
 sg13g2_nand2_1 _25411_ (.Y(_06568_),
    .A(\cpu.icache.r_tag[0][16] ),
    .B(net422));
 sg13g2_o21ai_1 _25412_ (.B1(_06568_),
    .Y(_02274_),
    .A1(net451),
    .A2(net421));
 sg13g2_nand2_1 _25413_ (.Y(_06569_),
    .A(\cpu.icache.r_tag[0][17] ),
    .B(net422));
 sg13g2_o21ai_1 _25414_ (.B1(_06569_),
    .Y(_02275_),
    .A1(_08918_),
    .A2(net421));
 sg13g2_nand2_1 _25415_ (.Y(_06570_),
    .A(\cpu.icache.r_tag[0][18] ),
    .B(_06453_));
 sg13g2_o21ai_1 _25416_ (.B1(_06570_),
    .Y(_02276_),
    .A1(net414),
    .A2(net421));
 sg13g2_nand2_1 _25417_ (.Y(_06571_),
    .A(\cpu.icache.r_tag[0][19] ),
    .B(net422));
 sg13g2_o21ai_1 _25418_ (.B1(_06571_),
    .Y(_02277_),
    .A1(net448),
    .A2(net421));
 sg13g2_buf_1 _25419_ (.A(_06451_),
    .X(_06572_));
 sg13g2_nand2_1 _25420_ (.Y(_06573_),
    .A(\cpu.icache.r_tag[0][20] ),
    .B(net420));
 sg13g2_o21ai_1 _25421_ (.B1(_06573_),
    .Y(_02278_),
    .A1(net412),
    .A2(net421));
 sg13g2_nand2_1 _25422_ (.Y(_06574_),
    .A(\cpu.icache.r_tag[0][21] ),
    .B(net420));
 sg13g2_o21ai_1 _25423_ (.B1(_06574_),
    .Y(_02279_),
    .A1(net411),
    .A2(_06565_));
 sg13g2_nand2_1 _25424_ (.Y(_06575_),
    .A(\cpu.icache.r_tag[0][22] ),
    .B(net420));
 sg13g2_o21ai_1 _25425_ (.B1(_06575_),
    .Y(_02280_),
    .A1(net449),
    .A2(_06565_));
 sg13g2_nand2_1 _25426_ (.Y(_06576_),
    .A(\cpu.icache.r_tag[0][23] ),
    .B(net420));
 sg13g2_o21ai_1 _25427_ (.B1(_06576_),
    .Y(_02281_),
    .A1(net500),
    .A2(net423));
 sg13g2_nand2_1 _25428_ (.Y(_06577_),
    .A(\cpu.icache.r_tag[0][6] ),
    .B(net420));
 sg13g2_o21ai_1 _25429_ (.B1(_06577_),
    .Y(_02282_),
    .A1(net980),
    .A2(net423));
 sg13g2_nand2_1 _25430_ (.Y(_06578_),
    .A(\cpu.icache.r_tag[0][7] ),
    .B(net420));
 sg13g2_o21ai_1 _25431_ (.B1(_06578_),
    .Y(_02283_),
    .A1(net939),
    .A2(net423));
 sg13g2_nand2_1 _25432_ (.Y(_06579_),
    .A(\cpu.icache.r_tag[0][8] ),
    .B(_06572_));
 sg13g2_o21ai_1 _25433_ (.B1(_06579_),
    .Y(_02284_),
    .A1(net940),
    .A2(net423));
 sg13g2_nand2_1 _25434_ (.Y(_06580_),
    .A(\cpu.icache.r_tag[0][9] ),
    .B(net420));
 sg13g2_o21ai_1 _25435_ (.B1(_06580_),
    .Y(_02285_),
    .A1(net974),
    .A2(net423));
 sg13g2_mux2_1 _25436_ (.A0(net978),
    .A1(\cpu.icache.r_tag[0][10] ),
    .S(_06453_),
    .X(_02286_));
 sg13g2_nand2_1 _25437_ (.Y(_06581_),
    .A(\cpu.icache.r_tag[0][11] ),
    .B(net420));
 sg13g2_o21ai_1 _25438_ (.B1(_06581_),
    .Y(_02287_),
    .A1(net979),
    .A2(net423));
 sg13g2_nand2_1 _25439_ (.Y(_06582_),
    .A(\cpu.icache.r_tag[0][12] ),
    .B(_06572_));
 sg13g2_o21ai_1 _25440_ (.B1(_06582_),
    .Y(_02288_),
    .A1(net349),
    .A2(net423));
 sg13g2_nand2_1 _25441_ (.Y(_06583_),
    .A(\cpu.icache.r_tag[0][13] ),
    .B(_06451_));
 sg13g2_o21ai_1 _25442_ (.B1(_06583_),
    .Y(_02289_),
    .A1(net415),
    .A2(_06452_));
 sg13g2_nand2_1 _25443_ (.Y(_06584_),
    .A(\cpu.icache.r_tag[0][14] ),
    .B(_06451_));
 sg13g2_o21ai_1 _25444_ (.B1(_06584_),
    .Y(_02290_),
    .A1(net410),
    .A2(_06452_));
 sg13g2_nor2b_1 _25445_ (.A(_06429_),
    .B_N(_06440_),
    .Y(_06585_));
 sg13g2_buf_1 _25446_ (.A(_06585_),
    .X(_06586_));
 sg13g2_nand2_1 _25447_ (.Y(_06587_),
    .A(_08591_),
    .B(_06586_));
 sg13g2_buf_1 _25448_ (.A(_06587_),
    .X(_06588_));
 sg13g2_buf_1 _25449_ (.A(net359),
    .X(_06589_));
 sg13g2_buf_1 _25450_ (.A(net359),
    .X(_06590_));
 sg13g2_nand2_1 _25451_ (.Y(_06591_),
    .A(\cpu.icache.r_tag[1][5] ),
    .B(net286));
 sg13g2_o21ai_1 _25452_ (.B1(_06591_),
    .Y(_02291_),
    .A1(net938),
    .A2(net287));
 sg13g2_buf_1 _25453_ (.A(_06588_),
    .X(_06592_));
 sg13g2_nand2_1 _25454_ (.Y(_06593_),
    .A(\cpu.icache.r_tag[1][15] ),
    .B(net285));
 sg13g2_o21ai_1 _25455_ (.B1(_06593_),
    .Y(_02292_),
    .A1(net450),
    .A2(net287));
 sg13g2_nand2_1 _25456_ (.Y(_06594_),
    .A(\cpu.icache.r_tag[1][16] ),
    .B(net285));
 sg13g2_o21ai_1 _25457_ (.B1(_06594_),
    .Y(_02293_),
    .A1(net451),
    .A2(net287));
 sg13g2_nand2_1 _25458_ (.Y(_06595_),
    .A(\cpu.icache.r_tag[1][17] ),
    .B(net285));
 sg13g2_o21ai_1 _25459_ (.B1(_06595_),
    .Y(_02294_),
    .A1(net413),
    .A2(net287));
 sg13g2_nand2_1 _25460_ (.Y(_06596_),
    .A(\cpu.icache.r_tag[1][18] ),
    .B(net285));
 sg13g2_o21ai_1 _25461_ (.B1(_06596_),
    .Y(_02295_),
    .A1(_08728_),
    .A2(net287));
 sg13g2_nand2_1 _25462_ (.Y(_06597_),
    .A(\cpu.icache.r_tag[1][19] ),
    .B(net285));
 sg13g2_o21ai_1 _25463_ (.B1(_06597_),
    .Y(_02296_),
    .A1(net448),
    .A2(net287));
 sg13g2_nand2_1 _25464_ (.Y(_06598_),
    .A(\cpu.icache.r_tag[1][20] ),
    .B(net285));
 sg13g2_o21ai_1 _25465_ (.B1(_06598_),
    .Y(_02297_),
    .A1(net412),
    .A2(net287));
 sg13g2_nand2_1 _25466_ (.Y(_06599_),
    .A(\cpu.icache.r_tag[1][21] ),
    .B(net285));
 sg13g2_o21ai_1 _25467_ (.B1(_06599_),
    .Y(_02298_),
    .A1(_08960_),
    .A2(net287));
 sg13g2_nand2_1 _25468_ (.Y(_06600_),
    .A(\cpu.icache.r_tag[1][22] ),
    .B(_06592_));
 sg13g2_o21ai_1 _25469_ (.B1(_06600_),
    .Y(_02299_),
    .A1(net449),
    .A2(_06589_));
 sg13g2_nand2_1 _25470_ (.Y(_06601_),
    .A(\cpu.icache.r_tag[1][23] ),
    .B(_06592_));
 sg13g2_o21ai_1 _25471_ (.B1(_06601_),
    .Y(_02300_),
    .A1(net500),
    .A2(_06589_));
 sg13g2_nand2_1 _25472_ (.Y(_06602_),
    .A(\cpu.icache.r_tag[1][6] ),
    .B(net285));
 sg13g2_o21ai_1 _25473_ (.B1(_06602_),
    .Y(_02301_),
    .A1(net980),
    .A2(_06590_));
 sg13g2_nand2_1 _25474_ (.Y(_06603_),
    .A(\cpu.icache.r_tag[1][7] ),
    .B(net359));
 sg13g2_o21ai_1 _25475_ (.B1(_06603_),
    .Y(_02302_),
    .A1(net939),
    .A2(net286));
 sg13g2_nand2_1 _25476_ (.Y(_06604_),
    .A(\cpu.icache.r_tag[1][8] ),
    .B(net359));
 sg13g2_o21ai_1 _25477_ (.B1(_06604_),
    .Y(_02303_),
    .A1(net940),
    .A2(net286));
 sg13g2_nand2_1 _25478_ (.Y(_06605_),
    .A(\cpu.icache.r_tag[1][9] ),
    .B(net359));
 sg13g2_o21ai_1 _25479_ (.B1(_06605_),
    .Y(_02304_),
    .A1(net974),
    .A2(net286));
 sg13g2_mux2_1 _25480_ (.A0(net978),
    .A1(\cpu.icache.r_tag[1][10] ),
    .S(net286),
    .X(_02305_));
 sg13g2_nand2_1 _25481_ (.Y(_06606_),
    .A(\cpu.icache.r_tag[1][11] ),
    .B(net359));
 sg13g2_o21ai_1 _25482_ (.B1(_06606_),
    .Y(_02306_),
    .A1(net979),
    .A2(net286));
 sg13g2_nand2_1 _25483_ (.Y(_06607_),
    .A(\cpu.icache.r_tag[1][12] ),
    .B(_06588_));
 sg13g2_o21ai_1 _25484_ (.B1(_06607_),
    .Y(_02307_),
    .A1(net349),
    .A2(_06590_));
 sg13g2_nand2_1 _25485_ (.Y(_06608_),
    .A(\cpu.icache.r_tag[1][13] ),
    .B(net359));
 sg13g2_o21ai_1 _25486_ (.B1(_06608_),
    .Y(_02308_),
    .A1(net415),
    .A2(net286));
 sg13g2_nand2_1 _25487_ (.Y(_06609_),
    .A(\cpu.icache.r_tag[1][14] ),
    .B(net359));
 sg13g2_o21ai_1 _25488_ (.B1(_06609_),
    .Y(_02309_),
    .A1(net410),
    .A2(net286));
 sg13g2_nand2_1 _25489_ (.Y(_06610_),
    .A(_08580_),
    .B(_06586_));
 sg13g2_buf_1 _25490_ (.A(_06610_),
    .X(_06611_));
 sg13g2_buf_1 _25491_ (.A(net419),
    .X(_06612_));
 sg13g2_buf_1 _25492_ (.A(net419),
    .X(_06613_));
 sg13g2_nand2_1 _25493_ (.Y(_06614_),
    .A(\cpu.icache.r_tag[2][5] ),
    .B(net357));
 sg13g2_o21ai_1 _25494_ (.B1(_06614_),
    .Y(_02310_),
    .A1(net938),
    .A2(_06612_));
 sg13g2_buf_1 _25495_ (.A(net419),
    .X(_06615_));
 sg13g2_nand2_1 _25496_ (.Y(_06616_),
    .A(\cpu.icache.r_tag[2][15] ),
    .B(net356));
 sg13g2_o21ai_1 _25497_ (.B1(_06616_),
    .Y(_02311_),
    .A1(net450),
    .A2(net358));
 sg13g2_nand2_1 _25498_ (.Y(_06617_),
    .A(\cpu.icache.r_tag[2][16] ),
    .B(net356));
 sg13g2_o21ai_1 _25499_ (.B1(_06617_),
    .Y(_02312_),
    .A1(net451),
    .A2(net358));
 sg13g2_nand2_1 _25500_ (.Y(_06618_),
    .A(\cpu.icache.r_tag[2][17] ),
    .B(net356));
 sg13g2_o21ai_1 _25501_ (.B1(_06618_),
    .Y(_02313_),
    .A1(net413),
    .A2(net358));
 sg13g2_nand2_1 _25502_ (.Y(_06619_),
    .A(\cpu.icache.r_tag[2][18] ),
    .B(net356));
 sg13g2_o21ai_1 _25503_ (.B1(_06619_),
    .Y(_02314_),
    .A1(net414),
    .A2(net358));
 sg13g2_nand2_1 _25504_ (.Y(_06620_),
    .A(\cpu.icache.r_tag[2][19] ),
    .B(_06615_));
 sg13g2_o21ai_1 _25505_ (.B1(_06620_),
    .Y(_02315_),
    .A1(net448),
    .A2(_06612_));
 sg13g2_nand2_1 _25506_ (.Y(_06621_),
    .A(\cpu.icache.r_tag[2][20] ),
    .B(net356));
 sg13g2_o21ai_1 _25507_ (.B1(_06621_),
    .Y(_02316_),
    .A1(net412),
    .A2(net358));
 sg13g2_nand2_1 _25508_ (.Y(_06622_),
    .A(\cpu.icache.r_tag[2][21] ),
    .B(net356));
 sg13g2_o21ai_1 _25509_ (.B1(_06622_),
    .Y(_02317_),
    .A1(net411),
    .A2(net358));
 sg13g2_nand2_1 _25510_ (.Y(_06623_),
    .A(\cpu.icache.r_tag[2][22] ),
    .B(net356));
 sg13g2_o21ai_1 _25511_ (.B1(_06623_),
    .Y(_02318_),
    .A1(net449),
    .A2(net358));
 sg13g2_nand2_1 _25512_ (.Y(_06624_),
    .A(\cpu.icache.r_tag[2][23] ),
    .B(net356));
 sg13g2_o21ai_1 _25513_ (.B1(_06624_),
    .Y(_02319_),
    .A1(net500),
    .A2(net358));
 sg13g2_nand2_1 _25514_ (.Y(_06625_),
    .A(\cpu.icache.r_tag[2][6] ),
    .B(_06615_));
 sg13g2_o21ai_1 _25515_ (.B1(_06625_),
    .Y(_02320_),
    .A1(net980),
    .A2(net357));
 sg13g2_nand2_1 _25516_ (.Y(_06626_),
    .A(\cpu.icache.r_tag[2][7] ),
    .B(_06611_));
 sg13g2_o21ai_1 _25517_ (.B1(_06626_),
    .Y(_02321_),
    .A1(net939),
    .A2(_06613_));
 sg13g2_nand2_1 _25518_ (.Y(_06627_),
    .A(\cpu.icache.r_tag[2][8] ),
    .B(net419));
 sg13g2_o21ai_1 _25519_ (.B1(_06627_),
    .Y(_02322_),
    .A1(net940),
    .A2(net357));
 sg13g2_nand2_1 _25520_ (.Y(_06628_),
    .A(\cpu.icache.r_tag[2][9] ),
    .B(net419));
 sg13g2_o21ai_1 _25521_ (.B1(_06628_),
    .Y(_02323_),
    .A1(net974),
    .A2(net357));
 sg13g2_mux2_1 _25522_ (.A0(net978),
    .A1(\cpu.icache.r_tag[2][10] ),
    .S(_06613_),
    .X(_02324_));
 sg13g2_nand2_1 _25523_ (.Y(_06629_),
    .A(\cpu.icache.r_tag[2][11] ),
    .B(_06611_));
 sg13g2_o21ai_1 _25524_ (.B1(_06629_),
    .Y(_02325_),
    .A1(net979),
    .A2(net357));
 sg13g2_nand2_1 _25525_ (.Y(_06630_),
    .A(\cpu.icache.r_tag[2][12] ),
    .B(net419));
 sg13g2_o21ai_1 _25526_ (.B1(_06630_),
    .Y(_02326_),
    .A1(net349),
    .A2(net357));
 sg13g2_nand2_1 _25527_ (.Y(_06631_),
    .A(\cpu.icache.r_tag[2][13] ),
    .B(net419));
 sg13g2_o21ai_1 _25528_ (.B1(_06631_),
    .Y(_02327_),
    .A1(net415),
    .A2(net357));
 sg13g2_nand2_1 _25529_ (.Y(_06632_),
    .A(\cpu.icache.r_tag[2][14] ),
    .B(net419));
 sg13g2_o21ai_1 _25530_ (.B1(_06632_),
    .Y(_02328_),
    .A1(net410),
    .A2(net357));
 sg13g2_buf_1 _25531_ (.A(_06515_),
    .X(_06633_));
 sg13g2_nand2_1 _25532_ (.Y(_06634_),
    .A(\cpu.icache.r_tag[3][5] ),
    .B(_06517_));
 sg13g2_o21ai_1 _25533_ (.B1(_06634_),
    .Y(_02329_),
    .A1(net938),
    .A2(_06633_));
 sg13g2_nand2_1 _25534_ (.Y(_06635_),
    .A(\cpu.icache.r_tag[3][15] ),
    .B(net288));
 sg13g2_o21ai_1 _25535_ (.B1(_06635_),
    .Y(_02330_),
    .A1(net450),
    .A2(net284));
 sg13g2_nand2_1 _25536_ (.Y(_06636_),
    .A(\cpu.icache.r_tag[3][16] ),
    .B(net288));
 sg13g2_o21ai_1 _25537_ (.B1(_06636_),
    .Y(_02331_),
    .A1(net451),
    .A2(net284));
 sg13g2_nand2_1 _25538_ (.Y(_06637_),
    .A(\cpu.icache.r_tag[3][17] ),
    .B(net288));
 sg13g2_o21ai_1 _25539_ (.B1(_06637_),
    .Y(_02332_),
    .A1(net413),
    .A2(net284));
 sg13g2_nand2_1 _25540_ (.Y(_06638_),
    .A(\cpu.icache.r_tag[3][18] ),
    .B(net288));
 sg13g2_o21ai_1 _25541_ (.B1(_06638_),
    .Y(_02333_),
    .A1(net414),
    .A2(net284));
 sg13g2_nand2_1 _25542_ (.Y(_06639_),
    .A(\cpu.icache.r_tag[3][19] ),
    .B(net288));
 sg13g2_o21ai_1 _25543_ (.B1(_06639_),
    .Y(_02334_),
    .A1(net448),
    .A2(net284));
 sg13g2_buf_1 _25544_ (.A(_06515_),
    .X(_06640_));
 sg13g2_nand2_1 _25545_ (.Y(_06641_),
    .A(\cpu.icache.r_tag[3][20] ),
    .B(net283));
 sg13g2_o21ai_1 _25546_ (.B1(_06641_),
    .Y(_02335_),
    .A1(net412),
    .A2(net284));
 sg13g2_nand2_1 _25547_ (.Y(_06642_),
    .A(\cpu.icache.r_tag[3][21] ),
    .B(net283));
 sg13g2_o21ai_1 _25548_ (.B1(_06642_),
    .Y(_02336_),
    .A1(net411),
    .A2(_06633_));
 sg13g2_nand2_1 _25549_ (.Y(_06643_),
    .A(\cpu.icache.r_tag[3][22] ),
    .B(_06640_));
 sg13g2_o21ai_1 _25550_ (.B1(_06643_),
    .Y(_02337_),
    .A1(net449),
    .A2(net284));
 sg13g2_nand2_1 _25551_ (.Y(_06644_),
    .A(\cpu.icache.r_tag[3][23] ),
    .B(net283));
 sg13g2_o21ai_1 _25552_ (.B1(_06644_),
    .Y(_02338_),
    .A1(net500),
    .A2(net289));
 sg13g2_nand2_1 _25553_ (.Y(_06645_),
    .A(\cpu.icache.r_tag[3][6] ),
    .B(net283));
 sg13g2_o21ai_1 _25554_ (.B1(_06645_),
    .Y(_02339_),
    .A1(net980),
    .A2(_06516_));
 sg13g2_nand2_1 _25555_ (.Y(_06646_),
    .A(\cpu.icache.r_tag[3][7] ),
    .B(net283));
 sg13g2_o21ai_1 _25556_ (.B1(_06646_),
    .Y(_02340_),
    .A1(net939),
    .A2(net289));
 sg13g2_nand2_1 _25557_ (.Y(_06647_),
    .A(\cpu.icache.r_tag[3][8] ),
    .B(net283));
 sg13g2_o21ai_1 _25558_ (.B1(_06647_),
    .Y(_02341_),
    .A1(net940),
    .A2(_06516_));
 sg13g2_nand2_1 _25559_ (.Y(_06648_),
    .A(\cpu.icache.r_tag[3][9] ),
    .B(net283));
 sg13g2_o21ai_1 _25560_ (.B1(_06648_),
    .Y(_02342_),
    .A1(net974),
    .A2(net289));
 sg13g2_mux2_1 _25561_ (.A0(net978),
    .A1(\cpu.icache.r_tag[3][10] ),
    .S(_06517_),
    .X(_02343_));
 sg13g2_nand2_1 _25562_ (.Y(_06649_),
    .A(\cpu.icache.r_tag[3][11] ),
    .B(net283));
 sg13g2_o21ai_1 _25563_ (.B1(_06649_),
    .Y(_02344_),
    .A1(net979),
    .A2(net289));
 sg13g2_nand2_1 _25564_ (.Y(_06650_),
    .A(\cpu.icache.r_tag[3][12] ),
    .B(_06640_));
 sg13g2_o21ai_1 _25565_ (.B1(_06650_),
    .Y(_02345_),
    .A1(net349),
    .A2(net289));
 sg13g2_nand2_1 _25566_ (.Y(_06651_),
    .A(\cpu.icache.r_tag[3][13] ),
    .B(_06515_));
 sg13g2_o21ai_1 _25567_ (.B1(_06651_),
    .Y(_02346_),
    .A1(net415),
    .A2(net289));
 sg13g2_nand2_1 _25568_ (.Y(_06652_),
    .A(\cpu.icache.r_tag[3][14] ),
    .B(_06515_));
 sg13g2_o21ai_1 _25569_ (.B1(_06652_),
    .Y(_02347_),
    .A1(net410),
    .A2(net289));
 sg13g2_nand2_1 _25570_ (.Y(_06653_),
    .A(_09007_),
    .B(_06586_));
 sg13g2_buf_1 _25571_ (.A(_06653_),
    .X(_06654_));
 sg13g2_buf_1 _25572_ (.A(net509),
    .X(_06655_));
 sg13g2_buf_1 _25573_ (.A(net509),
    .X(_06656_));
 sg13g2_nand2_1 _25574_ (.Y(_06657_),
    .A(\cpu.icache.r_tag[4][5] ),
    .B(_06656_));
 sg13g2_o21ai_1 _25575_ (.B1(_06657_),
    .Y(_02348_),
    .A1(net938),
    .A2(net461));
 sg13g2_buf_1 _25576_ (.A(net509),
    .X(_06658_));
 sg13g2_nand2_1 _25577_ (.Y(_06659_),
    .A(\cpu.icache.r_tag[4][15] ),
    .B(net459));
 sg13g2_o21ai_1 _25578_ (.B1(_06659_),
    .Y(_02349_),
    .A1(net450),
    .A2(net461));
 sg13g2_nand2_1 _25579_ (.Y(_06660_),
    .A(\cpu.icache.r_tag[4][16] ),
    .B(net459));
 sg13g2_o21ai_1 _25580_ (.B1(_06660_),
    .Y(_02350_),
    .A1(net451),
    .A2(net461));
 sg13g2_nand2_1 _25581_ (.Y(_06661_),
    .A(\cpu.icache.r_tag[4][17] ),
    .B(net459));
 sg13g2_o21ai_1 _25582_ (.B1(_06661_),
    .Y(_02351_),
    .A1(net413),
    .A2(net461));
 sg13g2_nand2_1 _25583_ (.Y(_06662_),
    .A(\cpu.icache.r_tag[4][18] ),
    .B(net459));
 sg13g2_o21ai_1 _25584_ (.B1(_06662_),
    .Y(_02352_),
    .A1(net414),
    .A2(net461));
 sg13g2_nand2_1 _25585_ (.Y(_06663_),
    .A(\cpu.icache.r_tag[4][19] ),
    .B(_06658_));
 sg13g2_o21ai_1 _25586_ (.B1(_06663_),
    .Y(_02353_),
    .A1(net448),
    .A2(_06655_));
 sg13g2_nand2_1 _25587_ (.Y(_06664_),
    .A(\cpu.icache.r_tag[4][20] ),
    .B(net459));
 sg13g2_o21ai_1 _25588_ (.B1(_06664_),
    .Y(_02354_),
    .A1(_08939_),
    .A2(net461));
 sg13g2_nand2_1 _25589_ (.Y(_06665_),
    .A(\cpu.icache.r_tag[4][21] ),
    .B(net459));
 sg13g2_o21ai_1 _25590_ (.B1(_06665_),
    .Y(_02355_),
    .A1(net411),
    .A2(net461));
 sg13g2_nand2_1 _25591_ (.Y(_06666_),
    .A(\cpu.icache.r_tag[4][22] ),
    .B(net459));
 sg13g2_o21ai_1 _25592_ (.B1(_06666_),
    .Y(_02356_),
    .A1(_08854_),
    .A2(net461));
 sg13g2_nand2_1 _25593_ (.Y(_06667_),
    .A(\cpu.icache.r_tag[4][23] ),
    .B(_06658_));
 sg13g2_o21ai_1 _25594_ (.B1(_06667_),
    .Y(_02357_),
    .A1(net500),
    .A2(_06655_));
 sg13g2_nand2_1 _25595_ (.Y(_06668_),
    .A(\cpu.icache.r_tag[4][6] ),
    .B(net459));
 sg13g2_o21ai_1 _25596_ (.B1(_06668_),
    .Y(_02358_),
    .A1(net980),
    .A2(net460));
 sg13g2_nand2_1 _25597_ (.Y(_06669_),
    .A(\cpu.icache.r_tag[4][7] ),
    .B(net509));
 sg13g2_o21ai_1 _25598_ (.B1(_06669_),
    .Y(_02359_),
    .A1(net939),
    .A2(net460));
 sg13g2_nand2_1 _25599_ (.Y(_06670_),
    .A(\cpu.icache.r_tag[4][8] ),
    .B(net509));
 sg13g2_o21ai_1 _25600_ (.B1(_06670_),
    .Y(_02360_),
    .A1(net940),
    .A2(net460));
 sg13g2_nand2_1 _25601_ (.Y(_06671_),
    .A(\cpu.icache.r_tag[4][9] ),
    .B(net509));
 sg13g2_o21ai_1 _25602_ (.B1(_06671_),
    .Y(_02361_),
    .A1(net974),
    .A2(net460));
 sg13g2_mux2_1 _25603_ (.A0(net978),
    .A1(\cpu.icache.r_tag[4][10] ),
    .S(net460),
    .X(_02362_));
 sg13g2_nand2_1 _25604_ (.Y(_06672_),
    .A(\cpu.icache.r_tag[4][11] ),
    .B(net509));
 sg13g2_o21ai_1 _25605_ (.B1(_06672_),
    .Y(_02363_),
    .A1(net979),
    .A2(net460));
 sg13g2_nand2_1 _25606_ (.Y(_06673_),
    .A(\cpu.icache.r_tag[4][12] ),
    .B(_06654_));
 sg13g2_o21ai_1 _25607_ (.B1(_06673_),
    .Y(_02364_),
    .A1(net349),
    .A2(net460));
 sg13g2_nand2_1 _25608_ (.Y(_06674_),
    .A(\cpu.icache.r_tag[4][13] ),
    .B(_06654_));
 sg13g2_o21ai_1 _25609_ (.B1(_06674_),
    .Y(_02365_),
    .A1(net415),
    .A2(_06656_));
 sg13g2_nand2_1 _25610_ (.Y(_06675_),
    .A(\cpu.icache.r_tag[4][14] ),
    .B(net509));
 sg13g2_o21ai_1 _25611_ (.B1(_06675_),
    .Y(_02366_),
    .A1(net410),
    .A2(net460));
 sg13g2_nand2_1 _25612_ (.Y(_06676_),
    .A(_08992_),
    .B(_06586_));
 sg13g2_buf_1 _25613_ (.A(_06676_),
    .X(_06677_));
 sg13g2_buf_1 _25614_ (.A(net418),
    .X(_06678_));
 sg13g2_buf_1 _25615_ (.A(net418),
    .X(_06679_));
 sg13g2_nand2_1 _25616_ (.Y(_06680_),
    .A(\cpu.icache.r_tag[5][5] ),
    .B(net354));
 sg13g2_o21ai_1 _25617_ (.B1(_06680_),
    .Y(_02367_),
    .A1(net938),
    .A2(net355));
 sg13g2_buf_1 _25618_ (.A(net418),
    .X(_06681_));
 sg13g2_nand2_1 _25619_ (.Y(_06682_),
    .A(\cpu.icache.r_tag[5][15] ),
    .B(net353));
 sg13g2_o21ai_1 _25620_ (.B1(_06682_),
    .Y(_02368_),
    .A1(net450),
    .A2(net355));
 sg13g2_nand2_1 _25621_ (.Y(_06683_),
    .A(\cpu.icache.r_tag[5][16] ),
    .B(net353));
 sg13g2_o21ai_1 _25622_ (.B1(_06683_),
    .Y(_02369_),
    .A1(net451),
    .A2(net355));
 sg13g2_nand2_1 _25623_ (.Y(_06684_),
    .A(\cpu.icache.r_tag[5][17] ),
    .B(net353));
 sg13g2_o21ai_1 _25624_ (.B1(_06684_),
    .Y(_02370_),
    .A1(net413),
    .A2(net355));
 sg13g2_nand2_1 _25625_ (.Y(_06685_),
    .A(\cpu.icache.r_tag[5][18] ),
    .B(net353));
 sg13g2_o21ai_1 _25626_ (.B1(_06685_),
    .Y(_02371_),
    .A1(net414),
    .A2(net355));
 sg13g2_nand2_1 _25627_ (.Y(_06686_),
    .A(\cpu.icache.r_tag[5][19] ),
    .B(net353));
 sg13g2_o21ai_1 _25628_ (.B1(_06686_),
    .Y(_02372_),
    .A1(net448),
    .A2(net355));
 sg13g2_nand2_1 _25629_ (.Y(_06687_),
    .A(\cpu.icache.r_tag[5][20] ),
    .B(net353));
 sg13g2_o21ai_1 _25630_ (.B1(_06687_),
    .Y(_02373_),
    .A1(net412),
    .A2(net355));
 sg13g2_nand2_1 _25631_ (.Y(_06688_),
    .A(\cpu.icache.r_tag[5][21] ),
    .B(_06681_));
 sg13g2_o21ai_1 _25632_ (.B1(_06688_),
    .Y(_02374_),
    .A1(net411),
    .A2(_06678_));
 sg13g2_nand2_1 _25633_ (.Y(_06689_),
    .A(\cpu.icache.r_tag[5][22] ),
    .B(_06681_));
 sg13g2_o21ai_1 _25634_ (.B1(_06689_),
    .Y(_02375_),
    .A1(net449),
    .A2(_06678_));
 sg13g2_nand2_1 _25635_ (.Y(_06690_),
    .A(\cpu.icache.r_tag[5][23] ),
    .B(net353));
 sg13g2_o21ai_1 _25636_ (.B1(_06690_),
    .Y(_02376_),
    .A1(net500),
    .A2(net355));
 sg13g2_nand2_1 _25637_ (.Y(_06691_),
    .A(\cpu.icache.r_tag[5][6] ),
    .B(net353));
 sg13g2_o21ai_1 _25638_ (.B1(_06691_),
    .Y(_02377_),
    .A1(net980),
    .A2(net354));
 sg13g2_nand2_1 _25639_ (.Y(_06692_),
    .A(\cpu.icache.r_tag[5][7] ),
    .B(net418));
 sg13g2_o21ai_1 _25640_ (.B1(_06692_),
    .Y(_02378_),
    .A1(net939),
    .A2(net354));
 sg13g2_nand2_1 _25641_ (.Y(_06693_),
    .A(\cpu.icache.r_tag[5][8] ),
    .B(net418));
 sg13g2_o21ai_1 _25642_ (.B1(_06693_),
    .Y(_02379_),
    .A1(net940),
    .A2(net354));
 sg13g2_nand2_1 _25643_ (.Y(_06694_),
    .A(\cpu.icache.r_tag[5][9] ),
    .B(net418));
 sg13g2_o21ai_1 _25644_ (.B1(_06694_),
    .Y(_02380_),
    .A1(net974),
    .A2(net354));
 sg13g2_mux2_1 _25645_ (.A0(net978),
    .A1(\cpu.icache.r_tag[5][10] ),
    .S(_06679_),
    .X(_02381_));
 sg13g2_nand2_1 _25646_ (.Y(_06695_),
    .A(\cpu.icache.r_tag[5][11] ),
    .B(net418));
 sg13g2_o21ai_1 _25647_ (.B1(_06695_),
    .Y(_02382_),
    .A1(net979),
    .A2(net354));
 sg13g2_nand2_1 _25648_ (.Y(_06696_),
    .A(\cpu.icache.r_tag[5][12] ),
    .B(_06677_));
 sg13g2_o21ai_1 _25649_ (.B1(_06696_),
    .Y(_02383_),
    .A1(net349),
    .A2(net354));
 sg13g2_nand2_1 _25650_ (.Y(_06697_),
    .A(\cpu.icache.r_tag[5][13] ),
    .B(_06677_));
 sg13g2_o21ai_1 _25651_ (.B1(_06697_),
    .Y(_02384_),
    .A1(net415),
    .A2(net354));
 sg13g2_nand2_1 _25652_ (.Y(_06698_),
    .A(\cpu.icache.r_tag[5][14] ),
    .B(net418));
 sg13g2_o21ai_1 _25653_ (.B1(_06698_),
    .Y(_02385_),
    .A1(net410),
    .A2(_06679_));
 sg13g2_nand2_1 _25654_ (.Y(_06699_),
    .A(_08667_),
    .B(_06586_));
 sg13g2_buf_1 _25655_ (.A(_06699_),
    .X(_06700_));
 sg13g2_buf_1 _25656_ (.A(net417),
    .X(_06701_));
 sg13g2_buf_1 _25657_ (.A(net417),
    .X(_06702_));
 sg13g2_nand2_1 _25658_ (.Y(_06703_),
    .A(\cpu.icache.r_tag[6][5] ),
    .B(net351));
 sg13g2_o21ai_1 _25659_ (.B1(_06703_),
    .Y(_02386_),
    .A1(net938),
    .A2(_06701_));
 sg13g2_buf_1 _25660_ (.A(net417),
    .X(_06704_));
 sg13g2_nand2_1 _25661_ (.Y(_06705_),
    .A(\cpu.icache.r_tag[6][15] ),
    .B(net350));
 sg13g2_o21ai_1 _25662_ (.B1(_06705_),
    .Y(_02387_),
    .A1(net450),
    .A2(net352));
 sg13g2_nand2_1 _25663_ (.Y(_06706_),
    .A(\cpu.icache.r_tag[6][16] ),
    .B(net350));
 sg13g2_o21ai_1 _25664_ (.B1(_06706_),
    .Y(_02388_),
    .A1(net451),
    .A2(net352));
 sg13g2_nand2_1 _25665_ (.Y(_06707_),
    .A(\cpu.icache.r_tag[6][17] ),
    .B(net350));
 sg13g2_o21ai_1 _25666_ (.B1(_06707_),
    .Y(_02389_),
    .A1(net413),
    .A2(net352));
 sg13g2_nand2_1 _25667_ (.Y(_06708_),
    .A(\cpu.icache.r_tag[6][18] ),
    .B(net350));
 sg13g2_o21ai_1 _25668_ (.B1(_06708_),
    .Y(_02390_),
    .A1(net414),
    .A2(net352));
 sg13g2_nand2_1 _25669_ (.Y(_06709_),
    .A(\cpu.icache.r_tag[6][19] ),
    .B(net350));
 sg13g2_o21ai_1 _25670_ (.B1(_06709_),
    .Y(_02391_),
    .A1(net448),
    .A2(_06701_));
 sg13g2_nand2_1 _25671_ (.Y(_06710_),
    .A(\cpu.icache.r_tag[6][20] ),
    .B(net350));
 sg13g2_o21ai_1 _25672_ (.B1(_06710_),
    .Y(_02392_),
    .A1(net412),
    .A2(net352));
 sg13g2_nand2_1 _25673_ (.Y(_06711_),
    .A(\cpu.icache.r_tag[6][21] ),
    .B(net350));
 sg13g2_o21ai_1 _25674_ (.B1(_06711_),
    .Y(_02393_),
    .A1(net411),
    .A2(net352));
 sg13g2_nand2_1 _25675_ (.Y(_06712_),
    .A(\cpu.icache.r_tag[6][22] ),
    .B(_06704_));
 sg13g2_o21ai_1 _25676_ (.B1(_06712_),
    .Y(_02394_),
    .A1(net449),
    .A2(net352));
 sg13g2_nand2_1 _25677_ (.Y(_06713_),
    .A(\cpu.icache.r_tag[6][23] ),
    .B(_06704_));
 sg13g2_o21ai_1 _25678_ (.B1(_06713_),
    .Y(_02395_),
    .A1(net500),
    .A2(net352));
 sg13g2_nand2_1 _25679_ (.Y(_06714_),
    .A(\cpu.icache.r_tag[6][6] ),
    .B(net350));
 sg13g2_o21ai_1 _25680_ (.B1(_06714_),
    .Y(_02396_),
    .A1(_04211_),
    .A2(net351));
 sg13g2_nand2_1 _25681_ (.Y(_06715_),
    .A(\cpu.icache.r_tag[6][7] ),
    .B(net417));
 sg13g2_o21ai_1 _25682_ (.B1(_06715_),
    .Y(_02397_),
    .A1(net939),
    .A2(_06702_));
 sg13g2_nand2_1 _25683_ (.Y(_06716_),
    .A(\cpu.icache.r_tag[6][8] ),
    .B(net417));
 sg13g2_o21ai_1 _25684_ (.B1(_06716_),
    .Y(_02398_),
    .A1(net940),
    .A2(net351));
 sg13g2_nand2_1 _25685_ (.Y(_06717_),
    .A(\cpu.icache.r_tag[6][9] ),
    .B(net417));
 sg13g2_o21ai_1 _25686_ (.B1(_06717_),
    .Y(_02399_),
    .A1(net974),
    .A2(net351));
 sg13g2_mux2_1 _25687_ (.A0(_04732_),
    .A1(\cpu.icache.r_tag[6][10] ),
    .S(net351),
    .X(_02400_));
 sg13g2_nand2_1 _25688_ (.Y(_06718_),
    .A(\cpu.icache.r_tag[6][11] ),
    .B(_06700_));
 sg13g2_o21ai_1 _25689_ (.B1(_06718_),
    .Y(_02401_),
    .A1(net979),
    .A2(_06702_));
 sg13g2_nand2_1 _25690_ (.Y(_06719_),
    .A(\cpu.icache.r_tag[6][12] ),
    .B(net417));
 sg13g2_o21ai_1 _25691_ (.B1(_06719_),
    .Y(_02402_),
    .A1(net349),
    .A2(net351));
 sg13g2_nand2_1 _25692_ (.Y(_06720_),
    .A(\cpu.icache.r_tag[6][13] ),
    .B(_06700_));
 sg13g2_o21ai_1 _25693_ (.B1(_06720_),
    .Y(_02403_),
    .A1(net415),
    .A2(net351));
 sg13g2_nand2_1 _25694_ (.Y(_06721_),
    .A(\cpu.icache.r_tag[6][14] ),
    .B(net417));
 sg13g2_o21ai_1 _25695_ (.B1(_06721_),
    .Y(_02404_),
    .A1(net410),
    .A2(net351));
 sg13g2_nand2_1 _25696_ (.Y(_06722_),
    .A(_08700_),
    .B(_06586_));
 sg13g2_buf_1 _25697_ (.A(_06722_),
    .X(_06723_));
 sg13g2_buf_1 _25698_ (.A(net508),
    .X(_06724_));
 sg13g2_buf_1 _25699_ (.A(net508),
    .X(_06725_));
 sg13g2_nand2_1 _25700_ (.Y(_06726_),
    .A(\cpu.icache.r_tag[7][5] ),
    .B(net457));
 sg13g2_o21ai_1 _25701_ (.B1(_06726_),
    .Y(_02405_),
    .A1(_08808_),
    .A2(net458));
 sg13g2_buf_1 _25702_ (.A(net508),
    .X(_06727_));
 sg13g2_nand2_1 _25703_ (.Y(_06728_),
    .A(\cpu.icache.r_tag[7][15] ),
    .B(net456));
 sg13g2_o21ai_1 _25704_ (.B1(_06728_),
    .Y(_02406_),
    .A1(_08698_),
    .A2(net458));
 sg13g2_nand2_1 _25705_ (.Y(_06729_),
    .A(\cpu.icache.r_tag[7][16] ),
    .B(net456));
 sg13g2_o21ai_1 _25706_ (.B1(_06729_),
    .Y(_02407_),
    .A1(net451),
    .A2(net458));
 sg13g2_nand2_1 _25707_ (.Y(_06730_),
    .A(\cpu.icache.r_tag[7][17] ),
    .B(net456));
 sg13g2_o21ai_1 _25708_ (.B1(_06730_),
    .Y(_02408_),
    .A1(net413),
    .A2(net458));
 sg13g2_nand2_1 _25709_ (.Y(_06731_),
    .A(\cpu.icache.r_tag[7][18] ),
    .B(_06727_));
 sg13g2_o21ai_1 _25710_ (.B1(_06731_),
    .Y(_02409_),
    .A1(net414),
    .A2(_06724_));
 sg13g2_nand2_1 _25711_ (.Y(_06732_),
    .A(\cpu.icache.r_tag[7][19] ),
    .B(net456));
 sg13g2_o21ai_1 _25712_ (.B1(_06732_),
    .Y(_02410_),
    .A1(_08896_),
    .A2(net458));
 sg13g2_nand2_1 _25713_ (.Y(_06733_),
    .A(\cpu.icache.r_tag[7][20] ),
    .B(net456));
 sg13g2_o21ai_1 _25714_ (.B1(_06733_),
    .Y(_02411_),
    .A1(net412),
    .A2(net458));
 sg13g2_nand2_1 _25715_ (.Y(_06734_),
    .A(\cpu.icache.r_tag[7][21] ),
    .B(net456));
 sg13g2_o21ai_1 _25716_ (.B1(_06734_),
    .Y(_02412_),
    .A1(net411),
    .A2(net458));
 sg13g2_nand2_1 _25717_ (.Y(_06735_),
    .A(\cpu.icache.r_tag[7][22] ),
    .B(net456));
 sg13g2_o21ai_1 _25718_ (.B1(_06735_),
    .Y(_02413_),
    .A1(net449),
    .A2(net458));
 sg13g2_nand2_1 _25719_ (.Y(_06736_),
    .A(\cpu.icache.r_tag[7][23] ),
    .B(_06727_));
 sg13g2_o21ai_1 _25720_ (.B1(_06736_),
    .Y(_02414_),
    .A1(net500),
    .A2(_06724_));
 sg13g2_nand2_1 _25721_ (.Y(_06737_),
    .A(\cpu.icache.r_tag[7][6] ),
    .B(net456));
 sg13g2_o21ai_1 _25722_ (.B1(_06737_),
    .Y(_02415_),
    .A1(_04211_),
    .A2(net457));
 sg13g2_nand2_1 _25723_ (.Y(_06738_),
    .A(\cpu.icache.r_tag[7][7] ),
    .B(net508));
 sg13g2_o21ai_1 _25724_ (.B1(_06738_),
    .Y(_02416_),
    .A1(_08779_),
    .A2(net457));
 sg13g2_nand2_1 _25725_ (.Y(_06739_),
    .A(\cpu.icache.r_tag[7][8] ),
    .B(net508));
 sg13g2_o21ai_1 _25726_ (.B1(_06739_),
    .Y(_02417_),
    .A1(_08759_),
    .A2(net457));
 sg13g2_nand2_1 _25727_ (.Y(_06740_),
    .A(\cpu.icache.r_tag[7][9] ),
    .B(net508));
 sg13g2_o21ai_1 _25728_ (.B1(_06740_),
    .Y(_02418_),
    .A1(_05748_),
    .A2(net457));
 sg13g2_mux2_1 _25729_ (.A0(_04732_),
    .A1(\cpu.icache.r_tag[7][10] ),
    .S(net457),
    .X(_02419_));
 sg13g2_nand2_1 _25730_ (.Y(_06741_),
    .A(\cpu.icache.r_tag[7][11] ),
    .B(_06723_));
 sg13g2_o21ai_1 _25731_ (.B1(_06741_),
    .Y(_02420_),
    .A1(_04278_),
    .A2(_06725_));
 sg13g2_nand2_1 _25732_ (.Y(_06742_),
    .A(\cpu.icache.r_tag[7][12] ),
    .B(net508));
 sg13g2_o21ai_1 _25733_ (.B1(_06742_),
    .Y(_02421_),
    .A1(_08558_),
    .A2(net457));
 sg13g2_nand2_1 _25734_ (.Y(_06743_),
    .A(\cpu.icache.r_tag[7][13] ),
    .B(net508));
 sg13g2_o21ai_1 _25735_ (.B1(_06743_),
    .Y(_02422_),
    .A1(_08634_),
    .A2(net457));
 sg13g2_nand2_1 _25736_ (.Y(_06744_),
    .A(\cpu.icache.r_tag[7][14] ),
    .B(_06723_));
 sg13g2_o21ai_1 _25737_ (.B1(_06744_),
    .Y(_02423_),
    .A1(_09158_),
    .A2(_06725_));
 sg13g2_buf_1 _25738_ (.A(_10128_),
    .X(_06745_));
 sg13g2_nand2_1 _25739_ (.Y(_06746_),
    .A(net124),
    .B(net652));
 sg13g2_buf_2 _25740_ (.A(_06746_),
    .X(_06747_));
 sg13g2_buf_1 _25741_ (.A(_06747_),
    .X(_06748_));
 sg13g2_mux2_1 _25742_ (.A0(net897),
    .A1(\cpu.intr.r_clock_cmp[0] ),
    .S(net80),
    .X(_02433_));
 sg13g2_mux2_1 _25743_ (.A0(_10312_),
    .A1(\cpu.intr.r_clock_cmp[10] ),
    .S(net80),
    .X(_02434_));
 sg13g2_mux2_1 _25744_ (.A0(_10319_),
    .A1(\cpu.intr.r_clock_cmp[11] ),
    .S(net80),
    .X(_02435_));
 sg13g2_mux2_1 _25745_ (.A0(_10324_),
    .A1(\cpu.intr.r_clock_cmp[12] ),
    .S(net80),
    .X(_02436_));
 sg13g2_mux2_1 _25746_ (.A0(_10326_),
    .A1(\cpu.intr.r_clock_cmp[13] ),
    .S(net80),
    .X(_02437_));
 sg13g2_mux2_1 _25747_ (.A0(_10339_),
    .A1(\cpu.intr.r_clock_cmp[14] ),
    .S(net80),
    .X(_02438_));
 sg13g2_mux2_1 _25748_ (.A0(_10344_),
    .A1(\cpu.intr.r_clock_cmp[15] ),
    .S(net80),
    .X(_02439_));
 sg13g2_nand2_1 _25749_ (.Y(_06749_),
    .A(net124),
    .B(net653));
 sg13g2_buf_2 _25750_ (.A(_06749_),
    .X(_06750_));
 sg13g2_buf_1 _25751_ (.A(_06750_),
    .X(_06751_));
 sg13g2_mux2_1 _25752_ (.A0(net897),
    .A1(\cpu.intr.r_clock_cmp[16] ),
    .S(_06751_),
    .X(_02440_));
 sg13g2_mux2_1 _25753_ (.A0(net918),
    .A1(\cpu.intr.r_clock_cmp[17] ),
    .S(net79),
    .X(_02441_));
 sg13g2_mux2_1 _25754_ (.A0(net917),
    .A1(\cpu.intr.r_clock_cmp[18] ),
    .S(net79),
    .X(_02442_));
 sg13g2_mux2_1 _25755_ (.A0(net1033),
    .A1(\cpu.intr.r_clock_cmp[19] ),
    .S(net79),
    .X(_02443_));
 sg13g2_mux2_1 _25756_ (.A0(net918),
    .A1(\cpu.intr.r_clock_cmp[1] ),
    .S(net80),
    .X(_02444_));
 sg13g2_mux2_1 _25757_ (.A0(net1032),
    .A1(\cpu.intr.r_clock_cmp[20] ),
    .S(net79),
    .X(_02445_));
 sg13g2_mux2_1 _25758_ (.A0(net916),
    .A1(\cpu.intr.r_clock_cmp[21] ),
    .S(net79),
    .X(_02446_));
 sg13g2_mux2_1 _25759_ (.A0(net1031),
    .A1(\cpu.intr.r_clock_cmp[22] ),
    .S(_06751_),
    .X(_02447_));
 sg13g2_mux2_1 _25760_ (.A0(net991),
    .A1(\cpu.intr.r_clock_cmp[23] ),
    .S(net79),
    .X(_02448_));
 sg13g2_mux2_1 _25761_ (.A0(_10302_),
    .A1(\cpu.intr.r_clock_cmp[24] ),
    .S(net79),
    .X(_02449_));
 sg13g2_mux2_1 _25762_ (.A0(_10307_),
    .A1(\cpu.intr.r_clock_cmp[25] ),
    .S(net79),
    .X(_02450_));
 sg13g2_mux2_1 _25763_ (.A0(_10312_),
    .A1(\cpu.intr.r_clock_cmp[26] ),
    .S(_06750_),
    .X(_02451_));
 sg13g2_mux2_1 _25764_ (.A0(_10319_),
    .A1(\cpu.intr.r_clock_cmp[27] ),
    .S(_06750_),
    .X(_02452_));
 sg13g2_mux2_1 _25765_ (.A0(_10324_),
    .A1(\cpu.intr.r_clock_cmp[28] ),
    .S(_06750_),
    .X(_02453_));
 sg13g2_mux2_1 _25766_ (.A0(_10326_),
    .A1(\cpu.intr.r_clock_cmp[29] ),
    .S(_06750_),
    .X(_02454_));
 sg13g2_mux2_1 _25767_ (.A0(net917),
    .A1(\cpu.intr.r_clock_cmp[2] ),
    .S(_06748_),
    .X(_02455_));
 sg13g2_mux2_1 _25768_ (.A0(_10339_),
    .A1(\cpu.intr.r_clock_cmp[30] ),
    .S(_06750_),
    .X(_02456_));
 sg13g2_mux2_1 _25769_ (.A0(_10344_),
    .A1(\cpu.intr.r_clock_cmp[31] ),
    .S(_06750_),
    .X(_02457_));
 sg13g2_mux2_1 _25770_ (.A0(net1033),
    .A1(\cpu.intr.r_clock_cmp[3] ),
    .S(_06748_),
    .X(_02458_));
 sg13g2_mux2_1 _25771_ (.A0(net1002),
    .A1(\cpu.intr.r_clock_cmp[4] ),
    .S(_06747_),
    .X(_02459_));
 sg13g2_mux2_1 _25772_ (.A0(net1001),
    .A1(\cpu.intr.r_clock_cmp[5] ),
    .S(_06747_),
    .X(_02460_));
 sg13g2_mux2_1 _25773_ (.A0(net1000),
    .A1(\cpu.intr.r_clock_cmp[6] ),
    .S(_06747_),
    .X(_02461_));
 sg13g2_mux2_1 _25774_ (.A0(net991),
    .A1(\cpu.intr.r_clock_cmp[7] ),
    .S(_06747_),
    .X(_02462_));
 sg13g2_mux2_1 _25775_ (.A0(_10302_),
    .A1(\cpu.intr.r_clock_cmp[8] ),
    .S(_06747_),
    .X(_02463_));
 sg13g2_mux2_1 _25776_ (.A0(_10307_),
    .A1(\cpu.intr.r_clock_cmp[9] ),
    .S(_06747_),
    .X(_02464_));
 sg13g2_nor4_1 _25777_ (.A(net542),
    .B(_09368_),
    .C(_10178_),
    .D(_10126_),
    .Y(_06752_));
 sg13g2_buf_2 _25778_ (.A(_06752_),
    .X(_06753_));
 sg13g2_buf_1 _25779_ (.A(_06753_),
    .X(_06754_));
 sg13g2_mux2_1 _25780_ (.A0(\cpu.intr.r_timer_reload[0] ),
    .A1(net897),
    .S(net123),
    .X(_02488_));
 sg13g2_mux2_1 _25781_ (.A0(\cpu.intr.r_timer_reload[10] ),
    .A1(_10312_),
    .S(net123),
    .X(_02489_));
 sg13g2_mux2_1 _25782_ (.A0(\cpu.intr.r_timer_reload[11] ),
    .A1(_10319_),
    .S(net123),
    .X(_02490_));
 sg13g2_mux2_1 _25783_ (.A0(\cpu.intr.r_timer_reload[12] ),
    .A1(_10324_),
    .S(net123),
    .X(_02491_));
 sg13g2_mux2_1 _25784_ (.A0(\cpu.intr.r_timer_reload[13] ),
    .A1(_10326_),
    .S(net123),
    .X(_02492_));
 sg13g2_mux2_1 _25785_ (.A0(\cpu.intr.r_timer_reload[14] ),
    .A1(_10339_),
    .S(net123),
    .X(_02493_));
 sg13g2_mux2_1 _25786_ (.A0(\cpu.intr.r_timer_reload[15] ),
    .A1(_10344_),
    .S(net123),
    .X(_02494_));
 sg13g2_o21ai_1 _25787_ (.B1(_10188_),
    .Y(_02495_),
    .A1(_10182_),
    .A2(_10181_));
 sg13g2_mux2_1 _25788_ (.A0(\cpu.intr.r_timer_reload[17] ),
    .A1(net918),
    .S(_10181_),
    .X(_02496_));
 sg13g2_inv_1 _25789_ (.Y(_06755_),
    .A(\cpu.intr.r_timer_reload[18] ));
 sg13g2_o21ai_1 _25790_ (.B1(_10203_),
    .Y(_02497_),
    .A1(_06755_),
    .A2(net133));
 sg13g2_inv_1 _25791_ (.Y(_06756_),
    .A(\cpu.intr.r_timer_reload[19] ));
 sg13g2_o21ai_1 _25792_ (.B1(_10210_),
    .Y(_02498_),
    .A1(_06756_),
    .A2(net133));
 sg13g2_mux2_1 _25793_ (.A0(\cpu.intr.r_timer_reload[1] ),
    .A1(net921),
    .S(_06754_),
    .X(_02499_));
 sg13g2_inv_1 _25794_ (.Y(_06757_),
    .A(\cpu.intr.r_timer_reload[20] ));
 sg13g2_o21ai_1 _25795_ (.B1(_10216_),
    .Y(_02500_),
    .A1(_06757_),
    .A2(net133));
 sg13g2_inv_1 _25796_ (.Y(_06758_),
    .A(\cpu.intr.r_timer_reload[21] ));
 sg13g2_o21ai_1 _25797_ (.B1(_10222_),
    .Y(_02501_),
    .A1(_06758_),
    .A2(net133));
 sg13g2_inv_1 _25798_ (.Y(_06759_),
    .A(\cpu.intr.r_timer_reload[22] ));
 sg13g2_o21ai_1 _25799_ (.B1(_10228_),
    .Y(_02502_),
    .A1(_06759_),
    .A2(net133));
 sg13g2_mux2_1 _25800_ (.A0(\cpu.intr.r_timer_reload[23] ),
    .A1(net991),
    .S(net148),
    .X(_02503_));
 sg13g2_mux2_1 _25801_ (.A0(\cpu.intr.r_timer_reload[2] ),
    .A1(net917),
    .S(net123),
    .X(_02504_));
 sg13g2_mux2_1 _25802_ (.A0(\cpu.intr.r_timer_reload[3] ),
    .A1(_12232_),
    .S(_06754_),
    .X(_02505_));
 sg13g2_mux2_1 _25803_ (.A0(\cpu.intr.r_timer_reload[4] ),
    .A1(net1002),
    .S(_06753_),
    .X(_02506_));
 sg13g2_mux2_1 _25804_ (.A0(\cpu.intr.r_timer_reload[5] ),
    .A1(net1001),
    .S(_06753_),
    .X(_02507_));
 sg13g2_mux2_1 _25805_ (.A0(\cpu.intr.r_timer_reload[6] ),
    .A1(net1000),
    .S(_06753_),
    .X(_02508_));
 sg13g2_mux2_1 _25806_ (.A0(\cpu.intr.r_timer_reload[7] ),
    .A1(net991),
    .S(_06753_),
    .X(_02509_));
 sg13g2_mux2_1 _25807_ (.A0(\cpu.intr.r_timer_reload[8] ),
    .A1(_10302_),
    .S(_06753_),
    .X(_02510_));
 sg13g2_mux2_1 _25808_ (.A0(\cpu.intr.r_timer_reload[9] ),
    .A1(_10307_),
    .S(_06753_),
    .X(_02511_));
 sg13g2_inv_1 _25809_ (.Y(_06760_),
    .A(_09941_));
 sg13g2_nor4_2 _25810_ (.A(_12008_),
    .B(_12023_),
    .C(_09960_),
    .Y(_06761_),
    .D(_12006_));
 sg13g2_nor3_2 _25811_ (.A(_12024_),
    .B(_12009_),
    .C(_12003_),
    .Y(_06762_));
 sg13g2_nand2_1 _25812_ (.Y(_06763_),
    .A(_06761_),
    .B(_06762_));
 sg13g2_nor4_1 _25813_ (.A(_09948_),
    .B(_09938_),
    .C(_09936_),
    .D(_06763_),
    .Y(_06764_));
 sg13g2_o21ai_1 _25814_ (.B1(_06764_),
    .Y(_06765_),
    .A1(_09982_),
    .A2(_09983_));
 sg13g2_buf_1 _25815_ (.A(_06765_),
    .X(_06766_));
 sg13g2_inv_1 _25816_ (.Y(_06767_),
    .A(_10034_));
 sg13g2_and2_1 _25817_ (.A(\cpu.qspi.r_read_delay[1][0] ),
    .B(_09975_),
    .X(_06768_));
 sg13g2_a221oi_1 _25818_ (.B2(\cpu.qspi.r_read_delay[0][0] ),
    .C1(_06768_),
    .B1(_09979_),
    .A1(\cpu.qspi.r_read_delay[2][0] ),
    .Y(_06769_),
    .A2(_09977_));
 sg13g2_or4_1 _25819_ (.A(_09947_),
    .B(_09959_),
    .C(net1047),
    .D(_09950_),
    .X(_06770_));
 sg13g2_buf_1 _25820_ (.A(_06770_),
    .X(_06771_));
 sg13g2_a221oi_1 _25821_ (.B2(_06771_),
    .C1(_09954_),
    .B1(_00183_),
    .A1(net1119),
    .Y(_06772_),
    .A2(_06760_));
 sg13g2_o21ai_1 _25822_ (.B1(_06772_),
    .Y(_06773_),
    .A1(_06767_),
    .A2(_06769_));
 sg13g2_nor2_1 _25823_ (.A(net28),
    .B(_06773_),
    .Y(_06774_));
 sg13g2_a21oi_1 _25824_ (.A1(_06760_),
    .A2(net28),
    .Y(_02512_),
    .B1(_06774_));
 sg13g2_inv_1 _25825_ (.Y(_06775_),
    .A(_09942_));
 sg13g2_a22oi_1 _25826_ (.Y(_06776_),
    .B1(_09975_),
    .B2(\cpu.qspi.r_read_delay[1][1] ),
    .A2(_09977_),
    .A1(\cpu.qspi.r_read_delay[2][1] ));
 sg13g2_nand2_1 _25827_ (.Y(_06777_),
    .A(\cpu.qspi.r_read_delay[0][1] ),
    .B(_09979_));
 sg13g2_a21oi_1 _25828_ (.A1(_06776_),
    .A2(_06777_),
    .Y(_06778_),
    .B1(_06767_));
 sg13g2_xnor2_1 _25829_ (.Y(_06779_),
    .A(_09941_),
    .B(_09942_));
 sg13g2_nor2_1 _25830_ (.A(net1119),
    .B(_06771_),
    .Y(_06780_));
 sg13g2_mux2_1 _25831_ (.A0(_06779_),
    .A1(_06767_),
    .S(_06780_),
    .X(_06781_));
 sg13g2_nor4_1 _25832_ (.A(_09954_),
    .B(_06766_),
    .C(_06778_),
    .D(_06781_),
    .Y(_06782_));
 sg13g2_a21oi_1 _25833_ (.A1(_06775_),
    .A2(_06766_),
    .Y(_02513_),
    .B1(_06782_));
 sg13g2_inv_1 _25834_ (.Y(_06783_),
    .A(_09943_));
 sg13g2_nor2_1 _25835_ (.A(_09941_),
    .B(_09942_),
    .Y(_06784_));
 sg13g2_xor2_1 _25836_ (.B(_06784_),
    .A(_00184_),
    .X(_06785_));
 sg13g2_mux2_1 _25837_ (.A0(_06771_),
    .A1(net788),
    .S(net1119),
    .X(_06786_));
 sg13g2_a22oi_1 _25838_ (.Y(_06787_),
    .B1(_06785_),
    .B2(_06786_),
    .A2(_06780_),
    .A1(_10034_));
 sg13g2_a22oi_1 _25839_ (.Y(_06788_),
    .B1(_09975_),
    .B2(\cpu.qspi.r_read_delay[1][2] ),
    .A2(_09977_),
    .A1(\cpu.qspi.r_read_delay[2][2] ));
 sg13g2_nand2_1 _25840_ (.Y(_06789_),
    .A(\cpu.qspi.r_read_delay[0][2] ),
    .B(_09979_));
 sg13g2_a21oi_1 _25841_ (.A1(_06788_),
    .A2(_06789_),
    .Y(_06790_),
    .B1(_06767_));
 sg13g2_nor4_1 _25842_ (.A(_09954_),
    .B(net28),
    .C(_06787_),
    .D(_06790_),
    .Y(_06791_));
 sg13g2_a21oi_1 _25843_ (.A1(_06783_),
    .A2(net28),
    .Y(_02514_),
    .B1(_06791_));
 sg13g2_nand2b_1 _25844_ (.Y(_06792_),
    .B(net1119),
    .A_N(_09940_));
 sg13g2_nand2b_1 _25845_ (.Y(_06793_),
    .B(_06792_),
    .A_N(_06771_));
 sg13g2_a22oi_1 _25846_ (.Y(_06794_),
    .B1(_09975_),
    .B2(\cpu.qspi.r_read_delay[1][3] ),
    .A2(_09977_),
    .A1(\cpu.qspi.r_read_delay[2][3] ));
 sg13g2_nand2_1 _25847_ (.Y(_06795_),
    .A(\cpu.qspi.r_read_delay[0][3] ),
    .B(_09979_));
 sg13g2_nand2_1 _25848_ (.Y(_06796_),
    .A(_06794_),
    .B(_06795_));
 sg13g2_a22oi_1 _25849_ (.Y(_06797_),
    .B1(_06796_),
    .B2(_10034_),
    .A2(_06793_),
    .A1(_09944_));
 sg13g2_a21oi_1 _25850_ (.A1(_06783_),
    .A2(_06784_),
    .Y(_06798_),
    .B1(_06780_));
 sg13g2_o21ai_1 _25851_ (.B1(\cpu.qspi.r_count[3] ),
    .Y(_06799_),
    .A1(net28),
    .A2(_06798_));
 sg13g2_o21ai_1 _25852_ (.B1(_06799_),
    .Y(_02515_),
    .A1(net28),
    .A2(_06797_));
 sg13g2_nand3_1 _25853_ (.B(_09944_),
    .C(_06771_),
    .A(_09940_),
    .Y(_06800_));
 sg13g2_or3_1 _25854_ (.A(_09940_),
    .B(_09944_),
    .C(_06780_),
    .X(_06801_));
 sg13g2_a21oi_1 _25855_ (.A1(_06800_),
    .A2(_06801_),
    .Y(_06802_),
    .B1(net28));
 sg13g2_a21o_1 _25856_ (.A2(net28),
    .A1(\cpu.qspi.r_count[4] ),
    .B1(_06802_),
    .X(_02516_));
 sg13g2_nand2_1 _25857_ (.Y(_06803_),
    .A(_10124_),
    .B(_06385_));
 sg13g2_buf_1 _25858_ (.A(_06803_),
    .X(_06804_));
 sg13g2_nor2_1 _25859_ (.A(_09353_),
    .B(net110),
    .Y(_06805_));
 sg13g2_buf_1 _25860_ (.A(_06805_),
    .X(_06806_));
 sg13g2_nand2_1 _25861_ (.Y(_06807_),
    .A(net893),
    .B(_06806_));
 sg13g2_nand3_1 _25862_ (.B(_10124_),
    .C(_06385_),
    .A(_09382_),
    .Y(_06808_));
 sg13g2_buf_1 _25863_ (.A(_06808_),
    .X(_06809_));
 sg13g2_nand2_1 _25864_ (.Y(_06810_),
    .A(\cpu.qspi.r_read_delay[0][0] ),
    .B(_06809_));
 sg13g2_a21oi_1 _25865_ (.A1(_06807_),
    .A2(_06810_),
    .Y(_02527_),
    .B1(net630));
 sg13g2_nand2_1 _25866_ (.Y(_06811_),
    .A(_12694_),
    .B(_06806_));
 sg13g2_nand2_1 _25867_ (.Y(_06812_),
    .A(\cpu.qspi.r_read_delay[0][1] ),
    .B(_06809_));
 sg13g2_buf_2 _25868_ (.A(net804),
    .X(_06813_));
 sg13g2_buf_1 _25869_ (.A(_06813_),
    .X(_06814_));
 sg13g2_a21oi_1 _25870_ (.A1(_06811_),
    .A2(_06812_),
    .Y(_02528_),
    .B1(net577));
 sg13g2_nand2_1 _25871_ (.Y(_06815_),
    .A(net892),
    .B(_06806_));
 sg13g2_nand2_1 _25872_ (.Y(_06816_),
    .A(\cpu.qspi.r_read_delay[0][2] ),
    .B(_06809_));
 sg13g2_nand3_1 _25873_ (.B(_06815_),
    .C(_06816_),
    .A(net650),
    .Y(_02529_));
 sg13g2_nand2_1 _25874_ (.Y(_06817_),
    .A(_12751_),
    .B(_06806_));
 sg13g2_nand2_1 _25875_ (.Y(_06818_),
    .A(\cpu.qspi.r_read_delay[0][3] ),
    .B(_06809_));
 sg13g2_a21oi_1 _25876_ (.A1(_06817_),
    .A2(_06818_),
    .Y(_02530_),
    .B1(net577));
 sg13g2_nor2_1 _25877_ (.A(_10252_),
    .B(_06804_),
    .Y(_06819_));
 sg13g2_nand2_1 _25878_ (.Y(_06820_),
    .A(_12807_),
    .B(_06819_));
 sg13g2_nand3_1 _25879_ (.B(net515),
    .C(_06385_),
    .A(_10124_),
    .Y(_06821_));
 sg13g2_buf_1 _25880_ (.A(_06821_),
    .X(_06822_));
 sg13g2_nand2_1 _25881_ (.Y(_06823_),
    .A(\cpu.qspi.r_read_delay[1][0] ),
    .B(_06822_));
 sg13g2_a21oi_1 _25882_ (.A1(_06820_),
    .A2(_06823_),
    .Y(_02531_),
    .B1(_06814_));
 sg13g2_buf_1 _25883_ (.A(_10194_),
    .X(_06824_));
 sg13g2_nand2_1 _25884_ (.Y(_06825_),
    .A(_06824_),
    .B(_06819_));
 sg13g2_nand2_1 _25885_ (.Y(_06826_),
    .A(\cpu.qspi.r_read_delay[1][1] ),
    .B(_06822_));
 sg13g2_a21oi_1 _25886_ (.A1(_06825_),
    .A2(_06826_),
    .Y(_02532_),
    .B1(net577));
 sg13g2_nand2_1 _25887_ (.Y(_06827_),
    .A(_12814_),
    .B(_06819_));
 sg13g2_nand2_1 _25888_ (.Y(_06828_),
    .A(\cpu.qspi.r_read_delay[1][2] ),
    .B(_06822_));
 sg13g2_nand3_1 _25889_ (.B(_06827_),
    .C(_06828_),
    .A(net650),
    .Y(_02533_));
 sg13g2_nand2_1 _25890_ (.Y(_06829_),
    .A(net986),
    .B(_06819_));
 sg13g2_nand2_1 _25891_ (.Y(_06830_),
    .A(\cpu.qspi.r_read_delay[1][3] ),
    .B(_06822_));
 sg13g2_a21oi_1 _25892_ (.A1(_06829_),
    .A2(_06830_),
    .Y(_02534_),
    .B1(net577));
 sg13g2_nor2_1 _25893_ (.A(_04936_),
    .B(net110),
    .Y(_06831_));
 sg13g2_buf_1 _25894_ (.A(_06831_),
    .X(_06832_));
 sg13g2_nand2_1 _25895_ (.Y(_06833_),
    .A(_10241_),
    .B(_06832_));
 sg13g2_or2_1 _25896_ (.X(_06834_),
    .B(net110),
    .A(_04936_));
 sg13g2_buf_1 _25897_ (.A(_06834_),
    .X(_06835_));
 sg13g2_nand2_1 _25898_ (.Y(_06836_),
    .A(\cpu.qspi.r_read_delay[2][0] ),
    .B(_06835_));
 sg13g2_a21oi_1 _25899_ (.A1(_06833_),
    .A2(_06836_),
    .Y(_02535_),
    .B1(net577));
 sg13g2_nand2_1 _25900_ (.Y(_06837_),
    .A(net966),
    .B(_06832_));
 sg13g2_nand2_1 _25901_ (.Y(_06838_),
    .A(\cpu.qspi.r_read_delay[2][1] ),
    .B(_06835_));
 sg13g2_a21oi_1 _25902_ (.A1(_06837_),
    .A2(_06838_),
    .Y(_02536_),
    .B1(net577));
 sg13g2_nand2_1 _25903_ (.Y(_06839_),
    .A(_12814_),
    .B(_06832_));
 sg13g2_nand2_1 _25904_ (.Y(_06840_),
    .A(\cpu.qspi.r_read_delay[2][2] ),
    .B(_06835_));
 sg13g2_nand3_1 _25905_ (.B(_06839_),
    .C(_06840_),
    .A(net650),
    .Y(_02537_));
 sg13g2_nand2_1 _25906_ (.Y(_06841_),
    .A(_12751_),
    .B(_06832_));
 sg13g2_nand2_1 _25907_ (.Y(_06842_),
    .A(\cpu.qspi.r_read_delay[2][3] ),
    .B(_06835_));
 sg13g2_a21oi_1 _25908_ (.A1(_06841_),
    .A2(_06842_),
    .Y(_02538_),
    .B1(net577));
 sg13g2_buf_1 _25909_ (.A(net802),
    .X(_06843_));
 sg13g2_nand2_1 _25910_ (.Y(_06844_),
    .A(_09499_),
    .B(_09924_));
 sg13g2_buf_1 _25911_ (.A(_06844_),
    .X(_06845_));
 sg13g2_mux2_1 _25912_ (.A0(net406),
    .A1(_09706_),
    .S(net122),
    .X(_06846_));
 sg13g2_nand2_1 _25913_ (.Y(_06847_),
    .A(net644),
    .B(_06846_));
 sg13g2_o21ai_1 _25914_ (.B1(_06847_),
    .Y(_06848_),
    .A1(net644),
    .A2(_08660_));
 sg13g2_buf_1 _25915_ (.A(net1069),
    .X(_06849_));
 sg13g2_mux2_1 _25916_ (.A0(_09866_),
    .A1(_09874_),
    .S(_06845_),
    .X(_06850_));
 sg13g2_nand2b_1 _25917_ (.Y(_06851_),
    .B(net831),
    .A_N(_11317_));
 sg13g2_o21ai_1 _25918_ (.B1(_06851_),
    .Y(_06852_),
    .A1(net831),
    .A2(_06850_));
 sg13g2_a21oi_1 _25919_ (.A1(_09960_),
    .A2(_09956_),
    .Y(_06853_),
    .B1(_12008_));
 sg13g2_buf_1 _25920_ (.A(_12106_),
    .X(_06854_));
 sg13g2_a22oi_1 _25921_ (.Y(_06855_),
    .B1(_05189_),
    .B2(_12130_),
    .A2(_05182_),
    .A1(_12105_));
 sg13g2_nand3_1 _25922_ (.B(net1009),
    .C(_04840_),
    .A(net1008),
    .Y(_06856_));
 sg13g2_o21ai_1 _25923_ (.B1(_06856_),
    .Y(_06857_),
    .A1(net1008),
    .A2(_06855_));
 sg13g2_nand3_1 _25924_ (.B(net1009),
    .C(_04876_),
    .A(net1008),
    .Y(_06858_));
 sg13g2_nand3b_1 _25925_ (.B(_12105_),
    .C(_05517_),
    .Y(_06859_),
    .A_N(net1008));
 sg13g2_a21oi_1 _25926_ (.A1(_06858_),
    .A2(_06859_),
    .Y(_06860_),
    .B1(_06854_));
 sg13g2_a21oi_1 _25927_ (.A1(net965),
    .A2(_06857_),
    .Y(_06861_),
    .B1(_06860_));
 sg13g2_and2_1 _25928_ (.A(net1008),
    .B(net1007),
    .X(_06862_));
 sg13g2_nand2_1 _25929_ (.Y(_06863_),
    .A(_12106_),
    .B(_04847_));
 sg13g2_o21ai_1 _25930_ (.B1(_06863_),
    .Y(_06864_),
    .A1(net965),
    .A2(_04859_));
 sg13g2_nor2b_1 _25931_ (.A(_12237_),
    .B_N(_12130_),
    .Y(_06865_));
 sg13g2_nor2_1 _25932_ (.A(_12105_),
    .B(_06865_),
    .Y(_06866_));
 sg13g2_a22oi_1 _25933_ (.Y(_06867_),
    .B1(_06866_),
    .B2(_05526_),
    .A2(_06864_),
    .A1(_06862_));
 sg13g2_a21o_1 _25934_ (.A2(_06867_),
    .A1(_06861_),
    .B1(_12010_),
    .X(_06868_));
 sg13g2_inv_1 _25935_ (.Y(_06869_),
    .A(_09939_));
 sg13g2_buf_1 _25936_ (.A(\cpu.qspi.r_state[0] ),
    .X(_06870_));
 sg13g2_nand2_1 _25937_ (.Y(_06871_),
    .A(net1127),
    .B(net1069));
 sg13g2_o21ai_1 _25938_ (.B1(_06871_),
    .Y(_06872_),
    .A1(net1069),
    .A2(_12062_));
 sg13g2_nor2_1 _25939_ (.A(_09959_),
    .B(_09950_),
    .Y(_06873_));
 sg13g2_and2_1 _25940_ (.A(_06762_),
    .B(_06873_),
    .X(_06874_));
 sg13g2_nor2b_1 _25941_ (.A(_09962_),
    .B_N(_06761_),
    .Y(_06875_));
 sg13g2_and4_1 _25942_ (.A(_12005_),
    .B(_00277_),
    .C(_06874_),
    .D(_06875_),
    .X(_06876_));
 sg13g2_buf_1 _25943_ (.A(_06876_),
    .X(_06877_));
 sg13g2_a221oi_1 _25944_ (.B2(_12003_),
    .C1(_06877_),
    .B1(_06872_),
    .A1(_06869_),
    .Y(_06878_),
    .A2(_06870_));
 sg13g2_buf_1 _25945_ (.A(_06844_),
    .X(_06879_));
 sg13g2_mux2_1 _25946_ (.A0(net403),
    .A1(_09776_),
    .S(net121),
    .X(_06880_));
 sg13g2_nor2_1 _25947_ (.A(net802),
    .B(_08558_),
    .Y(_06881_));
 sg13g2_a21oi_1 _25948_ (.A1(_09485_),
    .A2(_06880_),
    .Y(_06882_),
    .B1(_06881_));
 sg13g2_nand2b_1 _25949_ (.Y(_06883_),
    .B(_12009_),
    .A_N(_06882_));
 sg13g2_nand4_1 _25950_ (.B(_06868_),
    .C(_06878_),
    .A(_06853_),
    .Y(_06884_),
    .D(_06883_));
 sg13g2_a221oi_1 _25951_ (.B2(_12023_),
    .C1(_06884_),
    .B1(_06852_),
    .A1(_12024_),
    .Y(_06885_),
    .A2(_06848_));
 sg13g2_nand2_1 _25952_ (.Y(_06886_),
    .A(_09962_),
    .B(_09939_));
 sg13g2_nand3_1 _25953_ (.B(_00183_),
    .C(_06886_),
    .A(_06775_),
    .Y(_06887_));
 sg13g2_nor2_1 _25954_ (.A(net1047),
    .B(_09956_),
    .Y(_06888_));
 sg13g2_o21ai_1 _25955_ (.B1(_09943_),
    .Y(_06889_),
    .A1(_06887_),
    .A2(_06888_));
 sg13g2_nand3_1 _25956_ (.B(_09942_),
    .C(_06886_),
    .A(_06760_),
    .Y(_06890_));
 sg13g2_o21ai_1 _25957_ (.B1(_06890_),
    .Y(_06891_),
    .A1(_06760_),
    .A2(_06886_));
 sg13g2_nor2_1 _25958_ (.A(_09943_),
    .B(_06891_),
    .Y(_06892_));
 sg13g2_o21ai_1 _25959_ (.B1(_06892_),
    .Y(_06893_),
    .A1(net1047),
    .A2(_09942_));
 sg13g2_o21ai_1 _25960_ (.B1(_06893_),
    .Y(_06894_),
    .A1(_09942_),
    .A2(_06889_));
 sg13g2_nor3_1 _25961_ (.A(net1047),
    .B(_09941_),
    .C(_06889_),
    .Y(_06895_));
 sg13g2_o21ai_1 _25962_ (.B1(_09956_),
    .Y(_06896_),
    .A1(_06892_),
    .A2(_06895_));
 sg13g2_nand2b_1 _25963_ (.Y(_06897_),
    .B(_06896_),
    .A_N(_06894_));
 sg13g2_o21ai_1 _25964_ (.B1(_06897_),
    .Y(_06898_),
    .A1(_09959_),
    .A2(net1047));
 sg13g2_xnor2_1 _25965_ (.Y(_06899_),
    .A(_09957_),
    .B(_09982_));
 sg13g2_a22oi_1 _25966_ (.Y(_06900_),
    .B1(_06899_),
    .B2(_06877_),
    .A2(_06898_),
    .A1(_06885_));
 sg13g2_and2_1 _25967_ (.A(\cpu.qspi.r_mask[1] ),
    .B(_09975_),
    .X(_06901_));
 sg13g2_a221oi_1 _25968_ (.B2(\cpu.qspi.r_mask[0] ),
    .C1(_06901_),
    .B1(_09979_),
    .A1(\cpu.qspi.r_mask[2] ),
    .Y(_06902_),
    .A2(_09977_));
 sg13g2_nand2_1 _25969_ (.Y(_06903_),
    .A(_12008_),
    .B(_06902_));
 sg13g2_nor2_1 _25970_ (.A(net1119),
    .B(_09936_),
    .Y(_06904_));
 sg13g2_nor3_2 _25971_ (.A(_09947_),
    .B(_09948_),
    .C(_09938_),
    .Y(_06905_));
 sg13g2_nand4_1 _25972_ (.B(_06903_),
    .C(_06904_),
    .A(_06767_),
    .Y(_06906_),
    .D(_06905_));
 sg13g2_buf_2 _25973_ (.A(_06906_),
    .X(_06907_));
 sg13g2_mux2_1 _25974_ (.A0(_06900_),
    .A1(net11),
    .S(_06907_),
    .X(_02543_));
 sg13g2_nor3_1 _25975_ (.A(_09954_),
    .B(net1047),
    .C(_09964_),
    .Y(_06908_));
 sg13g2_nand4_1 _25976_ (.B(_06762_),
    .C(_06873_),
    .A(_06761_),
    .Y(_06909_),
    .D(_06908_));
 sg13g2_mux2_1 _25977_ (.A0(net408),
    .A1(_09594_),
    .S(net122),
    .X(_06910_));
 sg13g2_nand2_1 _25978_ (.Y(_06911_),
    .A(net644),
    .B(_06910_));
 sg13g2_o21ai_1 _25979_ (.B1(_06911_),
    .Y(_06912_),
    .A1(net644),
    .A2(_08918_));
 sg13g2_buf_1 _25980_ (.A(net1069),
    .X(_06913_));
 sg13g2_nand2_1 _25981_ (.Y(_06914_),
    .A(net830),
    .B(_11316_));
 sg13g2_mux2_1 _25982_ (.A0(_00237_),
    .A1(_09864_),
    .S(_06879_),
    .X(_06915_));
 sg13g2_nand2_1 _25983_ (.Y(_06916_),
    .A(net644),
    .B(_06915_));
 sg13g2_nand3_1 _25984_ (.B(_06914_),
    .C(_06916_),
    .A(_12023_),
    .Y(_06917_));
 sg13g2_nor2b_1 _25985_ (.A(_05228_),
    .B_N(_12130_),
    .Y(_06918_));
 sg13g2_inv_1 _25986_ (.Y(_06919_),
    .A(_12105_));
 sg13g2_nor3_1 _25987_ (.A(_12106_),
    .B(_06919_),
    .C(_05600_),
    .Y(_06920_));
 sg13g2_a21oi_1 _25988_ (.A1(_06854_),
    .A2(_06918_),
    .Y(_06921_),
    .B1(_06920_));
 sg13g2_nand2_1 _25989_ (.Y(_06922_),
    .A(_12106_),
    .B(_05307_));
 sg13g2_o21ai_1 _25990_ (.B1(_06922_),
    .Y(_06923_),
    .A1(net965),
    .A2(_05299_));
 sg13g2_nand3_1 _25991_ (.B(net1009),
    .C(_06923_),
    .A(net1008),
    .Y(_06924_));
 sg13g2_o21ai_1 _25992_ (.B1(_06924_),
    .Y(_06925_),
    .A1(_12177_),
    .A2(_06921_));
 sg13g2_nand2_1 _25993_ (.Y(_06926_),
    .A(_05592_),
    .B(_06866_));
 sg13g2_nand3_1 _25994_ (.B(_12134_),
    .C(_05293_),
    .A(net1007),
    .Y(_06927_));
 sg13g2_nand2_1 _25995_ (.Y(_06928_),
    .A(net1099),
    .B(_05318_));
 sg13g2_o21ai_1 _25996_ (.B1(_06928_),
    .Y(_06929_),
    .A1(net1008),
    .A2(_05220_));
 sg13g2_nand3_1 _25997_ (.B(net1007),
    .C(_06929_),
    .A(net965),
    .Y(_06930_));
 sg13g2_nand3_1 _25998_ (.B(_06927_),
    .C(_06930_),
    .A(_06926_),
    .Y(_06931_));
 sg13g2_o21ai_1 _25999_ (.B1(_09950_),
    .Y(_06932_),
    .A1(_06925_),
    .A2(_06931_));
 sg13g2_nand2_1 _26000_ (.Y(_06933_),
    .A(_09783_),
    .B(net121));
 sg13g2_o21ai_1 _26001_ (.B1(_06933_),
    .Y(_06934_),
    .A1(net402),
    .A2(net122));
 sg13g2_nand2b_1 _26002_ (.Y(_06935_),
    .B(net1069),
    .A_N(_08634_));
 sg13g2_o21ai_1 _26003_ (.B1(_06935_),
    .Y(_06936_),
    .A1(net830),
    .A2(_06934_));
 sg13g2_mux2_1 _26004_ (.A0(_04887_),
    .A1(_09846_),
    .S(net121),
    .X(_06937_));
 sg13g2_nand2_1 _26005_ (.Y(_06938_),
    .A(_09485_),
    .B(_06937_));
 sg13g2_o21ai_1 _26006_ (.B1(_06938_),
    .Y(_06939_),
    .A1(net802),
    .A2(_11401_));
 sg13g2_a22oi_1 _26007_ (.Y(_06940_),
    .B1(_06939_),
    .B2(_12003_),
    .A2(_06936_),
    .A1(_12009_));
 sg13g2_nand4_1 _26008_ (.B(_06917_),
    .C(_06932_),
    .A(_06853_),
    .Y(_06941_),
    .D(_06940_));
 sg13g2_a21oi_1 _26009_ (.A1(_12024_),
    .A2(_06912_),
    .Y(_06942_),
    .B1(_06941_));
 sg13g2_o21ai_1 _26010_ (.B1(_06942_),
    .Y(_06943_),
    .A1(_09982_),
    .A2(_06909_));
 sg13g2_mux2_1 _26011_ (.A0(_06943_),
    .A1(net12),
    .S(_06907_),
    .X(_02544_));
 sg13g2_nand2_1 _26012_ (.Y(_06944_),
    .A(net712),
    .B(_06913_));
 sg13g2_nand2_1 _26013_ (.Y(_06945_),
    .A(net802),
    .B(net475));
 sg13g2_a21oi_1 _26014_ (.A1(_06944_),
    .A2(_06945_),
    .Y(_06946_),
    .B1(_00185_));
 sg13g2_mux2_1 _26015_ (.A0(_05259_),
    .A1(_05124_),
    .S(net1099),
    .X(_06947_));
 sg13g2_nand2_1 _26016_ (.Y(_06948_),
    .A(net1099),
    .B(_05118_));
 sg13g2_o21ai_1 _26017_ (.B1(_06948_),
    .Y(_06949_),
    .A1(net1099),
    .A2(_05253_));
 sg13g2_a22oi_1 _26018_ (.Y(_06950_),
    .B1(_06949_),
    .B2(net1007),
    .A2(_06947_),
    .A1(net1009));
 sg13g2_a22oi_1 _26019_ (.Y(_06951_),
    .B1(_05388_),
    .B2(_12130_),
    .A2(_05380_),
    .A1(_12105_));
 sg13g2_a21oi_1 _26020_ (.A1(_12105_),
    .A2(_05695_),
    .Y(_06952_),
    .B1(net1099));
 sg13g2_a21oi_1 _26021_ (.A1(net1008),
    .A2(_06951_),
    .Y(_06953_),
    .B1(_06952_));
 sg13g2_nor2_1 _26022_ (.A(net965),
    .B(_06953_),
    .Y(_06954_));
 sg13g2_a21oi_1 _26023_ (.A1(net965),
    .A2(_06950_),
    .Y(_06955_),
    .B1(_06954_));
 sg13g2_a21oi_1 _26024_ (.A1(_05706_),
    .A2(_06866_),
    .Y(_06956_),
    .B1(_06955_));
 sg13g2_nor2_1 _26025_ (.A(_12010_),
    .B(_06956_),
    .Y(_06957_));
 sg13g2_nor4_1 _26026_ (.A(_12008_),
    .B(_06877_),
    .C(_06946_),
    .D(_06957_),
    .Y(_06958_));
 sg13g2_mux2_1 _26027_ (.A0(net405),
    .A1(_09728_),
    .S(net121),
    .X(_06959_));
 sg13g2_nand2_1 _26028_ (.Y(_06960_),
    .A(net644),
    .B(_06959_));
 sg13g2_o21ai_1 _26029_ (.B1(_06960_),
    .Y(_06961_),
    .A1(net644),
    .A2(_08728_));
 sg13g2_mux2_1 _26030_ (.A0(net409),
    .A1(_09538_),
    .S(net121),
    .X(_06962_));
 sg13g2_nor2_1 _26031_ (.A(net830),
    .B(_06962_),
    .Y(_06963_));
 sg13g2_a21oi_1 _26032_ (.A1(net831),
    .A2(_09158_),
    .Y(_06964_),
    .B1(_06963_));
 sg13g2_a22oi_1 _26033_ (.Y(_06965_),
    .B1(_06964_),
    .B2(_12009_),
    .A2(_06961_),
    .A1(_12024_));
 sg13g2_nor2_1 _26034_ (.A(_00231_),
    .B(_06879_),
    .Y(_06966_));
 sg13g2_a21o_1 _26035_ (.A2(net122),
    .A1(_09817_),
    .B1(_06966_),
    .X(_06967_));
 sg13g2_mux2_1 _26036_ (.A0(_11407_),
    .A1(_06967_),
    .S(_06843_),
    .X(_06968_));
 sg13g2_mux2_1 _26037_ (.A0(_00239_),
    .A1(_09825_),
    .S(net122),
    .X(_06969_));
 sg13g2_nand2_1 _26038_ (.Y(_06970_),
    .A(net830),
    .B(_11292_));
 sg13g2_o21ai_1 _26039_ (.B1(_06970_),
    .Y(_06971_),
    .A1(net831),
    .A2(_06969_));
 sg13g2_a22oi_1 _26040_ (.Y(_06972_),
    .B1(_06971_),
    .B2(_12023_),
    .A2(_06968_),
    .A1(_12003_));
 sg13g2_and3_1 _26041_ (.X(_06973_),
    .A(_06958_),
    .B(_06965_),
    .C(_06972_));
 sg13g2_inv_1 _26042_ (.Y(_06974_),
    .A(_09982_));
 sg13g2_a21oi_1 _26043_ (.A1(_09956_),
    .A2(_06974_),
    .Y(_06975_),
    .B1(_06909_));
 sg13g2_nor3_1 _26044_ (.A(_06907_),
    .B(_06973_),
    .C(_06975_),
    .Y(_06976_));
 sg13g2_a21o_1 _26045_ (.A2(_06907_),
    .A1(net13),
    .B1(_06976_),
    .X(_02545_));
 sg13g2_mux2_1 _26046_ (.A0(_00233_),
    .A1(_09855_),
    .S(_06845_),
    .X(_06977_));
 sg13g2_nand2_1 _26047_ (.Y(_06978_),
    .A(net830),
    .B(_11430_));
 sg13g2_o21ai_1 _26048_ (.B1(_06978_),
    .Y(_06979_),
    .A1(net831),
    .A2(_06977_));
 sg13g2_mux2_1 _26049_ (.A0(_09649_),
    .A1(_09631_),
    .S(net121),
    .X(_06980_));
 sg13g2_nor2_1 _26050_ (.A(net830),
    .B(_06980_),
    .Y(_06981_));
 sg13g2_a21oi_1 _26051_ (.A1(net831),
    .A2(_08698_),
    .Y(_06982_),
    .B1(_06981_));
 sg13g2_a22oi_1 _26052_ (.Y(_06983_),
    .B1(_06982_),
    .B2(_12009_),
    .A2(_06979_),
    .A1(_12003_));
 sg13g2_nand2_1 _26053_ (.Y(_06984_),
    .A(_09621_),
    .B(net121));
 sg13g2_o21ai_1 _26054_ (.B1(_06984_),
    .Y(_06985_),
    .A1(_09968_),
    .A2(net121));
 sg13g2_inv_1 _26055_ (.Y(_06986_),
    .A(_06985_));
 sg13g2_o21ai_1 _26056_ (.B1(_09969_),
    .Y(_06987_),
    .A1(net830),
    .A2(_06986_));
 sg13g2_nand4_1 _26057_ (.B(_09966_),
    .C(_12006_),
    .A(_09967_),
    .Y(_06988_),
    .D(_06987_));
 sg13g2_nor2_1 _26058_ (.A(net644),
    .B(_08896_),
    .Y(_06989_));
 sg13g2_nand2_1 _26059_ (.Y(_06990_),
    .A(_09677_),
    .B(net122));
 sg13g2_o21ai_1 _26060_ (.B1(_06990_),
    .Y(_06991_),
    .A1(_09666_),
    .A2(net122));
 sg13g2_nor2_1 _26061_ (.A(net831),
    .B(_06991_),
    .Y(_06992_));
 sg13g2_o21ai_1 _26062_ (.B1(_12024_),
    .Y(_06993_),
    .A1(_06989_),
    .A2(_06992_));
 sg13g2_mux2_1 _26063_ (.A0(_00241_),
    .A1(_09807_),
    .S(net122),
    .X(_06994_));
 sg13g2_nand2_1 _26064_ (.Y(_06995_),
    .A(net830),
    .B(_11273_));
 sg13g2_o21ai_1 _26065_ (.B1(_06995_),
    .Y(_06996_),
    .A1(_06913_),
    .A2(_06994_));
 sg13g2_mux4_1 _26066_ (.S0(net1099),
    .A0(_05090_),
    .A1(_05456_),
    .A2(_05084_),
    .A3(_05159_),
    .S1(net965),
    .X(_06997_));
 sg13g2_mux2_1 _26067_ (.A0(_05100_),
    .A1(_05151_),
    .S(net1099),
    .X(_06998_));
 sg13g2_a22oi_1 _26068_ (.Y(_06999_),
    .B1(_06998_),
    .B2(net965),
    .A2(_05449_),
    .A1(_12134_));
 sg13g2_nor2b_1 _26069_ (.A(_06999_),
    .B_N(net1009),
    .Y(_07000_));
 sg13g2_a221oi_1 _26070_ (.B2(net1007),
    .C1(_07000_),
    .B1(_06997_),
    .A1(_05075_),
    .Y(_07001_),
    .A2(_06866_));
 sg13g2_nand2_1 _26071_ (.Y(_07002_),
    .A(net711),
    .B(net1069));
 sg13g2_nand2_1 _26072_ (.Y(_07003_),
    .A(net802),
    .B(net437));
 sg13g2_a21oi_1 _26073_ (.A1(_07002_),
    .A2(_07003_),
    .Y(_07004_),
    .B1(_00185_));
 sg13g2_nor4_1 _26074_ (.A(_12008_),
    .B(_09960_),
    .C(_06877_),
    .D(_07004_),
    .Y(_07005_));
 sg13g2_o21ai_1 _26075_ (.B1(_07005_),
    .Y(_07006_),
    .A1(_12010_),
    .A2(_07001_));
 sg13g2_a21oi_1 _26076_ (.A1(_12023_),
    .A2(_06996_),
    .Y(_07007_),
    .B1(_07006_));
 sg13g2_and4_1 _26077_ (.A(_06983_),
    .B(_06988_),
    .C(_06993_),
    .D(_07007_),
    .X(_07008_));
 sg13g2_nor3_1 _26078_ (.A(_06907_),
    .B(_06975_),
    .C(_07008_),
    .Y(_07009_));
 sg13g2_a21o_1 _26079_ (.A2(_06907_),
    .A1(net14),
    .B1(_07009_),
    .X(_02546_));
 sg13g2_mux4_1 _26080_ (.S0(_05540_),
    .A0(_09304_),
    .A1(_09310_),
    .A2(_09299_),
    .A3(_09290_),
    .S1(_06397_),
    .X(_07010_));
 sg13g2_mux4_1 _26081_ (.S0(_05540_),
    .A0(_09288_),
    .A1(_09302_),
    .A2(_09308_),
    .A3(_09297_),
    .S1(_06397_),
    .X(_07011_));
 sg13g2_nor2b_1 _26082_ (.A(\cpu.gpio.r_spi_miso_src[1][2] ),
    .B_N(_07011_),
    .Y(_07012_));
 sg13g2_a21oi_1 _26083_ (.A1(\cpu.gpio.r_spi_miso_src[1][2] ),
    .A2(_07010_),
    .Y(_07013_),
    .B1(_07012_));
 sg13g2_mux4_1 _26084_ (.S0(_05540_),
    .A0(_09292_),
    .A1(_09313_),
    .A2(_09315_),
    .A3(_09294_),
    .S1(_06397_),
    .X(_07014_));
 sg13g2_nand3b_1 _26085_ (.B(\cpu.gpio.r_spi_miso_src[1][3] ),
    .C(_07014_),
    .Y(_07015_),
    .A_N(_00150_));
 sg13g2_o21ai_1 _26086_ (.B1(_07015_),
    .Y(_07016_),
    .A1(\cpu.gpio.r_spi_miso_src[1][3] ),
    .A2(_07013_));
 sg13g2_mux4_1 _26087_ (.S0(_04981_),
    .A0(_09304_),
    .A1(_09310_),
    .A2(_09299_),
    .A3(_09290_),
    .S1(_06396_),
    .X(_07017_));
 sg13g2_mux4_1 _26088_ (.S0(_04981_),
    .A0(_09288_),
    .A1(_09302_),
    .A2(_09308_),
    .A3(_09297_),
    .S1(_06396_),
    .X(_07018_));
 sg13g2_nor2b_1 _26089_ (.A(\cpu.gpio.r_spi_miso_src[0][2] ),
    .B_N(_07018_),
    .Y(_07019_));
 sg13g2_a21oi_1 _26090_ (.A1(\cpu.gpio.r_spi_miso_src[0][2] ),
    .A2(_07017_),
    .Y(_07020_),
    .B1(_07019_));
 sg13g2_mux4_1 _26091_ (.S0(_04981_),
    .A0(_09292_),
    .A1(_09313_),
    .A2(_09315_),
    .A3(_09294_),
    .S1(_06396_),
    .X(_07021_));
 sg13g2_nand3b_1 _26092_ (.B(\cpu.gpio.r_spi_miso_src[0][3] ),
    .C(_07021_),
    .Y(_07022_),
    .A_N(_00110_));
 sg13g2_o21ai_1 _26093_ (.B1(_07022_),
    .Y(_07023_),
    .A1(\cpu.gpio.r_spi_miso_src[0][3] ),
    .A2(_07020_));
 sg13g2_mux2_1 _26094_ (.A0(_07016_),
    .A1(_07023_),
    .S(_12045_),
    .X(_07024_));
 sg13g2_nor2_1 _26095_ (.A(net1123),
    .B(_12090_),
    .Y(_07025_));
 sg13g2_nor2b_1 _26096_ (.A(_09430_),
    .B_N(_09440_),
    .Y(_07026_));
 sg13g2_a22oi_1 _26097_ (.Y(_07027_),
    .B1(_07026_),
    .B2(net608),
    .A2(_07025_),
    .A1(_09430_));
 sg13g2_nor3_1 _26098_ (.A(net931),
    .B(net447),
    .C(_07027_),
    .Y(_07028_));
 sg13g2_buf_4 _26099_ (.X(_07029_),
    .A(_07028_));
 sg13g2_mux2_1 _26100_ (.A0(_09417_),
    .A1(_07024_),
    .S(_07029_),
    .X(_02586_));
 sg13g2_mux2_1 _26101_ (.A0(_09416_),
    .A1(_09417_),
    .S(_07029_),
    .X(_02587_));
 sg13g2_mux2_1 _26102_ (.A0(_09420_),
    .A1(_09416_),
    .S(_07029_),
    .X(_02588_));
 sg13g2_mux2_1 _26103_ (.A0(_09414_),
    .A1(_09420_),
    .S(_07029_),
    .X(_02589_));
 sg13g2_mux2_1 _26104_ (.A0(_09422_),
    .A1(_09414_),
    .S(_07029_),
    .X(_02590_));
 sg13g2_mux2_1 _26105_ (.A0(_09421_),
    .A1(_09422_),
    .S(_07029_),
    .X(_02591_));
 sg13g2_mux2_1 _26106_ (.A0(_09415_),
    .A1(_09421_),
    .S(_07029_),
    .X(_02592_));
 sg13g2_mux2_1 _26107_ (.A0(\cpu.spi.r_in[7] ),
    .A1(_09415_),
    .S(_07029_),
    .X(_02593_));
 sg13g2_buf_1 _26108_ (.A(_00225_),
    .X(_07030_));
 sg13g2_buf_1 _26109_ (.A(_07030_),
    .X(_07031_));
 sg13g2_nor2b_1 _26110_ (.A(net608),
    .B_N(_00223_),
    .Y(_07032_));
 sg13g2_buf_1 _26111_ (.A(net1124),
    .X(_07033_));
 sg13g2_o21ai_1 _26112_ (.B1(_07033_),
    .Y(_07034_),
    .A1(_07031_),
    .A2(_07032_));
 sg13g2_o21ai_1 _26113_ (.B1(_07034_),
    .Y(_07035_),
    .A1(_09432_),
    .A2(net1041));
 sg13g2_nand2_1 _26114_ (.Y(_07036_),
    .A(_12032_),
    .B(_07035_));
 sg13g2_nand2_1 _26115_ (.Y(_07037_),
    .A(_09394_),
    .B(_12090_));
 sg13g2_nor2_1 _26116_ (.A(net1124),
    .B(net898),
    .Y(_07038_));
 sg13g2_buf_2 _26117_ (.A(_07038_),
    .X(_07039_));
 sg13g2_a221oi_1 _26118_ (.B2(_12026_),
    .C1(_12095_),
    .B1(_07039_),
    .A1(_09436_),
    .Y(_07040_),
    .A2(_07037_));
 sg13g2_o21ai_1 _26119_ (.B1(_09383_),
    .Y(_07041_),
    .A1(_09377_),
    .A2(_09374_));
 sg13g2_and2_1 _26120_ (.A(_07040_),
    .B(_07041_),
    .X(_07042_));
 sg13g2_buf_4 _26121_ (.X(_07043_),
    .A(_07042_));
 sg13g2_mux2_1 _26122_ (.A0(\cpu.spi.r_out[0] ),
    .A1(_07036_),
    .S(_07043_),
    .X(_02601_));
 sg13g2_buf_1 _26123_ (.A(_09366_),
    .X(_07044_));
 sg13g2_mux2_1 _26124_ (.A0(_00178_),
    .A1(_00223_),
    .S(net608),
    .X(_07045_));
 sg13g2_a22oi_1 _26125_ (.Y(_07046_),
    .B1(_07039_),
    .B2(_10194_),
    .A2(net898),
    .A1(\cpu.spi.r_out[0] ));
 sg13g2_o21ai_1 _26126_ (.B1(_07046_),
    .Y(_07047_),
    .A1(net829),
    .A2(_07045_));
 sg13g2_mux2_1 _26127_ (.A0(\cpu.spi.r_out[1] ),
    .A1(_07047_),
    .S(_07043_),
    .X(_02602_));
 sg13g2_mux2_1 _26128_ (.A0(_00179_),
    .A1(_00178_),
    .S(net608),
    .X(_07048_));
 sg13g2_a22oi_1 _26129_ (.Y(_07049_),
    .B1(_07039_),
    .B2(net1039),
    .A2(net898),
    .A1(\cpu.spi.r_out[1] ));
 sg13g2_o21ai_1 _26130_ (.B1(_07049_),
    .Y(_07050_),
    .A1(net829),
    .A2(_07048_));
 sg13g2_mux2_1 _26131_ (.A0(\cpu.spi.r_out[2] ),
    .A1(_07050_),
    .S(_07043_),
    .X(_02603_));
 sg13g2_mux2_1 _26132_ (.A0(_00287_),
    .A1(_00179_),
    .S(net608),
    .X(_07051_));
 sg13g2_a22oi_1 _26133_ (.Y(_07052_),
    .B1(_07039_),
    .B2(net1116),
    .A2(net898),
    .A1(\cpu.spi.r_out[2] ));
 sg13g2_o21ai_1 _26134_ (.B1(_07052_),
    .Y(_07053_),
    .A1(net829),
    .A2(_07051_));
 sg13g2_mux2_1 _26135_ (.A0(\cpu.spi.r_out[3] ),
    .A1(_07053_),
    .S(_07043_),
    .X(_02604_));
 sg13g2_mux2_1 _26136_ (.A0(_00180_),
    .A1(_00287_),
    .S(net608),
    .X(_07054_));
 sg13g2_a22oi_1 _26137_ (.Y(_07055_),
    .B1(_07039_),
    .B2(_10214_),
    .A2(net898),
    .A1(\cpu.spi.r_out[3] ));
 sg13g2_o21ai_1 _26138_ (.B1(_07055_),
    .Y(_07056_),
    .A1(net829),
    .A2(_07054_));
 sg13g2_mux2_1 _26139_ (.A0(\cpu.spi.r_out[4] ),
    .A1(_07056_),
    .S(_07043_),
    .X(_02605_));
 sg13g2_mux2_1 _26140_ (.A0(_00181_),
    .A1(_00180_),
    .S(net608),
    .X(_07057_));
 sg13g2_a22oi_1 _26141_ (.Y(_07058_),
    .B1(_07039_),
    .B2(_10220_),
    .A2(net898),
    .A1(\cpu.spi.r_out[4] ));
 sg13g2_o21ai_1 _26142_ (.B1(_07058_),
    .Y(_07059_),
    .A1(net829),
    .A2(_07057_));
 sg13g2_mux2_1 _26143_ (.A0(\cpu.spi.r_out[5] ),
    .A1(_07059_),
    .S(_07043_),
    .X(_02606_));
 sg13g2_buf_1 _26144_ (.A(_00182_),
    .X(_07060_));
 sg13g2_mux2_1 _26145_ (.A0(_07060_),
    .A1(_00181_),
    .S(_12096_),
    .X(_07061_));
 sg13g2_a22oi_1 _26146_ (.Y(_07062_),
    .B1(_07039_),
    .B2(_10226_),
    .A2(net898),
    .A1(\cpu.spi.r_out[5] ));
 sg13g2_o21ai_1 _26147_ (.B1(_07062_),
    .Y(_07063_),
    .A1(_07044_),
    .A2(_07061_));
 sg13g2_mux2_1 _26148_ (.A0(\cpu.spi.r_out[6] ),
    .A1(_07063_),
    .S(_07043_),
    .X(_02607_));
 sg13g2_buf_1 _26149_ (.A(_00281_),
    .X(_07064_));
 sg13g2_mux2_1 _26150_ (.A0(_07064_),
    .A1(_07060_),
    .S(_12096_),
    .X(_07065_));
 sg13g2_a22oi_1 _26151_ (.Y(_07066_),
    .B1(_07039_),
    .B2(_10229_),
    .A2(_12080_),
    .A1(\cpu.spi.r_out[6] ));
 sg13g2_o21ai_1 _26152_ (.B1(_07066_),
    .Y(_07067_),
    .A1(_07044_),
    .A2(_07065_));
 sg13g2_mux2_1 _26153_ (.A0(\cpu.spi.r_out[7] ),
    .A1(_07067_),
    .S(_07043_),
    .X(_02608_));
 sg13g2_nand3_1 _26154_ (.B(net930),
    .C(_09448_),
    .A(_09377_),
    .Y(_07068_));
 sg13g2_buf_1 _26155_ (.A(_07068_),
    .X(_07069_));
 sg13g2_nand2_1 _26156_ (.Y(_07070_),
    .A(net900),
    .B(_07069_));
 sg13g2_o21ai_1 _26157_ (.B1(_07070_),
    .Y(_02611_),
    .A1(net656),
    .A2(_07069_));
 sg13g2_nand2_1 _26158_ (.Y(_07071_),
    .A(_12034_),
    .B(_07069_));
 sg13g2_o21ai_1 _26159_ (.B1(_07071_),
    .Y(_02612_),
    .A1(_02943_),
    .A2(_07069_));
 sg13g2_nand2b_1 _26160_ (.Y(_07072_),
    .B(_04905_),
    .A_N(_09370_));
 sg13g2_buf_4 _26161_ (.X(_07073_),
    .A(_07072_));
 sg13g2_mux2_1 _26162_ (.A0(net897),
    .A1(\cpu.spi.r_timeout[0] ),
    .S(_07073_),
    .X(_02616_));
 sg13g2_mux2_1 _26163_ (.A0(net918),
    .A1(\cpu.spi.r_timeout[1] ),
    .S(_07073_),
    .X(_02617_));
 sg13g2_mux2_1 _26164_ (.A0(_10264_),
    .A1(\cpu.spi.r_timeout[2] ),
    .S(_07073_),
    .X(_02618_));
 sg13g2_mux2_1 _26165_ (.A0(net1033),
    .A1(\cpu.spi.r_timeout[3] ),
    .S(_07073_),
    .X(_02619_));
 sg13g2_mux2_1 _26166_ (.A0(net1002),
    .A1(\cpu.spi.r_timeout[4] ),
    .S(_07073_),
    .X(_02620_));
 sg13g2_mux2_1 _26167_ (.A0(net1001),
    .A1(\cpu.spi.r_timeout[5] ),
    .S(_07073_),
    .X(_02621_));
 sg13g2_mux2_1 _26168_ (.A0(net1000),
    .A1(\cpu.spi.r_timeout[6] ),
    .S(_07073_),
    .X(_02622_));
 sg13g2_mux2_1 _26169_ (.A0(net991),
    .A1(\cpu.spi.r_timeout[7] ),
    .S(_07073_),
    .X(_02623_));
 sg13g2_nand2_1 _26170_ (.Y(_07074_),
    .A(net1124),
    .B(_09372_));
 sg13g2_inv_1 _26171_ (.Y(_07075_),
    .A(_09426_));
 sg13g2_nor2_1 _26172_ (.A(_09437_),
    .B(_07075_),
    .Y(_07076_));
 sg13g2_nor3_1 _26173_ (.A(_00226_),
    .B(_09397_),
    .C(_09426_),
    .Y(_07077_));
 sg13g2_nor3_1 _26174_ (.A(net497),
    .B(_07076_),
    .C(_07077_),
    .Y(_07078_));
 sg13g2_a21oi_1 _26175_ (.A1(_09437_),
    .A2(net497),
    .Y(_07079_),
    .B1(_07078_));
 sg13g2_nand3_1 _26176_ (.B(_09429_),
    .C(_07078_),
    .A(_09366_),
    .Y(_07080_));
 sg13g2_o21ai_1 _26177_ (.B1(_07080_),
    .Y(_07081_),
    .A1(_07074_),
    .A2(_07079_));
 sg13g2_nand2_1 _26178_ (.Y(_07082_),
    .A(net930),
    .B(_07081_));
 sg13g2_buf_2 _26179_ (.A(_07082_),
    .X(_07083_));
 sg13g2_buf_1 _26180_ (.A(_07083_),
    .X(_07084_));
 sg13g2_and2_1 _26181_ (.A(net963),
    .B(\cpu.spi.r_timeout[0] ),
    .X(_07085_));
 sg13g2_a21oi_1 _26182_ (.A1(net829),
    .A2(_00284_),
    .Y(_07086_),
    .B1(_07085_));
 sg13g2_nand2_1 _26183_ (.Y(_07087_),
    .A(_09399_),
    .B(net33));
 sg13g2_o21ai_1 _26184_ (.B1(_07087_),
    .Y(_02624_),
    .A1(net33),
    .A2(_07086_));
 sg13g2_nor3_1 _26185_ (.A(_09399_),
    .B(_09400_),
    .C(_07083_),
    .Y(_07088_));
 sg13g2_a21oi_1 _26186_ (.A1(_09399_),
    .A2(_09400_),
    .Y(_07089_),
    .B1(_07088_));
 sg13g2_nor2_1 _26187_ (.A(net829),
    .B(_07083_),
    .Y(_07090_));
 sg13g2_buf_2 _26188_ (.A(_07090_),
    .X(_07091_));
 sg13g2_a22oi_1 _26189_ (.Y(_07092_),
    .B1(_07091_),
    .B2(\cpu.spi.r_timeout[1] ),
    .A2(net33),
    .A1(_09400_));
 sg13g2_o21ai_1 _26190_ (.B1(_07092_),
    .Y(_02625_),
    .A1(net1049),
    .A2(_07089_));
 sg13g2_o21ai_1 _26191_ (.B1(\cpu.spi.r_timeout_count[2] ),
    .Y(_07093_),
    .A1(_09399_),
    .A2(_09400_));
 sg13g2_o21ai_1 _26192_ (.B1(_07093_),
    .Y(_07094_),
    .A1(_09402_),
    .A2(net33));
 sg13g2_nand2_1 _26193_ (.Y(_07095_),
    .A(net829),
    .B(_07094_));
 sg13g2_a22oi_1 _26194_ (.Y(_07096_),
    .B1(_07091_),
    .B2(\cpu.spi.r_timeout[2] ),
    .A2(net33),
    .A1(\cpu.spi.r_timeout_count[2] ));
 sg13g2_nand2_1 _26195_ (.Y(_02626_),
    .A(_07095_),
    .B(_07096_));
 sg13g2_nor2_1 _26196_ (.A(_09404_),
    .B(_07083_),
    .Y(_07097_));
 sg13g2_a21oi_1 _26197_ (.A1(\cpu.spi.r_timeout_count[3] ),
    .A2(_09402_),
    .Y(_07098_),
    .B1(_07097_));
 sg13g2_a22oi_1 _26198_ (.Y(_07099_),
    .B1(_07091_),
    .B2(\cpu.spi.r_timeout[3] ),
    .A2(_07084_),
    .A1(\cpu.spi.r_timeout_count[3] ));
 sg13g2_o21ai_1 _26199_ (.B1(_07099_),
    .Y(_02627_),
    .A1(net1049),
    .A2(_07098_));
 sg13g2_nor2_1 _26200_ (.A(_09406_),
    .B(_07083_),
    .Y(_07100_));
 sg13g2_a21oi_1 _26201_ (.A1(\cpu.spi.r_timeout_count[4] ),
    .A2(_09404_),
    .Y(_07101_),
    .B1(_07100_));
 sg13g2_a22oi_1 _26202_ (.Y(_07102_),
    .B1(_07091_),
    .B2(\cpu.spi.r_timeout[4] ),
    .A2(net33),
    .A1(\cpu.spi.r_timeout_count[4] ));
 sg13g2_o21ai_1 _26203_ (.B1(_07102_),
    .Y(_02628_),
    .A1(net1049),
    .A2(_07101_));
 sg13g2_nor2_1 _26204_ (.A(_09408_),
    .B(_07083_),
    .Y(_07103_));
 sg13g2_a21oi_1 _26205_ (.A1(\cpu.spi.r_timeout_count[5] ),
    .A2(_09406_),
    .Y(_07104_),
    .B1(_07103_));
 sg13g2_a22oi_1 _26206_ (.Y(_07105_),
    .B1(_07091_),
    .B2(\cpu.spi.r_timeout[5] ),
    .A2(_07084_),
    .A1(\cpu.spi.r_timeout_count[5] ));
 sg13g2_o21ai_1 _26207_ (.B1(_07105_),
    .Y(_02629_),
    .A1(net1049),
    .A2(_07104_));
 sg13g2_nor2_1 _26208_ (.A(_09410_),
    .B(_07083_),
    .Y(_07106_));
 sg13g2_a21oi_1 _26209_ (.A1(\cpu.spi.r_timeout_count[6] ),
    .A2(_09408_),
    .Y(_07107_),
    .B1(_07106_));
 sg13g2_a22oi_1 _26210_ (.Y(_07108_),
    .B1(_07091_),
    .B2(\cpu.spi.r_timeout[6] ),
    .A2(net33),
    .A1(\cpu.spi.r_timeout_count[6] ));
 sg13g2_o21ai_1 _26211_ (.B1(_07108_),
    .Y(_02630_),
    .A1(net1049),
    .A2(_07107_));
 sg13g2_nor3_1 _26212_ (.A(_09398_),
    .B(_09410_),
    .C(_07083_),
    .Y(_07109_));
 sg13g2_a21oi_1 _26213_ (.A1(_09398_),
    .A2(_09410_),
    .Y(_07110_),
    .B1(_07109_));
 sg13g2_a22oi_1 _26214_ (.Y(_07111_),
    .B1(_07091_),
    .B2(\cpu.spi.r_timeout[7] ),
    .A2(net33),
    .A1(_09398_));
 sg13g2_o21ai_1 _26215_ (.B1(_07111_),
    .Y(_02631_),
    .A1(net1049),
    .A2(_07110_));
 sg13g2_buf_1 _26216_ (.A(\cpu.uart.r_rcnt[0] ),
    .X(_07112_));
 sg13g2_nor2_1 _26217_ (.A(_07112_),
    .B(\cpu.uart.r_rcnt[1] ),
    .Y(_07113_));
 sg13g2_nand2_1 _26218_ (.Y(_07114_),
    .A(net348),
    .B(_07113_));
 sg13g2_nor2_1 _26219_ (.A(net931),
    .B(_07114_),
    .Y(_07115_));
 sg13g2_buf_1 _26220_ (.A(\cpu.uart.r_rstate[3] ),
    .X(_07116_));
 sg13g2_buf_1 _26221_ (.A(net1082),
    .X(_07117_));
 sg13g2_buf_1 _26222_ (.A(\cpu.uart.r_rstate[1] ),
    .X(_07118_));
 sg13g2_buf_1 _26223_ (.A(\cpu.uart.r_rstate[2] ),
    .X(_07119_));
 sg13g2_buf_1 _26224_ (.A(_07119_),
    .X(_07120_));
 sg13g2_nor2_2 _26225_ (.A(net1081),
    .B(net961),
    .Y(_07121_));
 sg13g2_buf_2 _26226_ (.A(\cpu.uart.r_rstate[0] ),
    .X(_07122_));
 sg13g2_inv_1 _26227_ (.Y(_07123_),
    .A(_07122_));
 sg13g2_nand3_1 _26228_ (.B(net962),
    .C(_07121_),
    .A(_07123_),
    .Y(_07124_));
 sg13g2_o21ai_1 _26229_ (.B1(_07124_),
    .Y(_07125_),
    .A1(net962),
    .A2(_07121_));
 sg13g2_and2_1 _26230_ (.A(_07115_),
    .B(_07125_),
    .X(_07126_));
 sg13g2_buf_2 _26231_ (.A(_07126_),
    .X(_07127_));
 sg13g2_mux2_1 _26232_ (.A0(\cpu.uart.r_ib[0] ),
    .A1(\cpu.uart.r_ib[1] ),
    .S(_07127_),
    .X(_02644_));
 sg13g2_mux2_1 _26233_ (.A0(\cpu.uart.r_ib[1] ),
    .A1(\cpu.uart.r_ib[2] ),
    .S(_07127_),
    .X(_02645_));
 sg13g2_mux2_1 _26234_ (.A0(\cpu.uart.r_ib[2] ),
    .A1(\cpu.uart.r_ib[3] ),
    .S(_07127_),
    .X(_02646_));
 sg13g2_mux2_1 _26235_ (.A0(\cpu.uart.r_ib[3] ),
    .A1(\cpu.uart.r_ib[4] ),
    .S(_07127_),
    .X(_02647_));
 sg13g2_mux2_1 _26236_ (.A0(\cpu.uart.r_ib[4] ),
    .A1(\cpu.uart.r_ib[5] ),
    .S(_07127_),
    .X(_02648_));
 sg13g2_mux2_1 _26237_ (.A0(\cpu.uart.r_ib[5] ),
    .A1(\cpu.uart.r_ib[6] ),
    .S(_07127_),
    .X(_02649_));
 sg13g2_xor2_1 _26238_ (.B(\cpu.uart.r_r ),
    .A(\cpu.uart.r_r_invert ),
    .X(_07128_));
 sg13g2_mux2_1 _26239_ (.A0(\cpu.uart.r_ib[6] ),
    .A1(_07128_),
    .S(_07127_),
    .X(_02650_));
 sg13g2_and4_1 _26240_ (.A(_07122_),
    .B(net962),
    .C(_07115_),
    .D(_07121_),
    .X(_07129_));
 sg13g2_buf_1 _26241_ (.A(_07129_),
    .X(_07130_));
 sg13g2_mux2_1 _26242_ (.A0(\cpu.uart.r_in[0] ),
    .A1(\cpu.uart.r_ib[0] ),
    .S(net154),
    .X(_02651_));
 sg13g2_mux2_1 _26243_ (.A0(\cpu.uart.r_in[1] ),
    .A1(\cpu.uart.r_ib[1] ),
    .S(net154),
    .X(_02652_));
 sg13g2_mux2_1 _26244_ (.A0(\cpu.uart.r_in[2] ),
    .A1(\cpu.uart.r_ib[2] ),
    .S(net154),
    .X(_02653_));
 sg13g2_mux2_1 _26245_ (.A0(\cpu.uart.r_in[3] ),
    .A1(\cpu.uart.r_ib[3] ),
    .S(net154),
    .X(_02654_));
 sg13g2_mux2_1 _26246_ (.A0(\cpu.uart.r_in[4] ),
    .A1(\cpu.uart.r_ib[4] ),
    .S(net154),
    .X(_02655_));
 sg13g2_mux2_1 _26247_ (.A0(\cpu.uart.r_in[5] ),
    .A1(\cpu.uart.r_ib[5] ),
    .S(net154),
    .X(_02656_));
 sg13g2_mux2_1 _26248_ (.A0(\cpu.uart.r_in[6] ),
    .A1(\cpu.uart.r_ib[6] ),
    .S(net154),
    .X(_02657_));
 sg13g2_mux2_1 _26249_ (.A0(\cpu.uart.r_in[7] ),
    .A1(_07128_),
    .S(net154),
    .X(_02658_));
 sg13g2_buf_2 _26250_ (.A(\cpu.uart.r_xstate[2] ),
    .X(_07131_));
 sg13g2_buf_1 _26251_ (.A(_07131_),
    .X(_07132_));
 sg13g2_buf_1 _26252_ (.A(\cpu.uart.r_xstate[3] ),
    .X(_07133_));
 sg13g2_buf_1 _26253_ (.A(_07133_),
    .X(_07134_));
 sg13g2_nor2_1 _26254_ (.A(net1056),
    .B(_09280_),
    .Y(_07135_));
 sg13g2_nand3_1 _26255_ (.B(_07135_),
    .C(_06385_),
    .A(_10123_),
    .Y(_07136_));
 sg13g2_buf_1 _26256_ (.A(_07136_),
    .X(_07137_));
 sg13g2_nor2_2 _26257_ (.A(_05564_),
    .B(_07137_),
    .Y(_07138_));
 sg13g2_buf_2 _26258_ (.A(\cpu.uart.r_xstate[1] ),
    .X(_07139_));
 sg13g2_buf_2 _26259_ (.A(\cpu.uart.r_xstate[0] ),
    .X(_07140_));
 sg13g2_nand2_1 _26260_ (.Y(_07141_),
    .A(_07139_),
    .B(_07140_));
 sg13g2_nor2_1 _26261_ (.A(_07138_),
    .B(_07141_),
    .Y(_07142_));
 sg13g2_buf_1 _26262_ (.A(_07140_),
    .X(_07143_));
 sg13g2_nand2b_1 _26263_ (.Y(_07144_),
    .B(_07138_),
    .A_N(_07143_));
 sg13g2_nor2_1 _26264_ (.A(_07139_),
    .B(net959),
    .Y(_07145_));
 sg13g2_a22oi_1 _26265_ (.Y(_07146_),
    .B1(_07144_),
    .B2(_07145_),
    .A2(_07142_),
    .A1(net959));
 sg13g2_nor2_1 _26266_ (.A(net960),
    .B(_07146_),
    .Y(_07147_));
 sg13g2_inv_2 _26267_ (.Y(_07148_),
    .A(_07133_));
 sg13g2_buf_1 _26268_ (.A(\cpu.uart.r_xcnt[0] ),
    .X(_07149_));
 sg13g2_nor2_1 _26269_ (.A(_07149_),
    .B(\cpu.uart.r_xcnt[1] ),
    .Y(_07150_));
 sg13g2_and2_1 _26270_ (.A(net348),
    .B(_07150_),
    .X(_07151_));
 sg13g2_buf_2 _26271_ (.A(_07151_),
    .X(_07152_));
 sg13g2_inv_2 _26272_ (.Y(_07153_),
    .A(_07139_));
 sg13g2_nor2_1 _26273_ (.A(_07148_),
    .B(_07152_),
    .Y(_07154_));
 sg13g2_a21oi_1 _26274_ (.A1(_07143_),
    .A2(net959),
    .Y(_07155_),
    .B1(_07153_));
 sg13g2_a21oi_1 _26275_ (.A1(_07153_),
    .A2(_07154_),
    .Y(_07156_),
    .B1(_07155_));
 sg13g2_inv_1 _26276_ (.Y(_07157_),
    .A(_07131_));
 sg13g2_a22oi_1 _26277_ (.Y(_07158_),
    .B1(_07156_),
    .B2(_07157_),
    .A2(_07152_),
    .A1(_07148_));
 sg13g2_nor3_1 _26278_ (.A(net931),
    .B(_07147_),
    .C(_07158_),
    .Y(_07159_));
 sg13g2_buf_2 _26279_ (.A(_07159_),
    .X(_07160_));
 sg13g2_buf_1 _26280_ (.A(_07160_),
    .X(_07161_));
 sg13g2_nor2_1 _26281_ (.A(_07139_),
    .B(_07131_),
    .Y(_07162_));
 sg13g2_xnor2_1 _26282_ (.Y(_07163_),
    .A(net959),
    .B(_07162_));
 sg13g2_buf_2 _26283_ (.A(_07163_),
    .X(_07164_));
 sg13g2_buf_1 _26284_ (.A(_07164_),
    .X(_07165_));
 sg13g2_nor2b_1 _26285_ (.A(net643),
    .B_N(_10186_),
    .Y(_07166_));
 sg13g2_a21oi_1 _26286_ (.A1(\cpu.uart.r_out[1] ),
    .A2(net643),
    .Y(_07167_),
    .B1(_07166_));
 sg13g2_nor2_1 _26287_ (.A(\cpu.uart.r_out[0] ),
    .B(net30),
    .Y(_07168_));
 sg13g2_a21oi_1 _26288_ (.A1(net30),
    .A2(_07167_),
    .Y(_02659_),
    .B1(_07168_));
 sg13g2_nor2b_1 _26289_ (.A(net643),
    .B_N(_10194_),
    .Y(_07169_));
 sg13g2_a21oi_1 _26290_ (.A1(\cpu.uart.r_out[2] ),
    .A2(net643),
    .Y(_07170_),
    .B1(_07169_));
 sg13g2_nor2_1 _26291_ (.A(\cpu.uart.r_out[1] ),
    .B(_07161_),
    .Y(_07171_));
 sg13g2_a21oi_1 _26292_ (.A1(net30),
    .A2(_07170_),
    .Y(_02660_),
    .B1(_07171_));
 sg13g2_nor2b_1 _26293_ (.A(_07164_),
    .B_N(net1039),
    .Y(_07172_));
 sg13g2_a21oi_1 _26294_ (.A1(\cpu.uart.r_out[3] ),
    .A2(net643),
    .Y(_07173_),
    .B1(_07172_));
 sg13g2_nor2_1 _26295_ (.A(\cpu.uart.r_out[2] ),
    .B(_07160_),
    .Y(_07174_));
 sg13g2_a21oi_1 _26296_ (.A1(net30),
    .A2(_07173_),
    .Y(_02661_),
    .B1(_07174_));
 sg13g2_nor2b_1 _26297_ (.A(_07164_),
    .B_N(net1116),
    .Y(_07175_));
 sg13g2_a21oi_1 _26298_ (.A1(\cpu.uart.r_out[4] ),
    .A2(net643),
    .Y(_07176_),
    .B1(_07175_));
 sg13g2_nor2_1 _26299_ (.A(\cpu.uart.r_out[3] ),
    .B(_07160_),
    .Y(_07177_));
 sg13g2_a21oi_1 _26300_ (.A1(net30),
    .A2(_07176_),
    .Y(_02662_),
    .B1(_07177_));
 sg13g2_nor2b_1 _26301_ (.A(_07164_),
    .B_N(_10214_),
    .Y(_07178_));
 sg13g2_a21oi_1 _26302_ (.A1(\cpu.uart.r_out[5] ),
    .A2(_07165_),
    .Y(_07179_),
    .B1(_07178_));
 sg13g2_nor2_1 _26303_ (.A(\cpu.uart.r_out[4] ),
    .B(_07160_),
    .Y(_07180_));
 sg13g2_a21oi_1 _26304_ (.A1(net30),
    .A2(_07179_),
    .Y(_02663_),
    .B1(_07180_));
 sg13g2_nor2b_1 _26305_ (.A(_07164_),
    .B_N(_10220_),
    .Y(_07181_));
 sg13g2_a21oi_1 _26306_ (.A1(\cpu.uart.r_out[6] ),
    .A2(_07165_),
    .Y(_07182_),
    .B1(_07181_));
 sg13g2_nor2_1 _26307_ (.A(\cpu.uart.r_out[5] ),
    .B(_07160_),
    .Y(_07183_));
 sg13g2_a21oi_1 _26308_ (.A1(_07161_),
    .A2(_07182_),
    .Y(_02664_),
    .B1(_07183_));
 sg13g2_nor2b_1 _26309_ (.A(_07164_),
    .B_N(_10226_),
    .Y(_07184_));
 sg13g2_a21oi_1 _26310_ (.A1(\cpu.uart.r_out[7] ),
    .A2(net643),
    .Y(_07185_),
    .B1(_07184_));
 sg13g2_nor2_1 _26311_ (.A(\cpu.uart.r_out[6] ),
    .B(_07160_),
    .Y(_07186_));
 sg13g2_a21oi_1 _26312_ (.A1(net30),
    .A2(_07185_),
    .Y(_02665_),
    .B1(_07186_));
 sg13g2_nor2_1 _26313_ (.A(_07064_),
    .B(net643),
    .Y(_07187_));
 sg13g2_mux2_1 _26314_ (.A0(\cpu.uart.r_out[7] ),
    .A1(_07187_),
    .S(net30),
    .X(_02666_));
 sg13g2_nand2b_1 _26315_ (.Y(_07188_),
    .B(_10086_),
    .A_N(_10047_));
 sg13g2_nor3_1 _26316_ (.A(net1081),
    .B(_07119_),
    .C(net1082),
    .Y(_07189_));
 sg13g2_a22oi_1 _26317_ (.Y(_07190_),
    .B1(_07188_),
    .B2(_07189_),
    .A2(net1082),
    .A1(net1081));
 sg13g2_nor4_1 _26318_ (.A(_07122_),
    .B(\cpu.uart.r_rstate[1] ),
    .C(_07119_),
    .D(_07116_),
    .Y(_07191_));
 sg13g2_a21o_1 _26319_ (.A2(_07188_),
    .A1(net1081),
    .B1(_07119_),
    .X(_07192_));
 sg13g2_a22oi_1 _26320_ (.Y(_07193_),
    .B1(_07192_),
    .B2(net1082),
    .A2(_07191_),
    .A1(_07128_));
 sg13g2_o21ai_1 _26321_ (.B1(_07193_),
    .Y(_07194_),
    .A1(_07123_),
    .A2(_07190_));
 sg13g2_nor2_1 _26322_ (.A(_07123_),
    .B(net1081),
    .Y(_07195_));
 sg13g2_nor2b_1 _26323_ (.A(net1082),
    .B_N(_07128_),
    .Y(_07196_));
 sg13g2_nand2_1 _26324_ (.Y(_07197_),
    .A(net1081),
    .B(net1082));
 sg13g2_nor2_1 _26325_ (.A(_07122_),
    .B(_07197_),
    .Y(_07198_));
 sg13g2_a21oi_1 _26326_ (.A1(_07195_),
    .A2(_07196_),
    .Y(_07199_),
    .B1(_07198_));
 sg13g2_nor3_1 _26327_ (.A(net961),
    .B(_07114_),
    .C(_07199_),
    .Y(_07200_));
 sg13g2_xor2_1 _26328_ (.B(_07121_),
    .A(net962),
    .X(_07201_));
 sg13g2_o21ai_1 _26329_ (.B1(net930),
    .Y(_07202_),
    .A1(net348),
    .A2(_07201_));
 sg13g2_nor3_1 _26330_ (.A(_07194_),
    .B(_07200_),
    .C(_07202_),
    .Y(_07203_));
 sg13g2_and2_1 _26331_ (.A(_07122_),
    .B(net1081),
    .X(_07204_));
 sg13g2_buf_1 _26332_ (.A(_07204_),
    .X(_07205_));
 sg13g2_o21ai_1 _26333_ (.B1(net962),
    .Y(_07206_),
    .A1(_07120_),
    .A2(_07205_));
 sg13g2_nor2b_1 _26334_ (.A(_07191_),
    .B_N(_07206_),
    .Y(_07207_));
 sg13g2_and2_1 _26335_ (.A(_07203_),
    .B(_07207_),
    .X(_07208_));
 sg13g2_nor2_1 _26336_ (.A(_07112_),
    .B(_07203_),
    .Y(_07209_));
 sg13g2_a21oi_1 _26337_ (.A1(_07112_),
    .A2(_07208_),
    .Y(_02669_),
    .B1(_07209_));
 sg13g2_nand2_1 _26338_ (.Y(_07210_),
    .A(_07112_),
    .B(_07207_));
 sg13g2_inv_1 _26339_ (.Y(_07211_),
    .A(\cpu.uart.r_rcnt[1] ));
 sg13g2_a21oi_1 _26340_ (.A1(_07203_),
    .A2(_07210_),
    .Y(_07212_),
    .B1(_07211_));
 sg13g2_a21o_1 _26341_ (.A2(_07208_),
    .A1(_07113_),
    .B1(_07212_),
    .X(_02670_));
 sg13g2_nor3_2 _26342_ (.A(_07153_),
    .B(_07148_),
    .C(_07131_),
    .Y(_07213_));
 sg13g2_nor2_1 _26343_ (.A(_07148_),
    .B(net960),
    .Y(_07214_));
 sg13g2_nand2_1 _26344_ (.Y(_07215_),
    .A(_07148_),
    .B(_07131_));
 sg13g2_nor2_1 _26345_ (.A(_07139_),
    .B(_07140_),
    .Y(_07216_));
 sg13g2_nand2_1 _26346_ (.Y(_07217_),
    .A(_07215_),
    .B(_07216_));
 sg13g2_nor2_1 _26347_ (.A(_07214_),
    .B(_07217_),
    .Y(_07218_));
 sg13g2_nor3_1 _26348_ (.A(net931),
    .B(_07213_),
    .C(_07218_),
    .Y(_07219_));
 sg13g2_nand2_1 _26349_ (.Y(_07220_),
    .A(\cpu.uart.r_out[0] ),
    .B(_07164_));
 sg13g2_xor2_1 _26350_ (.B(_07220_),
    .A(\cpu.uart.r_x_invert ),
    .X(_07221_));
 sg13g2_nor2_1 _26351_ (.A(_00280_),
    .B(_07219_),
    .Y(_07222_));
 sg13g2_a21oi_1 _26352_ (.A1(_07219_),
    .A2(_07221_),
    .Y(_07223_),
    .B1(_07222_));
 sg13g2_buf_1 _26353_ (.A(\cpu.gpio.genblk1[3].srcs_o[1] ),
    .X(_07224_));
 sg13g2_nand2_1 _26354_ (.Y(_07225_),
    .A(_07133_),
    .B(_07131_));
 sg13g2_o21ai_1 _26355_ (.B1(_07225_),
    .Y(_07226_),
    .A1(net959),
    .A2(net348));
 sg13g2_nand2b_1 _26356_ (.Y(_07227_),
    .B(_07162_),
    .A_N(_07152_));
 sg13g2_o21ai_1 _26357_ (.B1(_07227_),
    .Y(_07228_),
    .A1(_07153_),
    .A2(_07157_));
 sg13g2_a21o_1 _26358_ (.A2(_07133_),
    .A1(_07140_),
    .B1(_07153_),
    .X(_07229_));
 sg13g2_a21oi_1 _26359_ (.A1(_07229_),
    .A2(_07215_),
    .Y(_07230_),
    .B1(_07152_));
 sg13g2_a221oi_1 _26360_ (.B2(_07134_),
    .C1(_07230_),
    .B1(_07228_),
    .A1(_07140_),
    .Y(_07231_),
    .A2(_07226_));
 sg13g2_nand3_1 _26361_ (.B(_07138_),
    .C(_07213_),
    .A(net958),
    .Y(_07232_));
 sg13g2_buf_1 _26362_ (.A(_07232_),
    .X(_07233_));
 sg13g2_a21oi_1 _26363_ (.A1(_07231_),
    .A2(_07233_),
    .Y(_07234_),
    .B1(net804));
 sg13g2_mux2_1 _26364_ (.A0(_07223_),
    .A1(net1080),
    .S(_07234_),
    .X(_02675_));
 sg13g2_a21oi_1 _26365_ (.A1(_07140_),
    .A2(_07150_),
    .Y(_07235_),
    .B1(_07132_));
 sg13g2_o21ai_1 _26366_ (.B1(_07132_),
    .Y(_07236_),
    .A1(_07140_),
    .A2(_07150_));
 sg13g2_o21ai_1 _26367_ (.B1(_07236_),
    .Y(_07237_),
    .A1(_07153_),
    .A2(_07235_));
 sg13g2_nand2_1 _26368_ (.Y(_07238_),
    .A(_07134_),
    .B(_07237_));
 sg13g2_nor3_1 _26369_ (.A(_07139_),
    .B(net959),
    .C(_07131_),
    .Y(_07239_));
 sg13g2_nand2b_1 _26370_ (.Y(_07240_),
    .B(_07239_),
    .A_N(_07140_));
 sg13g2_nand4_1 _26371_ (.B(_10058_),
    .C(_07238_),
    .A(net930),
    .Y(_07241_),
    .D(_07240_));
 sg13g2_nor2b_1 _26372_ (.A(_07241_),
    .B_N(_07233_),
    .Y(_07242_));
 sg13g2_nor2_1 _26373_ (.A(_07225_),
    .B(_07216_),
    .Y(_07243_));
 sg13g2_nor2_1 _26374_ (.A(_07239_),
    .B(_07243_),
    .Y(_07244_));
 sg13g2_nand2_1 _26375_ (.Y(_07245_),
    .A(_07242_),
    .B(_07244_));
 sg13g2_nor2b_1 _26376_ (.A(_07149_),
    .B_N(_07242_),
    .Y(_07246_));
 sg13g2_a21oi_1 _26377_ (.A1(_07149_),
    .A2(_07245_),
    .Y(_07247_),
    .B1(_07246_));
 sg13g2_inv_1 _26378_ (.Y(_02678_),
    .A(_07247_));
 sg13g2_nand2_1 _26379_ (.Y(_07248_),
    .A(_07149_),
    .B(_07244_));
 sg13g2_nand2_1 _26380_ (.Y(_07249_),
    .A(_07242_),
    .B(_07248_));
 sg13g2_o21ai_1 _26381_ (.B1(\cpu.uart.r_xcnt[1] ),
    .Y(_07250_),
    .A1(_07149_),
    .A2(_07245_));
 sg13g2_o21ai_1 _26382_ (.B1(_07250_),
    .Y(_02679_),
    .A1(\cpu.uart.r_xcnt[1] ),
    .A2(_07249_));
 sg13g2_nand3_1 _26383_ (.B(net444),
    .C(net124),
    .A(net620),
    .Y(_07251_));
 sg13g2_buf_2 _26384_ (.A(_07251_),
    .X(_07252_));
 sg13g2_buf_1 _26385_ (.A(_07252_),
    .X(_07253_));
 sg13g2_nand2_1 _26386_ (.Y(_07254_),
    .A(_10128_),
    .B(net399));
 sg13g2_buf_1 _26387_ (.A(_07254_),
    .X(_07255_));
 sg13g2_buf_1 _26388_ (.A(net109),
    .X(_07256_));
 sg13g2_buf_1 _26389_ (.A(net109),
    .X(_07257_));
 sg13g2_nand4_1 _26390_ (.B(_10333_),
    .C(_10341_),
    .A(_10327_),
    .Y(_07258_),
    .D(_04954_));
 sg13g2_buf_1 _26391_ (.A(_07258_),
    .X(_07259_));
 sg13g2_nor2_1 _26392_ (.A(_10336_),
    .B(_07259_),
    .Y(_07260_));
 sg13g2_nand2_1 _26393_ (.Y(_07261_),
    .A(net94),
    .B(_07260_));
 sg13g2_o21ai_1 _26394_ (.B1(_07261_),
    .Y(_07262_),
    .A1(net1041),
    .A2(_07256_));
 sg13g2_nand3_1 _26395_ (.B(_10333_),
    .C(_10341_),
    .A(_10327_),
    .Y(_07263_));
 sg13g2_o21ai_1 _26396_ (.B1(net94),
    .Y(_07264_),
    .A1(_10336_),
    .A2(_07263_));
 sg13g2_a21oi_1 _26397_ (.A1(_07252_),
    .A2(_07264_),
    .Y(_07265_),
    .B1(_04954_));
 sg13g2_a21oi_1 _26398_ (.A1(net78),
    .A2(_07262_),
    .Y(_02465_),
    .B1(_07265_));
 sg13g2_inv_1 _26399_ (.Y(_07266_),
    .A(_05360_));
 sg13g2_nor3_2 _26400_ (.A(_07266_),
    .B(_10336_),
    .C(_07259_),
    .Y(_07267_));
 sg13g2_nand2_1 _26401_ (.Y(_07268_),
    .A(net94),
    .B(_07267_));
 sg13g2_o21ai_1 _26402_ (.B1(_07268_),
    .Y(_07269_),
    .A1(net1040),
    .A2(net95));
 sg13g2_buf_1 _26403_ (.A(_07252_),
    .X(_07270_));
 sg13g2_o21ai_1 _26404_ (.B1(net77),
    .Y(_07271_),
    .A1(net104),
    .A2(_07260_));
 sg13g2_a22oi_1 _26405_ (.Y(_02466_),
    .B1(_07271_),
    .B2(_07266_),
    .A2(_07269_),
    .A1(net78));
 sg13g2_nand3_1 _26406_ (.B(_07255_),
    .C(_07267_),
    .A(_05416_),
    .Y(_07272_));
 sg13g2_o21ai_1 _26407_ (.B1(_07272_),
    .Y(_07273_),
    .A1(net1039),
    .A2(net95));
 sg13g2_o21ai_1 _26408_ (.B1(net77),
    .Y(_07274_),
    .A1(net104),
    .A2(_07267_));
 sg13g2_inv_1 _26409_ (.Y(_07275_),
    .A(_05416_));
 sg13g2_a22oi_1 _26410_ (.Y(_02467_),
    .B1(_07274_),
    .B2(_07275_),
    .A2(_07273_),
    .A1(net78));
 sg13g2_nand2_1 _26411_ (.Y(_07276_),
    .A(_05360_),
    .B(_05416_));
 sg13g2_nor4_1 _26412_ (.A(_10328_),
    .B(_10329_),
    .C(_07259_),
    .D(_07276_),
    .Y(_07277_));
 sg13g2_nand2_1 _26413_ (.Y(_07278_),
    .A(_05488_),
    .B(_07277_));
 sg13g2_inv_1 _26414_ (.Y(_07279_),
    .A(_07278_));
 sg13g2_nand2_1 _26415_ (.Y(_07280_),
    .A(net109),
    .B(_07279_));
 sg13g2_o21ai_1 _26416_ (.B1(_07280_),
    .Y(_07281_),
    .A1(net1116),
    .A2(net95));
 sg13g2_o21ai_1 _26417_ (.B1(_07270_),
    .Y(_07282_),
    .A1(net104),
    .A2(_07277_));
 sg13g2_inv_1 _26418_ (.Y(_07283_),
    .A(_05488_));
 sg13g2_a22oi_1 _26419_ (.Y(_02468_),
    .B1(_07282_),
    .B2(_07283_),
    .A2(_07281_),
    .A1(net78));
 sg13g2_nand3_1 _26420_ (.B(_05488_),
    .C(_07267_),
    .A(_05416_),
    .Y(_07284_));
 sg13g2_buf_1 _26421_ (.A(_07284_),
    .X(_07285_));
 sg13g2_nor2_1 _26422_ (.A(_10258_),
    .B(_07285_),
    .Y(_07286_));
 sg13g2_nand2_1 _26423_ (.Y(_07287_),
    .A(_05559_),
    .B(_07286_));
 sg13g2_o21ai_1 _26424_ (.B1(_07287_),
    .Y(_07288_),
    .A1(net1037),
    .A2(net95));
 sg13g2_nand2_1 _26425_ (.Y(_07289_),
    .A(_07257_),
    .B(_07285_));
 sg13g2_a21oi_1 _26426_ (.A1(_07252_),
    .A2(_07289_),
    .Y(_07290_),
    .B1(_05559_));
 sg13g2_a21oi_1 _26427_ (.A1(net78),
    .A2(_07288_),
    .Y(_02469_),
    .B1(_07290_));
 sg13g2_nand2_1 _26428_ (.Y(_07291_),
    .A(_05559_),
    .B(_05623_));
 sg13g2_nand2b_1 _26429_ (.Y(_07292_),
    .B(_10276_),
    .A_N(_10220_));
 sg13g2_o21ai_1 _26430_ (.B1(_07292_),
    .Y(_07293_),
    .A1(_07280_),
    .A2(_07291_));
 sg13g2_a21o_1 _26431_ (.A2(_07279_),
    .A1(_05559_),
    .B1(_10258_),
    .X(_07294_));
 sg13g2_a21oi_1 _26432_ (.A1(_07252_),
    .A2(_07294_),
    .Y(_07295_),
    .B1(_05623_));
 sg13g2_a21oi_1 _26433_ (.A1(_07253_),
    .A2(_07293_),
    .Y(_02470_),
    .B1(_07295_));
 sg13g2_nand4_1 _26434_ (.B(_05623_),
    .C(_05655_),
    .A(_05559_),
    .Y(_07296_),
    .D(_07286_));
 sg13g2_o21ai_1 _26435_ (.B1(_07296_),
    .Y(_07297_),
    .A1(net1035),
    .A2(_07256_));
 sg13g2_o21ai_1 _26436_ (.B1(_07257_),
    .Y(_07298_),
    .A1(_07285_),
    .A2(_07291_));
 sg13g2_a21oi_1 _26437_ (.A1(_07252_),
    .A2(_07298_),
    .Y(_07299_),
    .B1(_05655_));
 sg13g2_a21oi_1 _26438_ (.A1(_07253_),
    .A2(_07297_),
    .Y(_02471_),
    .B1(_07299_));
 sg13g2_nand3_1 _26439_ (.B(_05623_),
    .C(_05655_),
    .A(_05559_),
    .Y(_07300_));
 sg13g2_buf_1 _26440_ (.A(_07300_),
    .X(_07301_));
 sg13g2_nor2_1 _26441_ (.A(_07278_),
    .B(_07301_),
    .Y(_07302_));
 sg13g2_nand3_1 _26442_ (.B(_07255_),
    .C(_07302_),
    .A(_05037_),
    .Y(_07303_));
 sg13g2_o21ai_1 _26443_ (.B1(_07303_),
    .Y(_07304_),
    .A1(_10229_),
    .A2(net95));
 sg13g2_o21ai_1 _26444_ (.B1(_07270_),
    .Y(_07305_),
    .A1(net104),
    .A2(_07302_));
 sg13g2_inv_1 _26445_ (.Y(_07306_),
    .A(_05037_));
 sg13g2_a22oi_1 _26446_ (.Y(_02472_),
    .B1(_07305_),
    .B2(_07306_),
    .A2(_07304_),
    .A1(net78));
 sg13g2_inv_1 _26447_ (.Y(_07307_),
    .A(_05725_));
 sg13g2_or2_1 _26448_ (.X(_07308_),
    .B(_07301_),
    .A(_07306_));
 sg13g2_buf_1 _26449_ (.A(_07308_),
    .X(_07309_));
 sg13g2_nor3_2 _26450_ (.A(_07307_),
    .B(_07285_),
    .C(_07309_),
    .Y(_07310_));
 sg13g2_nand2_1 _26451_ (.Y(_07311_),
    .A(net94),
    .B(_07310_));
 sg13g2_o21ai_1 _26452_ (.B1(_07311_),
    .Y(_07312_),
    .A1(_10302_),
    .A2(net95));
 sg13g2_nor2_1 _26453_ (.A(_07285_),
    .B(_07309_),
    .Y(_07313_));
 sg13g2_o21ai_1 _26454_ (.B1(net77),
    .Y(_07314_),
    .A1(net104),
    .A2(_07313_));
 sg13g2_a22oi_1 _26455_ (.Y(_02473_),
    .B1(_07314_),
    .B2(_07307_),
    .A2(_07312_),
    .A1(net77));
 sg13g2_nand3_1 _26456_ (.B(net109),
    .C(_07310_),
    .A(_05739_),
    .Y(_07315_));
 sg13g2_o21ai_1 _26457_ (.B1(_07315_),
    .Y(_07316_),
    .A1(_10307_),
    .A2(net94));
 sg13g2_o21ai_1 _26458_ (.B1(net77),
    .Y(_07317_),
    .A1(net104),
    .A2(_07310_));
 sg13g2_inv_1 _26459_ (.Y(_07318_),
    .A(_05739_));
 sg13g2_a22oi_1 _26460_ (.Y(_02474_),
    .B1(_07317_),
    .B2(_07318_),
    .A2(_07316_),
    .A1(net77));
 sg13g2_nand4_1 _26461_ (.B(_05133_),
    .C(net109),
    .A(_05739_),
    .Y(_07319_),
    .D(_07310_));
 sg13g2_o21ai_1 _26462_ (.B1(_07319_),
    .Y(_07320_),
    .A1(_10312_),
    .A2(net95));
 sg13g2_a21o_1 _26463_ (.A2(_07310_),
    .A1(_05739_),
    .B1(_10258_),
    .X(_07321_));
 sg13g2_a21oi_1 _26464_ (.A1(_07252_),
    .A2(_07321_),
    .Y(_07322_),
    .B1(_05133_));
 sg13g2_a21oi_1 _26465_ (.A1(net78),
    .A2(_07320_),
    .Y(_02475_),
    .B1(_07322_));
 sg13g2_nand3_1 _26466_ (.B(_05739_),
    .C(_05133_),
    .A(_05725_),
    .Y(_07323_));
 sg13g2_nor4_2 _26467_ (.A(_07306_),
    .B(_07278_),
    .C(_07301_),
    .Y(_07324_),
    .D(_07323_));
 sg13g2_nand3_1 _26468_ (.B(net109),
    .C(_07324_),
    .A(_05164_),
    .Y(_07325_));
 sg13g2_o21ai_1 _26469_ (.B1(_07325_),
    .Y(_07326_),
    .A1(_10319_),
    .A2(net94));
 sg13g2_o21ai_1 _26470_ (.B1(net77),
    .Y(_07327_),
    .A1(net104),
    .A2(_07324_));
 sg13g2_inv_1 _26471_ (.Y(_07328_),
    .A(_05164_));
 sg13g2_a22oi_1 _26472_ (.Y(_02476_),
    .B1(_07327_),
    .B2(_07328_),
    .A2(_07326_),
    .A1(net77));
 sg13g2_nand3_1 _26473_ (.B(_05488_),
    .C(_07267_),
    .A(_05416_),
    .Y(_07329_));
 sg13g2_nor4_1 _26474_ (.A(_07307_),
    .B(_07318_),
    .C(_07329_),
    .D(_07309_),
    .Y(_07330_));
 sg13g2_nand3_1 _26475_ (.B(_05164_),
    .C(_07330_),
    .A(_05133_),
    .Y(_07331_));
 sg13g2_nor3_1 _26476_ (.A(_05194_),
    .B(net103),
    .C(_07331_),
    .Y(_07332_));
 sg13g2_a21oi_1 _26477_ (.A1(_10324_),
    .A2(net103),
    .Y(_07333_),
    .B1(_07332_));
 sg13g2_and2_1 _26478_ (.A(net109),
    .B(_07331_),
    .X(_07334_));
 sg13g2_o21ai_1 _26479_ (.B1(_05194_),
    .Y(_07335_),
    .A1(net72),
    .A2(_07334_));
 sg13g2_o21ai_1 _26480_ (.B1(_07335_),
    .Y(_02477_),
    .A1(net73),
    .A2(_07333_));
 sg13g2_and3_1 _26481_ (.X(_07336_),
    .A(_05164_),
    .B(_05194_),
    .C(_05208_));
 sg13g2_buf_1 _26482_ (.A(_07336_),
    .X(_07337_));
 sg13g2_nand3_1 _26483_ (.B(_07324_),
    .C(_07337_),
    .A(net94),
    .Y(_07338_));
 sg13g2_o21ai_1 _26484_ (.B1(_07338_),
    .Y(_07339_),
    .A1(_10326_),
    .A2(net95));
 sg13g2_nand3_1 _26485_ (.B(_05194_),
    .C(_07324_),
    .A(_05164_),
    .Y(_07340_));
 sg13g2_nand2_1 _26486_ (.Y(_07341_),
    .A(net94),
    .B(_07340_));
 sg13g2_a21oi_1 _26487_ (.A1(_07252_),
    .A2(_07341_),
    .Y(_07342_),
    .B1(_05208_));
 sg13g2_a21oi_1 _26488_ (.A1(net78),
    .A2(_07339_),
    .Y(_02478_),
    .B1(_07342_));
 sg13g2_nand3_1 _26489_ (.B(_07330_),
    .C(_07337_),
    .A(_05133_),
    .Y(_07343_));
 sg13g2_nor3_1 _26490_ (.A(_05241_),
    .B(_10258_),
    .C(_07343_),
    .Y(_07344_));
 sg13g2_a21oi_1 _26491_ (.A1(_10339_),
    .A2(net103),
    .Y(_07345_),
    .B1(_07344_));
 sg13g2_and2_1 _26492_ (.A(net109),
    .B(_07343_),
    .X(_07346_));
 sg13g2_o21ai_1 _26493_ (.B1(_05241_),
    .Y(_07347_),
    .A1(net72),
    .A2(_07346_));
 sg13g2_o21ai_1 _26494_ (.B1(_07347_),
    .Y(_02479_),
    .A1(net73),
    .A2(_07345_));
 sg13g2_nand3_1 _26495_ (.B(_07324_),
    .C(_07337_),
    .A(_05241_),
    .Y(_07348_));
 sg13g2_nor3_1 _26496_ (.A(_05275_),
    .B(_10258_),
    .C(_07348_),
    .Y(_07349_));
 sg13g2_a21oi_1 _26497_ (.A1(_10344_),
    .A2(net103),
    .Y(_07350_),
    .B1(_07349_));
 sg13g2_and2_1 _26498_ (.A(_10238_),
    .B(_07348_),
    .X(_07351_));
 sg13g2_o21ai_1 _26499_ (.B1(_05275_),
    .Y(_07352_),
    .A1(net72),
    .A2(_07351_));
 sg13g2_o21ai_1 _26500_ (.B1(_07352_),
    .Y(_02480_),
    .A1(net73),
    .A2(_07350_));
 sg13g2_nor2_1 _26501_ (.A(\cpu.r_clk_invert ),
    .B(net707),
    .Y(_07353_));
 sg13g2_a21oi_1 _26502_ (.A1(_09290_),
    .A2(net705),
    .Y(_02547_),
    .B1(_07353_));
 sg13g2_nand2b_1 _26503_ (.Y(_07354_),
    .B(net803),
    .A_N(\cpu.d_flush_all ));
 sg13g2_buf_2 _26504_ (.A(_07354_),
    .X(_07355_));
 sg13g2_nor2b_1 _26505_ (.A(\cpu.dcache.r_valid[0] ),
    .B_N(net440),
    .Y(_07356_));
 sg13g2_nand4_1 _26506_ (.B(_02926_),
    .C(_12208_),
    .A(_09486_),
    .Y(_07357_),
    .D(_12108_));
 sg13g2_buf_2 _26507_ (.A(_07357_),
    .X(_07358_));
 sg13g2_nor2_1 _26508_ (.A(net607),
    .B(_07358_),
    .Y(_07359_));
 sg13g2_nor3_1 _26509_ (.A(_07355_),
    .B(_07356_),
    .C(_07359_),
    .Y(_00741_));
 sg13g2_nor2_1 _26510_ (.A(\cpu.dcache.r_valid[1] ),
    .B(net483),
    .Y(_07360_));
 sg13g2_nor2_1 _26511_ (.A(net661),
    .B(_07358_),
    .Y(_07361_));
 sg13g2_nor3_1 _26512_ (.A(_07355_),
    .B(_07360_),
    .C(_07361_),
    .Y(_00742_));
 sg13g2_nor2_1 _26513_ (.A(\cpu.dcache.r_valid[2] ),
    .B(net481),
    .Y(_07362_));
 sg13g2_nor2_1 _26514_ (.A(net606),
    .B(_07358_),
    .Y(_07363_));
 sg13g2_nor3_1 _26515_ (.A(_07355_),
    .B(_07362_),
    .C(_07363_),
    .Y(_00743_));
 sg13g2_nor2_1 _26516_ (.A(\cpu.dcache.r_valid[3] ),
    .B(net197),
    .Y(_07364_));
 sg13g2_nor2_1 _26517_ (.A(net271),
    .B(_07358_),
    .Y(_07365_));
 sg13g2_nor3_1 _26518_ (.A(_07355_),
    .B(_07364_),
    .C(_07365_),
    .Y(_00744_));
 sg13g2_inv_1 _26519_ (.Y(_07366_),
    .A(\cpu.dcache.r_valid[4] ));
 sg13g2_inv_1 _26520_ (.Y(_07367_),
    .A(_07358_));
 sg13g2_a221oi_1 _26521_ (.B2(net444),
    .C1(_07355_),
    .B1(_07367_),
    .A1(_07366_),
    .Y(_00745_),
    .A2(net386));
 sg13g2_nor2_1 _26522_ (.A(\cpu.dcache.r_valid[5] ),
    .B(_12840_),
    .Y(_07368_));
 sg13g2_nor2_1 _26523_ (.A(_12771_),
    .B(_07358_),
    .Y(_07369_));
 sg13g2_nor3_1 _26524_ (.A(_07355_),
    .B(_07368_),
    .C(_07369_),
    .Y(_00746_));
 sg13g2_nor2_1 _26525_ (.A(\cpu.dcache.r_valid[6] ),
    .B(_02791_),
    .Y(_07370_));
 sg13g2_nor2_1 _26526_ (.A(_02722_),
    .B(_07358_),
    .Y(_07371_));
 sg13g2_nor3_1 _26527_ (.A(_07355_),
    .B(_07370_),
    .C(_07371_),
    .Y(_00747_));
 sg13g2_nor2_1 _26528_ (.A(\cpu.dcache.r_valid[7] ),
    .B(net227),
    .Y(_07372_));
 sg13g2_nor2_1 _26529_ (.A(_02833_),
    .B(_07358_),
    .Y(_07373_));
 sg13g2_nor3_1 _26530_ (.A(_07355_),
    .B(_07372_),
    .C(_07373_),
    .Y(_00748_));
 sg13g2_nor2_1 _26531_ (.A(net1114),
    .B(net1113),
    .Y(_07374_));
 sg13g2_nand3_1 _26532_ (.B(_07374_),
    .C(_04746_),
    .A(_10355_),
    .Y(_07375_));
 sg13g2_buf_1 _26533_ (.A(_07375_),
    .X(_07376_));
 sg13g2_nand2_1 _26534_ (.Y(_07377_),
    .A(_08397_),
    .B(net576));
 sg13g2_o21ai_1 _26535_ (.B1(_07377_),
    .Y(_07378_),
    .A1(net656),
    .A2(net576));
 sg13g2_and3_1 _26536_ (.X(_00797_),
    .A(net214),
    .B(_09445_),
    .C(_07378_));
 sg13g2_and4_1 _26537_ (.A(net745),
    .B(_10962_),
    .C(\cpu.dec.do_flush_all ),
    .D(net666),
    .X(_00930_));
 sg13g2_and4_1 _26538_ (.A(net745),
    .B(_10796_),
    .C(\cpu.dec.do_flush_all ),
    .D(net666),
    .X(_00948_));
 sg13g2_nand2_1 _26539_ (.Y(_07379_),
    .A(net666),
    .B(_03498_));
 sg13g2_nor2_1 _26540_ (.A(_06849_),
    .B(net666),
    .Y(_07380_));
 sg13g2_a21oi_1 _26541_ (.A1(_05790_),
    .A2(_07379_),
    .Y(_07381_),
    .B1(_07380_));
 sg13g2_nor2_1 _26542_ (.A(_11678_),
    .B(_11281_),
    .Y(_07382_));
 sg13g2_nand3_1 _26543_ (.B(net666),
    .C(_07382_),
    .A(net745),
    .Y(_07383_));
 sg13g2_mux2_1 _26544_ (.A0(_10789_),
    .A1(_09285_),
    .S(_07383_),
    .X(_07384_));
 sg13g2_nor2_1 _26545_ (.A(_11541_),
    .B(net576),
    .Y(_07385_));
 sg13g2_a21oi_1 _26546_ (.A1(net576),
    .A2(_07384_),
    .Y(_07386_),
    .B1(_07385_));
 sg13g2_nor3_1 _26547_ (.A(net707),
    .B(_07381_),
    .C(_07386_),
    .Y(_00949_));
 sg13g2_nor2_1 _26548_ (.A(_08390_),
    .B(_00298_),
    .Y(_07387_));
 sg13g2_nand2_1 _26549_ (.Y(_07388_),
    .A(_08392_),
    .B(net666));
 sg13g2_nor2_1 _26550_ (.A(_00310_),
    .B(_07388_),
    .Y(_07389_));
 sg13g2_nand2_1 _26551_ (.Y(_07390_),
    .A(_09486_),
    .B(_09498_));
 sg13g2_o21ai_1 _26552_ (.B1(_07390_),
    .Y(_07391_),
    .A1(_09385_),
    .A2(net663));
 sg13g2_nor2_1 _26553_ (.A(_11693_),
    .B(_07391_),
    .Y(_07392_));
 sg13g2_o21ai_1 _26554_ (.B1(_09443_),
    .Y(_07393_),
    .A1(net957),
    .A2(_07392_));
 sg13g2_inv_1 _26555_ (.Y(_07394_),
    .A(_07393_));
 sg13g2_o21ai_1 _26556_ (.B1(_07394_),
    .Y(_07395_),
    .A1(_08390_),
    .A2(_07389_));
 sg13g2_a21oi_1 _26557_ (.A1(_04814_),
    .A2(_07387_),
    .Y(_01068_),
    .B1(_07395_));
 sg13g2_o21ai_1 _26558_ (.B1(_07389_),
    .Y(_07396_),
    .A1(_11680_),
    .A2(_04814_));
 sg13g2_a21oi_1 _26559_ (.A1(_08416_),
    .A2(_07396_),
    .Y(_01069_),
    .B1(_07393_));
 sg13g2_inv_1 _26560_ (.Y(_07397_),
    .A(\cpu.icache.r_valid[0] ));
 sg13g2_nand2b_1 _26561_ (.Y(_07398_),
    .B(_09444_),
    .A_N(\cpu.ex.i_flush_all ));
 sg13g2_buf_2 _26562_ (.A(_07398_),
    .X(_07399_));
 sg13g2_a21oi_1 _26563_ (.A1(_07397_),
    .A2(net421),
    .Y(_02424_),
    .B1(_07399_));
 sg13g2_nor2_1 _26564_ (.A(\cpu.icache.r_valid[1] ),
    .B(_06484_),
    .Y(_07400_));
 sg13g2_nor2_1 _26565_ (.A(_07399_),
    .B(_07400_),
    .Y(_02425_));
 sg13g2_nor2_1 _26566_ (.A(\cpu.icache.r_valid[2] ),
    .B(_06501_),
    .Y(_07401_));
 sg13g2_nor2_1 _26567_ (.A(_07399_),
    .B(_07401_),
    .Y(_02426_));
 sg13g2_inv_1 _26568_ (.Y(_07402_),
    .A(\cpu.icache.r_valid[3] ));
 sg13g2_a21oi_1 _26569_ (.A1(_07402_),
    .A2(net284),
    .Y(_02427_),
    .B1(_07399_));
 sg13g2_nor2_1 _26570_ (.A(\cpu.icache.r_valid[4] ),
    .B(_06527_),
    .Y(_07403_));
 sg13g2_nor2_1 _26571_ (.A(_07399_),
    .B(_07403_),
    .Y(_02428_));
 sg13g2_inv_1 _26572_ (.Y(_07404_),
    .A(\cpu.icache.r_valid[5] ));
 sg13g2_a21oi_1 _26573_ (.A1(_07404_),
    .A2(_06536_),
    .Y(_02429_),
    .B1(_07399_));
 sg13g2_nor2_1 _26574_ (.A(\cpu.icache.r_valid[6] ),
    .B(_06551_),
    .Y(_07405_));
 sg13g2_nor2_1 _26575_ (.A(_07399_),
    .B(_07405_),
    .Y(_02430_));
 sg13g2_nor2_1 _26576_ (.A(\cpu.icache.r_valid[7] ),
    .B(_06562_),
    .Y(_07406_));
 sg13g2_nor2_1 _26577_ (.A(_07399_),
    .B(_07406_),
    .Y(_02431_));
 sg13g2_nand3_1 _26578_ (.B(net124),
    .C(_04930_),
    .A(net1116),
    .Y(_07407_));
 sg13g2_nand2_1 _26579_ (.Y(_07408_),
    .A(_09326_),
    .B(_07407_));
 sg13g2_nand3_1 _26580_ (.B(_06745_),
    .C(_04934_),
    .A(net1038),
    .Y(_07409_));
 sg13g2_a21oi_1 _26581_ (.A1(_07408_),
    .A2(_07409_),
    .Y(_00317_),
    .B1(net577));
 sg13g2_nor2_1 _26582_ (.A(_02926_),
    .B(net1100),
    .Y(_07410_));
 sg13g2_nor2b_1 _26583_ (.A(_07410_),
    .B_N(_00315_),
    .Y(_00586_));
 sg13g2_nor2_1 _26584_ (.A(_12134_),
    .B(_12178_),
    .Y(_07411_));
 sg13g2_nor2_1 _26585_ (.A(_07410_),
    .B(_07411_),
    .Y(_00587_));
 sg13g2_xor2_1 _26586_ (.B(_12108_),
    .A(_12131_),
    .X(_07412_));
 sg13g2_nor2_1 _26587_ (.A(_07410_),
    .B(_07412_),
    .Y(_00588_));
 sg13g2_nor2_1 _26588_ (.A(_12656_),
    .B(net576),
    .Y(_07413_));
 sg13g2_a21oi_1 _26589_ (.A1(_08531_),
    .A2(net576),
    .Y(_07414_),
    .B1(_07413_));
 sg13g2_nor2_1 _26590_ (.A(net631),
    .B(_07414_),
    .Y(_00798_));
 sg13g2_nand2_1 _26591_ (.Y(_07415_),
    .A(_08500_),
    .B(net666));
 sg13g2_a21oi_2 _26592_ (.B1(net215),
    .Y(_07416_),
    .A2(_07415_),
    .A1(_11671_));
 sg13g2_nor2b_1 _26593_ (.A(net745),
    .B_N(_07416_),
    .Y(_07417_));
 sg13g2_nand3b_1 _26594_ (.B(_04139_),
    .C(_07382_),
    .Y(_07418_),
    .A_N(_10964_));
 sg13g2_a21oi_1 _26595_ (.A1(net745),
    .A2(_07418_),
    .Y(_07419_),
    .B1(_09386_));
 sg13g2_nor2_1 _26596_ (.A(_03687_),
    .B(_07419_),
    .Y(_07420_));
 sg13g2_nor2_1 _26597_ (.A(_10964_),
    .B(_07420_),
    .Y(_07421_));
 sg13g2_a21oi_1 _26598_ (.A1(_11541_),
    .A2(_07420_),
    .Y(_07422_),
    .B1(_07421_));
 sg13g2_nor2_1 _26599_ (.A(_07416_),
    .B(_07422_),
    .Y(_07423_));
 sg13g2_o21ai_1 _26600_ (.B1(_09990_),
    .Y(_00799_),
    .A1(_07417_),
    .A2(_07423_));
 sg13g2_mux2_1 _26601_ (.A0(net983),
    .A1(_11029_),
    .S(net576),
    .X(_07424_));
 sg13g2_and2_1 _26602_ (.A(_12004_),
    .B(_07424_),
    .X(_00800_));
 sg13g2_nor2_1 _26603_ (.A(_06843_),
    .B(_09998_),
    .Y(_07425_));
 sg13g2_nor2_1 _26604_ (.A(net957),
    .B(_07392_),
    .Y(_07426_));
 sg13g2_nor4_1 _26605_ (.A(\cpu.ex.r_branch_stall ),
    .B(_11669_),
    .C(_03373_),
    .D(_07388_),
    .Y(_07427_));
 sg13g2_nor3_1 _26606_ (.A(_10364_),
    .B(_07426_),
    .C(_07427_),
    .Y(_07428_));
 sg13g2_nand2_1 _26607_ (.Y(_07429_),
    .A(_08500_),
    .B(_11675_));
 sg13g2_o21ai_1 _26608_ (.B1(_04828_),
    .Y(_07430_),
    .A1(_07428_),
    .A2(_07429_));
 sg13g2_nor2_1 _26609_ (.A(_06849_),
    .B(_07430_),
    .Y(_07431_));
 sg13g2_o21ai_1 _26610_ (.B1(_09990_),
    .Y(_00946_),
    .A1(_07425_),
    .A2(_07431_));
 sg13g2_nand2_1 _26611_ (.Y(_07432_),
    .A(_09486_),
    .B(_09457_));
 sg13g2_nand3_1 _26612_ (.B(\cpu.dec.do_flush_write ),
    .C(_04139_),
    .A(net745),
    .Y(_07433_));
 sg13g2_a21oi_1 _26613_ (.A1(_07432_),
    .A2(_07433_),
    .Y(_00947_),
    .B1(_06814_));
 sg13g2_nand2_1 _26614_ (.Y(_07434_),
    .A(\cpu.dec.io ),
    .B(_04139_));
 sg13g2_nand2_1 _26615_ (.Y(_07435_),
    .A(net891),
    .B(_09457_));
 sg13g2_buf_1 _26616_ (.A(_06813_),
    .X(_07436_));
 sg13g2_a21oi_1 _26617_ (.A1(_07434_),
    .A2(_07435_),
    .Y(_00950_),
    .B1(net575));
 sg13g2_and2_1 _26618_ (.A(_09286_),
    .B(_07416_),
    .X(_07437_));
 sg13g2_nand2_1 _26619_ (.Y(_07438_),
    .A(_10789_),
    .B(net576));
 sg13g2_o21ai_1 _26620_ (.B1(_07438_),
    .Y(_07439_),
    .A1(net620),
    .A2(_07376_));
 sg13g2_nor2_1 _26621_ (.A(_07416_),
    .B(_07439_),
    .Y(_07440_));
 sg13g2_nor3_1 _26622_ (.A(net707),
    .B(_07437_),
    .C(_07440_),
    .Y(_00997_));
 sg13g2_a22oi_1 _26623_ (.Y(_07441_),
    .B1(_11695_),
    .B2(net1053),
    .A2(_04139_),
    .A1(_11669_));
 sg13g2_nor2_1 _26624_ (.A(_09390_),
    .B(_07441_),
    .Y(_00998_));
 sg13g2_and2_1 _26625_ (.A(_11541_),
    .B(_05802_),
    .X(_07442_));
 sg13g2_buf_1 _26626_ (.A(_07442_),
    .X(_07443_));
 sg13g2_mux2_1 _26627_ (.A0(_10930_),
    .A1(net437),
    .S(_07443_),
    .X(_07444_));
 sg13g2_nand2_1 _26628_ (.Y(_07445_),
    .A(_05790_),
    .B(_07444_));
 sg13g2_a21oi_1 _26629_ (.A1(_11671_),
    .A2(_07445_),
    .Y(_01074_),
    .B1(net575));
 sg13g2_mux2_1 _26630_ (.A0(net1016),
    .A1(_09349_),
    .S(_07443_),
    .X(_07446_));
 sg13g2_nand2_1 _26631_ (.Y(_07447_),
    .A(net214),
    .B(_07446_));
 sg13g2_o21ai_1 _26632_ (.B1(_07447_),
    .Y(_07448_),
    .A1(net796),
    .A2(net214));
 sg13g2_nor2_1 _26633_ (.A(_09390_),
    .B(_07448_),
    .Y(_01075_));
 sg13g2_inv_1 _26634_ (.Y(_07449_),
    .A(_08525_));
 sg13g2_mux2_1 _26635_ (.A0(\cpu.ex.mmu_read[1] ),
    .A1(_10246_),
    .S(_07443_),
    .X(_07450_));
 sg13g2_nand2b_1 _26636_ (.Y(_07451_),
    .B(_07450_),
    .A_N(_08431_));
 sg13g2_a21oi_1 _26637_ (.A1(_07449_),
    .A2(_07451_),
    .Y(_01076_),
    .B1(net575));
 sg13g2_buf_1 _26638_ (.A(net707),
    .X(_07452_));
 sg13g2_nor2_1 _26639_ (.A(net1024),
    .B(net1109),
    .Y(_07453_));
 sg13g2_nand3_1 _26640_ (.B(net1083),
    .C(_07453_),
    .A(_05837_),
    .Y(_07454_));
 sg13g2_nor3_2 _26641_ (.A(net970),
    .B(_05815_),
    .C(_07454_),
    .Y(_07455_));
 sg13g2_nor2b_1 _26642_ (.A(_00257_),
    .B_N(_05800_),
    .Y(_07456_));
 sg13g2_nand2b_1 _26643_ (.Y(_07457_),
    .B(net1052),
    .A_N(_00255_));
 sg13g2_inv_1 _26644_ (.Y(_07458_),
    .A(\cpu.dec.do_inv_mmu ));
 sg13g2_nor2_1 _26645_ (.A(_07458_),
    .B(_05797_),
    .Y(_07459_));
 sg13g2_buf_2 _26646_ (.A(_07459_),
    .X(_07460_));
 sg13g2_a21oi_1 _26647_ (.A1(_07456_),
    .A2(_07457_),
    .Y(_07461_),
    .B1(_07460_));
 sg13g2_nor3_2 _26648_ (.A(_08431_),
    .B(_08525_),
    .C(_07461_),
    .Y(_07462_));
 sg13g2_nand2_1 _26649_ (.Y(_07463_),
    .A(_05799_),
    .B(_07462_));
 sg13g2_buf_1 _26650_ (.A(_07463_),
    .X(_07464_));
 sg13g2_nor3_1 _26651_ (.A(_07458_),
    .B(_10962_),
    .C(_05797_),
    .Y(_07465_));
 sg13g2_nor2b_1 _26652_ (.A(_07465_),
    .B_N(_07462_),
    .Y(_07466_));
 sg13g2_buf_2 _26653_ (.A(_07466_),
    .X(_07467_));
 sg13g2_o21ai_1 _26654_ (.B1(_07467_),
    .Y(_07468_),
    .A1(_07455_),
    .A2(net213));
 sg13g2_nor2_1 _26655_ (.A(net620),
    .B(_07463_),
    .Y(_07469_));
 sg13g2_buf_1 _26656_ (.A(_07469_),
    .X(_07470_));
 sg13g2_a22oi_1 _26657_ (.Y(_07471_),
    .B1(_07470_),
    .B2(_07455_),
    .A2(_07468_),
    .A1(\cpu.genblk1.mmu.r_valid_d[0] ));
 sg13g2_nor2_1 _26658_ (.A(net574),
    .B(_07471_),
    .Y(_01077_));
 sg13g2_nor2_2 _26659_ (.A(net975),
    .B(_05860_),
    .Y(_07472_));
 sg13g2_nand2_1 _26660_ (.Y(_07473_),
    .A(_00288_),
    .B(_07453_));
 sg13g2_nand2_1 _26661_ (.Y(_07474_),
    .A(net971),
    .B(_07473_));
 sg13g2_o21ai_1 _26662_ (.B1(_07474_),
    .Y(_07475_),
    .A1(_05810_),
    .A2(_07454_));
 sg13g2_nor4_1 _26663_ (.A(net1016),
    .B(_05815_),
    .C(net971),
    .D(_07473_),
    .Y(_07476_));
 sg13g2_a21o_1 _26664_ (.A2(_07475_),
    .A1(net1016),
    .B1(_07476_),
    .X(_07477_));
 sg13g2_buf_1 _26665_ (.A(_07477_),
    .X(_07478_));
 sg13g2_inv_1 _26666_ (.Y(_07479_),
    .A(net455));
 sg13g2_nor2_1 _26667_ (.A(net213),
    .B(_07479_),
    .Y(_07480_));
 sg13g2_buf_1 _26668_ (.A(net213),
    .X(_07481_));
 sg13g2_buf_1 _26669_ (.A(_07467_),
    .X(_07482_));
 sg13g2_o21ai_1 _26670_ (.B1(net186),
    .Y(_07483_),
    .A1(_05862_),
    .A2(net187));
 sg13g2_a22oi_1 _26671_ (.Y(_07484_),
    .B1(_07483_),
    .B2(\cpu.genblk1.mmu.r_valid_d[10] ),
    .A2(_07480_),
    .A1(_07472_));
 sg13g2_nor2_1 _26672_ (.A(net574),
    .B(_07484_),
    .Y(_01078_));
 sg13g2_o21ai_1 _26673_ (.B1(net186),
    .Y(_07485_),
    .A1(_05871_),
    .A2(net187));
 sg13g2_a22oi_1 _26674_ (.Y(_07486_),
    .B1(_07485_),
    .B2(\cpu.genblk1.mmu.r_valid_d[11] ),
    .A2(net188),
    .A1(_05871_));
 sg13g2_nor2_1 _26675_ (.A(_07452_),
    .B(_07486_),
    .Y(_01079_));
 sg13g2_nand2_1 _26676_ (.Y(_07487_),
    .A(net1109),
    .B(_12152_));
 sg13g2_nor3_1 _26677_ (.A(net973),
    .B(net1024),
    .C(_07487_),
    .Y(_07488_));
 sg13g2_buf_2 _26678_ (.A(_07488_),
    .X(_07489_));
 sg13g2_nor2_1 _26679_ (.A(net1109),
    .B(_05827_),
    .Y(_07490_));
 sg13g2_a21oi_1 _26680_ (.A1(net972),
    .A2(_05817_),
    .Y(_07491_),
    .B1(_07490_));
 sg13g2_nor2b_1 _26681_ (.A(_07491_),
    .B_N(net1083),
    .Y(_07492_));
 sg13g2_and2_1 _26682_ (.A(net455),
    .B(_07492_),
    .X(_07493_));
 sg13g2_o21ai_1 _26683_ (.B1(net186),
    .Y(_07494_),
    .A1(net187),
    .A2(_07493_));
 sg13g2_a22oi_1 _26684_ (.Y(_07495_),
    .B1(_07494_),
    .B2(\cpu.genblk1.mmu.r_valid_d[12] ),
    .A2(_07489_),
    .A1(_07480_));
 sg13g2_nor2_1 _26685_ (.A(net574),
    .B(_07495_),
    .Y(_01080_));
 sg13g2_nor4_2 _26686_ (.A(_05810_),
    .B(_10542_),
    .C(net870),
    .Y(_07496_),
    .D(_07479_));
 sg13g2_o21ai_1 _26687_ (.B1(net186),
    .Y(_07497_),
    .A1(net187),
    .A2(_07496_));
 sg13g2_a22oi_1 _26688_ (.Y(_07498_),
    .B1(_07497_),
    .B2(\cpu.genblk1.mmu.r_valid_d[13] ),
    .A2(_07496_),
    .A1(net188));
 sg13g2_nor2_1 _26689_ (.A(_07452_),
    .B(_07498_),
    .Y(_01081_));
 sg13g2_inv_1 _26690_ (.Y(_07499_),
    .A(_05858_));
 sg13g2_nor2_1 _26691_ (.A(_07499_),
    .B(_07487_),
    .Y(_07500_));
 sg13g2_buf_2 _26692_ (.A(_07500_),
    .X(_07501_));
 sg13g2_nor2_1 _26693_ (.A(_05823_),
    .B(_07499_),
    .Y(_07502_));
 sg13g2_and2_1 _26694_ (.A(net455),
    .B(_07502_),
    .X(_07503_));
 sg13g2_o21ai_1 _26695_ (.B1(net186),
    .Y(_07504_),
    .A1(net187),
    .A2(_07503_));
 sg13g2_a22oi_1 _26696_ (.Y(_07505_),
    .B1(_07504_),
    .B2(\cpu.genblk1.mmu.r_valid_d[14] ),
    .A2(_07501_),
    .A1(_07480_));
 sg13g2_nor2_1 _26697_ (.A(net574),
    .B(_07505_),
    .Y(_01082_));
 sg13g2_and2_1 _26698_ (.A(_05828_),
    .B(net455),
    .X(_07506_));
 sg13g2_buf_1 _26699_ (.A(_07506_),
    .X(_07507_));
 sg13g2_o21ai_1 _26700_ (.B1(net186),
    .Y(_07508_),
    .A1(net187),
    .A2(_07507_));
 sg13g2_a22oi_1 _26701_ (.Y(_07509_),
    .B1(_07508_),
    .B2(\cpu.genblk1.mmu.r_valid_d[15] ),
    .A2(_07507_),
    .A1(net188));
 sg13g2_nor2_1 _26702_ (.A(net574),
    .B(_07509_),
    .Y(_01083_));
 sg13g2_nor3_1 _26703_ (.A(_07458_),
    .B(_10805_),
    .C(_05797_),
    .Y(_07510_));
 sg13g2_nor2b_1 _26704_ (.A(_07510_),
    .B_N(_07462_),
    .Y(_07511_));
 sg13g2_buf_2 _26705_ (.A(_07511_),
    .X(_07512_));
 sg13g2_nor2_1 _26706_ (.A(_05847_),
    .B(_05902_),
    .Y(_07513_));
 sg13g2_o21ai_1 _26707_ (.B1(_05803_),
    .Y(_07514_),
    .A1(_05828_),
    .A2(_07513_));
 sg13g2_o21ai_1 _26708_ (.B1(_05799_),
    .Y(_07515_),
    .A1(_07479_),
    .A2(_07514_));
 sg13g2_nand2_1 _26709_ (.Y(_07516_),
    .A(_07512_),
    .B(_07515_));
 sg13g2_a21oi_1 _26710_ (.A1(_05803_),
    .A2(_05847_),
    .Y(_07517_),
    .B1(_05311_));
 sg13g2_nor2b_1 _26711_ (.A(_05902_),
    .B_N(_07517_),
    .Y(_07518_));
 sg13g2_buf_1 _26712_ (.A(_07518_),
    .X(_07519_));
 sg13g2_and3_1 _26713_ (.X(_07520_),
    .A(_05799_),
    .B(net455),
    .C(_07519_));
 sg13g2_buf_1 _26714_ (.A(_07512_),
    .X(_07521_));
 sg13g2_a22oi_1 _26715_ (.Y(_07522_),
    .B1(_07520_),
    .B2(net185),
    .A2(_07516_),
    .A1(\cpu.genblk1.mmu.r_valid_d[16] ));
 sg13g2_nor2_1 _26716_ (.A(net574),
    .B(_07522_),
    .Y(_01084_));
 sg13g2_nor3_2 _26717_ (.A(_05810_),
    .B(net1024),
    .C(net972),
    .Y(_07523_));
 sg13g2_nor4_1 _26718_ (.A(net970),
    .B(net973),
    .C(_05836_),
    .D(net1083),
    .Y(_07524_));
 sg13g2_a21oi_1 _26719_ (.A1(net1083),
    .A2(_06207_),
    .Y(_07525_),
    .B1(_07524_));
 sg13g2_nand2b_1 _26720_ (.Y(_07526_),
    .B(_10483_),
    .A_N(net1083));
 sg13g2_a21oi_1 _26721_ (.A1(_07453_),
    .A2(_07526_),
    .Y(_07527_),
    .B1(_05836_));
 sg13g2_nand2_1 _26722_ (.Y(_07528_),
    .A(_05846_),
    .B(_07527_));
 sg13g2_o21ai_1 _26723_ (.B1(_07528_),
    .Y(_07529_),
    .A1(_06108_),
    .A2(_07525_));
 sg13g2_buf_2 _26724_ (.A(_07529_),
    .X(_07530_));
 sg13g2_and2_1 _26725_ (.A(_07523_),
    .B(_07530_),
    .X(_07531_));
 sg13g2_buf_1 _26726_ (.A(_07531_),
    .X(_07532_));
 sg13g2_and2_1 _26727_ (.A(_05799_),
    .B(_07462_),
    .X(_07533_));
 sg13g2_buf_1 _26728_ (.A(_07533_),
    .X(_07534_));
 sg13g2_and2_1 _26729_ (.A(net542),
    .B(_07534_),
    .X(_07535_));
 sg13g2_buf_2 _26730_ (.A(_07535_),
    .X(_07536_));
 sg13g2_buf_1 _26731_ (.A(_07460_),
    .X(_07537_));
 sg13g2_o21ai_1 _26732_ (.B1(net185),
    .Y(_07538_),
    .A1(net507),
    .A2(_07532_));
 sg13g2_a22oi_1 _26733_ (.Y(_07539_),
    .B1(_07538_),
    .B2(\cpu.genblk1.mmu.r_valid_d[17] ),
    .A2(_07536_),
    .A1(_07532_));
 sg13g2_nor2_1 _26734_ (.A(net574),
    .B(_07539_),
    .Y(_01085_));
 sg13g2_buf_1 _26735_ (.A(_07460_),
    .X(_07540_));
 sg13g2_o21ai_1 _26736_ (.B1(_07512_),
    .Y(_07541_),
    .A1(_07540_),
    .A2(_05910_));
 sg13g2_and2_1 _26737_ (.A(_07530_),
    .B(_07534_),
    .X(_07542_));
 sg13g2_buf_1 _26738_ (.A(_07542_),
    .X(_07543_));
 sg13g2_a22oi_1 _26739_ (.Y(_07544_),
    .B1(_07543_),
    .B2(_07472_),
    .A2(_07541_),
    .A1(\cpu.genblk1.mmu.r_valid_d[18] ));
 sg13g2_nor2_1 _26740_ (.A(net574),
    .B(_07544_),
    .Y(_01086_));
 sg13g2_buf_1 _26741_ (.A(_09389_),
    .X(_07545_));
 sg13g2_o21ai_1 _26742_ (.B1(net185),
    .Y(_07546_),
    .A1(net507),
    .A2(_05918_));
 sg13g2_a22oi_1 _26743_ (.Y(_07547_),
    .B1(_07546_),
    .B2(\cpu.genblk1.mmu.r_valid_d[19] ),
    .A2(_07536_),
    .A1(_05918_));
 sg13g2_nor2_1 _26744_ (.A(net573),
    .B(_07547_),
    .Y(_01087_));
 sg13g2_nor3_1 _26745_ (.A(net973),
    .B(net1083),
    .C(_05901_),
    .Y(_07548_));
 sg13g2_a21oi_1 _26746_ (.A1(net1083),
    .A2(_05877_),
    .Y(_07549_),
    .B1(_07548_));
 sg13g2_nand2_1 _26747_ (.Y(_07550_),
    .A(net1016),
    .B(_07527_));
 sg13g2_o21ai_1 _26748_ (.B1(_07550_),
    .Y(_07551_),
    .A1(_06108_),
    .A2(_07549_));
 sg13g2_buf_2 _26749_ (.A(_07551_),
    .X(_07552_));
 sg13g2_and2_1 _26750_ (.A(_07523_),
    .B(_07552_),
    .X(_07553_));
 sg13g2_buf_1 _26751_ (.A(_07553_),
    .X(_07554_));
 sg13g2_o21ai_1 _26752_ (.B1(net186),
    .Y(_07555_),
    .A1(net213),
    .A2(_07554_));
 sg13g2_a22oi_1 _26753_ (.Y(_07556_),
    .B1(_07555_),
    .B2(\cpu.genblk1.mmu.r_valid_d[1] ),
    .A2(_07554_),
    .A1(net188));
 sg13g2_nor2_1 _26754_ (.A(_07545_),
    .B(_07556_),
    .Y(_01088_));
 sg13g2_and2_1 _26755_ (.A(_07492_),
    .B(_07530_),
    .X(_07557_));
 sg13g2_o21ai_1 _26756_ (.B1(net185),
    .Y(_07558_),
    .A1(net507),
    .A2(_07557_));
 sg13g2_a22oi_1 _26757_ (.Y(_07559_),
    .B1(_07558_),
    .B2(\cpu.genblk1.mmu.r_valid_d[20] ),
    .A2(_07543_),
    .A1(_07489_));
 sg13g2_nor2_1 _26758_ (.A(net573),
    .B(_07559_),
    .Y(_01089_));
 sg13g2_nand3_1 _26759_ (.B(_05884_),
    .C(_07530_),
    .A(net972),
    .Y(_07560_));
 sg13g2_inv_1 _26760_ (.Y(_07561_),
    .A(_07560_));
 sg13g2_o21ai_1 _26761_ (.B1(net185),
    .Y(_07562_),
    .A1(net507),
    .A2(_07561_));
 sg13g2_a22oi_1 _26762_ (.Y(_07563_),
    .B1(_07562_),
    .B2(\cpu.genblk1.mmu.r_valid_d[21] ),
    .A2(_07561_),
    .A1(_07536_));
 sg13g2_nor2_1 _26763_ (.A(net573),
    .B(_07563_),
    .Y(_01090_));
 sg13g2_nor3_1 _26764_ (.A(net870),
    .B(_07499_),
    .C(_07528_),
    .Y(_07564_));
 sg13g2_o21ai_1 _26765_ (.B1(net185),
    .Y(_07565_),
    .A1(net507),
    .A2(_07564_));
 sg13g2_a22oi_1 _26766_ (.Y(_07566_),
    .B1(_07565_),
    .B2(\cpu.genblk1.mmu.r_valid_d[22] ),
    .A2(_07543_),
    .A1(_07501_));
 sg13g2_nor2_1 _26767_ (.A(net573),
    .B(_07566_),
    .Y(_01091_));
 sg13g2_nor3_2 _26768_ (.A(net1016),
    .B(_05810_),
    .C(_06004_),
    .Y(_07567_));
 sg13g2_o21ai_1 _26769_ (.B1(net185),
    .Y(_07568_),
    .A1(net507),
    .A2(_07567_));
 sg13g2_a22oi_1 _26770_ (.Y(_07569_),
    .B1(_07568_),
    .B2(\cpu.genblk1.mmu.r_valid_d[23] ),
    .A2(_07567_),
    .A1(_07536_));
 sg13g2_nor2_1 _26771_ (.A(net573),
    .B(_07569_),
    .Y(_01092_));
 sg13g2_nor2b_1 _26772_ (.A(_07514_),
    .B_N(_07530_),
    .Y(_07570_));
 sg13g2_o21ai_1 _26773_ (.B1(_07512_),
    .Y(_07571_),
    .A1(net506),
    .A2(_07570_));
 sg13g2_nand2_1 _26774_ (.Y(_07572_),
    .A(\cpu.genblk1.mmu.r_valid_d[24] ),
    .B(_07571_));
 sg13g2_nand3_1 _26775_ (.B(_07530_),
    .C(_07534_),
    .A(_07519_),
    .Y(_07573_));
 sg13g2_a21oi_1 _26776_ (.A1(_07572_),
    .A2(_07573_),
    .Y(_01093_),
    .B1(net575));
 sg13g2_a21o_1 _26777_ (.A2(_07475_),
    .A1(net970),
    .B1(_07455_),
    .X(_07574_));
 sg13g2_buf_1 _26778_ (.A(_07574_),
    .X(_07575_));
 sg13g2_and2_1 _26779_ (.A(_07523_),
    .B(net454),
    .X(_07576_));
 sg13g2_buf_1 _26780_ (.A(_07576_),
    .X(_07577_));
 sg13g2_o21ai_1 _26781_ (.B1(_07521_),
    .Y(_07578_),
    .A1(_07537_),
    .A2(_07577_));
 sg13g2_a22oi_1 _26782_ (.Y(_07579_),
    .B1(_07578_),
    .B2(\cpu.genblk1.mmu.r_valid_d[25] ),
    .A2(_07577_),
    .A1(_07536_));
 sg13g2_nor2_1 _26783_ (.A(net573),
    .B(_07579_),
    .Y(_01094_));
 sg13g2_o21ai_1 _26784_ (.B1(_07512_),
    .Y(_07580_),
    .A1(_07460_),
    .A2(_05956_));
 sg13g2_and2_1 _26785_ (.A(_07534_),
    .B(net454),
    .X(_07581_));
 sg13g2_buf_1 _26786_ (.A(_07581_),
    .X(_07582_));
 sg13g2_a22oi_1 _26787_ (.Y(_07583_),
    .B1(_07582_),
    .B2(_07472_),
    .A2(_07580_),
    .A1(\cpu.genblk1.mmu.r_valid_d[26] ));
 sg13g2_nor2_1 _26788_ (.A(net573),
    .B(_07583_),
    .Y(_01095_));
 sg13g2_o21ai_1 _26789_ (.B1(_07521_),
    .Y(_07584_),
    .A1(net507),
    .A2(_05961_));
 sg13g2_a22oi_1 _26790_ (.Y(_07585_),
    .B1(_07584_),
    .B2(\cpu.genblk1.mmu.r_valid_d[27] ),
    .A2(_07536_),
    .A1(_05961_));
 sg13g2_nor2_1 _26791_ (.A(_07545_),
    .B(_07585_),
    .Y(_01096_));
 sg13g2_and2_1 _26792_ (.A(_07492_),
    .B(_07575_),
    .X(_07586_));
 sg13g2_o21ai_1 _26793_ (.B1(_07512_),
    .Y(_07587_),
    .A1(net507),
    .A2(_07586_));
 sg13g2_a22oi_1 _26794_ (.Y(_07588_),
    .B1(_07587_),
    .B2(\cpu.genblk1.mmu.r_valid_d[28] ),
    .A2(_07582_),
    .A1(_07489_));
 sg13g2_nor2_1 _26795_ (.A(net573),
    .B(_07588_),
    .Y(_01097_));
 sg13g2_buf_1 _26796_ (.A(_09389_),
    .X(_07589_));
 sg13g2_and3_1 _26797_ (.X(_07590_),
    .A(net972),
    .B(_05884_),
    .C(net454));
 sg13g2_buf_1 _26798_ (.A(_07590_),
    .X(_07591_));
 sg13g2_o21ai_1 _26799_ (.B1(_07512_),
    .Y(_07592_),
    .A1(_07537_),
    .A2(_07591_));
 sg13g2_a22oi_1 _26800_ (.Y(_07593_),
    .B1(_07592_),
    .B2(\cpu.genblk1.mmu.r_valid_d[29] ),
    .A2(_07591_),
    .A1(_07536_));
 sg13g2_nor2_1 _26801_ (.A(net572),
    .B(_07593_),
    .Y(_01098_));
 sg13g2_inv_1 _26802_ (.Y(_07594_),
    .A(_07552_));
 sg13g2_nor2_1 _26803_ (.A(_05860_),
    .B(_07594_),
    .Y(_07595_));
 sg13g2_o21ai_1 _26804_ (.B1(_07467_),
    .Y(_07596_),
    .A1(_07464_),
    .A2(_07595_));
 sg13g2_nor3_1 _26805_ (.A(_05311_),
    .B(_05860_),
    .C(_07594_),
    .Y(_07597_));
 sg13g2_inv_1 _26806_ (.Y(_07598_),
    .A(_07481_));
 sg13g2_a22oi_1 _26807_ (.Y(_07599_),
    .B1(_07597_),
    .B2(_07598_),
    .A2(_07596_),
    .A1(\cpu.genblk1.mmu.r_valid_d[2] ));
 sg13g2_nor2_1 _26808_ (.A(net572),
    .B(_07599_),
    .Y(_01099_));
 sg13g2_a21oi_1 _26809_ (.A1(_07502_),
    .A2(net454),
    .Y(_07600_),
    .B1(_07460_));
 sg13g2_nand2b_1 _26810_ (.Y(_07601_),
    .B(net185),
    .A_N(_07600_));
 sg13g2_a22oi_1 _26811_ (.Y(_07602_),
    .B1(_07601_),
    .B2(\cpu.genblk1.mmu.r_valid_d[30] ),
    .A2(_07582_),
    .A1(_07501_));
 sg13g2_nor2_1 _26812_ (.A(net572),
    .B(_07602_),
    .Y(_01100_));
 sg13g2_and2_1 _26813_ (.A(_05828_),
    .B(net454),
    .X(_07603_));
 sg13g2_buf_1 _26814_ (.A(_07603_),
    .X(_07604_));
 sg13g2_o21ai_1 _26815_ (.B1(_07512_),
    .Y(_07605_),
    .A1(_07540_),
    .A2(_07604_));
 sg13g2_a22oi_1 _26816_ (.Y(_07606_),
    .B1(_07605_),
    .B2(\cpu.genblk1.mmu.r_valid_d[31] ),
    .A2(_07604_),
    .A1(_07536_));
 sg13g2_nor2_1 _26817_ (.A(net572),
    .B(_07606_),
    .Y(_01101_));
 sg13g2_and2_1 _26818_ (.A(_07490_),
    .B(_07552_),
    .X(_07607_));
 sg13g2_buf_1 _26819_ (.A(_07607_),
    .X(_07608_));
 sg13g2_o21ai_1 _26820_ (.B1(_07482_),
    .Y(_07609_),
    .A1(net213),
    .A2(_07608_));
 sg13g2_a22oi_1 _26821_ (.Y(_07610_),
    .B1(_07609_),
    .B2(\cpu.genblk1.mmu.r_valid_d[3] ),
    .A2(_07608_),
    .A1(net188));
 sg13g2_nor2_1 _26822_ (.A(net572),
    .B(_07610_),
    .Y(_01102_));
 sg13g2_nor2_1 _26823_ (.A(_07464_),
    .B(_07594_),
    .Y(_07611_));
 sg13g2_and2_1 _26824_ (.A(_07492_),
    .B(_07552_),
    .X(_07612_));
 sg13g2_o21ai_1 _26825_ (.B1(_07482_),
    .Y(_07613_),
    .A1(net213),
    .A2(_07612_));
 sg13g2_a22oi_1 _26826_ (.Y(_07614_),
    .B1(_07613_),
    .B2(\cpu.genblk1.mmu.r_valid_d[4] ),
    .A2(_07611_),
    .A1(_07489_));
 sg13g2_nor2_1 _26827_ (.A(net572),
    .B(_07614_),
    .Y(_01103_));
 sg13g2_o21ai_1 _26828_ (.B1(net186),
    .Y(_07615_),
    .A1(_05999_),
    .A2(net187));
 sg13g2_a22oi_1 _26829_ (.Y(_07616_),
    .B1(_07615_),
    .B2(\cpu.genblk1.mmu.r_valid_d[5] ),
    .A2(net188),
    .A1(_05999_));
 sg13g2_nor2_1 _26830_ (.A(net572),
    .B(_07616_),
    .Y(_01104_));
 sg13g2_o21ai_1 _26831_ (.B1(_07467_),
    .Y(_07617_),
    .A1(_06005_),
    .A2(net187));
 sg13g2_a22oi_1 _26832_ (.Y(_07618_),
    .B1(_07617_),
    .B2(\cpu.genblk1.mmu.r_valid_d[6] ),
    .A2(_07611_),
    .A1(_07501_));
 sg13g2_nor2_1 _26833_ (.A(_07589_),
    .B(_07618_),
    .Y(_01105_));
 sg13g2_o21ai_1 _26834_ (.B1(_07467_),
    .Y(_07619_),
    .A1(_06010_),
    .A2(_07481_));
 sg13g2_a22oi_1 _26835_ (.Y(_07620_),
    .B1(_07619_),
    .B2(\cpu.genblk1.mmu.r_valid_d[7] ),
    .A2(net188),
    .A1(_06010_));
 sg13g2_nor2_1 _26836_ (.A(_07589_),
    .B(_07620_),
    .Y(_01106_));
 sg13g2_nor2_1 _26837_ (.A(_07514_),
    .B(_07594_),
    .Y(_07621_));
 sg13g2_o21ai_1 _26838_ (.B1(_07467_),
    .Y(_07622_),
    .A1(net213),
    .A2(_07621_));
 sg13g2_a22oi_1 _26839_ (.Y(_07623_),
    .B1(_07622_),
    .B2(\cpu.genblk1.mmu.r_valid_d[8] ),
    .A2(_07611_),
    .A1(_07519_));
 sg13g2_nor2_1 _26840_ (.A(net572),
    .B(_07623_),
    .Y(_01107_));
 sg13g2_buf_1 _26841_ (.A(_06813_),
    .X(_07624_));
 sg13g2_and2_1 _26842_ (.A(net455),
    .B(_07523_),
    .X(_07625_));
 sg13g2_buf_1 _26843_ (.A(_07625_),
    .X(_07626_));
 sg13g2_o21ai_1 _26844_ (.B1(_07467_),
    .Y(_07627_),
    .A1(net213),
    .A2(_07626_));
 sg13g2_a22oi_1 _26845_ (.Y(_07628_),
    .B1(_07627_),
    .B2(\cpu.genblk1.mmu.r_valid_d[9] ),
    .A2(_07626_),
    .A1(net188));
 sg13g2_nor2_1 _26846_ (.A(_07624_),
    .B(_07628_),
    .Y(_01108_));
 sg13g2_nand2_1 _26847_ (.Y(_07629_),
    .A(net1052),
    .B(_00255_));
 sg13g2_a21oi_1 _26848_ (.A1(_07456_),
    .A2(_07629_),
    .Y(_07630_),
    .B1(_07460_));
 sg13g2_nor3_2 _26849_ (.A(_08431_),
    .B(_08525_),
    .C(_07630_),
    .Y(_07631_));
 sg13g2_nand2_1 _26850_ (.Y(_07632_),
    .A(_05799_),
    .B(_07631_));
 sg13g2_buf_1 _26851_ (.A(_07632_),
    .X(_07633_));
 sg13g2_nor3_1 _26852_ (.A(_07458_),
    .B(_10796_),
    .C(_05795_),
    .Y(_07634_));
 sg13g2_nor2b_1 _26853_ (.A(_07634_),
    .B_N(_07631_),
    .Y(_07635_));
 sg13g2_buf_2 _26854_ (.A(_07635_),
    .X(_07636_));
 sg13g2_o21ai_1 _26855_ (.B1(_07636_),
    .Y(_07637_),
    .A1(_07455_),
    .A2(_07633_));
 sg13g2_nor2_1 _26856_ (.A(_10172_),
    .B(_07633_),
    .Y(_07638_));
 sg13g2_buf_1 _26857_ (.A(_07638_),
    .X(_07639_));
 sg13g2_a22oi_1 _26858_ (.Y(_07640_),
    .B1(net153),
    .B2(_07455_),
    .A2(_07637_),
    .A1(\cpu.genblk1.mmu.r_valid_i[0] ));
 sg13g2_nor2_1 _26859_ (.A(net571),
    .B(_07640_),
    .Y(_01109_));
 sg13g2_and2_1 _26860_ (.A(_05799_),
    .B(_07631_),
    .X(_07641_));
 sg13g2_buf_1 _26861_ (.A(_07641_),
    .X(_07642_));
 sg13g2_and2_1 _26862_ (.A(_07472_),
    .B(_07642_),
    .X(_07643_));
 sg13g2_buf_1 _26863_ (.A(_07643_),
    .X(_07644_));
 sg13g2_buf_1 _26864_ (.A(_07633_),
    .X(_07645_));
 sg13g2_buf_1 _26865_ (.A(_07636_),
    .X(_07646_));
 sg13g2_o21ai_1 _26866_ (.B1(net183),
    .Y(_07647_),
    .A1(_05862_),
    .A2(net184));
 sg13g2_a22oi_1 _26867_ (.Y(_07648_),
    .B1(_07647_),
    .B2(\cpu.genblk1.mmu.r_valid_i[10] ),
    .A2(_07644_),
    .A1(net455));
 sg13g2_nor2_1 _26868_ (.A(net571),
    .B(_07648_),
    .Y(_01110_));
 sg13g2_o21ai_1 _26869_ (.B1(net183),
    .Y(_07649_),
    .A1(_05871_),
    .A2(net184));
 sg13g2_a22oi_1 _26870_ (.Y(_07650_),
    .B1(_07649_),
    .B2(\cpu.genblk1.mmu.r_valid_i[11] ),
    .A2(_07639_),
    .A1(_05871_));
 sg13g2_nor2_1 _26871_ (.A(net571),
    .B(_07650_),
    .Y(_01111_));
 sg13g2_and2_1 _26872_ (.A(_07489_),
    .B(_07642_),
    .X(_07651_));
 sg13g2_buf_1 _26873_ (.A(_07651_),
    .X(_07652_));
 sg13g2_o21ai_1 _26874_ (.B1(_07646_),
    .Y(_07653_),
    .A1(_07493_),
    .A2(net184));
 sg13g2_a22oi_1 _26875_ (.Y(_07654_),
    .B1(_07653_),
    .B2(\cpu.genblk1.mmu.r_valid_i[12] ),
    .A2(_07652_),
    .A1(_07478_));
 sg13g2_nor2_1 _26876_ (.A(_07624_),
    .B(_07654_),
    .Y(_01112_));
 sg13g2_o21ai_1 _26877_ (.B1(net183),
    .Y(_07655_),
    .A1(_07496_),
    .A2(net184));
 sg13g2_a22oi_1 _26878_ (.Y(_07656_),
    .B1(_07655_),
    .B2(\cpu.genblk1.mmu.r_valid_i[13] ),
    .A2(net153),
    .A1(_07496_));
 sg13g2_nor2_1 _26879_ (.A(net571),
    .B(_07656_),
    .Y(_01113_));
 sg13g2_and2_1 _26880_ (.A(_07501_),
    .B(_07642_),
    .X(_07657_));
 sg13g2_o21ai_1 _26881_ (.B1(_07646_),
    .Y(_07658_),
    .A1(_07503_),
    .A2(net184));
 sg13g2_a22oi_1 _26882_ (.Y(_07659_),
    .B1(_07658_),
    .B2(\cpu.genblk1.mmu.r_valid_i[14] ),
    .A2(_07657_),
    .A1(net455));
 sg13g2_nor2_1 _26883_ (.A(net571),
    .B(_07659_),
    .Y(_01114_));
 sg13g2_o21ai_1 _26884_ (.B1(net183),
    .Y(_07660_),
    .A1(_07507_),
    .A2(_07645_));
 sg13g2_a22oi_1 _26885_ (.Y(_07661_),
    .B1(_07660_),
    .B2(\cpu.genblk1.mmu.r_valid_i[15] ),
    .A2(net153),
    .A1(_07507_));
 sg13g2_nor2_1 _26886_ (.A(net571),
    .B(_07661_),
    .Y(_01115_));
 sg13g2_nor3_1 _26887_ (.A(_07458_),
    .B(_10937_),
    .C(_05797_),
    .Y(_07662_));
 sg13g2_nor2b_1 _26888_ (.A(_07662_),
    .B_N(_07631_),
    .Y(_07663_));
 sg13g2_buf_2 _26889_ (.A(_07663_),
    .X(_07664_));
 sg13g2_buf_1 _26890_ (.A(_07664_),
    .X(_07665_));
 sg13g2_nand2_1 _26891_ (.Y(_07666_),
    .A(_07515_),
    .B(net182));
 sg13g2_a22oi_1 _26892_ (.Y(_07667_),
    .B1(_07666_),
    .B2(\cpu.genblk1.mmu.r_valid_i[16] ),
    .A2(_07665_),
    .A1(_07520_));
 sg13g2_nor2_1 _26893_ (.A(net571),
    .B(_07667_),
    .Y(_01116_));
 sg13g2_o21ai_1 _26894_ (.B1(_07664_),
    .Y(_07668_),
    .A1(_07460_),
    .A2(_07532_));
 sg13g2_inv_1 _26895_ (.Y(_07669_),
    .A(_07664_));
 sg13g2_nor3_1 _26896_ (.A(_10172_),
    .B(_07460_),
    .C(_07669_),
    .Y(_07670_));
 sg13g2_buf_1 _26897_ (.A(_07670_),
    .X(_07671_));
 sg13g2_a22oi_1 _26898_ (.Y(_07672_),
    .B1(_07671_),
    .B2(_07532_),
    .A2(_07668_),
    .A1(\cpu.genblk1.mmu.r_valid_i[17] ));
 sg13g2_nor2_1 _26899_ (.A(net571),
    .B(_07672_),
    .Y(_01117_));
 sg13g2_buf_1 _26900_ (.A(_06813_),
    .X(_07673_));
 sg13g2_o21ai_1 _26901_ (.B1(net182),
    .Y(_07674_),
    .A1(net506),
    .A2(_05910_));
 sg13g2_a22oi_1 _26902_ (.Y(_07675_),
    .B1(_07674_),
    .B2(\cpu.genblk1.mmu.r_valid_i[18] ),
    .A2(_07644_),
    .A1(_07530_));
 sg13g2_nor2_1 _26903_ (.A(_07673_),
    .B(_07675_),
    .Y(_01118_));
 sg13g2_o21ai_1 _26904_ (.B1(net182),
    .Y(_07676_),
    .A1(net506),
    .A2(_05918_));
 sg13g2_a22oi_1 _26905_ (.Y(_07677_),
    .B1(_07676_),
    .B2(\cpu.genblk1.mmu.r_valid_i[19] ),
    .A2(_07671_),
    .A1(_05918_));
 sg13g2_nor2_1 _26906_ (.A(net570),
    .B(_07677_),
    .Y(_01119_));
 sg13g2_o21ai_1 _26907_ (.B1(net183),
    .Y(_07678_),
    .A1(_07554_),
    .A2(_07645_));
 sg13g2_a22oi_1 _26908_ (.Y(_07679_),
    .B1(_07678_),
    .B2(\cpu.genblk1.mmu.r_valid_i[1] ),
    .A2(net153),
    .A1(_07554_));
 sg13g2_nor2_1 _26909_ (.A(net570),
    .B(_07679_),
    .Y(_01120_));
 sg13g2_and2_1 _26910_ (.A(_07530_),
    .B(_07642_),
    .X(_07680_));
 sg13g2_buf_1 _26911_ (.A(_07680_),
    .X(_07681_));
 sg13g2_o21ai_1 _26912_ (.B1(_07665_),
    .Y(_07682_),
    .A1(_07557_),
    .A2(net184));
 sg13g2_a22oi_1 _26913_ (.Y(_07683_),
    .B1(_07682_),
    .B2(\cpu.genblk1.mmu.r_valid_i[20] ),
    .A2(_07681_),
    .A1(_07489_));
 sg13g2_nor2_1 _26914_ (.A(net570),
    .B(_07683_),
    .Y(_01121_));
 sg13g2_o21ai_1 _26915_ (.B1(net182),
    .Y(_07684_),
    .A1(net506),
    .A2(_07561_));
 sg13g2_a22oi_1 _26916_ (.Y(_07685_),
    .B1(_07684_),
    .B2(\cpu.genblk1.mmu.r_valid_i[21] ),
    .A2(_07671_),
    .A1(_07561_));
 sg13g2_nor2_1 _26917_ (.A(net570),
    .B(_07685_),
    .Y(_01122_));
 sg13g2_o21ai_1 _26918_ (.B1(net182),
    .Y(_07686_),
    .A1(_07564_),
    .A2(net184));
 sg13g2_a22oi_1 _26919_ (.Y(_07687_),
    .B1(_07686_),
    .B2(\cpu.genblk1.mmu.r_valid_i[22] ),
    .A2(_07681_),
    .A1(_07501_));
 sg13g2_nor2_1 _26920_ (.A(net570),
    .B(_07687_),
    .Y(_01123_));
 sg13g2_o21ai_1 _26921_ (.B1(net182),
    .Y(_07688_),
    .A1(net506),
    .A2(_07567_));
 sg13g2_a22oi_1 _26922_ (.Y(_07689_),
    .B1(_07688_),
    .B2(\cpu.genblk1.mmu.r_valid_i[23] ),
    .A2(_07671_),
    .A1(_07567_));
 sg13g2_nor2_1 _26923_ (.A(net570),
    .B(_07689_),
    .Y(_01124_));
 sg13g2_o21ai_1 _26924_ (.B1(net182),
    .Y(_07690_),
    .A1(_07570_),
    .A2(net184));
 sg13g2_a22oi_1 _26925_ (.Y(_07691_),
    .B1(_07690_),
    .B2(\cpu.genblk1.mmu.r_valid_i[24] ),
    .A2(_07681_),
    .A1(_07519_));
 sg13g2_nor2_1 _26926_ (.A(_07673_),
    .B(_07691_),
    .Y(_01125_));
 sg13g2_o21ai_1 _26927_ (.B1(net182),
    .Y(_07692_),
    .A1(net506),
    .A2(_07577_));
 sg13g2_a22oi_1 _26928_ (.Y(_07693_),
    .B1(_07692_),
    .B2(\cpu.genblk1.mmu.r_valid_i[25] ),
    .A2(_07671_),
    .A1(_07577_));
 sg13g2_nor2_1 _26929_ (.A(net570),
    .B(_07693_),
    .Y(_01126_));
 sg13g2_o21ai_1 _26930_ (.B1(_07664_),
    .Y(_07694_),
    .A1(net506),
    .A2(_05956_));
 sg13g2_a22oi_1 _26931_ (.Y(_07695_),
    .B1(_07694_),
    .B2(\cpu.genblk1.mmu.r_valid_i[26] ),
    .A2(_07644_),
    .A1(net454));
 sg13g2_nor2_1 _26932_ (.A(net570),
    .B(_07695_),
    .Y(_01127_));
 sg13g2_buf_1 _26933_ (.A(_06813_),
    .X(_07696_));
 sg13g2_o21ai_1 _26934_ (.B1(_07664_),
    .Y(_07697_),
    .A1(net506),
    .A2(_05961_));
 sg13g2_a22oi_1 _26935_ (.Y(_07698_),
    .B1(_07697_),
    .B2(\cpu.genblk1.mmu.r_valid_i[27] ),
    .A2(_07671_),
    .A1(_05961_));
 sg13g2_nor2_1 _26936_ (.A(net569),
    .B(_07698_),
    .Y(_01128_));
 sg13g2_buf_1 _26937_ (.A(_07633_),
    .X(_07699_));
 sg13g2_o21ai_1 _26938_ (.B1(_07664_),
    .Y(_07700_),
    .A1(_07586_),
    .A2(net181));
 sg13g2_a22oi_1 _26939_ (.Y(_07701_),
    .B1(_07700_),
    .B2(\cpu.genblk1.mmu.r_valid_i[28] ),
    .A2(_07652_),
    .A1(net454));
 sg13g2_nor2_1 _26940_ (.A(net569),
    .B(_07701_),
    .Y(_01129_));
 sg13g2_o21ai_1 _26941_ (.B1(_07664_),
    .Y(_07702_),
    .A1(_07591_),
    .A2(net181));
 sg13g2_a22oi_1 _26942_ (.Y(_07703_),
    .B1(_07702_),
    .B2(\cpu.genblk1.mmu.r_valid_i[29] ),
    .A2(net153),
    .A1(_07591_));
 sg13g2_nor2_1 _26943_ (.A(net569),
    .B(_07703_),
    .Y(_01130_));
 sg13g2_o21ai_1 _26944_ (.B1(net183),
    .Y(_07704_),
    .A1(_07595_),
    .A2(_07699_));
 sg13g2_a22oi_1 _26945_ (.Y(_07705_),
    .B1(_07704_),
    .B2(\cpu.genblk1.mmu.r_valid_i[2] ),
    .A2(_07642_),
    .A1(_07597_));
 sg13g2_nor2_1 _26946_ (.A(net569),
    .B(_07705_),
    .Y(_01131_));
 sg13g2_nand4_1 _26947_ (.B(_07501_),
    .C(net454),
    .A(_05799_),
    .Y(_07706_),
    .D(_07631_));
 sg13g2_o21ai_1 _26948_ (.B1(\cpu.genblk1.mmu.r_valid_i[30] ),
    .Y(_07707_),
    .A1(_07600_),
    .A2(_07669_));
 sg13g2_a21oi_1 _26949_ (.A1(_07706_),
    .A2(_07707_),
    .Y(_01132_),
    .B1(net575));
 sg13g2_o21ai_1 _26950_ (.B1(_07664_),
    .Y(_07708_),
    .A1(_07604_),
    .A2(net181));
 sg13g2_a22oi_1 _26951_ (.Y(_07709_),
    .B1(_07708_),
    .B2(\cpu.genblk1.mmu.r_valid_i[31] ),
    .A2(net153),
    .A1(_07604_));
 sg13g2_nor2_1 _26952_ (.A(net569),
    .B(_07709_),
    .Y(_01133_));
 sg13g2_o21ai_1 _26953_ (.B1(net183),
    .Y(_07710_),
    .A1(_07608_),
    .A2(net181));
 sg13g2_a22oi_1 _26954_ (.Y(_07711_),
    .B1(_07710_),
    .B2(\cpu.genblk1.mmu.r_valid_i[3] ),
    .A2(_07639_),
    .A1(_07608_));
 sg13g2_nor2_1 _26955_ (.A(_07696_),
    .B(_07711_),
    .Y(_01134_));
 sg13g2_o21ai_1 _26956_ (.B1(net183),
    .Y(_07712_),
    .A1(_07612_),
    .A2(_07699_));
 sg13g2_a22oi_1 _26957_ (.Y(_07713_),
    .B1(_07712_),
    .B2(\cpu.genblk1.mmu.r_valid_i[4] ),
    .A2(_07652_),
    .A1(_07552_));
 sg13g2_nor2_1 _26958_ (.A(net569),
    .B(_07713_),
    .Y(_01135_));
 sg13g2_o21ai_1 _26959_ (.B1(_07636_),
    .Y(_07714_),
    .A1(_05999_),
    .A2(net181));
 sg13g2_a22oi_1 _26960_ (.Y(_07715_),
    .B1(_07714_),
    .B2(\cpu.genblk1.mmu.r_valid_i[5] ),
    .A2(net153),
    .A1(_05999_));
 sg13g2_nor2_1 _26961_ (.A(_07696_),
    .B(_07715_),
    .Y(_01136_));
 sg13g2_nand3_1 _26962_ (.B(_07552_),
    .C(_07642_),
    .A(_07501_),
    .Y(_07716_));
 sg13g2_o21ai_1 _26963_ (.B1(_07636_),
    .Y(_07717_),
    .A1(_06005_),
    .A2(_07633_));
 sg13g2_nand2_1 _26964_ (.Y(_07718_),
    .A(\cpu.genblk1.mmu.r_valid_i[6] ),
    .B(_07717_));
 sg13g2_a21oi_1 _26965_ (.A1(_07716_),
    .A2(_07718_),
    .Y(_01137_),
    .B1(_07436_));
 sg13g2_o21ai_1 _26966_ (.B1(_07636_),
    .Y(_07719_),
    .A1(_06010_),
    .A2(net181));
 sg13g2_a22oi_1 _26967_ (.Y(_07720_),
    .B1(_07719_),
    .B2(\cpu.genblk1.mmu.r_valid_i[7] ),
    .A2(net153),
    .A1(_06010_));
 sg13g2_nor2_1 _26968_ (.A(net569),
    .B(_07720_),
    .Y(_01138_));
 sg13g2_o21ai_1 _26969_ (.B1(_07636_),
    .Y(_07721_),
    .A1(_07621_),
    .A2(net181));
 sg13g2_nand2_1 _26970_ (.Y(_07722_),
    .A(\cpu.genblk1.mmu.r_valid_i[8] ),
    .B(_07721_));
 sg13g2_nand3_1 _26971_ (.B(_07552_),
    .C(_07642_),
    .A(_07519_),
    .Y(_07723_));
 sg13g2_a21oi_1 _26972_ (.A1(_07722_),
    .A2(_07723_),
    .Y(_01139_),
    .B1(_07436_));
 sg13g2_o21ai_1 _26973_ (.B1(_07636_),
    .Y(_07724_),
    .A1(_07626_),
    .A2(net181));
 sg13g2_a22oi_1 _26974_ (.Y(_07725_),
    .B1(_07724_),
    .B2(\cpu.genblk1.mmu.r_valid_i[9] ),
    .A2(_07638_),
    .A1(_07626_));
 sg13g2_nor2_1 _26975_ (.A(net569),
    .B(_07725_),
    .Y(_01140_));
 sg13g2_nor3_1 _26976_ (.A(_12066_),
    .B(_04994_),
    .C(_06387_),
    .Y(_07726_));
 sg13g2_buf_2 _26977_ (.A(_07726_),
    .X(_07727_));
 sg13g2_nand2_1 _26978_ (.Y(_07728_),
    .A(_10241_),
    .B(_07727_));
 sg13g2_nand4_1 _26979_ (.B(_09866_),
    .C(_04996_),
    .A(net983),
    .Y(_07729_),
    .D(_06385_));
 sg13g2_buf_2 _26980_ (.A(_07729_),
    .X(_07730_));
 sg13g2_nand2_1 _26981_ (.Y(_07731_),
    .A(_09287_),
    .B(_07730_));
 sg13g2_a21oi_1 _26982_ (.A1(_07728_),
    .A2(_07731_),
    .Y(_01941_),
    .B1(net575));
 sg13g2_nand2_1 _26983_ (.Y(_07732_),
    .A(_06824_),
    .B(_07727_));
 sg13g2_nand2_1 _26984_ (.Y(_07733_),
    .A(_09301_),
    .B(_07730_));
 sg13g2_a21oi_1 _26985_ (.A1(_07732_),
    .A2(_07733_),
    .Y(_01942_),
    .B1(net575));
 sg13g2_nand2_1 _26986_ (.Y(_07734_),
    .A(net892),
    .B(_07727_));
 sg13g2_nand2_1 _26987_ (.Y(_07735_),
    .A(_09307_),
    .B(_07730_));
 sg13g2_a21oi_1 _26988_ (.A1(_07734_),
    .A2(_07735_),
    .Y(_01943_),
    .B1(net575));
 sg13g2_nand2_1 _26989_ (.Y(_07736_),
    .A(net1038),
    .B(_07727_));
 sg13g2_nand2_1 _26990_ (.Y(_07737_),
    .A(_09296_),
    .B(_07730_));
 sg13g2_buf_1 _26991_ (.A(_06813_),
    .X(_07738_));
 sg13g2_a21oi_1 _26992_ (.A1(_07736_),
    .A2(_07737_),
    .Y(_01944_),
    .B1(net568));
 sg13g2_nand2_1 _26993_ (.Y(_07739_),
    .A(_10215_),
    .B(_07727_));
 sg13g2_nand2_1 _26994_ (.Y(_07740_),
    .A(_09303_),
    .B(_07730_));
 sg13g2_a21oi_1 _26995_ (.A1(_07739_),
    .A2(_07740_),
    .Y(_01945_),
    .B1(net568));
 sg13g2_nand2_1 _26996_ (.Y(_07741_),
    .A(_10221_),
    .B(_07727_));
 sg13g2_nand2_1 _26997_ (.Y(_07742_),
    .A(_09309_),
    .B(_07730_));
 sg13g2_a21oi_1 _26998_ (.A1(_07741_),
    .A2(_07742_),
    .Y(_01946_),
    .B1(net568));
 sg13g2_nand2_1 _26999_ (.Y(_07743_),
    .A(_10227_),
    .B(_07727_));
 sg13g2_nand2_1 _27000_ (.Y(_07744_),
    .A(_09298_),
    .B(_07730_));
 sg13g2_a21oi_1 _27001_ (.A1(_07743_),
    .A2(_07744_),
    .Y(_01947_),
    .B1(net568));
 sg13g2_nand2_1 _27002_ (.Y(_07745_),
    .A(net985),
    .B(_07727_));
 sg13g2_nand2_1 _27003_ (.Y(_07746_),
    .A(_09289_),
    .B(_07730_));
 sg13g2_a21oi_1 _27004_ (.A1(_07745_),
    .A2(_07746_),
    .Y(_01948_),
    .B1(net568));
 sg13g2_nor3_1 _27005_ (.A(_12066_),
    .B(_04883_),
    .C(_06387_),
    .Y(_07747_));
 sg13g2_buf_2 _27006_ (.A(_07747_),
    .X(_07748_));
 sg13g2_nand2_1 _27007_ (.Y(_07749_),
    .A(net1037),
    .B(_07748_));
 sg13g2_nand2b_1 _27008_ (.Y(_07750_),
    .B(\cpu.gpio.r_enable_io[4] ),
    .A_N(_07748_));
 sg13g2_a21oi_1 _27009_ (.A1(_07749_),
    .A2(_07750_),
    .Y(_01949_),
    .B1(net568));
 sg13g2_nand2_1 _27010_ (.Y(_07751_),
    .A(net1036),
    .B(_07748_));
 sg13g2_nand2b_1 _27011_ (.Y(_07752_),
    .B(_09312_),
    .A_N(_07748_));
 sg13g2_a21oi_1 _27012_ (.A1(_07751_),
    .A2(_07752_),
    .Y(_01950_),
    .B1(net568));
 sg13g2_nand2_1 _27013_ (.Y(_07753_),
    .A(_10227_),
    .B(_07748_));
 sg13g2_nand2b_1 _27014_ (.Y(_07754_),
    .B(_09314_),
    .A_N(_07748_));
 sg13g2_a21oi_1 _27015_ (.A1(_07753_),
    .A2(_07754_),
    .Y(_01951_),
    .B1(net568));
 sg13g2_nand2_1 _27016_ (.Y(_07755_),
    .A(_02785_),
    .B(_07748_));
 sg13g2_nand2b_1 _27017_ (.Y(_07756_),
    .B(_09293_),
    .A_N(_07748_));
 sg13g2_a21oi_1 _27018_ (.A1(_07755_),
    .A2(_07756_),
    .Y(_01952_),
    .B1(_07738_));
 sg13g2_nor4_1 _27019_ (.A(net542),
    .B(net872),
    .C(_09836_),
    .D(_06387_),
    .Y(_07757_));
 sg13g2_buf_2 _27020_ (.A(_07757_),
    .X(_07758_));
 sg13g2_nand2_1 _27021_ (.Y(_07759_),
    .A(_10215_),
    .B(_07758_));
 sg13g2_nand2b_1 _27022_ (.Y(_07760_),
    .B(net7),
    .A_N(_07758_));
 sg13g2_a21oi_1 _27023_ (.A1(_07759_),
    .A2(_07760_),
    .Y(_01953_),
    .B1(_07738_));
 sg13g2_nand2_1 _27024_ (.Y(_07761_),
    .A(_10221_),
    .B(_07758_));
 sg13g2_nand2b_1 _27025_ (.Y(_07762_),
    .B(net8),
    .A_N(_07758_));
 sg13g2_buf_1 _27026_ (.A(_09452_),
    .X(_07763_));
 sg13g2_a21oi_1 _27027_ (.A1(_07761_),
    .A2(_07762_),
    .Y(_01954_),
    .B1(net567));
 sg13g2_nand2_1 _27028_ (.Y(_07764_),
    .A(net1035),
    .B(_07758_));
 sg13g2_nand2b_1 _27029_ (.Y(_07765_),
    .B(net9),
    .A_N(_07758_));
 sg13g2_a21oi_1 _27030_ (.A1(_07764_),
    .A2(_07765_),
    .Y(_01955_),
    .B1(net567));
 sg13g2_nand2_1 _27031_ (.Y(_07766_),
    .A(net985),
    .B(_07758_));
 sg13g2_nand2b_1 _27032_ (.Y(_07767_),
    .B(net10),
    .A_N(_07758_));
 sg13g2_a21oi_1 _27033_ (.A1(_07766_),
    .A2(_07767_),
    .Y(_01956_),
    .B1(net567));
 sg13g2_nor2_1 _27034_ (.A(net343),
    .B(net96),
    .Y(_07768_));
 sg13g2_nand2_1 _27035_ (.Y(_07769_),
    .A(net893),
    .B(_07768_));
 sg13g2_o21ai_1 _27036_ (.B1(_05000_),
    .Y(_07770_),
    .A1(net343),
    .A2(net96));
 sg13g2_nand3_1 _27037_ (.B(_07769_),
    .C(_07770_),
    .A(net650),
    .Y(_02002_));
 sg13g2_nand2_1 _27038_ (.Y(_07771_),
    .A(net966),
    .B(_07768_));
 sg13g2_buf_1 _27039_ (.A(\cpu.gpio.r_src_o[6][1] ),
    .X(_07772_));
 sg13g2_o21ai_1 _27040_ (.B1(_07772_),
    .Y(_07773_),
    .A1(net343),
    .A2(net96));
 sg13g2_a21oi_1 _27041_ (.A1(_07771_),
    .A2(_07773_),
    .Y(_02003_),
    .B1(net567));
 sg13g2_nand2_1 _27042_ (.Y(_07774_),
    .A(_10202_),
    .B(_07768_));
 sg13g2_o21ai_1 _27043_ (.B1(\cpu.gpio.r_src_o[6][2] ),
    .Y(_07775_),
    .A1(net343),
    .A2(net96));
 sg13g2_a21oi_1 _27044_ (.A1(_07774_),
    .A2(_07775_),
    .Y(_02004_),
    .B1(net567));
 sg13g2_nand2_1 _27045_ (.Y(_07776_),
    .A(_10209_),
    .B(_07768_));
 sg13g2_o21ai_1 _27046_ (.B1(\cpu.gpio.r_src_o[6][3] ),
    .Y(_07777_),
    .A1(net343),
    .A2(net96));
 sg13g2_a21oi_1 _27047_ (.A1(_07776_),
    .A2(_07777_),
    .Y(_02005_),
    .B1(net567));
 sg13g2_nor2_1 _27048_ (.A(_05346_),
    .B(net96),
    .Y(_07778_));
 sg13g2_nand2_1 _27049_ (.Y(_07779_),
    .A(net919),
    .B(_07778_));
 sg13g2_o21ai_1 _27050_ (.B1(_04998_),
    .Y(_07780_),
    .A1(_05346_),
    .A2(net96));
 sg13g2_a21oi_1 _27051_ (.A1(_07779_),
    .A2(_07780_),
    .Y(_02010_),
    .B1(net567));
 sg13g2_nand2_1 _27052_ (.Y(_07781_),
    .A(net966),
    .B(_07778_));
 sg13g2_o21ai_1 _27053_ (.B1(\cpu.gpio.r_uart_rx_src[1] ),
    .Y(_07782_),
    .A1(_05346_),
    .A2(_06404_));
 sg13g2_a21oi_1 _27054_ (.A1(_07781_),
    .A2(_07782_),
    .Y(_02011_),
    .B1(net567));
 sg13g2_nand2_1 _27055_ (.Y(_07783_),
    .A(_10202_),
    .B(_07778_));
 sg13g2_o21ai_1 _27056_ (.B1(\cpu.gpio.r_uart_rx_src[2] ),
    .Y(_07784_),
    .A1(_05346_),
    .A2(_06404_));
 sg13g2_a21oi_1 _27057_ (.A1(_07783_),
    .A2(_07784_),
    .Y(_02012_),
    .B1(_07763_));
 sg13g2_and2_1 _27058_ (.A(\cpu.i_wstrobe_d ),
    .B(_00316_),
    .X(_02269_));
 sg13g2_nor2_1 _27059_ (.A(_06422_),
    .B(_06434_),
    .Y(_07785_));
 sg13g2_nor2_1 _27060_ (.A(_06448_),
    .B(_07785_),
    .Y(_02270_));
 sg13g2_xor2_1 _27061_ (.B(_06429_),
    .A(\cpu.icache.r_offset[2] ),
    .X(_07786_));
 sg13g2_nor2_1 _27062_ (.A(_06448_),
    .B(_07786_),
    .Y(_02271_));
 sg13g2_buf_1 _27063_ (.A(_06813_),
    .X(_07787_));
 sg13g2_nand4_1 _27064_ (.B(_10194_),
    .C(net124),
    .A(net437),
    .Y(_07788_),
    .D(_04891_));
 sg13g2_xnor2_1 _27065_ (.Y(_07789_),
    .A(\cpu.intr.r_clock_cmp[3] ),
    .B(_10270_));
 sg13g2_xnor2_1 _27066_ (.Y(_07790_),
    .A(\cpu.intr.r_clock_cmp[0] ),
    .B(_10260_));
 sg13g2_xnor2_1 _27067_ (.Y(_07791_),
    .A(\cpu.intr.r_clock_cmp[20] ),
    .B(_05559_));
 sg13g2_xnor2_1 _27068_ (.Y(_07792_),
    .A(\cpu.intr.r_clock_cmp[17] ),
    .B(_05360_));
 sg13g2_nand4_1 _27069_ (.B(_07790_),
    .C(_07791_),
    .A(_07789_),
    .Y(_07793_),
    .D(_07792_));
 sg13g2_xnor2_1 _27070_ (.Y(_07794_),
    .A(\cpu.intr.r_clock_cmp[31] ),
    .B(_05275_));
 sg13g2_xnor2_1 _27071_ (.Y(_07795_),
    .A(\cpu.intr.r_clock_cmp[2] ),
    .B(_10265_));
 sg13g2_xnor2_1 _27072_ (.Y(_07796_),
    .A(\cpu.intr.r_clock_cmp[25] ),
    .B(_05739_));
 sg13g2_xnor2_1 _27073_ (.Y(_07797_),
    .A(\cpu.intr.r_clock_cmp[23] ),
    .B(_05037_));
 sg13g2_nand4_1 _27074_ (.B(_07795_),
    .C(_07796_),
    .A(_07794_),
    .Y(_07798_),
    .D(_07797_));
 sg13g2_xnor2_1 _27075_ (.Y(_07799_),
    .A(\cpu.intr.r_clock_cmp[8] ),
    .B(_10297_));
 sg13g2_xnor2_1 _27076_ (.Y(_07800_),
    .A(\cpu.intr.r_clock_cmp[19] ),
    .B(_05488_));
 sg13g2_xnor2_1 _27077_ (.Y(_07801_),
    .A(\cpu.intr.r_clock_cmp[6] ),
    .B(_10289_));
 sg13g2_xnor2_1 _27078_ (.Y(_07802_),
    .A(\cpu.intr.r_clock_cmp[29] ),
    .B(_05208_));
 sg13g2_nand4_1 _27079_ (.B(_07800_),
    .C(_07801_),
    .A(_07799_),
    .Y(_07803_),
    .D(_07802_));
 sg13g2_xnor2_1 _27080_ (.Y(_07804_),
    .A(\cpu.intr.r_clock_cmp[27] ),
    .B(_05164_));
 sg13g2_xnor2_1 _27081_ (.Y(_07805_),
    .A(\cpu.intr.r_clock_cmp[14] ),
    .B(_10333_));
 sg13g2_xnor2_1 _27082_ (.Y(_07806_),
    .A(\cpu.intr.r_clock_cmp[12] ),
    .B(_10321_));
 sg13g2_xnor2_1 _27083_ (.Y(_07807_),
    .A(\cpu.intr.r_clock_cmp[18] ),
    .B(_05416_));
 sg13g2_nand4_1 _27084_ (.B(_07805_),
    .C(_07806_),
    .A(_07804_),
    .Y(_07808_),
    .D(_07807_));
 sg13g2_nor4_1 _27085_ (.A(_07793_),
    .B(_07798_),
    .C(_07803_),
    .D(_07808_),
    .Y(_07809_));
 sg13g2_xnor2_1 _27086_ (.Y(_07810_),
    .A(\cpu.intr.r_clock_cmp[16] ),
    .B(_04954_));
 sg13g2_xnor2_1 _27087_ (.Y(_07811_),
    .A(\cpu.intr.r_clock_cmp[30] ),
    .B(_05241_));
 sg13g2_xnor2_1 _27088_ (.Y(_07812_),
    .A(\cpu.intr.r_clock_cmp[21] ),
    .B(_05623_));
 sg13g2_xnor2_1 _27089_ (.Y(_07813_),
    .A(\cpu.intr.r_clock_cmp[15] ),
    .B(_10341_));
 sg13g2_nand4_1 _27090_ (.B(_07811_),
    .C(_07812_),
    .A(_07810_),
    .Y(_07814_),
    .D(_07813_));
 sg13g2_xnor2_1 _27091_ (.Y(_07815_),
    .A(\cpu.intr.r_clock_cmp[5] ),
    .B(_10283_));
 sg13g2_xnor2_1 _27092_ (.Y(_07816_),
    .A(\cpu.intr.r_clock_cmp[26] ),
    .B(_05133_));
 sg13g2_xnor2_1 _27093_ (.Y(_07817_),
    .A(\cpu.intr.r_clock_cmp[22] ),
    .B(_05655_));
 sg13g2_xnor2_1 _27094_ (.Y(_07818_),
    .A(\cpu.intr.r_clock_cmp[10] ),
    .B(_10309_));
 sg13g2_nand4_1 _27095_ (.B(_07816_),
    .C(_07817_),
    .A(_07815_),
    .Y(_07819_),
    .D(_07818_));
 sg13g2_xnor2_1 _27096_ (.Y(_07820_),
    .A(\cpu.intr.r_clock_cmp[7] ),
    .B(_10293_));
 sg13g2_xnor2_1 _27097_ (.Y(_07821_),
    .A(\cpu.intr.r_clock_cmp[11] ),
    .B(_10314_));
 sg13g2_xnor2_1 _27098_ (.Y(_07822_),
    .A(\cpu.intr.r_clock_cmp[24] ),
    .B(_05725_));
 sg13g2_xnor2_1 _27099_ (.Y(_07823_),
    .A(\cpu.intr.r_clock_cmp[4] ),
    .B(_10277_));
 sg13g2_nand4_1 _27100_ (.B(_07821_),
    .C(_07822_),
    .A(_07820_),
    .Y(_07824_),
    .D(_07823_));
 sg13g2_xnor2_1 _27101_ (.Y(_07825_),
    .A(\cpu.intr.r_clock_cmp[1] ),
    .B(_10261_));
 sg13g2_xnor2_1 _27102_ (.Y(_07826_),
    .A(\cpu.intr.r_clock_cmp[13] ),
    .B(_10327_));
 sg13g2_xnor2_1 _27103_ (.Y(_07827_),
    .A(\cpu.intr.r_clock_cmp[28] ),
    .B(_05194_));
 sg13g2_xnor2_1 _27104_ (.Y(_07828_),
    .A(\cpu.intr.r_clock_cmp[9] ),
    .B(_10304_));
 sg13g2_nand4_1 _27105_ (.B(_07826_),
    .C(_07827_),
    .A(_07825_),
    .Y(_07829_),
    .D(_07828_));
 sg13g2_nor4_1 _27106_ (.A(_07814_),
    .B(_07819_),
    .C(_07824_),
    .D(_07829_),
    .Y(_07830_));
 sg13g2_nor2_1 _27107_ (.A(net542),
    .B(_07788_),
    .Y(_07831_));
 sg13g2_a221oi_1 _27108_ (.B2(_07830_),
    .C1(_07831_),
    .B1(_07809_),
    .A1(\cpu.intr.r_clock ),
    .Y(_07832_),
    .A2(_07788_));
 sg13g2_nor2_1 _27109_ (.A(_07787_),
    .B(_07832_),
    .Y(_02432_));
 sg13g2_and2_1 _27110_ (.A(net124),
    .B(net382),
    .X(_07833_));
 sg13g2_buf_1 _27111_ (.A(_07833_),
    .X(_07834_));
 sg13g2_nand2_1 _27112_ (.Y(_07835_),
    .A(net919),
    .B(_07834_));
 sg13g2_nand2_1 _27113_ (.Y(_07836_),
    .A(net124),
    .B(net382));
 sg13g2_buf_1 _27114_ (.A(_07836_),
    .X(_07837_));
 sg13g2_nand2_1 _27115_ (.Y(_07838_),
    .A(\cpu.intr.r_enable[0] ),
    .B(_07837_));
 sg13g2_a21oi_1 _27116_ (.A1(_07835_),
    .A2(_07838_),
    .Y(_02481_),
    .B1(_07763_));
 sg13g2_nand2_1 _27117_ (.Y(_07839_),
    .A(net966),
    .B(_07834_));
 sg13g2_nand2_1 _27118_ (.Y(_07840_),
    .A(_09325_),
    .B(_07837_));
 sg13g2_buf_1 _27119_ (.A(_09452_),
    .X(_07841_));
 sg13g2_a21oi_1 _27120_ (.A1(_07839_),
    .A2(_07840_),
    .Y(_02482_),
    .B1(net565));
 sg13g2_nand2_1 _27121_ (.Y(_07842_),
    .A(net920),
    .B(_07834_));
 sg13g2_nand2_1 _27122_ (.Y(_07843_),
    .A(\cpu.intr.r_enable[2] ),
    .B(_07837_));
 sg13g2_a21oi_1 _27123_ (.A1(_07842_),
    .A2(_07843_),
    .Y(_02483_),
    .B1(net565));
 sg13g2_nand2_1 _27124_ (.Y(_07844_),
    .A(net1038),
    .B(_07834_));
 sg13g2_nand2_1 _27125_ (.Y(_07845_),
    .A(\cpu.intr.r_enable[3] ),
    .B(_07837_));
 sg13g2_a21oi_1 _27126_ (.A1(_07844_),
    .A2(_07845_),
    .Y(_02484_),
    .B1(_07841_));
 sg13g2_nand2_1 _27127_ (.Y(_07846_),
    .A(net1037),
    .B(_07834_));
 sg13g2_nand2_1 _27128_ (.Y(_07847_),
    .A(_09318_),
    .B(_07837_));
 sg13g2_a21oi_1 _27129_ (.A1(_07846_),
    .A2(_07847_),
    .Y(_02485_),
    .B1(net565));
 sg13g2_nand2_1 _27130_ (.Y(_07848_),
    .A(net1036),
    .B(_07834_));
 sg13g2_nand2_1 _27131_ (.Y(_07849_),
    .A(_09323_),
    .B(_07837_));
 sg13g2_a21oi_1 _27132_ (.A1(_07848_),
    .A2(_07849_),
    .Y(_02486_),
    .B1(_07841_));
 sg13g2_nand3_1 _27133_ (.B(net124),
    .C(_04930_),
    .A(net1039),
    .Y(_07850_));
 sg13g2_nand3_1 _27134_ (.B(_06745_),
    .C(_04934_),
    .A(_10200_),
    .Y(_07851_));
 sg13g2_nand2_1 _27135_ (.Y(_07852_),
    .A(_10114_),
    .B(_07851_));
 sg13g2_a21oi_1 _27136_ (.A1(_09321_),
    .A2(_07850_),
    .Y(_07853_),
    .B1(_07852_));
 sg13g2_nor2_1 _27137_ (.A(_07787_),
    .B(_07853_),
    .Y(_02487_));
 sg13g2_nand3_1 _27138_ (.B(_06762_),
    .C(_06873_),
    .A(_06767_),
    .Y(_07854_));
 sg13g2_nor2_1 _27139_ (.A(_09954_),
    .B(_07854_),
    .Y(_07855_));
 sg13g2_nand4_1 _27140_ (.B(_06904_),
    .C(_06875_),
    .A(_09986_),
    .Y(_07856_),
    .D(_07855_));
 sg13g2_buf_1 _27141_ (.A(_07856_),
    .X(_07857_));
 sg13g2_o21ai_1 _27142_ (.B1(net803),
    .Y(_07858_),
    .A1(_06905_),
    .A2(_07857_));
 sg13g2_nor2_1 _27143_ (.A(_09964_),
    .B(_09979_),
    .Y(_07859_));
 sg13g2_o21ai_1 _27144_ (.B1(net19),
    .Y(_07860_),
    .A1(_07857_),
    .A2(_07859_));
 sg13g2_nand2b_1 _27145_ (.Y(_02517_),
    .B(_07860_),
    .A_N(_07858_));
 sg13g2_nand3_1 _27146_ (.B(_09964_),
    .C(_06870_),
    .A(_09939_),
    .Y(_07861_));
 sg13g2_a21o_1 _27147_ (.A2(_07861_),
    .A1(_06905_),
    .B1(_07857_),
    .X(_07862_));
 sg13g2_nand2_1 _27148_ (.Y(_07863_),
    .A(_00277_),
    .B(_06905_));
 sg13g2_nor2_1 _27149_ (.A(_09975_),
    .B(_07863_),
    .Y(_07864_));
 sg13g2_o21ai_1 _27150_ (.B1(net20),
    .Y(_07865_),
    .A1(_07857_),
    .A2(_07864_));
 sg13g2_nand3_1 _27151_ (.B(_07862_),
    .C(_07865_),
    .A(net650),
    .Y(_02518_));
 sg13g2_nor2_1 _27152_ (.A(_09964_),
    .B(_09977_),
    .Y(_07866_));
 sg13g2_buf_1 _27153_ (.A(\cpu.gpio.genblk1[3].srcs_o[11] ),
    .X(_07867_));
 sg13g2_o21ai_1 _27154_ (.B1(_07867_),
    .Y(_07868_),
    .A1(_07857_),
    .A2(_07866_));
 sg13g2_nand2b_1 _27155_ (.Y(_02519_),
    .B(_07868_),
    .A_N(_07858_));
 sg13g2_nor4_1 _27156_ (.A(\cpu.qspi.r_state[17] ),
    .B(_09947_),
    .C(_09963_),
    .D(_06870_),
    .Y(_07869_));
 sg13g2_nand2_1 _27157_ (.Y(_07870_),
    .A(_06761_),
    .B(_07869_));
 sg13g2_nor4_1 _27158_ (.A(_09948_),
    .B(_09987_),
    .C(_07854_),
    .D(_07870_),
    .Y(_07871_));
 sg13g2_a21oi_1 _27159_ (.A1(_12005_),
    .A2(_07871_),
    .Y(_07872_),
    .B1(_09939_));
 sg13g2_nor2_1 _27160_ (.A(net566),
    .B(_07872_),
    .Y(_02520_));
 sg13g2_nand2_1 _27161_ (.Y(_07873_),
    .A(_02785_),
    .B(_06806_));
 sg13g2_nand2_1 _27162_ (.Y(_07874_),
    .A(\cpu.qspi.r_mask[0] ),
    .B(_06809_));
 sg13g2_a21oi_1 _27163_ (.A1(_07873_),
    .A2(_07874_),
    .Y(_02521_),
    .B1(net565));
 sg13g2_nor4_1 _27164_ (.A(net975),
    .B(_07064_),
    .C(_04960_),
    .D(net110),
    .Y(_07875_));
 sg13g2_a21oi_1 _27165_ (.A1(\cpu.qspi.r_mask[1] ),
    .A2(_06822_),
    .Y(_07876_),
    .B1(_07875_));
 sg13g2_nand2_1 _27166_ (.Y(_02522_),
    .A(net685),
    .B(_07876_));
 sg13g2_nor2_1 _27167_ (.A(_07064_),
    .B(_06835_),
    .Y(_07877_));
 sg13g2_a21oi_1 _27168_ (.A1(\cpu.qspi.r_mask[2] ),
    .A2(_06835_),
    .Y(_07878_),
    .B1(_07877_));
 sg13g2_nor2_1 _27169_ (.A(net566),
    .B(_07878_),
    .Y(_02523_));
 sg13g2_nand2_1 _27170_ (.Y(_07879_),
    .A(\cpu.qspi.r_quad[0] ),
    .B(_06809_));
 sg13g2_nand2_1 _27171_ (.Y(_07880_),
    .A(net1035),
    .B(_06806_));
 sg13g2_nand3_1 _27172_ (.B(_07879_),
    .C(_07880_),
    .A(net650),
    .Y(_02524_));
 sg13g2_nor4_1 _27173_ (.A(net975),
    .B(_07060_),
    .C(_04960_),
    .D(net110),
    .Y(_07881_));
 sg13g2_a21oi_1 _27174_ (.A1(\cpu.qspi.r_quad[1] ),
    .A2(_06822_),
    .Y(_07882_),
    .B1(_07881_));
 sg13g2_nor2_1 _27175_ (.A(net566),
    .B(_07882_),
    .Y(_02525_));
 sg13g2_nand2_1 _27176_ (.Y(_07883_),
    .A(_07060_),
    .B(_06832_));
 sg13g2_o21ai_1 _27177_ (.B1(_07883_),
    .Y(_07884_),
    .A1(\cpu.qspi.r_quad[2] ),
    .A2(_06832_));
 sg13g2_nand2_1 _27178_ (.Y(_02526_),
    .A(net685),
    .B(_07884_));
 sg13g2_nor2_1 _27179_ (.A(_04903_),
    .B(net110),
    .Y(_07885_));
 sg13g2_nand2_1 _27180_ (.Y(_07886_),
    .A(_12807_),
    .B(_07885_));
 sg13g2_o21ai_1 _27181_ (.B1(_09967_),
    .Y(_07887_),
    .A1(_04903_),
    .A2(net110));
 sg13g2_nand3_1 _27182_ (.B(_07886_),
    .C(_07887_),
    .A(net650),
    .Y(_02539_));
 sg13g2_nand2_1 _27183_ (.Y(_07888_),
    .A(_12694_),
    .B(_07885_));
 sg13g2_o21ai_1 _27184_ (.B1(\cpu.qspi.r_rom_mode[1] ),
    .Y(_07889_),
    .A1(_04903_),
    .A2(net110));
 sg13g2_nand3_1 _27185_ (.B(_07888_),
    .C(_07889_),
    .A(net650),
    .Y(_02540_));
 sg13g2_nand2b_1 _27186_ (.Y(_07890_),
    .B(_12008_),
    .A_N(_06902_));
 sg13g2_nor4_1 _27187_ (.A(_12023_),
    .B(_09947_),
    .C(_09963_),
    .D(_09960_),
    .Y(_07891_));
 sg13g2_nand4_1 _27188_ (.B(_07855_),
    .C(_07890_),
    .A(_09937_),
    .Y(_07892_),
    .D(_07891_));
 sg13g2_buf_1 _27189_ (.A(_07892_),
    .X(_07893_));
 sg13g2_nor2b_1 _27190_ (.A(net3),
    .B_N(_07893_),
    .Y(_07894_));
 sg13g2_nor4_1 _27191_ (.A(_12008_),
    .B(_09948_),
    .C(_09938_),
    .D(net1119),
    .Y(_07895_));
 sg13g2_nor4_1 _27192_ (.A(_12006_),
    .B(_06870_),
    .C(_07893_),
    .D(_07895_),
    .Y(_07896_));
 sg13g2_nor3_1 _27193_ (.A(net707),
    .B(_07894_),
    .C(_07896_),
    .Y(_02541_));
 sg13g2_nor2b_1 _27194_ (.A(net6),
    .B_N(_07893_),
    .Y(_07897_));
 sg13g2_nand2b_1 _27195_ (.Y(_07898_),
    .B(_07895_),
    .A_N(_06870_));
 sg13g2_o21ai_1 _27196_ (.B1(_12007_),
    .Y(_07899_),
    .A1(_09982_),
    .A2(_07898_));
 sg13g2_nor2_1 _27197_ (.A(_07893_),
    .B(_07899_),
    .Y(_07900_));
 sg13g2_nor3_1 _27198_ (.A(net707),
    .B(_07897_),
    .C(_07900_),
    .Y(_02542_));
 sg13g2_nand2b_1 _27199_ (.Y(_07901_),
    .B(net758),
    .A_N(_09370_));
 sg13g2_nor3_1 _27200_ (.A(_09377_),
    .B(net1124),
    .C(_09429_),
    .Y(_07902_));
 sg13g2_a221oi_1 _27201_ (.B2(net1050),
    .C1(_07902_),
    .B1(_09276_),
    .A1(net1124),
    .Y(_07903_),
    .A2(_07901_));
 sg13g2_buf_1 _27202_ (.A(_07903_),
    .X(_07904_));
 sg13g2_nand3_1 _27203_ (.B(net1050),
    .C(_07904_),
    .A(_09395_),
    .Y(_07905_));
 sg13g2_o21ai_1 _27204_ (.B1(_07905_),
    .Y(_07906_),
    .A1(_09395_),
    .A2(_07904_));
 sg13g2_nand2_1 _27205_ (.Y(_02548_),
    .A(net685),
    .B(_07906_));
 sg13g2_nand2_1 _27206_ (.Y(_07907_),
    .A(_09395_),
    .B(_12031_));
 sg13g2_a21oi_1 _27207_ (.A1(_07904_),
    .A2(_07907_),
    .Y(_07908_),
    .B1(_09396_));
 sg13g2_inv_1 _27208_ (.Y(_07909_),
    .A(_09395_));
 sg13g2_and4_1 _27209_ (.A(_07909_),
    .B(_09396_),
    .C(_12031_),
    .D(_07904_),
    .X(_07910_));
 sg13g2_o21ai_1 _27210_ (.B1(net685),
    .Y(_02549_),
    .A1(_07908_),
    .A2(_07910_));
 sg13g2_nor2_1 _27211_ (.A(_09395_),
    .B(_09396_),
    .Y(_07911_));
 sg13g2_or2_1 _27212_ (.X(_07912_),
    .B(_07911_),
    .A(_00226_));
 sg13g2_a21oi_1 _27213_ (.A1(_07904_),
    .A2(_07912_),
    .Y(_07913_),
    .B1(\cpu.spi.r_bits[2] ));
 sg13g2_and4_1 _27214_ (.A(\cpu.spi.r_bits[2] ),
    .B(_12031_),
    .C(_07911_),
    .D(_07904_),
    .X(_07914_));
 sg13g2_o21ai_1 _27215_ (.B1(net685),
    .Y(_02550_),
    .A1(_07913_),
    .A2(_07914_));
 sg13g2_nor3_2 _27216_ (.A(net899),
    .B(_04890_),
    .C(_09370_),
    .Y(_07915_));
 sg13g2_and2_1 _27217_ (.A(net760),
    .B(_07915_),
    .X(_07916_));
 sg13g2_buf_1 _27218_ (.A(_07916_),
    .X(_07917_));
 sg13g2_nand2_1 _27219_ (.Y(_07918_),
    .A(net515),
    .B(_07917_));
 sg13g2_buf_2 _27220_ (.A(_07918_),
    .X(_07919_));
 sg13g2_nand2_1 _27221_ (.Y(_07920_),
    .A(\cpu.spi.r_clk_count[0][0] ),
    .B(_07919_));
 sg13g2_and2_1 _27222_ (.A(net515),
    .B(_07917_),
    .X(_07921_));
 sg13g2_buf_2 _27223_ (.A(_07921_),
    .X(_07922_));
 sg13g2_nand2_1 _27224_ (.Y(_07923_),
    .A(net919),
    .B(_07922_));
 sg13g2_a21oi_1 _27225_ (.A1(_07920_),
    .A2(_07923_),
    .Y(_02551_),
    .B1(net565));
 sg13g2_nand2_1 _27226_ (.Y(_07924_),
    .A(\cpu.spi.r_clk_count[0][1] ),
    .B(_07919_));
 sg13g2_nand2_1 _27227_ (.Y(_07925_),
    .A(net966),
    .B(_07922_));
 sg13g2_a21oi_1 _27228_ (.A1(_07924_),
    .A2(_07925_),
    .Y(_02552_),
    .B1(net565));
 sg13g2_nand2_1 _27229_ (.Y(_07926_),
    .A(\cpu.spi.r_clk_count[0][2] ),
    .B(_07919_));
 sg13g2_nand2_1 _27230_ (.Y(_07927_),
    .A(net920),
    .B(_07922_));
 sg13g2_a21oi_1 _27231_ (.A1(_07926_),
    .A2(_07927_),
    .Y(_02553_),
    .B1(net565));
 sg13g2_nand2_1 _27232_ (.Y(_07928_),
    .A(\cpu.spi.r_clk_count[0][3] ),
    .B(_07919_));
 sg13g2_nand2_1 _27233_ (.Y(_07929_),
    .A(net1038),
    .B(_07922_));
 sg13g2_a21oi_1 _27234_ (.A1(_07928_),
    .A2(_07929_),
    .Y(_02554_),
    .B1(net565));
 sg13g2_nand2_1 _27235_ (.Y(_07930_),
    .A(\cpu.spi.r_clk_count[0][4] ),
    .B(_07919_));
 sg13g2_nand2_1 _27236_ (.Y(_07931_),
    .A(net1037),
    .B(_07922_));
 sg13g2_buf_1 _27237_ (.A(_09452_),
    .X(_07932_));
 sg13g2_a21oi_1 _27238_ (.A1(_07930_),
    .A2(_07931_),
    .Y(_02555_),
    .B1(net564));
 sg13g2_nand2_1 _27239_ (.Y(_07933_),
    .A(\cpu.spi.r_clk_count[0][5] ),
    .B(_07919_));
 sg13g2_nand2_1 _27240_ (.Y(_07934_),
    .A(net1036),
    .B(_07922_));
 sg13g2_a21oi_1 _27241_ (.A1(_07933_),
    .A2(_07934_),
    .Y(_02556_),
    .B1(net564));
 sg13g2_nand2_1 _27242_ (.Y(_07935_),
    .A(\cpu.spi.r_clk_count[0][6] ),
    .B(_07919_));
 sg13g2_nand2_1 _27243_ (.Y(_07936_),
    .A(net1035),
    .B(_07922_));
 sg13g2_a21oi_1 _27244_ (.A1(_07935_),
    .A2(_07936_),
    .Y(_02557_),
    .B1(net564));
 sg13g2_nand2_1 _27245_ (.Y(_07937_),
    .A(\cpu.spi.r_clk_count[0][7] ),
    .B(_07919_));
 sg13g2_nand2_1 _27246_ (.Y(_07938_),
    .A(net985),
    .B(_07922_));
 sg13g2_a21oi_1 _27247_ (.A1(_07937_),
    .A2(_07938_),
    .Y(_02558_),
    .B1(net564));
 sg13g2_nand3_1 _27248_ (.B(net515),
    .C(_07915_),
    .A(net524),
    .Y(_07939_));
 sg13g2_buf_2 _27249_ (.A(_07939_),
    .X(_07940_));
 sg13g2_nand2_1 _27250_ (.Y(_07941_),
    .A(\cpu.spi.r_clk_count[1][0] ),
    .B(_07940_));
 sg13g2_and3_1 _27251_ (.X(_07942_),
    .A(net524),
    .B(net515),
    .C(_07915_));
 sg13g2_buf_2 _27252_ (.A(_07942_),
    .X(_07943_));
 sg13g2_nand2_1 _27253_ (.Y(_07944_),
    .A(net919),
    .B(_07943_));
 sg13g2_a21oi_1 _27254_ (.A1(_07941_),
    .A2(_07944_),
    .Y(_02559_),
    .B1(net564));
 sg13g2_nand2_1 _27255_ (.Y(_07945_),
    .A(\cpu.spi.r_clk_count[1][1] ),
    .B(_07940_));
 sg13g2_nand2_1 _27256_ (.Y(_07946_),
    .A(net1040),
    .B(_07943_));
 sg13g2_a21oi_1 _27257_ (.A1(_07945_),
    .A2(_07946_),
    .Y(_02560_),
    .B1(_07932_));
 sg13g2_nand2_1 _27258_ (.Y(_07947_),
    .A(\cpu.spi.r_clk_count[1][2] ),
    .B(_07940_));
 sg13g2_nand2_1 _27259_ (.Y(_07948_),
    .A(net920),
    .B(_07943_));
 sg13g2_a21oi_1 _27260_ (.A1(_07947_),
    .A2(_07948_),
    .Y(_02561_),
    .B1(_07932_));
 sg13g2_nand2_1 _27261_ (.Y(_07949_),
    .A(\cpu.spi.r_clk_count[1][3] ),
    .B(_07940_));
 sg13g2_nand2_1 _27262_ (.Y(_07950_),
    .A(net1038),
    .B(_07943_));
 sg13g2_a21oi_1 _27263_ (.A1(_07949_),
    .A2(_07950_),
    .Y(_02562_),
    .B1(net564));
 sg13g2_nand2_1 _27264_ (.Y(_07951_),
    .A(\cpu.spi.r_clk_count[1][4] ),
    .B(_07940_));
 sg13g2_nand2_1 _27265_ (.Y(_07952_),
    .A(net1037),
    .B(_07943_));
 sg13g2_a21oi_1 _27266_ (.A1(_07951_),
    .A2(_07952_),
    .Y(_02563_),
    .B1(net564));
 sg13g2_nand2_1 _27267_ (.Y(_07953_),
    .A(\cpu.spi.r_clk_count[1][5] ),
    .B(_07940_));
 sg13g2_nand2_1 _27268_ (.Y(_07954_),
    .A(net1036),
    .B(_07943_));
 sg13g2_a21oi_1 _27269_ (.A1(_07953_),
    .A2(_07954_),
    .Y(_02564_),
    .B1(net564));
 sg13g2_nand2_1 _27270_ (.Y(_07955_),
    .A(\cpu.spi.r_clk_count[1][6] ),
    .B(_07940_));
 sg13g2_nand2_1 _27271_ (.Y(_07956_),
    .A(net1035),
    .B(_07943_));
 sg13g2_buf_1 _27272_ (.A(_09452_),
    .X(_07957_));
 sg13g2_a21oi_1 _27273_ (.A1(_07955_),
    .A2(_07956_),
    .Y(_02565_),
    .B1(net563));
 sg13g2_nand2_1 _27274_ (.Y(_07958_),
    .A(\cpu.spi.r_clk_count[1][7] ),
    .B(_07940_));
 sg13g2_nand2_1 _27275_ (.Y(_07959_),
    .A(net985),
    .B(_07943_));
 sg13g2_a21oi_1 _27276_ (.A1(_07958_),
    .A2(_07959_),
    .Y(_02566_),
    .B1(net563));
 sg13g2_nand2_1 _27277_ (.Y(_07960_),
    .A(_12058_),
    .B(net760));
 sg13g2_nor3_1 _27278_ (.A(_04890_),
    .B(_09370_),
    .C(_07960_),
    .Y(_07961_));
 sg13g2_buf_1 _27279_ (.A(_07961_),
    .X(_07962_));
 sg13g2_nand2_1 _27280_ (.Y(_07963_),
    .A(net515),
    .B(_07962_));
 sg13g2_buf_2 _27281_ (.A(_07963_),
    .X(_07964_));
 sg13g2_nand2_1 _27282_ (.Y(_07965_),
    .A(_04916_),
    .B(_07964_));
 sg13g2_and2_1 _27283_ (.A(net515),
    .B(_07962_),
    .X(_07966_));
 sg13g2_buf_2 _27284_ (.A(_07966_),
    .X(_07967_));
 sg13g2_nand2_1 _27285_ (.Y(_07968_),
    .A(net919),
    .B(_07967_));
 sg13g2_a21oi_1 _27286_ (.A1(_07965_),
    .A2(_07968_),
    .Y(_02567_),
    .B1(net563));
 sg13g2_nand2_1 _27287_ (.Y(_07969_),
    .A(_05326_),
    .B(_07964_));
 sg13g2_nand2_1 _27288_ (.Y(_07970_),
    .A(net1040),
    .B(_07967_));
 sg13g2_a21oi_1 _27289_ (.A1(_07969_),
    .A2(_07970_),
    .Y(_02568_),
    .B1(net563));
 sg13g2_nand2_1 _27290_ (.Y(_07971_),
    .A(_05394_),
    .B(_07964_));
 sg13g2_nand2_1 _27291_ (.Y(_07972_),
    .A(net920),
    .B(_07967_));
 sg13g2_a21oi_1 _27292_ (.A1(_07971_),
    .A2(_07972_),
    .Y(_02569_),
    .B1(_07957_));
 sg13g2_nand2_1 _27293_ (.Y(_07973_),
    .A(_05479_),
    .B(_07964_));
 sg13g2_nand2_1 _27294_ (.Y(_07974_),
    .A(net1038),
    .B(_07967_));
 sg13g2_a21oi_1 _27295_ (.A1(_07973_),
    .A2(_07974_),
    .Y(_02570_),
    .B1(net563));
 sg13g2_nand2_1 _27296_ (.Y(_07975_),
    .A(_05570_),
    .B(_07964_));
 sg13g2_nand2_1 _27297_ (.Y(_07976_),
    .A(net1037),
    .B(_07967_));
 sg13g2_a21oi_1 _27298_ (.A1(_07975_),
    .A2(_07976_),
    .Y(_02571_),
    .B1(net563));
 sg13g2_nand2_1 _27299_ (.Y(_07977_),
    .A(_05610_),
    .B(_07964_));
 sg13g2_nand2_1 _27300_ (.Y(_07978_),
    .A(net1036),
    .B(_07967_));
 sg13g2_a21oi_1 _27301_ (.A1(_07977_),
    .A2(_07978_),
    .Y(_02572_),
    .B1(net563));
 sg13g2_nand2_1 _27302_ (.Y(_07979_),
    .A(_05683_),
    .B(_07964_));
 sg13g2_nand2_1 _27303_ (.Y(_07980_),
    .A(net1035),
    .B(_07967_));
 sg13g2_a21oi_1 _27304_ (.A1(_07979_),
    .A2(_07980_),
    .Y(_02573_),
    .B1(net563));
 sg13g2_nand2_1 _27305_ (.Y(_07981_),
    .A(_05022_),
    .B(_07964_));
 sg13g2_nand2_1 _27306_ (.Y(_07982_),
    .A(net985),
    .B(_07967_));
 sg13g2_a21oi_1 _27307_ (.A1(_07981_),
    .A2(_07982_),
    .Y(_02574_),
    .B1(_07957_));
 sg13g2_nand2_1 _27308_ (.Y(_07983_),
    .A(_09377_),
    .B(_09383_));
 sg13g2_o21ai_1 _27309_ (.B1(_09374_),
    .Y(_07984_),
    .A1(_09393_),
    .A2(_09364_));
 sg13g2_nor2_1 _27310_ (.A(_09375_),
    .B(\cpu.spi.r_state[5] ),
    .Y(_07985_));
 sg13g2_and2_1 _27311_ (.A(_12027_),
    .B(_07985_),
    .X(_07986_));
 sg13g2_buf_1 _27312_ (.A(_07986_),
    .X(_07987_));
 sg13g2_nand2_1 _27313_ (.Y(_07988_),
    .A(_07030_),
    .B(_07987_));
 sg13g2_buf_2 _27314_ (.A(_07988_),
    .X(_07989_));
 sg13g2_inv_1 _27315_ (.Y(_07990_),
    .A(_07989_));
 sg13g2_nand2_1 _27316_ (.Y(_07991_),
    .A(_12026_),
    .B(_07990_));
 sg13g2_nand3b_1 _27317_ (.B(_09372_),
    .C(_09275_),
    .Y(_07992_),
    .A_N(net964));
 sg13g2_nand4_1 _27318_ (.B(_07984_),
    .C(_07991_),
    .A(_07983_),
    .Y(_07993_),
    .D(_07992_));
 sg13g2_buf_1 _27319_ (.A(_07993_),
    .X(_07994_));
 sg13g2_buf_1 _27320_ (.A(_07994_),
    .X(_07995_));
 sg13g2_nand2b_1 _27321_ (.Y(_07996_),
    .B(net609),
    .A_N(\cpu.spi.r_clk_count[0][0] ));
 sg13g2_o21ai_1 _27322_ (.B1(_07996_),
    .Y(_07997_),
    .A1(net610),
    .A2(_04916_));
 sg13g2_mux2_1 _27323_ (.A0(\cpu.spi.r_clk_count[0][0] ),
    .A1(\cpu.spi.r_clk_count[1][0] ),
    .S(net609),
    .X(_07998_));
 sg13g2_nor2_1 _27324_ (.A(net664),
    .B(_07998_),
    .Y(_07999_));
 sg13g2_a21oi_1 _27325_ (.A1(net659),
    .A2(_07997_),
    .Y(_08000_),
    .B1(_07999_));
 sg13g2_nor2_1 _27326_ (.A(_07989_),
    .B(_08000_),
    .Y(_08001_));
 sg13g2_buf_1 _27327_ (.A(_07987_),
    .X(_08002_));
 sg13g2_buf_1 _27328_ (.A(net1012),
    .X(_08003_));
 sg13g2_nand2_1 _27329_ (.Y(_08004_),
    .A(net1014),
    .B(_00313_));
 sg13g2_o21ai_1 _27330_ (.B1(_08004_),
    .Y(_08005_),
    .A1(net828),
    .A2(_04911_));
 sg13g2_nor2_1 _27331_ (.A(net1012),
    .B(_04916_),
    .Y(_08006_));
 sg13g2_a21oi_1 _27332_ (.A1(_12038_),
    .A2(_00314_),
    .Y(_08007_),
    .B1(_08006_));
 sg13g2_nand2_1 _27333_ (.Y(_08008_),
    .A(net1013),
    .B(_08007_));
 sg13g2_o21ai_1 _27334_ (.B1(_08008_),
    .Y(_08009_),
    .A1(net1013),
    .A2(_08005_));
 sg13g2_nand2_1 _27335_ (.Y(_08010_),
    .A(_09433_),
    .B(_08009_));
 sg13g2_o21ai_1 _27336_ (.B1(_08010_),
    .Y(_08011_),
    .A1(_09267_),
    .A2(net90));
 sg13g2_nor2_1 _27337_ (.A(net447),
    .B(_08009_),
    .Y(_08012_));
 sg13g2_nor3_1 _27338_ (.A(_09267_),
    .B(net642),
    .C(_08012_),
    .Y(_08013_));
 sg13g2_a221oi_1 _27339_ (.B2(net963),
    .C1(_08013_),
    .B1(_08011_),
    .A1(net964),
    .Y(_08014_),
    .A2(net642));
 sg13g2_nor3_1 _27340_ (.A(_07994_),
    .B(_08001_),
    .C(_08014_),
    .Y(_08015_));
 sg13g2_a21oi_1 _27341_ (.A1(_09267_),
    .A2(net31),
    .Y(_08016_),
    .B1(_08015_));
 sg13g2_nor2_1 _27342_ (.A(net566),
    .B(_08016_),
    .Y(_02575_));
 sg13g2_mux2_1 _27343_ (.A0(\cpu.spi.r_clk_count[0][1] ),
    .A1(\cpu.spi.r_clk_count[1][1] ),
    .S(_12059_),
    .X(_08017_));
 sg13g2_nand2_1 _27344_ (.Y(_08018_),
    .A(net760),
    .B(_05326_));
 sg13g2_nand2_1 _27345_ (.Y(_08019_),
    .A(net665),
    .B(\cpu.spi.r_clk_count[0][1] ));
 sg13g2_nand3_1 _27346_ (.B(_08018_),
    .C(_08019_),
    .A(net761),
    .Y(_08020_));
 sg13g2_o21ai_1 _27347_ (.B1(_08020_),
    .Y(_08021_),
    .A1(net761),
    .A2(_08017_));
 sg13g2_nand2_1 _27348_ (.Y(_08022_),
    .A(_07990_),
    .B(_08021_));
 sg13g2_nand3_1 _27349_ (.B(_09374_),
    .C(_08022_),
    .A(_09267_),
    .Y(_08023_));
 sg13g2_nand2b_1 _27350_ (.Y(_08024_),
    .B(_08023_),
    .A_N(_07994_));
 sg13g2_nor2_1 _27351_ (.A(net828),
    .B(_05326_),
    .Y(_08025_));
 sg13g2_a21oi_1 _27352_ (.A1(net900),
    .A2(_00095_),
    .Y(_08026_),
    .B1(_08025_));
 sg13g2_nand2_1 _27353_ (.Y(_08027_),
    .A(net1014),
    .B(_00094_));
 sg13g2_o21ai_1 _27354_ (.B1(_08027_),
    .Y(_08028_),
    .A1(net828),
    .A2(_05328_));
 sg13g2_nor2_1 _27355_ (.A(_12040_),
    .B(_08028_),
    .Y(_08029_));
 sg13g2_a21oi_1 _27356_ (.A1(net1015),
    .A2(_08026_),
    .Y(_08030_),
    .B1(_08029_));
 sg13g2_nor2_1 _27357_ (.A(net107),
    .B(_09269_),
    .Y(_08031_));
 sg13g2_a21oi_1 _27358_ (.A1(net90),
    .A2(_08030_),
    .Y(_08032_),
    .B1(_08031_));
 sg13g2_nand2_1 _27359_ (.Y(_08033_),
    .A(_09267_),
    .B(_09268_));
 sg13g2_or2_1 _27360_ (.X(_08034_),
    .B(_09268_),
    .A(_09267_));
 sg13g2_a221oi_1 _27361_ (.B2(_08034_),
    .C1(_08002_),
    .B1(_08033_),
    .A1(net446),
    .Y(_08035_),
    .A2(_08030_));
 sg13g2_a221oi_1 _27362_ (.B2(net963),
    .C1(_08035_),
    .B1(_08032_),
    .A1(net964),
    .Y(_08036_),
    .A2(net642));
 sg13g2_nor2_1 _27363_ (.A(_07994_),
    .B(_08036_),
    .Y(_08037_));
 sg13g2_a22oi_1 _27364_ (.Y(_08038_),
    .B1(_08037_),
    .B2(_08022_),
    .A2(_08024_),
    .A1(_09268_));
 sg13g2_nor2_1 _27365_ (.A(net566),
    .B(_08038_),
    .Y(_02576_));
 sg13g2_nand2_1 _27366_ (.Y(_08039_),
    .A(\cpu.spi.r_count[2] ),
    .B(net31));
 sg13g2_nand2b_1 _27367_ (.Y(_08040_),
    .B(net610),
    .A_N(\cpu.spi.r_clk_count[0][2] ));
 sg13g2_o21ai_1 _27368_ (.B1(_08040_),
    .Y(_08041_),
    .A1(net610),
    .A2(_05394_));
 sg13g2_mux2_1 _27369_ (.A0(\cpu.spi.r_clk_count[0][2] ),
    .A1(\cpu.spi.r_clk_count[1][2] ),
    .S(net609),
    .X(_08042_));
 sg13g2_nor2_1 _27370_ (.A(net664),
    .B(_08042_),
    .Y(_08043_));
 sg13g2_a21oi_1 _27371_ (.A1(net659),
    .A2(_08041_),
    .Y(_08044_),
    .B1(_08043_));
 sg13g2_nor2_1 _27372_ (.A(_07989_),
    .B(_08044_),
    .Y(_08045_));
 sg13g2_nor2_1 _27373_ (.A(net900),
    .B(_05394_),
    .Y(_08046_));
 sg13g2_a21oi_1 _27374_ (.A1(net900),
    .A2(_00105_),
    .Y(_08047_),
    .B1(_08046_));
 sg13g2_nand2_1 _27375_ (.Y(_08048_),
    .A(net1014),
    .B(_00104_));
 sg13g2_o21ai_1 _27376_ (.B1(_08048_),
    .Y(_08049_),
    .A1(_08003_),
    .A2(_05393_));
 sg13g2_nor2_1 _27377_ (.A(net1015),
    .B(_08049_),
    .Y(_08050_));
 sg13g2_a21oi_1 _27378_ (.A1(net1015),
    .A2(_08047_),
    .Y(_08051_),
    .B1(_08050_));
 sg13g2_xnor2_1 _27379_ (.Y(_08052_),
    .A(\cpu.spi.r_count[2] ),
    .B(_08034_));
 sg13g2_nor2_1 _27380_ (.A(net107),
    .B(_08052_),
    .Y(_08053_));
 sg13g2_a21oi_1 _27381_ (.A1(net90),
    .A2(_08051_),
    .Y(_08054_),
    .B1(_08053_));
 sg13g2_inv_1 _27382_ (.Y(_08055_),
    .A(_07987_));
 sg13g2_nand2_1 _27383_ (.Y(_08056_),
    .A(_08055_),
    .B(_08052_));
 sg13g2_a21oi_1 _27384_ (.A1(net446),
    .A2(_08051_),
    .Y(_08057_),
    .B1(_08056_));
 sg13g2_a221oi_1 _27385_ (.B2(_07033_),
    .C1(_08057_),
    .B1(_08054_),
    .A1(net964),
    .Y(_08058_),
    .A2(_08002_));
 sg13g2_or3_1 _27386_ (.A(net31),
    .B(_08045_),
    .C(_08058_),
    .X(_08059_));
 sg13g2_buf_1 _27387_ (.A(_09452_),
    .X(_08060_));
 sg13g2_a21oi_1 _27388_ (.A1(_08039_),
    .A2(_08059_),
    .Y(_02577_),
    .B1(net562));
 sg13g2_nand2b_1 _27389_ (.Y(_08061_),
    .B(net609),
    .A_N(\cpu.spi.r_clk_count[0][3] ));
 sg13g2_o21ai_1 _27390_ (.B1(_08061_),
    .Y(_08062_),
    .A1(net610),
    .A2(_05479_));
 sg13g2_mux2_1 _27391_ (.A0(\cpu.spi.r_clk_count[0][3] ),
    .A1(\cpu.spi.r_clk_count[1][3] ),
    .S(net665),
    .X(_08063_));
 sg13g2_nor2_1 _27392_ (.A(net664),
    .B(_08063_),
    .Y(_08064_));
 sg13g2_a21oi_1 _27393_ (.A1(net659),
    .A2(_08062_),
    .Y(_08065_),
    .B1(_08064_));
 sg13g2_nor2_1 _27394_ (.A(_07989_),
    .B(_08065_),
    .Y(_08066_));
 sg13g2_xor2_1 _27395_ (.B(_09270_),
    .A(_09266_),
    .X(_08067_));
 sg13g2_nand2_1 _27396_ (.Y(_08068_),
    .A(net1012),
    .B(_00114_));
 sg13g2_o21ai_1 _27397_ (.B1(_08068_),
    .Y(_08069_),
    .A1(net828),
    .A2(_05478_));
 sg13g2_nor2_1 _27398_ (.A(net1012),
    .B(_05479_),
    .Y(_08070_));
 sg13g2_a21oi_1 _27399_ (.A1(net1014),
    .A2(_00115_),
    .Y(_08071_),
    .B1(_08070_));
 sg13g2_nand2_1 _27400_ (.Y(_08072_),
    .A(net1013),
    .B(_08071_));
 sg13g2_o21ai_1 _27401_ (.B1(_08072_),
    .Y(_08073_),
    .A1(net1013),
    .A2(_08069_));
 sg13g2_nand2_1 _27402_ (.Y(_08074_),
    .A(net107),
    .B(_08073_));
 sg13g2_o21ai_1 _27403_ (.B1(_08074_),
    .Y(_08075_),
    .A1(net90),
    .A2(_08067_));
 sg13g2_nor2_1 _27404_ (.A(net497),
    .B(_08073_),
    .Y(_08076_));
 sg13g2_nor3_1 _27405_ (.A(net642),
    .B(_08067_),
    .C(_08076_),
    .Y(_08077_));
 sg13g2_a221oi_1 _27406_ (.B2(net963),
    .C1(_08077_),
    .B1(_08075_),
    .A1(net964),
    .Y(_08078_),
    .A2(net642));
 sg13g2_nor3_1 _27407_ (.A(_07994_),
    .B(_08066_),
    .C(_08078_),
    .Y(_08079_));
 sg13g2_a21oi_1 _27408_ (.A1(_09266_),
    .A2(net31),
    .Y(_08080_),
    .B1(_08079_));
 sg13g2_nor2_1 _27409_ (.A(net566),
    .B(_08080_),
    .Y(_02578_));
 sg13g2_nand2b_1 _27410_ (.Y(_08081_),
    .B(net609),
    .A_N(\cpu.spi.r_clk_count[0][4] ));
 sg13g2_o21ai_1 _27411_ (.B1(_08081_),
    .Y(_08082_),
    .A1(net610),
    .A2(_05570_));
 sg13g2_mux2_1 _27412_ (.A0(\cpu.spi.r_clk_count[0][4] ),
    .A1(\cpu.spi.r_clk_count[1][4] ),
    .S(net665),
    .X(_08083_));
 sg13g2_nor2_1 _27413_ (.A(net664),
    .B(_08083_),
    .Y(_08084_));
 sg13g2_a21oi_1 _27414_ (.A1(net659),
    .A2(_08082_),
    .Y(_08085_),
    .B1(_08084_));
 sg13g2_nor2_1 _27415_ (.A(_07989_),
    .B(_08085_),
    .Y(_08086_));
 sg13g2_nor2_1 _27416_ (.A(_09266_),
    .B(_09270_),
    .Y(_08087_));
 sg13g2_xnor2_1 _27417_ (.Y(_08088_),
    .A(\cpu.spi.r_count[4] ),
    .B(_08087_));
 sg13g2_nand2_1 _27418_ (.Y(_08089_),
    .A(net1012),
    .B(_00125_));
 sg13g2_o21ai_1 _27419_ (.B1(_08089_),
    .Y(_08090_),
    .A1(net828),
    .A2(_05569_));
 sg13g2_nor2_1 _27420_ (.A(net1012),
    .B(_05570_),
    .Y(_08091_));
 sg13g2_a21oi_1 _27421_ (.A1(net1014),
    .A2(_00126_),
    .Y(_08092_),
    .B1(_08091_));
 sg13g2_nand2_1 _27422_ (.Y(_08093_),
    .A(net1013),
    .B(_08092_));
 sg13g2_o21ai_1 _27423_ (.B1(_08093_),
    .Y(_08094_),
    .A1(net1013),
    .A2(_08090_));
 sg13g2_nand2_1 _27424_ (.Y(_08095_),
    .A(net107),
    .B(_08094_));
 sg13g2_o21ai_1 _27425_ (.B1(_08095_),
    .Y(_08096_),
    .A1(net90),
    .A2(_08088_));
 sg13g2_nor2_1 _27426_ (.A(net497),
    .B(_08094_),
    .Y(_08097_));
 sg13g2_nor3_1 _27427_ (.A(_07987_),
    .B(_08088_),
    .C(_08097_),
    .Y(_08098_));
 sg13g2_a221oi_1 _27428_ (.B2(net963),
    .C1(_08098_),
    .B1(_08096_),
    .A1(net964),
    .Y(_08099_),
    .A2(net642));
 sg13g2_nor3_1 _27429_ (.A(_07994_),
    .B(_08086_),
    .C(_08099_),
    .Y(_08100_));
 sg13g2_a21oi_1 _27430_ (.A1(\cpu.spi.r_count[4] ),
    .A2(_07995_),
    .Y(_08101_),
    .B1(_08100_));
 sg13g2_nor2_1 _27431_ (.A(net566),
    .B(_08101_),
    .Y(_02579_));
 sg13g2_nand2b_1 _27432_ (.Y(_08102_),
    .B(net609),
    .A_N(\cpu.spi.r_clk_count[0][5] ));
 sg13g2_o21ai_1 _27433_ (.B1(_08102_),
    .Y(_08103_),
    .A1(net610),
    .A2(_05610_));
 sg13g2_mux2_1 _27434_ (.A0(\cpu.spi.r_clk_count[0][5] ),
    .A1(\cpu.spi.r_clk_count[1][5] ),
    .S(net665),
    .X(_08104_));
 sg13g2_nor2_1 _27435_ (.A(net761),
    .B(_08104_),
    .Y(_08105_));
 sg13g2_a21oi_1 _27436_ (.A1(net659),
    .A2(_08103_),
    .Y(_08106_),
    .B1(_08105_));
 sg13g2_nor2_1 _27437_ (.A(_07989_),
    .B(_08106_),
    .Y(_08107_));
 sg13g2_xnor2_1 _27438_ (.Y(_08108_),
    .A(\cpu.spi.r_count[5] ),
    .B(_09271_));
 sg13g2_mux2_1 _27439_ (.A0(_00133_),
    .A1(_00132_),
    .S(net1014),
    .X(_08109_));
 sg13g2_nor2_1 _27440_ (.A(net1012),
    .B(_05610_),
    .Y(_08110_));
 sg13g2_a21oi_1 _27441_ (.A1(net1014),
    .A2(_00133_),
    .Y(_08111_),
    .B1(_08110_));
 sg13g2_nand2_1 _27442_ (.Y(_08112_),
    .A(net1013),
    .B(_08111_));
 sg13g2_o21ai_1 _27443_ (.B1(_08112_),
    .Y(_08113_),
    .A1(net1013),
    .A2(_08109_));
 sg13g2_nand2_1 _27444_ (.Y(_08114_),
    .A(net107),
    .B(_08113_));
 sg13g2_o21ai_1 _27445_ (.B1(_08114_),
    .Y(_08115_),
    .A1(net90),
    .A2(_08108_));
 sg13g2_nor2_1 _27446_ (.A(net497),
    .B(_08113_),
    .Y(_08116_));
 sg13g2_nor3_1 _27447_ (.A(_07987_),
    .B(_08116_),
    .C(_08108_),
    .Y(_08117_));
 sg13g2_a221oi_1 _27448_ (.B2(net963),
    .C1(_08117_),
    .B1(_08115_),
    .A1(net964),
    .Y(_08118_),
    .A2(net642));
 sg13g2_nor3_1 _27449_ (.A(_07994_),
    .B(_08107_),
    .C(_08118_),
    .Y(_08119_));
 sg13g2_a21oi_1 _27450_ (.A1(\cpu.spi.r_count[5] ),
    .A2(_07995_),
    .Y(_08120_),
    .B1(_08119_));
 sg13g2_nor2_1 _27451_ (.A(net566),
    .B(_08120_),
    .Y(_02580_));
 sg13g2_nand2_1 _27452_ (.Y(_08121_),
    .A(\cpu.spi.r_count[6] ),
    .B(net31));
 sg13g2_nand2b_1 _27453_ (.Y(_08122_),
    .B(net609),
    .A_N(\cpu.spi.r_clk_count[0][6] ));
 sg13g2_o21ai_1 _27454_ (.B1(_08122_),
    .Y(_08123_),
    .A1(net610),
    .A2(_05683_));
 sg13g2_mux2_1 _27455_ (.A0(\cpu.spi.r_clk_count[0][6] ),
    .A1(\cpu.spi.r_clk_count[1][6] ),
    .S(net609),
    .X(_08124_));
 sg13g2_nor2_1 _27456_ (.A(net664),
    .B(_08124_),
    .Y(_08125_));
 sg13g2_a21oi_1 _27457_ (.A1(net659),
    .A2(_08123_),
    .Y(_08126_),
    .B1(_08125_));
 sg13g2_nor2_1 _27458_ (.A(_07989_),
    .B(_08126_),
    .Y(_08127_));
 sg13g2_nor2_1 _27459_ (.A(net828),
    .B(_05683_),
    .Y(_08128_));
 sg13g2_a21oi_1 _27460_ (.A1(net900),
    .A2(_00145_),
    .Y(_08129_),
    .B1(_08128_));
 sg13g2_mux2_1 _27461_ (.A0(_00145_),
    .A1(_00144_),
    .S(net828),
    .X(_08130_));
 sg13g2_nor2_1 _27462_ (.A(net1015),
    .B(_08130_),
    .Y(_08131_));
 sg13g2_a21oi_1 _27463_ (.A1(net1015),
    .A2(_08129_),
    .Y(_08132_),
    .B1(_08131_));
 sg13g2_xor2_1 _27464_ (.B(_09272_),
    .A(\cpu.spi.r_count[6] ),
    .X(_08133_));
 sg13g2_nor2_1 _27465_ (.A(net107),
    .B(_08133_),
    .Y(_08134_));
 sg13g2_a21oi_1 _27466_ (.A1(net90),
    .A2(_08132_),
    .Y(_08135_),
    .B1(_08134_));
 sg13g2_nand2_1 _27467_ (.Y(_08136_),
    .A(_08055_),
    .B(_08133_));
 sg13g2_a21oi_1 _27468_ (.A1(net446),
    .A2(_08132_),
    .Y(_08137_),
    .B1(_08136_));
 sg13g2_a221oi_1 _27469_ (.B2(net963),
    .C1(_08137_),
    .B1(_08135_),
    .A1(net964),
    .Y(_08138_),
    .A2(net642));
 sg13g2_or3_1 _27470_ (.A(net31),
    .B(_08127_),
    .C(_08138_),
    .X(_08139_));
 sg13g2_a21oi_1 _27471_ (.A1(_08121_),
    .A2(_08139_),
    .Y(_02581_),
    .B1(net562));
 sg13g2_nor2_1 _27472_ (.A(net828),
    .B(_05022_),
    .Y(_08140_));
 sg13g2_a21oi_1 _27473_ (.A1(net900),
    .A2(_00157_),
    .Y(_08141_),
    .B1(_08140_));
 sg13g2_mux2_1 _27474_ (.A0(_00157_),
    .A1(_00156_),
    .S(net1014),
    .X(_08142_));
 sg13g2_nor2_1 _27475_ (.A(net1015),
    .B(_08142_),
    .Y(_08143_));
 sg13g2_a21oi_1 _27476_ (.A1(net1015),
    .A2(_08141_),
    .Y(_08144_),
    .B1(_08143_));
 sg13g2_nand2_1 _27477_ (.Y(_08145_),
    .A(net90),
    .B(_08144_));
 sg13g2_nand2b_1 _27478_ (.Y(_08146_),
    .B(_09265_),
    .A_N(_09273_));
 sg13g2_nand3_1 _27479_ (.B(net447),
    .C(_08146_),
    .A(_07901_),
    .Y(_08147_));
 sg13g2_nand4_1 _27480_ (.B(_07989_),
    .C(_08145_),
    .A(net963),
    .Y(_08148_),
    .D(_08147_));
 sg13g2_and2_1 _27481_ (.A(net665),
    .B(\cpu.spi.r_clk_count[1][7] ),
    .X(_08149_));
 sg13g2_a21oi_1 _27482_ (.A1(net760),
    .A2(\cpu.spi.r_clk_count[0][7] ),
    .Y(_08150_),
    .B1(_08149_));
 sg13g2_mux2_1 _27483_ (.A0(_05022_),
    .A1(\cpu.spi.r_clk_count[0][7] ),
    .S(net665),
    .X(_08151_));
 sg13g2_nand2_1 _27484_ (.Y(_08152_),
    .A(net761),
    .B(_08151_));
 sg13g2_o21ai_1 _27485_ (.B1(_08152_),
    .Y(_08153_),
    .A1(net664),
    .A2(_08150_));
 sg13g2_o21ai_1 _27486_ (.B1(_08146_),
    .Y(_08154_),
    .A1(net447),
    .A2(_08144_));
 sg13g2_a22oi_1 _27487_ (.Y(_08155_),
    .B1(_08154_),
    .B2(_08055_),
    .A2(_08153_),
    .A1(_07990_));
 sg13g2_a21oi_1 _27488_ (.A1(_08148_),
    .A2(_08155_),
    .Y(_08156_),
    .B1(net31));
 sg13g2_a21oi_1 _27489_ (.A1(_09265_),
    .A2(net31),
    .Y(_08157_),
    .B1(_08156_));
 sg13g2_nor2_1 _27490_ (.A(_09453_),
    .B(_08157_),
    .Y(_02582_));
 sg13g2_buf_1 _27491_ (.A(\cpu.gpio.genblk1[3].srcs_o[6] ),
    .X(_08158_));
 sg13g2_inv_1 _27492_ (.Y(_08159_),
    .A(net1078));
 sg13g2_nor2_1 _27493_ (.A(_09433_),
    .B(_09391_),
    .Y(_08160_));
 sg13g2_inv_1 _27494_ (.Y(_08161_),
    .A(_09375_));
 sg13g2_nand2_1 _27495_ (.Y(_08162_),
    .A(_08161_),
    .B(_09366_));
 sg13g2_nand2_1 _27496_ (.Y(_08163_),
    .A(net446),
    .B(_08162_));
 sg13g2_nor3_1 _27497_ (.A(_09436_),
    .B(_09393_),
    .C(_08162_),
    .Y(_08164_));
 sg13g2_a21oi_1 _27498_ (.A1(_12033_),
    .A2(_08003_),
    .Y(_08165_),
    .B1(_09275_));
 sg13g2_nor3_1 _27499_ (.A(_00278_),
    .B(_08164_),
    .C(_08165_),
    .Y(_08166_));
 sg13g2_a21oi_1 _27500_ (.A1(_00278_),
    .A2(_08163_),
    .Y(_08167_),
    .B1(_08166_));
 sg13g2_o21ai_1 _27501_ (.B1(_08167_),
    .Y(_08168_),
    .A1(_07031_),
    .A2(_08160_));
 sg13g2_nor3_1 _27502_ (.A(_12034_),
    .B(net900),
    .C(_08168_),
    .Y(_08169_));
 sg13g2_inv_1 _27503_ (.Y(_08170_),
    .A(_08168_));
 sg13g2_a21oi_1 _27504_ (.A1(_08162_),
    .A2(_08170_),
    .Y(_08171_),
    .B1(net804));
 sg13g2_o21ai_1 _27505_ (.B1(_08171_),
    .Y(_02583_),
    .A1(_08159_),
    .A2(_08169_));
 sg13g2_buf_1 _27506_ (.A(\cpu.gpio.genblk1[3].srcs_o[7] ),
    .X(_08172_));
 sg13g2_nand3_1 _27507_ (.B(_12051_),
    .C(_08170_),
    .A(_12048_),
    .Y(_08173_));
 sg13g2_nand2_1 _27508_ (.Y(_08174_),
    .A(net1077),
    .B(_08173_));
 sg13g2_nand2_1 _27509_ (.Y(_02584_),
    .A(_08171_),
    .B(_08174_));
 sg13g2_buf_1 _27510_ (.A(\cpu.gpio.genblk1[3].srcs_o[8] ),
    .X(_08175_));
 sg13g2_inv_1 _27511_ (.Y(_08176_),
    .A(net1076));
 sg13g2_nor3_1 _27512_ (.A(_12048_),
    .B(_12051_),
    .C(_08168_),
    .Y(_08177_));
 sg13g2_o21ai_1 _27513_ (.B1(_08171_),
    .Y(_02585_),
    .A1(_08176_),
    .A2(_08177_));
 sg13g2_a21o_1 _27514_ (.A2(_09427_),
    .A1(_09429_),
    .B1(_07902_),
    .X(_08178_));
 sg13g2_buf_1 _27515_ (.A(_08178_),
    .X(_08179_));
 sg13g2_or2_1 _27516_ (.X(_08180_),
    .B(_09364_),
    .A(_07030_));
 sg13g2_o21ai_1 _27517_ (.B1(_07983_),
    .Y(_08181_),
    .A1(net107),
    .A2(_08180_));
 sg13g2_or3_1 _27518_ (.A(_09437_),
    .B(_08179_),
    .C(_08181_),
    .X(_08182_));
 sg13g2_o21ai_1 _27519_ (.B1(_09322_),
    .Y(_08183_),
    .A1(_08179_),
    .A2(_08181_));
 sg13g2_a21oi_1 _27520_ (.A1(_08182_),
    .A2(_08183_),
    .Y(_02594_),
    .B1(net562));
 sg13g2_nand2_2 _27521_ (.Y(_08184_),
    .A(net632),
    .B(_07917_));
 sg13g2_mux2_1 _27522_ (.A0(net1041),
    .A1(\cpu.spi.r_mode[0][0] ),
    .S(_08184_),
    .X(_08185_));
 sg13g2_and2_1 _27523_ (.A(net667),
    .B(_08185_),
    .X(_02595_));
 sg13g2_mux2_1 _27524_ (.A0(net1040),
    .A1(_12049_),
    .S(_08184_),
    .X(_08186_));
 sg13g2_and2_1 _27525_ (.A(net667),
    .B(_08186_),
    .X(_02596_));
 sg13g2_nand3_1 _27526_ (.B(net632),
    .C(_07915_),
    .A(_12067_),
    .Y(_08187_));
 sg13g2_buf_1 _27527_ (.A(_08187_),
    .X(_08188_));
 sg13g2_mux2_1 _27528_ (.A0(net1041),
    .A1(\cpu.spi.r_mode[1][0] ),
    .S(_08188_),
    .X(_08189_));
 sg13g2_and2_1 _27529_ (.A(net667),
    .B(_08189_),
    .X(_02597_));
 sg13g2_mux2_1 _27530_ (.A0(net1040),
    .A1(_12050_),
    .S(_08188_),
    .X(_08190_));
 sg13g2_and2_1 _27531_ (.A(net667),
    .B(_08190_),
    .X(_02598_));
 sg13g2_nand3_1 _27532_ (.B(net632),
    .C(_07962_),
    .A(net1041),
    .Y(_08191_));
 sg13g2_nand2_1 _27533_ (.Y(_08192_),
    .A(net632),
    .B(_07962_));
 sg13g2_nand2_1 _27534_ (.Y(_08193_),
    .A(\cpu.spi.r_mode[2][0] ),
    .B(_08192_));
 sg13g2_a21oi_1 _27535_ (.A1(_08191_),
    .A2(_08193_),
    .Y(_02599_),
    .B1(net562));
 sg13g2_nand3_1 _27536_ (.B(net632),
    .C(_07962_),
    .A(net1040),
    .Y(_08194_));
 sg13g2_nand2_1 _27537_ (.Y(_08195_),
    .A(_12054_),
    .B(_08192_));
 sg13g2_a21oi_1 _27538_ (.A1(_08194_),
    .A2(_08195_),
    .Y(_02600_),
    .B1(_08060_));
 sg13g2_a221oi_1 _27539_ (.B2(_08161_),
    .C1(_08181_),
    .B1(_07902_),
    .A1(net1050),
    .Y(_08196_),
    .A2(_09427_));
 sg13g2_nor2_1 _27540_ (.A(_09375_),
    .B(_09374_),
    .Y(_08197_));
 sg13g2_a22oi_1 _27541_ (.Y(_08198_),
    .B1(_08196_),
    .B2(_08197_),
    .A2(net447),
    .A1(_04899_));
 sg13g2_nor2_1 _27542_ (.A(net1050),
    .B(_08198_),
    .Y(_08199_));
 sg13g2_nor2_1 _27543_ (.A(\cpu.spi.r_ready ),
    .B(_08196_),
    .Y(_08200_));
 sg13g2_o21ai_1 _27544_ (.B1(net685),
    .Y(_02609_),
    .A1(_08199_),
    .A2(_08200_));
 sg13g2_nor4_1 _27545_ (.A(net437),
    .B(net632),
    .C(_09370_),
    .D(_08179_),
    .Y(_08201_));
 sg13g2_a21o_1 _27546_ (.A2(_07901_),
    .A1(_09411_),
    .B1(_08201_),
    .X(_08202_));
 sg13g2_a22oi_1 _27547_ (.Y(_08203_),
    .B1(_08202_),
    .B2(net1049),
    .A2(_08179_),
    .A1(_09411_));
 sg13g2_nor2_1 _27548_ (.A(net630),
    .B(_08203_),
    .Y(_02610_));
 sg13g2_mux2_1 _27549_ (.A0(net1039),
    .A1(\cpu.spi.r_src[0] ),
    .S(_08184_),
    .X(_08204_));
 sg13g2_and2_1 _27550_ (.A(net667),
    .B(_08204_),
    .X(_02613_));
 sg13g2_mux2_1 _27551_ (.A0(net1039),
    .A1(\cpu.spi.r_src[1] ),
    .S(_08188_),
    .X(_08205_));
 sg13g2_and2_1 _27552_ (.A(net667),
    .B(_08205_),
    .X(_02614_));
 sg13g2_nand3_1 _27553_ (.B(net632),
    .C(_07962_),
    .A(net920),
    .Y(_08206_));
 sg13g2_nand2_1 _27554_ (.Y(_08207_),
    .A(_12035_),
    .B(_08192_));
 sg13g2_a21oi_1 _27555_ (.A1(_08206_),
    .A2(_08207_),
    .Y(_02615_),
    .B1(_08060_));
 sg13g2_buf_1 _27556_ (.A(_07137_),
    .X(_08208_));
 sg13g2_nor2_1 _27557_ (.A(_04994_),
    .B(net93),
    .Y(_08209_));
 sg13g2_buf_2 _27558_ (.A(_08209_),
    .X(_08210_));
 sg13g2_nand2_1 _27559_ (.Y(_08211_),
    .A(net893),
    .B(_08210_));
 sg13g2_inv_1 _27560_ (.Y(_08212_),
    .A(_07137_));
 sg13g2_nand2_1 _27561_ (.Y(_08213_),
    .A(net429),
    .B(_08212_));
 sg13g2_buf_2 _27562_ (.A(_08213_),
    .X(_08214_));
 sg13g2_nand2_1 _27563_ (.Y(_08215_),
    .A(\cpu.uart.r_div_value[0] ),
    .B(_08214_));
 sg13g2_nand3_1 _27564_ (.B(_08211_),
    .C(_08215_),
    .A(net667),
    .Y(_02632_));
 sg13g2_nor2_1 _27565_ (.A(_04883_),
    .B(net93),
    .Y(_08216_));
 sg13g2_nand2_1 _27566_ (.Y(_08217_),
    .A(net920),
    .B(_08216_));
 sg13g2_o21ai_1 _27567_ (.B1(_10080_),
    .Y(_08218_),
    .A1(_04883_),
    .A2(net93));
 sg13g2_a21oi_1 _27568_ (.A1(_08217_),
    .A2(_08218_),
    .Y(_02633_),
    .B1(net562));
 sg13g2_nand2_1 _27569_ (.Y(_08219_),
    .A(net1038),
    .B(_08216_));
 sg13g2_o21ai_1 _27570_ (.B1(\cpu.uart.r_div_value[11] ),
    .Y(_08220_),
    .A1(_04883_),
    .A2(net93));
 sg13g2_a21oi_1 _27571_ (.A1(_08219_),
    .A2(_08220_),
    .Y(_02634_),
    .B1(net562));
 sg13g2_nand2_1 _27572_ (.Y(_08221_),
    .A(net966),
    .B(_08210_));
 sg13g2_nand2_1 _27573_ (.Y(_08222_),
    .A(\cpu.uart.r_div_value[1] ),
    .B(_08214_));
 sg13g2_a21oi_1 _27574_ (.A1(_08221_),
    .A2(_08222_),
    .Y(_02635_),
    .B1(net562));
 sg13g2_nand2_1 _27575_ (.Y(_08223_),
    .A(net920),
    .B(_08210_));
 sg13g2_nand2_1 _27576_ (.Y(_08224_),
    .A(\cpu.uart.r_div_value[2] ),
    .B(_08214_));
 sg13g2_a21oi_1 _27577_ (.A1(_08223_),
    .A2(_08224_),
    .Y(_02636_),
    .B1(net562));
 sg13g2_nand2_1 _27578_ (.Y(_08225_),
    .A(net1038),
    .B(_08210_));
 sg13g2_nand2_1 _27579_ (.Y(_08226_),
    .A(\cpu.uart.r_div_value[3] ),
    .B(_08214_));
 sg13g2_buf_1 _27580_ (.A(_09452_),
    .X(_08227_));
 sg13g2_a21oi_1 _27581_ (.A1(_08225_),
    .A2(_08226_),
    .Y(_02637_),
    .B1(net561));
 sg13g2_nand2_1 _27582_ (.Y(_08228_),
    .A(net1037),
    .B(_08210_));
 sg13g2_nand2_1 _27583_ (.Y(_08229_),
    .A(\cpu.uart.r_div_value[4] ),
    .B(_08214_));
 sg13g2_a21oi_1 _27584_ (.A1(_08228_),
    .A2(_08229_),
    .Y(_02638_),
    .B1(net561));
 sg13g2_nand2_1 _27585_ (.Y(_08230_),
    .A(net1036),
    .B(_08210_));
 sg13g2_nand2_1 _27586_ (.Y(_08231_),
    .A(\cpu.uart.r_div_value[5] ),
    .B(_08214_));
 sg13g2_a21oi_1 _27587_ (.A1(_08230_),
    .A2(_08231_),
    .Y(_02639_),
    .B1(net561));
 sg13g2_nand2_1 _27588_ (.Y(_08232_),
    .A(net1035),
    .B(_08210_));
 sg13g2_nand2_1 _27589_ (.Y(_08233_),
    .A(\cpu.uart.r_div_value[6] ),
    .B(_08214_));
 sg13g2_a21oi_1 _27590_ (.A1(_08232_),
    .A2(_08233_),
    .Y(_02640_),
    .B1(net561));
 sg13g2_nand2_1 _27591_ (.Y(_08234_),
    .A(net985),
    .B(_08210_));
 sg13g2_nand2_1 _27592_ (.Y(_08235_),
    .A(\cpu.uart.r_div_value[7] ),
    .B(_08214_));
 sg13g2_a21oi_1 _27593_ (.A1(_08234_),
    .A2(_08235_),
    .Y(_02641_),
    .B1(_08227_));
 sg13g2_nand2_1 _27594_ (.Y(_08236_),
    .A(net919),
    .B(_08216_));
 sg13g2_o21ai_1 _27595_ (.B1(\cpu.uart.r_div_value[8] ),
    .Y(_08237_),
    .A1(_04883_),
    .A2(net93));
 sg13g2_a21oi_1 _27596_ (.A1(_08236_),
    .A2(_08237_),
    .Y(_02642_),
    .B1(net561));
 sg13g2_nand2_1 _27597_ (.Y(_08238_),
    .A(net966),
    .B(_08216_));
 sg13g2_o21ai_1 _27598_ (.B1(\cpu.uart.r_div_value[9] ),
    .Y(_08239_),
    .A1(_04883_),
    .A2(net93));
 sg13g2_a21oi_1 _27599_ (.A1(_08238_),
    .A2(_08239_),
    .Y(_02643_),
    .B1(net561));
 sg13g2_nand3_1 _27600_ (.B(net382),
    .C(_08212_),
    .A(net1040),
    .Y(_08240_));
 sg13g2_nor4_1 _27601_ (.A(net984),
    .B(net1056),
    .C(net983),
    .D(_07960_),
    .Y(_08241_));
 sg13g2_nand4_1 _27602_ (.B(_09337_),
    .C(_09354_),
    .A(_08502_),
    .Y(_08242_),
    .D(_08241_));
 sg13g2_nand4_1 _27603_ (.B(net706),
    .C(_08240_),
    .A(_09329_),
    .Y(_08243_),
    .D(_08242_));
 sg13g2_nand2b_1 _27604_ (.Y(_02667_),
    .B(_08243_),
    .A_N(_07130_));
 sg13g2_nor2_1 _27605_ (.A(_05058_),
    .B(net93),
    .Y(_08244_));
 sg13g2_nand2_1 _27606_ (.Y(_08245_),
    .A(net966),
    .B(_08244_));
 sg13g2_o21ai_1 _27607_ (.B1(\cpu.uart.r_r_invert ),
    .Y(_08246_),
    .A1(_05058_),
    .A2(net93));
 sg13g2_a21oi_1 _27608_ (.A1(_08245_),
    .A2(_08246_),
    .Y(_02668_),
    .B1(net561));
 sg13g2_a21oi_1 _27609_ (.A1(_07122_),
    .A2(net348),
    .Y(_08247_),
    .B1(net1082));
 sg13g2_a21oi_1 _27610_ (.A1(_07123_),
    .A2(net348),
    .Y(_08248_),
    .B1(_07197_));
 sg13g2_a221oi_1 _27611_ (.B2(_08247_),
    .C1(_08248_),
    .B1(_07121_),
    .A1(net961),
    .Y(_08249_),
    .A2(net1082));
 sg13g2_a21oi_1 _27612_ (.A1(_07114_),
    .A2(_08249_),
    .Y(_08250_),
    .B1(_07194_));
 sg13g2_buf_2 _27613_ (.A(_08250_),
    .X(_08251_));
 sg13g2_o21ai_1 _27614_ (.B1(_08251_),
    .Y(_08252_),
    .A1(net961),
    .A2(_07197_));
 sg13g2_xnor2_1 _27615_ (.Y(_08253_),
    .A(_07123_),
    .B(_08252_));
 sg13g2_nor2_1 _27616_ (.A(net630),
    .B(_08253_),
    .Y(_02671_));
 sg13g2_o21ai_1 _27617_ (.B1(_08251_),
    .Y(_08254_),
    .A1(_07122_),
    .A2(net962));
 sg13g2_nand2_1 _27618_ (.Y(_08255_),
    .A(net1081),
    .B(_08254_));
 sg13g2_nand2b_1 _27619_ (.Y(_08256_),
    .B(net961),
    .A_N(net962));
 sg13g2_o21ai_1 _27620_ (.B1(_08256_),
    .Y(_08257_),
    .A1(net961),
    .A2(_07196_));
 sg13g2_nand3_1 _27621_ (.B(_08251_),
    .C(_08257_),
    .A(_07195_),
    .Y(_08258_));
 sg13g2_a21oi_1 _27622_ (.A1(_08255_),
    .A2(_08258_),
    .Y(_02672_),
    .B1(_08227_));
 sg13g2_nand2_1 _27623_ (.Y(_08259_),
    .A(_07122_),
    .B(_07118_));
 sg13g2_nor3_1 _27624_ (.A(net961),
    .B(_07117_),
    .C(_08259_),
    .Y(_08260_));
 sg13g2_o21ai_1 _27625_ (.B1(_08251_),
    .Y(_08261_),
    .A1(_07117_),
    .A2(_07205_));
 sg13g2_a22oi_1 _27626_ (.Y(_08262_),
    .B1(_08261_),
    .B2(_07120_),
    .A2(_08260_),
    .A1(_08251_));
 sg13g2_nor2_1 _27627_ (.A(net630),
    .B(_08262_),
    .Y(_02673_));
 sg13g2_a21oi_1 _27628_ (.A1(_07205_),
    .A2(_08251_),
    .Y(_08263_),
    .B1(net962));
 sg13g2_nor2b_1 _27629_ (.A(net961),
    .B_N(_07118_),
    .Y(_08264_));
 sg13g2_a21oi_1 _27630_ (.A1(_08251_),
    .A2(_08264_),
    .Y(_08265_),
    .B1(_06813_));
 sg13g2_nor2b_1 _27631_ (.A(_08263_),
    .B_N(_08265_),
    .Y(_02674_));
 sg13g2_nor2b_1 _27632_ (.A(net958),
    .B_N(_07213_),
    .Y(_08266_));
 sg13g2_o21ai_1 _27633_ (.B1(_08266_),
    .Y(_08267_),
    .A1(_09328_),
    .A2(_07152_));
 sg13g2_o21ai_1 _27634_ (.B1(_10252_),
    .Y(_08268_),
    .A1(_00223_),
    .A2(_04936_));
 sg13g2_nor2b_1 _27635_ (.A(_07240_),
    .B_N(_08268_),
    .Y(_08269_));
 sg13g2_a21o_1 _27636_ (.A2(net382),
    .A1(_10186_),
    .B1(net381),
    .X(_08270_));
 sg13g2_a22oi_1 _27637_ (.Y(_08271_),
    .B1(_08270_),
    .B2(_07213_),
    .A2(_08269_),
    .A1(net586));
 sg13g2_o21ai_1 _27638_ (.B1(_09328_),
    .Y(_08272_),
    .A1(_08208_),
    .A2(_08271_));
 sg13g2_a21oi_1 _27639_ (.A1(_08267_),
    .A2(_08272_),
    .Y(_02676_),
    .B1(net561));
 sg13g2_nand2_1 _27640_ (.Y(_08273_),
    .A(net919),
    .B(_08244_));
 sg13g2_o21ai_1 _27641_ (.B1(\cpu.uart.r_x_invert ),
    .Y(_08274_),
    .A1(_05058_),
    .A2(_08208_));
 sg13g2_a21oi_1 _27642_ (.A1(_08273_),
    .A2(_08274_),
    .Y(_02677_),
    .B1(net705));
 sg13g2_mux2_1 _27643_ (.A0(_07142_),
    .A1(_07216_),
    .S(net960),
    .X(_08275_));
 sg13g2_o21ai_1 _27644_ (.B1(_07231_),
    .Y(_08276_),
    .A1(_07138_),
    .A2(_07240_));
 sg13g2_a21oi_2 _27645_ (.B1(_08276_),
    .Y(_08277_),
    .A2(_08275_),
    .A1(_07154_));
 sg13g2_nand4_1 _27646_ (.B(_07138_),
    .C(_07152_),
    .A(net958),
    .Y(_08278_),
    .D(_07213_));
 sg13g2_nand4_1 _27647_ (.B(_07225_),
    .C(_08277_),
    .A(net958),
    .Y(_08279_),
    .D(_08278_));
 sg13g2_o21ai_1 _27648_ (.B1(_08279_),
    .Y(_08280_),
    .A1(net958),
    .A2(_08277_));
 sg13g2_nor2_1 _27649_ (.A(net630),
    .B(_08280_),
    .Y(_02680_));
 sg13g2_a21o_1 _27650_ (.A2(_08275_),
    .A1(_07154_),
    .B1(_08276_),
    .X(_08281_));
 sg13g2_buf_1 _27651_ (.A(_08281_),
    .X(_08282_));
 sg13g2_a21oi_1 _27652_ (.A1(net959),
    .A2(net960),
    .Y(_08283_),
    .B1(net958));
 sg13g2_o21ai_1 _27653_ (.B1(_07139_),
    .Y(_08284_),
    .A1(_08282_),
    .A2(_08283_));
 sg13g2_nand4_1 _27654_ (.B(net958),
    .C(_07225_),
    .A(_07153_),
    .Y(_08285_),
    .D(_08277_));
 sg13g2_a21oi_1 _27655_ (.A1(_08284_),
    .A2(_08285_),
    .Y(_02681_),
    .B1(net705));
 sg13g2_nor3_1 _27656_ (.A(net960),
    .B(_07141_),
    .C(_08282_),
    .Y(_08286_));
 sg13g2_and2_1 _27657_ (.A(net960),
    .B(_07141_),
    .X(_08287_));
 sg13g2_o21ai_1 _27658_ (.B1(_07148_),
    .Y(_08288_),
    .A1(_08286_),
    .A2(_08287_));
 sg13g2_nor2_1 _27659_ (.A(_07152_),
    .B(_07233_),
    .Y(_08289_));
 sg13g2_a21oi_1 _27660_ (.A1(net960),
    .A2(_08282_),
    .Y(_08290_),
    .B1(_08289_));
 sg13g2_a21oi_1 _27661_ (.A1(_08288_),
    .A2(_08290_),
    .Y(_02682_),
    .B1(net705));
 sg13g2_a21oi_1 _27662_ (.A1(_07139_),
    .A2(net958),
    .Y(_08291_),
    .B1(net960));
 sg13g2_o21ai_1 _27663_ (.B1(net959),
    .Y(_08292_),
    .A1(_08282_),
    .A2(_08291_));
 sg13g2_nor2_1 _27664_ (.A(_07141_),
    .B(_07215_),
    .Y(_08293_));
 sg13g2_o21ai_1 _27665_ (.B1(_08277_),
    .Y(_08294_),
    .A1(_08289_),
    .A2(_08293_));
 sg13g2_a21oi_1 _27666_ (.A1(_08292_),
    .A2(_08294_),
    .Y(_02683_),
    .B1(net705));
 sg13g2_nand2b_1 _27667_ (.Y(\cpu.ex.genblk3.c_supmode ),
    .B(_07419_),
    .A_N(_07416_));
 sg13g2_nand2_1 _27668_ (.Y(_08295_),
    .A(_09989_),
    .B(_07871_));
 sg13g2_o21ai_1 _27669_ (.B1(_09953_),
    .Y(\cpu.qspi.c_rstrobe_d ),
    .A1(_09956_),
    .A2(_08295_));
 sg13g2_nor4_1 _27670_ (.A(_09948_),
    .B(_09938_),
    .C(net788),
    .D(_07870_),
    .Y(_08296_));
 sg13g2_a22oi_1 _27671_ (.Y(_08297_),
    .B1(_07855_),
    .B2(_08296_),
    .A2(net788),
    .A1(_09947_));
 sg13g2_nor2_1 _27672_ (.A(net831),
    .B(_08297_),
    .Y(\cpu.qspi.c_wstrobe_d ));
 sg13g2_nor2_1 _27673_ (.A(_00189_),
    .B(_08297_),
    .Y(\cpu.qspi.c_wstrobe_i ));
 sg13g2_mux4_1 _27674_ (.S0(_04998_),
    .A0(_09288_),
    .A1(_09302_),
    .A2(_09308_),
    .A3(_09297_),
    .S1(\cpu.gpio.r_uart_rx_src[1] ),
    .X(_08298_));
 sg13g2_mux4_1 _27675_ (.S0(_04998_),
    .A0(_09304_),
    .A1(_09310_),
    .A2(_09299_),
    .A3(_09290_),
    .S1(\cpu.gpio.r_uart_rx_src[1] ),
    .X(_08299_));
 sg13g2_mux2_1 _27676_ (.A0(_08298_),
    .A1(_08299_),
    .S(\cpu.gpio.r_uart_rx_src[2] ),
    .X(\cpu.gpio.uart_rx ));
 sg13g2_mux4_1 _27677_ (.S0(_04989_),
    .A0(net1104),
    .A1(net1105),
    .A2(net1078),
    .A3(net1077),
    .S1(_05342_),
    .X(_08300_));
 sg13g2_mux4_1 _27678_ (.S0(_04989_),
    .A0(\cpu.gpio.genblk2[4].srcs_io[0] ),
    .A1(net1080),
    .A2(net1102),
    .A3(net1103),
    .S1(_05342_),
    .X(_08301_));
 sg13g2_nor2b_1 _27679_ (.A(_05404_),
    .B_N(_08301_),
    .Y(_08302_));
 sg13g2_a21oi_1 _27680_ (.A1(_05404_),
    .A2(_08300_),
    .Y(_08303_),
    .B1(_08302_));
 sg13g2_nand2b_1 _27681_ (.Y(_08304_),
    .B(net1076),
    .A_N(_04989_));
 sg13g2_nand3_1 _27682_ (.B(_05342_),
    .C(net1079),
    .A(_04989_),
    .Y(_08305_));
 sg13g2_o21ai_1 _27683_ (.B1(_08305_),
    .Y(_08306_),
    .A1(_05342_),
    .A2(_08304_));
 sg13g2_nand3_1 _27684_ (.B(_00187_),
    .C(_08306_),
    .A(_05465_),
    .Y(_08307_));
 sg13g2_o21ai_1 _27685_ (.B1(_08307_),
    .Y(net15),
    .A1(_05465_),
    .A2(_08303_));
 sg13g2_mux4_1 _27686_ (.S0(_05544_),
    .A0(net1104),
    .A1(net1105),
    .A2(net1078),
    .A3(net1077),
    .S1(_05639_),
    .X(_08308_));
 sg13g2_mux4_1 _27687_ (.S0(_05544_),
    .A0(\cpu.gpio.genblk2[5].srcs_io[0] ),
    .A1(net1080),
    .A2(net1102),
    .A3(net1103),
    .S1(_05639_),
    .X(_08309_));
 sg13g2_nor2b_1 _27688_ (.A(_05671_),
    .B_N(_08309_),
    .Y(_08310_));
 sg13g2_a21oi_1 _27689_ (.A1(_05671_),
    .A2(_08308_),
    .Y(_08311_),
    .B1(_08310_));
 sg13g2_nand2b_1 _27690_ (.Y(_08312_),
    .B(net1076),
    .A_N(_05544_));
 sg13g2_nand3_1 _27691_ (.B(_05639_),
    .C(net1079),
    .A(_05544_),
    .Y(_08313_));
 sg13g2_o21ai_1 _27692_ (.B1(_08313_),
    .Y(_08314_),
    .A1(_05639_),
    .A2(_08312_));
 sg13g2_nand3_1 _27693_ (.B(_00186_),
    .C(_08314_),
    .A(_05053_),
    .Y(_08315_));
 sg13g2_o21ai_1 _27694_ (.B1(_08315_),
    .Y(net16),
    .A1(_05053_),
    .A2(_08311_));
 sg13g2_mux4_1 _27695_ (.S0(_05006_),
    .A0(net1104),
    .A1(net1105),
    .A2(net1078),
    .A3(net1077),
    .S1(_06402_),
    .X(_08316_));
 sg13g2_mux4_1 _27696_ (.S0(_05006_),
    .A0(\cpu.gpio.genblk2[6].srcs_io[0] ),
    .A1(net1080),
    .A2(net1102),
    .A3(net1103),
    .S1(_06402_),
    .X(_08317_));
 sg13g2_nor2b_1 _27697_ (.A(\cpu.gpio.r_src_io[6][2] ),
    .B_N(_08317_),
    .Y(_08318_));
 sg13g2_a21oi_1 _27698_ (.A1(\cpu.gpio.r_src_io[6][2] ),
    .A2(_08316_),
    .Y(_08319_),
    .B1(_08318_));
 sg13g2_nand2b_1 _27699_ (.Y(_08320_),
    .B(net1076),
    .A_N(_05006_));
 sg13g2_nand3_1 _27700_ (.B(net1079),
    .C(_06402_),
    .A(_05006_),
    .Y(_08321_));
 sg13g2_o21ai_1 _27701_ (.B1(_08321_),
    .Y(_08322_),
    .A1(_06402_),
    .A2(_08320_));
 sg13g2_nand3_1 _27702_ (.B(\cpu.gpio.r_src_io[6][3] ),
    .C(_08322_),
    .A(_00106_),
    .Y(_08323_));
 sg13g2_o21ai_1 _27703_ (.B1(_08323_),
    .Y(net17),
    .A1(\cpu.gpio.r_src_io[6][3] ),
    .A2(_08319_));
 sg13g2_mux4_1 _27704_ (.S0(_05547_),
    .A0(net1104),
    .A1(net1105),
    .A2(net1078),
    .A3(net1077),
    .S1(_06403_),
    .X(_08324_));
 sg13g2_mux4_1 _27705_ (.S0(_05547_),
    .A0(\cpu.gpio.genblk2[7].srcs_io[0] ),
    .A1(net1080),
    .A2(net1102),
    .A3(net1103),
    .S1(_06403_),
    .X(_08325_));
 sg13g2_nor2b_1 _27706_ (.A(\cpu.gpio.r_src_io[7][2] ),
    .B_N(_08325_),
    .Y(_08326_));
 sg13g2_a21oi_1 _27707_ (.A1(\cpu.gpio.r_src_io[7][2] ),
    .A2(_08324_),
    .Y(_08327_),
    .B1(_08326_));
 sg13g2_nand2b_1 _27708_ (.Y(_08328_),
    .B(net1076),
    .A_N(_05547_));
 sg13g2_nand3_1 _27709_ (.B(net1079),
    .C(_06403_),
    .A(_05547_),
    .Y(_08329_));
 sg13g2_o21ai_1 _27710_ (.B1(_08329_),
    .Y(_08330_),
    .A1(_06403_),
    .A2(_08328_));
 sg13g2_nand3_1 _27711_ (.B(\cpu.gpio.r_src_io[7][3] ),
    .C(_08330_),
    .A(_00146_),
    .Y(_08331_));
 sg13g2_o21ai_1 _27712_ (.B1(_08331_),
    .Y(net18),
    .A1(\cpu.gpio.r_src_io[7][3] ),
    .A2(_08327_));
 sg13g2_xor2_1 _27713_ (.B(clknet_leaf_77_clk),
    .A(\cpu.r_clk_invert ),
    .X(net21));
 sg13g2_mux4_1 _27714_ (.S0(_05541_),
    .A0(net1104),
    .A1(net1105),
    .A2(net1078),
    .A3(net1077),
    .S1(_06406_),
    .X(_08332_));
 sg13g2_mux4_1 _27715_ (.S0(_05541_),
    .A0(\cpu.gpio.genblk1[3].srcs_o[0] ),
    .A1(net1080),
    .A2(net1102),
    .A3(net1103),
    .S1(_06406_),
    .X(_08333_));
 sg13g2_nor2b_1 _27716_ (.A(\cpu.gpio.r_src_o[3][2] ),
    .B_N(_08333_),
    .Y(_08334_));
 sg13g2_a21oi_1 _27717_ (.A1(\cpu.gpio.r_src_o[3][2] ),
    .A2(_08332_),
    .Y(_08335_),
    .B1(_08334_));
 sg13g2_nand2b_1 _27718_ (.Y(_08336_),
    .B(_08175_),
    .A_N(_05541_));
 sg13g2_nand3_1 _27719_ (.B(net1079),
    .C(_06406_),
    .A(_05541_),
    .Y(_08337_));
 sg13g2_o21ai_1 _27720_ (.B1(_08337_),
    .Y(_08338_),
    .A1(_06406_),
    .A2(_08336_));
 sg13g2_nand3_1 _27721_ (.B(\cpu.gpio.r_src_o[3][3] ),
    .C(_08338_),
    .A(_00149_),
    .Y(_08339_));
 sg13g2_o21ai_1 _27722_ (.B1(_08339_),
    .Y(net22),
    .A1(\cpu.gpio.r_src_o[3][3] ),
    .A2(_08335_));
 sg13g2_mux4_1 _27723_ (.S0(_04984_),
    .A0(net1104),
    .A1(net1105),
    .A2(_08158_),
    .A3(net1077),
    .S1(_06409_),
    .X(_08340_));
 sg13g2_mux4_1 _27724_ (.S0(_04984_),
    .A0(\cpu.gpio.genblk1[4].srcs_o[0] ),
    .A1(net1080),
    .A2(_12101_),
    .A3(_12085_),
    .S1(_06409_),
    .X(_08341_));
 sg13g2_nor2b_1 _27725_ (.A(\cpu.gpio.r_src_o[4][2] ),
    .B_N(_08341_),
    .Y(_08342_));
 sg13g2_a21oi_1 _27726_ (.A1(\cpu.gpio.r_src_o[4][2] ),
    .A2(_08340_),
    .Y(_08343_),
    .B1(_08342_));
 sg13g2_nand2b_1 _27727_ (.Y(_08344_),
    .B(net1076),
    .A_N(_04984_));
 sg13g2_nand3_1 _27728_ (.B(net1079),
    .C(_06409_),
    .A(_04984_),
    .Y(_08345_));
 sg13g2_o21ai_1 _27729_ (.B1(_08345_),
    .Y(_08346_),
    .A1(_06409_),
    .A2(_08344_));
 sg13g2_nand3_1 _27730_ (.B(\cpu.gpio.r_src_o[4][3] ),
    .C(_08346_),
    .A(_00108_),
    .Y(_08347_));
 sg13g2_o21ai_1 _27731_ (.B1(_08347_),
    .Y(net23),
    .A1(\cpu.gpio.r_src_o[4][3] ),
    .A2(_08343_));
 sg13g2_mux4_1 _27732_ (.S0(_05534_),
    .A0(_12083_),
    .A1(_12076_),
    .A2(_08158_),
    .A3(_08172_),
    .S1(_06410_),
    .X(_08348_));
 sg13g2_mux4_1 _27733_ (.S0(_05534_),
    .A0(\cpu.gpio.genblk1[5].srcs_o[0] ),
    .A1(net1080),
    .A2(net1102),
    .A3(net1103),
    .S1(_06410_),
    .X(_08349_));
 sg13g2_nor2b_1 _27734_ (.A(\cpu.gpio.r_src_o[5][2] ),
    .B_N(_08349_),
    .Y(_08350_));
 sg13g2_a21oi_1 _27735_ (.A1(\cpu.gpio.r_src_o[5][2] ),
    .A2(_08348_),
    .Y(_08351_),
    .B1(_08350_));
 sg13g2_nand2b_1 _27736_ (.Y(_08352_),
    .B(_08175_),
    .A_N(_05534_));
 sg13g2_nand3_1 _27737_ (.B(net1079),
    .C(_06410_),
    .A(_05534_),
    .Y(_08353_));
 sg13g2_o21ai_1 _27738_ (.B1(_08353_),
    .Y(_08354_),
    .A1(_06410_),
    .A2(_08352_));
 sg13g2_nand3_1 _27739_ (.B(\cpu.gpio.r_src_o[5][3] ),
    .C(_08354_),
    .A(_00148_),
    .Y(_08355_));
 sg13g2_o21ai_1 _27740_ (.B1(_08355_),
    .Y(net24),
    .A1(\cpu.gpio.r_src_o[5][3] ),
    .A2(_08351_));
 sg13g2_mux4_1 _27741_ (.S0(_05000_),
    .A0(_12083_),
    .A1(_12076_),
    .A2(net1078),
    .A3(_08172_),
    .S1(_07772_),
    .X(_08356_));
 sg13g2_mux4_1 _27742_ (.S0(_05000_),
    .A0(\cpu.gpio.genblk1[6].srcs_o[0] ),
    .A1(_07224_),
    .A2(_12101_),
    .A3(_12085_),
    .S1(_07772_),
    .X(_08357_));
 sg13g2_nor2b_1 _27743_ (.A(\cpu.gpio.r_src_o[6][2] ),
    .B_N(_08357_),
    .Y(_08358_));
 sg13g2_a21oi_1 _27744_ (.A1(\cpu.gpio.r_src_o[6][2] ),
    .A2(_08356_),
    .Y(_08359_),
    .B1(_08358_));
 sg13g2_nand2b_1 _27745_ (.Y(_08360_),
    .B(net1076),
    .A_N(_05000_));
 sg13g2_nand3_1 _27746_ (.B(_07867_),
    .C(_07772_),
    .A(_05000_),
    .Y(_08361_));
 sg13g2_o21ai_1 _27747_ (.B1(_08361_),
    .Y(_08362_),
    .A1(_07772_),
    .A2(_08360_));
 sg13g2_nand3_1 _27748_ (.B(\cpu.gpio.r_src_o[6][3] ),
    .C(_08362_),
    .A(_00107_),
    .Y(_08363_));
 sg13g2_o21ai_1 _27749_ (.B1(_08363_),
    .Y(net25),
    .A1(\cpu.gpio.r_src_o[6][3] ),
    .A2(_08359_));
 sg13g2_mux4_1 _27750_ (.S0(_05545_),
    .A0(net1104),
    .A1(net1105),
    .A2(net1078),
    .A3(net1077),
    .S1(_06412_),
    .X(_08364_));
 sg13g2_mux4_1 _27751_ (.S0(_05545_),
    .A0(\cpu.gpio.genblk1[7].srcs_o[0] ),
    .A1(_07224_),
    .A2(net1102),
    .A3(net1103),
    .S1(_06412_),
    .X(_08365_));
 sg13g2_nor2b_1 _27752_ (.A(\cpu.gpio.r_src_o[7][2] ),
    .B_N(_08365_),
    .Y(_08366_));
 sg13g2_a21oi_1 _27753_ (.A1(\cpu.gpio.r_src_o[7][2] ),
    .A2(_08364_),
    .Y(_08367_),
    .B1(_08366_));
 sg13g2_nand2b_1 _27754_ (.Y(_08368_),
    .B(net1076),
    .A_N(_05545_));
 sg13g2_nand3_1 _27755_ (.B(net1079),
    .C(_06412_),
    .A(_05545_),
    .Y(_08369_));
 sg13g2_o21ai_1 _27756_ (.B1(_08369_),
    .Y(_08370_),
    .A1(_06412_),
    .A2(_08368_));
 sg13g2_nand3_1 _27757_ (.B(\cpu.gpio.r_src_o[7][3] ),
    .C(_08370_),
    .A(_00147_),
    .Y(_08371_));
 sg13g2_o21ai_1 _27758_ (.B1(_08371_),
    .Y(net26),
    .A1(\cpu.gpio.r_src_o[7][3] ),
    .A2(_08367_));
 sg13g2_dfrbp_1 _27759_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1136),
    .D(_00317_),
    .Q_N(_15004_),
    .Q(\cpu.intr.r_swi ));
 sg13g2_dfrbp_1 _27760_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1137),
    .D(_00318_),
    .Q_N(_15003_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[5] ));
 sg13g2_dfrbp_1 _27761_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1138),
    .D(_00319_),
    .Q_N(_15002_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[4] ));
 sg13g2_dfrbp_1 _27762_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1139),
    .D(_00320_),
    .Q_N(_15001_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[3] ));
 sg13g2_dfrbp_1 _27763_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1140),
    .D(_00321_),
    .Q_N(_15000_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[2] ));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_1 _27765_ (.A(net6),
    .X(net4));
 sg13g2_buf_1 _27766_ (.A(net6),
    .X(net5));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1141),
    .D(_00322_),
    .Q_N(_14999_),
    .Q(\cpu.dcache.r_data[0][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1142),
    .D(_00323_),
    .Q_N(_00103_),
    .Q(\cpu.dcache.r_data[0][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1143),
    .D(_00324_),
    .Q_N(_00113_),
    .Q(\cpu.dcache.r_data[0][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1144),
    .D(_00325_),
    .Q_N(_00124_),
    .Q(\cpu.dcache.r_data[0][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1145),
    .D(_00326_),
    .Q_N(_00131_),
    .Q(\cpu.dcache.r_data[0][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1146),
    .D(_00327_),
    .Q_N(_00143_),
    .Q(\cpu.dcache.r_data[0][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1147),
    .D(_00328_),
    .Q_N(_00155_),
    .Q(\cpu.dcache.r_data[0][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1148),
    .D(_00329_),
    .Q_N(_14998_),
    .Q(\cpu.dcache.r_data[0][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1149),
    .D(_00330_),
    .Q_N(_00091_),
    .Q(\cpu.dcache.r_data[0][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1150),
    .D(_00331_),
    .Q_N(_00101_),
    .Q(\cpu.dcache.r_data[0][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][19]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1151),
    .D(_00332_),
    .Q_N(_00111_),
    .Q(\cpu.dcache.r_data[0][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1152),
    .D(_00333_),
    .Q_N(_14997_),
    .Q(\cpu.dcache.r_data[0][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][20]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1153),
    .D(_00334_),
    .Q_N(_00122_),
    .Q(\cpu.dcache.r_data[0][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][21]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1154),
    .D(_00335_),
    .Q_N(_00129_),
    .Q(\cpu.dcache.r_data[0][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][22]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1155),
    .D(_00336_),
    .Q_N(_00141_),
    .Q(\cpu.dcache.r_data[0][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][23]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1156),
    .D(_00337_),
    .Q_N(_00153_),
    .Q(\cpu.dcache.r_data[0][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][24]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1157),
    .D(_00338_),
    .Q_N(_00311_),
    .Q(\cpu.dcache.r_data[0][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][25]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1158),
    .D(_00339_),
    .Q_N(_00092_),
    .Q(\cpu.dcache.r_data[0][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][26]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1159),
    .D(_00340_),
    .Q_N(_00102_),
    .Q(\cpu.dcache.r_data[0][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][27]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1160),
    .D(_00341_),
    .Q_N(_00112_),
    .Q(\cpu.dcache.r_data[0][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][28]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1161),
    .D(_00342_),
    .Q_N(_00123_),
    .Q(\cpu.dcache.r_data[0][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][29]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1162),
    .D(_00343_),
    .Q_N(_00130_),
    .Q(\cpu.dcache.r_data[0][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1163),
    .D(_00344_),
    .Q_N(_14996_),
    .Q(\cpu.dcache.r_data[0][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][30]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1164),
    .D(_00345_),
    .Q_N(_00142_),
    .Q(\cpu.dcache.r_data[0][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][31]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1165),
    .D(_00346_),
    .Q_N(_00154_),
    .Q(\cpu.dcache.r_data[0][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1166),
    .D(_00347_),
    .Q_N(_14995_),
    .Q(\cpu.dcache.r_data[0][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1167),
    .D(_00348_),
    .Q_N(_00121_),
    .Q(\cpu.dcache.r_data[0][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1168),
    .D(_00349_),
    .Q_N(_00128_),
    .Q(\cpu.dcache.r_data[0][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1169),
    .D(_00350_),
    .Q_N(_00140_),
    .Q(\cpu.dcache.r_data[0][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1170),
    .D(_00351_),
    .Q_N(_00152_),
    .Q(\cpu.dcache.r_data[0][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1171),
    .D(_00352_),
    .Q_N(_00312_),
    .Q(\cpu.dcache.r_data[0][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1172),
    .D(_00353_),
    .Q_N(_00093_),
    .Q(\cpu.dcache.r_data[0][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1173),
    .D(_00354_),
    .Q_N(_14994_),
    .Q(\cpu.dcache.r_data[1][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1174),
    .D(_00355_),
    .Q_N(_14993_),
    .Q(\cpu.dcache.r_data[1][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1175),
    .D(_00356_),
    .Q_N(_14992_),
    .Q(\cpu.dcache.r_data[1][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1176),
    .D(_00357_),
    .Q_N(_14991_),
    .Q(\cpu.dcache.r_data[1][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1177),
    .D(_00358_),
    .Q_N(_14990_),
    .Q(\cpu.dcache.r_data[1][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1178),
    .D(_00359_),
    .Q_N(_14989_),
    .Q(\cpu.dcache.r_data[1][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1179),
    .D(_00360_),
    .Q_N(_14988_),
    .Q(\cpu.dcache.r_data[1][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1180),
    .D(_00361_),
    .Q_N(_14987_),
    .Q(\cpu.dcache.r_data[1][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1181),
    .D(_00362_),
    .Q_N(_14986_),
    .Q(\cpu.dcache.r_data[1][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1182),
    .D(_00363_),
    .Q_N(_14985_),
    .Q(\cpu.dcache.r_data[1][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][19]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1183),
    .D(_00364_),
    .Q_N(_14984_),
    .Q(\cpu.dcache.r_data[1][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1184),
    .D(_00365_),
    .Q_N(_14983_),
    .Q(\cpu.dcache.r_data[1][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][20]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1185),
    .D(_00366_),
    .Q_N(_14982_),
    .Q(\cpu.dcache.r_data[1][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][21]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1186),
    .D(_00367_),
    .Q_N(_14981_),
    .Q(\cpu.dcache.r_data[1][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][22]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1187),
    .D(_00368_),
    .Q_N(_14980_),
    .Q(\cpu.dcache.r_data[1][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][23]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1188),
    .D(_00369_),
    .Q_N(_14979_),
    .Q(\cpu.dcache.r_data[1][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][24]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1189),
    .D(_00370_),
    .Q_N(_14978_),
    .Q(\cpu.dcache.r_data[1][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][25]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1190),
    .D(_00371_),
    .Q_N(_14977_),
    .Q(\cpu.dcache.r_data[1][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][26]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1191),
    .D(_00372_),
    .Q_N(_14976_),
    .Q(\cpu.dcache.r_data[1][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][27]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1192),
    .D(_00373_),
    .Q_N(_14975_),
    .Q(\cpu.dcache.r_data[1][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][28]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1193),
    .D(_00374_),
    .Q_N(_14974_),
    .Q(\cpu.dcache.r_data[1][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][29]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1194),
    .D(_00375_),
    .Q_N(_14973_),
    .Q(\cpu.dcache.r_data[1][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1195),
    .D(_00376_),
    .Q_N(_14972_),
    .Q(\cpu.dcache.r_data[1][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][30]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1196),
    .D(_00377_),
    .Q_N(_14971_),
    .Q(\cpu.dcache.r_data[1][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][31]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1197),
    .D(_00378_),
    .Q_N(_14970_),
    .Q(\cpu.dcache.r_data[1][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1198),
    .D(_00379_),
    .Q_N(_14969_),
    .Q(\cpu.dcache.r_data[1][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1199),
    .D(_00380_),
    .Q_N(_14968_),
    .Q(\cpu.dcache.r_data[1][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1200),
    .D(_00381_),
    .Q_N(_14967_),
    .Q(\cpu.dcache.r_data[1][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1201),
    .D(_00382_),
    .Q_N(_14966_),
    .Q(\cpu.dcache.r_data[1][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1202),
    .D(_00383_),
    .Q_N(_14965_),
    .Q(\cpu.dcache.r_data[1][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1203),
    .D(_00384_),
    .Q_N(_14964_),
    .Q(\cpu.dcache.r_data[1][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1204),
    .D(_00385_),
    .Q_N(_14963_),
    .Q(\cpu.dcache.r_data[1][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1205),
    .D(_00386_),
    .Q_N(_14962_),
    .Q(\cpu.dcache.r_data[2][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1206),
    .D(_00387_),
    .Q_N(_14961_),
    .Q(\cpu.dcache.r_data[2][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1207),
    .D(_00388_),
    .Q_N(_14960_),
    .Q(\cpu.dcache.r_data[2][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1208),
    .D(_00389_),
    .Q_N(_14959_),
    .Q(\cpu.dcache.r_data[2][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1209),
    .D(_00390_),
    .Q_N(_14958_),
    .Q(\cpu.dcache.r_data[2][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1210),
    .D(_00391_),
    .Q_N(_14957_),
    .Q(\cpu.dcache.r_data[2][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1211),
    .D(_00392_),
    .Q_N(_14956_),
    .Q(\cpu.dcache.r_data[2][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1212),
    .D(_00393_),
    .Q_N(_14955_),
    .Q(\cpu.dcache.r_data[2][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1213),
    .D(_00394_),
    .Q_N(_14954_),
    .Q(\cpu.dcache.r_data[2][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1214),
    .D(_00395_),
    .Q_N(_14953_),
    .Q(\cpu.dcache.r_data[2][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][19]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1215),
    .D(_00396_),
    .Q_N(_14952_),
    .Q(\cpu.dcache.r_data[2][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1216),
    .D(_00397_),
    .Q_N(_14951_),
    .Q(\cpu.dcache.r_data[2][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][20]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1217),
    .D(_00398_),
    .Q_N(_14950_),
    .Q(\cpu.dcache.r_data[2][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][21]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1218),
    .D(_00399_),
    .Q_N(_14949_),
    .Q(\cpu.dcache.r_data[2][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][22]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1219),
    .D(_00400_),
    .Q_N(_14948_),
    .Q(\cpu.dcache.r_data[2][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][23]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1220),
    .D(_00401_),
    .Q_N(_14947_),
    .Q(\cpu.dcache.r_data[2][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][24]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1221),
    .D(_00402_),
    .Q_N(_14946_),
    .Q(\cpu.dcache.r_data[2][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][25]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1222),
    .D(_00403_),
    .Q_N(_14945_),
    .Q(\cpu.dcache.r_data[2][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][26]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1223),
    .D(_00404_),
    .Q_N(_14944_),
    .Q(\cpu.dcache.r_data[2][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][27]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1224),
    .D(_00405_),
    .Q_N(_14943_),
    .Q(\cpu.dcache.r_data[2][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][28]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1225),
    .D(_00406_),
    .Q_N(_14942_),
    .Q(\cpu.dcache.r_data[2][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][29]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1226),
    .D(_00407_),
    .Q_N(_14941_),
    .Q(\cpu.dcache.r_data[2][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1227),
    .D(_00408_),
    .Q_N(_14940_),
    .Q(\cpu.dcache.r_data[2][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][30]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1228),
    .D(_00409_),
    .Q_N(_14939_),
    .Q(\cpu.dcache.r_data[2][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][31]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1229),
    .D(_00410_),
    .Q_N(_14938_),
    .Q(\cpu.dcache.r_data[2][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1230),
    .D(_00411_),
    .Q_N(_14937_),
    .Q(\cpu.dcache.r_data[2][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1231),
    .D(_00412_),
    .Q_N(_14936_),
    .Q(\cpu.dcache.r_data[2][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1232),
    .D(_00413_),
    .Q_N(_14935_),
    .Q(\cpu.dcache.r_data[2][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1233),
    .D(_00414_),
    .Q_N(_14934_),
    .Q(\cpu.dcache.r_data[2][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1234),
    .D(_00415_),
    .Q_N(_14933_),
    .Q(\cpu.dcache.r_data[2][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1235),
    .D(_00416_),
    .Q_N(_14932_),
    .Q(\cpu.dcache.r_data[2][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1236),
    .D(_00417_),
    .Q_N(_14931_),
    .Q(\cpu.dcache.r_data[2][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1237),
    .D(_00418_),
    .Q_N(_14930_),
    .Q(\cpu.dcache.r_data[3][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1238),
    .D(_00419_),
    .Q_N(_14929_),
    .Q(\cpu.dcache.r_data[3][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1239),
    .D(_00420_),
    .Q_N(_14928_),
    .Q(\cpu.dcache.r_data[3][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1240),
    .D(_00421_),
    .Q_N(_14927_),
    .Q(\cpu.dcache.r_data[3][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1241),
    .D(_00422_),
    .Q_N(_14926_),
    .Q(\cpu.dcache.r_data[3][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1242),
    .D(_00423_),
    .Q_N(_14925_),
    .Q(\cpu.dcache.r_data[3][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1243),
    .D(_00424_),
    .Q_N(_14924_),
    .Q(\cpu.dcache.r_data[3][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1244),
    .D(_00425_),
    .Q_N(_14923_),
    .Q(\cpu.dcache.r_data[3][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1245),
    .D(_00426_),
    .Q_N(_14922_),
    .Q(\cpu.dcache.r_data[3][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1246),
    .D(_00427_),
    .Q_N(_14921_),
    .Q(\cpu.dcache.r_data[3][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][19]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1247),
    .D(_00428_),
    .Q_N(_14920_),
    .Q(\cpu.dcache.r_data[3][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1248),
    .D(_00429_),
    .Q_N(_14919_),
    .Q(\cpu.dcache.r_data[3][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][20]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1249),
    .D(_00430_),
    .Q_N(_14918_),
    .Q(\cpu.dcache.r_data[3][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][21]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1250),
    .D(_00431_),
    .Q_N(_14917_),
    .Q(\cpu.dcache.r_data[3][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][22]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1251),
    .D(_00432_),
    .Q_N(_14916_),
    .Q(\cpu.dcache.r_data[3][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][23]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1252),
    .D(_00433_),
    .Q_N(_14915_),
    .Q(\cpu.dcache.r_data[3][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][24]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1253),
    .D(_00434_),
    .Q_N(_14914_),
    .Q(\cpu.dcache.r_data[3][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][25]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1254),
    .D(_00435_),
    .Q_N(_14913_),
    .Q(\cpu.dcache.r_data[3][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][26]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1255),
    .D(_00436_),
    .Q_N(_14912_),
    .Q(\cpu.dcache.r_data[3][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][27]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1256),
    .D(_00437_),
    .Q_N(_14911_),
    .Q(\cpu.dcache.r_data[3][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][28]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1257),
    .D(_00438_),
    .Q_N(_14910_),
    .Q(\cpu.dcache.r_data[3][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][29]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1258),
    .D(_00439_),
    .Q_N(_14909_),
    .Q(\cpu.dcache.r_data[3][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1259),
    .D(_00440_),
    .Q_N(_14908_),
    .Q(\cpu.dcache.r_data[3][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][30]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1260),
    .D(_00441_),
    .Q_N(_14907_),
    .Q(\cpu.dcache.r_data[3][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][31]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1261),
    .D(_00442_),
    .Q_N(_14906_),
    .Q(\cpu.dcache.r_data[3][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1262),
    .D(_00443_),
    .Q_N(_14905_),
    .Q(\cpu.dcache.r_data[3][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1263),
    .D(_00444_),
    .Q_N(_14904_),
    .Q(\cpu.dcache.r_data[3][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1264),
    .D(_00445_),
    .Q_N(_14903_),
    .Q(\cpu.dcache.r_data[3][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1265),
    .D(_00446_),
    .Q_N(_14902_),
    .Q(\cpu.dcache.r_data[3][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1266),
    .D(_00447_),
    .Q_N(_14901_),
    .Q(\cpu.dcache.r_data[3][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1267),
    .D(_00448_),
    .Q_N(_14900_),
    .Q(\cpu.dcache.r_data[3][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1268),
    .D(_00449_),
    .Q_N(_14899_),
    .Q(\cpu.dcache.r_data[3][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1269),
    .D(_00450_),
    .Q_N(_14898_),
    .Q(\cpu.dcache.r_data[4][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1270),
    .D(_00451_),
    .Q_N(_14897_),
    .Q(\cpu.dcache.r_data[4][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1271),
    .D(_00452_),
    .Q_N(_14896_),
    .Q(\cpu.dcache.r_data[4][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1272),
    .D(_00453_),
    .Q_N(_14895_),
    .Q(\cpu.dcache.r_data[4][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1273),
    .D(_00454_),
    .Q_N(_14894_),
    .Q(\cpu.dcache.r_data[4][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1274),
    .D(_00455_),
    .Q_N(_14893_),
    .Q(\cpu.dcache.r_data[4][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1275),
    .D(_00456_),
    .Q_N(_14892_),
    .Q(\cpu.dcache.r_data[4][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1276),
    .D(_00457_),
    .Q_N(_14891_),
    .Q(\cpu.dcache.r_data[4][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1277),
    .D(_00458_),
    .Q_N(_14890_),
    .Q(\cpu.dcache.r_data[4][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1278),
    .D(_00459_),
    .Q_N(_14889_),
    .Q(\cpu.dcache.r_data[4][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][19]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1279),
    .D(_00460_),
    .Q_N(_14888_),
    .Q(\cpu.dcache.r_data[4][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1280),
    .D(_00461_),
    .Q_N(_14887_),
    .Q(\cpu.dcache.r_data[4][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][20]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1281),
    .D(_00462_),
    .Q_N(_14886_),
    .Q(\cpu.dcache.r_data[4][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][21]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1282),
    .D(_00463_),
    .Q_N(_14885_),
    .Q(\cpu.dcache.r_data[4][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][22]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1283),
    .D(_00464_),
    .Q_N(_14884_),
    .Q(\cpu.dcache.r_data[4][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][23]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1284),
    .D(_00465_),
    .Q_N(_14883_),
    .Q(\cpu.dcache.r_data[4][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][24]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1285),
    .D(_00466_),
    .Q_N(_14882_),
    .Q(\cpu.dcache.r_data[4][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][25]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1286),
    .D(_00467_),
    .Q_N(_14881_),
    .Q(\cpu.dcache.r_data[4][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][26]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1287),
    .D(_00468_),
    .Q_N(_14880_),
    .Q(\cpu.dcache.r_data[4][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][27]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1288),
    .D(_00469_),
    .Q_N(_14879_),
    .Q(\cpu.dcache.r_data[4][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][28]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1289),
    .D(_00470_),
    .Q_N(_14878_),
    .Q(\cpu.dcache.r_data[4][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][29]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1290),
    .D(_00471_),
    .Q_N(_14877_),
    .Q(\cpu.dcache.r_data[4][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1291),
    .D(_00472_),
    .Q_N(_14876_),
    .Q(\cpu.dcache.r_data[4][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][30]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1292),
    .D(_00473_),
    .Q_N(_14875_),
    .Q(\cpu.dcache.r_data[4][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][31]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1293),
    .D(_00474_),
    .Q_N(_14874_),
    .Q(\cpu.dcache.r_data[4][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1294),
    .D(_00475_),
    .Q_N(_14873_),
    .Q(\cpu.dcache.r_data[4][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1295),
    .D(_00476_),
    .Q_N(_14872_),
    .Q(\cpu.dcache.r_data[4][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1296),
    .D(_00477_),
    .Q_N(_14871_),
    .Q(\cpu.dcache.r_data[4][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1297),
    .D(_00478_),
    .Q_N(_14870_),
    .Q(\cpu.dcache.r_data[4][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1298),
    .D(_00479_),
    .Q_N(_14869_),
    .Q(\cpu.dcache.r_data[4][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1299),
    .D(_00480_),
    .Q_N(_14868_),
    .Q(\cpu.dcache.r_data[4][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1300),
    .D(_00481_),
    .Q_N(_14867_),
    .Q(\cpu.dcache.r_data[4][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1301),
    .D(_00482_),
    .Q_N(_14866_),
    .Q(\cpu.dcache.r_data[5][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1302),
    .D(_00483_),
    .Q_N(_14865_),
    .Q(\cpu.dcache.r_data[5][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1303),
    .D(_00484_),
    .Q_N(_14864_),
    .Q(\cpu.dcache.r_data[5][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1304),
    .D(_00485_),
    .Q_N(_14863_),
    .Q(\cpu.dcache.r_data[5][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1305),
    .D(_00486_),
    .Q_N(_14862_),
    .Q(\cpu.dcache.r_data[5][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1306),
    .D(_00487_),
    .Q_N(_14861_),
    .Q(\cpu.dcache.r_data[5][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1307),
    .D(_00488_),
    .Q_N(_14860_),
    .Q(\cpu.dcache.r_data[5][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1308),
    .D(_00489_),
    .Q_N(_14859_),
    .Q(\cpu.dcache.r_data[5][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1309),
    .D(_00490_),
    .Q_N(_14858_),
    .Q(\cpu.dcache.r_data[5][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1310),
    .D(_00491_),
    .Q_N(_14857_),
    .Q(\cpu.dcache.r_data[5][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][19]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1311),
    .D(_00492_),
    .Q_N(_14856_),
    .Q(\cpu.dcache.r_data[5][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1312),
    .D(_00493_),
    .Q_N(_14855_),
    .Q(\cpu.dcache.r_data[5][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][20]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1313),
    .D(_00494_),
    .Q_N(_14854_),
    .Q(\cpu.dcache.r_data[5][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][21]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1314),
    .D(_00495_),
    .Q_N(_14853_),
    .Q(\cpu.dcache.r_data[5][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][22]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1315),
    .D(_00496_),
    .Q_N(_14852_),
    .Q(\cpu.dcache.r_data[5][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][23]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1316),
    .D(_00497_),
    .Q_N(_14851_),
    .Q(\cpu.dcache.r_data[5][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][24]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1317),
    .D(_00498_),
    .Q_N(_14850_),
    .Q(\cpu.dcache.r_data[5][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][25]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1318),
    .D(_00499_),
    .Q_N(_14849_),
    .Q(\cpu.dcache.r_data[5][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][26]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1319),
    .D(_00500_),
    .Q_N(_14848_),
    .Q(\cpu.dcache.r_data[5][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][27]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1320),
    .D(_00501_),
    .Q_N(_14847_),
    .Q(\cpu.dcache.r_data[5][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][28]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1321),
    .D(_00502_),
    .Q_N(_14846_),
    .Q(\cpu.dcache.r_data[5][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][29]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1322),
    .D(_00503_),
    .Q_N(_14845_),
    .Q(\cpu.dcache.r_data[5][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1323),
    .D(_00504_),
    .Q_N(_14844_),
    .Q(\cpu.dcache.r_data[5][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][30]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1324),
    .D(_00505_),
    .Q_N(_14843_),
    .Q(\cpu.dcache.r_data[5][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][31]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1325),
    .D(_00506_),
    .Q_N(_14842_),
    .Q(\cpu.dcache.r_data[5][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1326),
    .D(_00507_),
    .Q_N(_14841_),
    .Q(\cpu.dcache.r_data[5][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1327),
    .D(_00508_),
    .Q_N(_14840_),
    .Q(\cpu.dcache.r_data[5][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1328),
    .D(_00509_),
    .Q_N(_14839_),
    .Q(\cpu.dcache.r_data[5][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1329),
    .D(_00510_),
    .Q_N(_14838_),
    .Q(\cpu.dcache.r_data[5][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1330),
    .D(_00511_),
    .Q_N(_14837_),
    .Q(\cpu.dcache.r_data[5][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1331),
    .D(_00512_),
    .Q_N(_14836_),
    .Q(\cpu.dcache.r_data[5][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1332),
    .D(_00513_),
    .Q_N(_14835_),
    .Q(\cpu.dcache.r_data[5][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1333),
    .D(_00514_),
    .Q_N(_14834_),
    .Q(\cpu.dcache.r_data[6][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1334),
    .D(_00515_),
    .Q_N(_14833_),
    .Q(\cpu.dcache.r_data[6][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1335),
    .D(_00516_),
    .Q_N(_14832_),
    .Q(\cpu.dcache.r_data[6][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1336),
    .D(_00517_),
    .Q_N(_14831_),
    .Q(\cpu.dcache.r_data[6][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1337),
    .D(_00518_),
    .Q_N(_14830_),
    .Q(\cpu.dcache.r_data[6][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1338),
    .D(_00519_),
    .Q_N(_14829_),
    .Q(\cpu.dcache.r_data[6][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1339),
    .D(_00520_),
    .Q_N(_14828_),
    .Q(\cpu.dcache.r_data[6][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1340),
    .D(_00521_),
    .Q_N(_14827_),
    .Q(\cpu.dcache.r_data[6][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1341),
    .D(_00522_),
    .Q_N(_14826_),
    .Q(\cpu.dcache.r_data[6][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1342),
    .D(_00523_),
    .Q_N(_14825_),
    .Q(\cpu.dcache.r_data[6][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][19]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1343),
    .D(_00524_),
    .Q_N(_14824_),
    .Q(\cpu.dcache.r_data[6][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1344),
    .D(_00525_),
    .Q_N(_14823_),
    .Q(\cpu.dcache.r_data[6][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][20]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1345),
    .D(_00526_),
    .Q_N(_14822_),
    .Q(\cpu.dcache.r_data[6][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][21]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1346),
    .D(_00527_),
    .Q_N(_14821_),
    .Q(\cpu.dcache.r_data[6][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][22]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1347),
    .D(_00528_),
    .Q_N(_14820_),
    .Q(\cpu.dcache.r_data[6][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][23]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1348),
    .D(_00529_),
    .Q_N(_14819_),
    .Q(\cpu.dcache.r_data[6][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][24]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1349),
    .D(_00530_),
    .Q_N(_14818_),
    .Q(\cpu.dcache.r_data[6][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][25]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1350),
    .D(_00531_),
    .Q_N(_14817_),
    .Q(\cpu.dcache.r_data[6][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][26]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1351),
    .D(_00532_),
    .Q_N(_14816_),
    .Q(\cpu.dcache.r_data[6][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][27]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1352),
    .D(_00533_),
    .Q_N(_14815_),
    .Q(\cpu.dcache.r_data[6][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][28]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1353),
    .D(_00534_),
    .Q_N(_14814_),
    .Q(\cpu.dcache.r_data[6][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][29]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1354),
    .D(_00535_),
    .Q_N(_14813_),
    .Q(\cpu.dcache.r_data[6][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1355),
    .D(_00536_),
    .Q_N(_14812_),
    .Q(\cpu.dcache.r_data[6][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][30]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1356),
    .D(_00537_),
    .Q_N(_14811_),
    .Q(\cpu.dcache.r_data[6][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][31]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1357),
    .D(_00538_),
    .Q_N(_14810_),
    .Q(\cpu.dcache.r_data[6][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1358),
    .D(_00539_),
    .Q_N(_14809_),
    .Q(\cpu.dcache.r_data[6][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1359),
    .D(_00540_),
    .Q_N(_14808_),
    .Q(\cpu.dcache.r_data[6][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1360),
    .D(_00541_),
    .Q_N(_14807_),
    .Q(\cpu.dcache.r_data[6][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1361),
    .D(_00542_),
    .Q_N(_14806_),
    .Q(\cpu.dcache.r_data[6][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1362),
    .D(_00543_),
    .Q_N(_14805_),
    .Q(\cpu.dcache.r_data[6][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1363),
    .D(_00544_),
    .Q_N(_14804_),
    .Q(\cpu.dcache.r_data[6][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1364),
    .D(_00545_),
    .Q_N(_14803_),
    .Q(\cpu.dcache.r_data[6][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1365),
    .D(_00546_),
    .Q_N(_14802_),
    .Q(\cpu.dcache.r_data[7][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1366),
    .D(_00547_),
    .Q_N(_14801_),
    .Q(\cpu.dcache.r_data[7][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1367),
    .D(_00548_),
    .Q_N(_14800_),
    .Q(\cpu.dcache.r_data[7][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1368),
    .D(_00549_),
    .Q_N(_14799_),
    .Q(\cpu.dcache.r_data[7][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1369),
    .D(_00550_),
    .Q_N(_14798_),
    .Q(\cpu.dcache.r_data[7][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1370),
    .D(_00551_),
    .Q_N(_14797_),
    .Q(\cpu.dcache.r_data[7][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1371),
    .D(_00552_),
    .Q_N(_14796_),
    .Q(\cpu.dcache.r_data[7][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1372),
    .D(_00553_),
    .Q_N(_14795_),
    .Q(\cpu.dcache.r_data[7][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1373),
    .D(_00554_),
    .Q_N(_14794_),
    .Q(\cpu.dcache.r_data[7][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1374),
    .D(_00555_),
    .Q_N(_14793_),
    .Q(\cpu.dcache.r_data[7][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][19]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1375),
    .D(_00556_),
    .Q_N(_14792_),
    .Q(\cpu.dcache.r_data[7][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1376),
    .D(_00557_),
    .Q_N(_14791_),
    .Q(\cpu.dcache.r_data[7][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][20]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1377),
    .D(_00558_),
    .Q_N(_14790_),
    .Q(\cpu.dcache.r_data[7][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][21]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1378),
    .D(_00559_),
    .Q_N(_14789_),
    .Q(\cpu.dcache.r_data[7][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][22]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1379),
    .D(_00560_),
    .Q_N(_14788_),
    .Q(\cpu.dcache.r_data[7][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][23]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1380),
    .D(_00561_),
    .Q_N(_14787_),
    .Q(\cpu.dcache.r_data[7][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][24]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1381),
    .D(_00562_),
    .Q_N(_14786_),
    .Q(\cpu.dcache.r_data[7][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][25]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1382),
    .D(_00563_),
    .Q_N(_14785_),
    .Q(\cpu.dcache.r_data[7][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][26]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1383),
    .D(_00564_),
    .Q_N(_14784_),
    .Q(\cpu.dcache.r_data[7][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][27]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1384),
    .D(_00565_),
    .Q_N(_14783_),
    .Q(\cpu.dcache.r_data[7][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][28]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1385),
    .D(_00566_),
    .Q_N(_14782_),
    .Q(\cpu.dcache.r_data[7][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][29]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1386),
    .D(_00567_),
    .Q_N(_14781_),
    .Q(\cpu.dcache.r_data[7][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1387),
    .D(_00568_),
    .Q_N(_14780_),
    .Q(\cpu.dcache.r_data[7][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][30]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1388),
    .D(_00569_),
    .Q_N(_14779_),
    .Q(\cpu.dcache.r_data[7][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][31]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1389),
    .D(_00570_),
    .Q_N(_14778_),
    .Q(\cpu.dcache.r_data[7][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1390),
    .D(_00571_),
    .Q_N(_14777_),
    .Q(\cpu.dcache.r_data[7][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1391),
    .D(_00572_),
    .Q_N(_14776_),
    .Q(\cpu.dcache.r_data[7][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1392),
    .D(_00573_),
    .Q_N(_14775_),
    .Q(\cpu.dcache.r_data[7][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1393),
    .D(_00574_),
    .Q_N(_14774_),
    .Q(\cpu.dcache.r_data[7][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1394),
    .D(_00575_),
    .Q_N(_14773_),
    .Q(\cpu.dcache.r_data[7][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1395),
    .D(_00576_),
    .Q_N(_14772_),
    .Q(\cpu.dcache.r_data[7][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1396),
    .D(_00577_),
    .Q_N(_14771_),
    .Q(\cpu.dcache.r_data[7][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[0]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1397),
    .D(_00578_),
    .Q_N(_14770_),
    .Q(\cpu.dcache.r_dirty[0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[1]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1398),
    .D(_00579_),
    .Q_N(_14769_),
    .Q(\cpu.dcache.r_dirty[1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[2]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1399),
    .D(_00580_),
    .Q_N(_14768_),
    .Q(\cpu.dcache.r_dirty[2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[3]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1400),
    .D(_00581_),
    .Q_N(_14767_),
    .Q(\cpu.dcache.r_dirty[3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[4]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1401),
    .D(_00582_),
    .Q_N(_14766_),
    .Q(\cpu.dcache.r_dirty[4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[5]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1402),
    .D(_00583_),
    .Q_N(_14765_),
    .Q(\cpu.dcache.r_dirty[5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[6]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1403),
    .D(_00584_),
    .Q_N(_14764_),
    .Q(\cpu.dcache.r_dirty[6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[7]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1404),
    .D(_00585_),
    .Q_N(_14763_),
    .Q(\cpu.dcache.r_dirty[7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_offset[0]$_SDFF_PN0_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1405),
    .D(_00586_),
    .Q_N(_00315_),
    .Q(\cpu.dcache.r_offset[0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_offset[1]$_SDFF_PN0_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1406),
    .D(_00587_),
    .Q_N(_14762_),
    .Q(\cpu.dcache.r_offset[1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_offset[2]$_SDFF_PN0_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1407),
    .D(_00588_),
    .Q_N(_00276_),
    .Q(\cpu.dcache.r_offset[2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1408),
    .D(_00589_),
    .Q_N(_00230_),
    .Q(\cpu.dcache.r_tag[0][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1409),
    .D(_00590_),
    .Q_N(_00246_),
    .Q(\cpu.dcache.r_tag[0][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1410),
    .D(_00591_),
    .Q_N(_00247_),
    .Q(\cpu.dcache.r_tag[0][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1411),
    .D(_00592_),
    .Q_N(_00248_),
    .Q(\cpu.dcache.r_tag[0][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1412),
    .D(_00593_),
    .Q_N(_00249_),
    .Q(\cpu.dcache.r_tag[0][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1413),
    .D(_00594_),
    .Q_N(_00250_),
    .Q(\cpu.dcache.r_tag[0][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1414),
    .D(_00595_),
    .Q_N(_14761_),
    .Q(\cpu.dcache.r_tag[0][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1415),
    .D(_00596_),
    .Q_N(_14760_),
    .Q(\cpu.dcache.r_tag[0][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1416),
    .D(_00597_),
    .Q_N(_14759_),
    .Q(\cpu.dcache.r_tag[0][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1417),
    .D(_00598_),
    .Q_N(_00251_),
    .Q(\cpu.dcache.r_tag[0][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1418),
    .D(_00599_),
    .Q_N(_00232_),
    .Q(\cpu.dcache.r_tag[0][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1419),
    .D(_00600_),
    .Q_N(_00234_),
    .Q(\cpu.dcache.r_tag[0][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1420),
    .D(_00601_),
    .Q_N(_00236_),
    .Q(\cpu.dcache.r_tag[0][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1421),
    .D(_00602_),
    .Q_N(_00238_),
    .Q(\cpu.dcache.r_tag[0][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1422),
    .D(_00603_),
    .Q_N(_00240_),
    .Q(\cpu.dcache.r_tag[0][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1423),
    .D(_00604_),
    .Q_N(_00242_),
    .Q(\cpu.dcache.r_tag[0][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1424),
    .D(_00605_),
    .Q_N(_00243_),
    .Q(\cpu.dcache.r_tag[0][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1425),
    .D(_00606_),
    .Q_N(_00244_),
    .Q(\cpu.dcache.r_tag[0][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1426),
    .D(_00607_),
    .Q_N(_00245_),
    .Q(\cpu.dcache.r_tag[0][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1427),
    .D(_00608_),
    .Q_N(_14758_),
    .Q(\cpu.dcache.r_tag[1][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1428),
    .D(_00609_),
    .Q_N(_14757_),
    .Q(\cpu.dcache.r_tag[1][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1429),
    .D(_00610_),
    .Q_N(_14756_),
    .Q(\cpu.dcache.r_tag[1][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1430),
    .D(_00611_),
    .Q_N(_14755_),
    .Q(\cpu.dcache.r_tag[1][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1431),
    .D(_00612_),
    .Q_N(_14754_),
    .Q(\cpu.dcache.r_tag[1][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1432),
    .D(_00613_),
    .Q_N(_14753_),
    .Q(\cpu.dcache.r_tag[1][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1433),
    .D(_00614_),
    .Q_N(_14752_),
    .Q(\cpu.dcache.r_tag[1][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1434),
    .D(_00615_),
    .Q_N(_14751_),
    .Q(\cpu.dcache.r_tag[1][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1435),
    .D(_00616_),
    .Q_N(_14750_),
    .Q(\cpu.dcache.r_tag[1][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1436),
    .D(_00617_),
    .Q_N(_14749_),
    .Q(\cpu.dcache.r_tag[1][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1437),
    .D(_00618_),
    .Q_N(_14748_),
    .Q(\cpu.dcache.r_tag[1][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1438),
    .D(_00619_),
    .Q_N(_14747_),
    .Q(\cpu.dcache.r_tag[1][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1439),
    .D(_00620_),
    .Q_N(_14746_),
    .Q(\cpu.dcache.r_tag[1][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1440),
    .D(_00621_),
    .Q_N(_14745_),
    .Q(\cpu.dcache.r_tag[1][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1441),
    .D(_00622_),
    .Q_N(_14744_),
    .Q(\cpu.dcache.r_tag[1][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1442),
    .D(_00623_),
    .Q_N(_14743_),
    .Q(\cpu.dcache.r_tag[1][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1443),
    .D(_00624_),
    .Q_N(_14742_),
    .Q(\cpu.dcache.r_tag[1][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1444),
    .D(_00625_),
    .Q_N(_14741_),
    .Q(\cpu.dcache.r_tag[1][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1445),
    .D(_00626_),
    .Q_N(_14740_),
    .Q(\cpu.dcache.r_tag[1][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1446),
    .D(_00627_),
    .Q_N(_14739_),
    .Q(\cpu.dcache.r_tag[2][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1447),
    .D(_00628_),
    .Q_N(_14738_),
    .Q(\cpu.dcache.r_tag[2][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1448),
    .D(_00629_),
    .Q_N(_14737_),
    .Q(\cpu.dcache.r_tag[2][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1449),
    .D(_00630_),
    .Q_N(_14736_),
    .Q(\cpu.dcache.r_tag[2][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1450),
    .D(_00631_),
    .Q_N(_14735_),
    .Q(\cpu.dcache.r_tag[2][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1451),
    .D(_00632_),
    .Q_N(_14734_),
    .Q(\cpu.dcache.r_tag[2][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1452),
    .D(_00633_),
    .Q_N(_14733_),
    .Q(\cpu.dcache.r_tag[2][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1453),
    .D(_00634_),
    .Q_N(_14732_),
    .Q(\cpu.dcache.r_tag[2][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1454),
    .D(_00635_),
    .Q_N(_14731_),
    .Q(\cpu.dcache.r_tag[2][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1455),
    .D(_00636_),
    .Q_N(_14730_),
    .Q(\cpu.dcache.r_tag[2][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1456),
    .D(_00637_),
    .Q_N(_14729_),
    .Q(\cpu.dcache.r_tag[2][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1457),
    .D(_00638_),
    .Q_N(_14728_),
    .Q(\cpu.dcache.r_tag[2][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1458),
    .D(_00639_),
    .Q_N(_14727_),
    .Q(\cpu.dcache.r_tag[2][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1459),
    .D(_00640_),
    .Q_N(_14726_),
    .Q(\cpu.dcache.r_tag[2][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1460),
    .D(_00641_),
    .Q_N(_14725_),
    .Q(\cpu.dcache.r_tag[2][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1461),
    .D(_00642_),
    .Q_N(_14724_),
    .Q(\cpu.dcache.r_tag[2][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1462),
    .D(_00643_),
    .Q_N(_14723_),
    .Q(\cpu.dcache.r_tag[2][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1463),
    .D(_00644_),
    .Q_N(_14722_),
    .Q(\cpu.dcache.r_tag[2][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1464),
    .D(_00645_),
    .Q_N(_14721_),
    .Q(\cpu.dcache.r_tag[2][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1465),
    .D(_00646_),
    .Q_N(_14720_),
    .Q(\cpu.dcache.r_tag[3][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1466),
    .D(_00647_),
    .Q_N(_14719_),
    .Q(\cpu.dcache.r_tag[3][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1467),
    .D(_00648_),
    .Q_N(_14718_),
    .Q(\cpu.dcache.r_tag[3][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1468),
    .D(_00649_),
    .Q_N(_14717_),
    .Q(\cpu.dcache.r_tag[3][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1469),
    .D(_00650_),
    .Q_N(_14716_),
    .Q(\cpu.dcache.r_tag[3][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1470),
    .D(_00651_),
    .Q_N(_14715_),
    .Q(\cpu.dcache.r_tag[3][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1471),
    .D(_00652_),
    .Q_N(_14714_),
    .Q(\cpu.dcache.r_tag[3][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1472),
    .D(_00653_),
    .Q_N(_14713_),
    .Q(\cpu.dcache.r_tag[3][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1473),
    .D(_00654_),
    .Q_N(_14712_),
    .Q(\cpu.dcache.r_tag[3][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1474),
    .D(_00655_),
    .Q_N(_14711_),
    .Q(\cpu.dcache.r_tag[3][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1475),
    .D(_00656_),
    .Q_N(_14710_),
    .Q(\cpu.dcache.r_tag[3][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1476),
    .D(_00657_),
    .Q_N(_14709_),
    .Q(\cpu.dcache.r_tag[3][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1477),
    .D(_00658_),
    .Q_N(_14708_),
    .Q(\cpu.dcache.r_tag[3][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1478),
    .D(_00659_),
    .Q_N(_14707_),
    .Q(\cpu.dcache.r_tag[3][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1479),
    .D(_00660_),
    .Q_N(_14706_),
    .Q(\cpu.dcache.r_tag[3][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1480),
    .D(_00661_),
    .Q_N(_14705_),
    .Q(\cpu.dcache.r_tag[3][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1481),
    .D(_00662_),
    .Q_N(_14704_),
    .Q(\cpu.dcache.r_tag[3][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1482),
    .D(_00663_),
    .Q_N(_14703_),
    .Q(\cpu.dcache.r_tag[3][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1483),
    .D(_00664_),
    .Q_N(_14702_),
    .Q(\cpu.dcache.r_tag[3][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1484),
    .D(_00665_),
    .Q_N(_14701_),
    .Q(\cpu.dcache.r_tag[4][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1485),
    .D(_00666_),
    .Q_N(_14700_),
    .Q(\cpu.dcache.r_tag[4][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1486),
    .D(_00667_),
    .Q_N(_14699_),
    .Q(\cpu.dcache.r_tag[4][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1487),
    .D(_00668_),
    .Q_N(_14698_),
    .Q(\cpu.dcache.r_tag[4][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1488),
    .D(_00669_),
    .Q_N(_14697_),
    .Q(\cpu.dcache.r_tag[4][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1489),
    .D(_00670_),
    .Q_N(_14696_),
    .Q(\cpu.dcache.r_tag[4][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1490),
    .D(_00671_),
    .Q_N(_14695_),
    .Q(\cpu.dcache.r_tag[4][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1491),
    .D(_00672_),
    .Q_N(_14694_),
    .Q(\cpu.dcache.r_tag[4][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1492),
    .D(_00673_),
    .Q_N(_14693_),
    .Q(\cpu.dcache.r_tag[4][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1493),
    .D(_00674_),
    .Q_N(_14692_),
    .Q(\cpu.dcache.r_tag[4][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1494),
    .D(_00675_),
    .Q_N(_14691_),
    .Q(\cpu.dcache.r_tag[4][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1495),
    .D(_00676_),
    .Q_N(_14690_),
    .Q(\cpu.dcache.r_tag[4][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1496),
    .D(_00677_),
    .Q_N(_14689_),
    .Q(\cpu.dcache.r_tag[4][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1497),
    .D(_00678_),
    .Q_N(_14688_),
    .Q(\cpu.dcache.r_tag[4][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1498),
    .D(_00679_),
    .Q_N(_14687_),
    .Q(\cpu.dcache.r_tag[4][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1499),
    .D(_00680_),
    .Q_N(_14686_),
    .Q(\cpu.dcache.r_tag[4][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1500),
    .D(_00681_),
    .Q_N(_14685_),
    .Q(\cpu.dcache.r_tag[4][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1501),
    .D(_00682_),
    .Q_N(_14684_),
    .Q(\cpu.dcache.r_tag[4][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1502),
    .D(_00683_),
    .Q_N(_14683_),
    .Q(\cpu.dcache.r_tag[4][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1503),
    .D(_00684_),
    .Q_N(_14682_),
    .Q(\cpu.dcache.r_tag[5][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1504),
    .D(_00685_),
    .Q_N(_14681_),
    .Q(\cpu.dcache.r_tag[5][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1505),
    .D(_00686_),
    .Q_N(_14680_),
    .Q(\cpu.dcache.r_tag[5][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1506),
    .D(_00687_),
    .Q_N(_14679_),
    .Q(\cpu.dcache.r_tag[5][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1507),
    .D(_00688_),
    .Q_N(_14678_),
    .Q(\cpu.dcache.r_tag[5][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1508),
    .D(_00689_),
    .Q_N(_14677_),
    .Q(\cpu.dcache.r_tag[5][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1509),
    .D(_00690_),
    .Q_N(_14676_),
    .Q(\cpu.dcache.r_tag[5][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1510),
    .D(_00691_),
    .Q_N(_14675_),
    .Q(\cpu.dcache.r_tag[5][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1511),
    .D(_00692_),
    .Q_N(_14674_),
    .Q(\cpu.dcache.r_tag[5][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1512),
    .D(_00693_),
    .Q_N(_14673_),
    .Q(\cpu.dcache.r_tag[5][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1513),
    .D(_00694_),
    .Q_N(_14672_),
    .Q(\cpu.dcache.r_tag[5][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1514),
    .D(_00695_),
    .Q_N(_14671_),
    .Q(\cpu.dcache.r_tag[5][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1515),
    .D(_00696_),
    .Q_N(_14670_),
    .Q(\cpu.dcache.r_tag[5][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1516),
    .D(_00697_),
    .Q_N(_14669_),
    .Q(\cpu.dcache.r_tag[5][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1517),
    .D(_00698_),
    .Q_N(_14668_),
    .Q(\cpu.dcache.r_tag[5][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1518),
    .D(_00699_),
    .Q_N(_14667_),
    .Q(\cpu.dcache.r_tag[5][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1519),
    .D(_00700_),
    .Q_N(_14666_),
    .Q(\cpu.dcache.r_tag[5][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1520),
    .D(_00701_),
    .Q_N(_14665_),
    .Q(\cpu.dcache.r_tag[5][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1521),
    .D(_00702_),
    .Q_N(_14664_),
    .Q(\cpu.dcache.r_tag[5][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1522),
    .D(_00703_),
    .Q_N(_14663_),
    .Q(\cpu.dcache.r_tag[6][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1523),
    .D(_00704_),
    .Q_N(_14662_),
    .Q(\cpu.dcache.r_tag[6][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1524),
    .D(_00705_),
    .Q_N(_14661_),
    .Q(\cpu.dcache.r_tag[6][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1525),
    .D(_00706_),
    .Q_N(_14660_),
    .Q(\cpu.dcache.r_tag[6][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1526),
    .D(_00707_),
    .Q_N(_14659_),
    .Q(\cpu.dcache.r_tag[6][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1527),
    .D(_00708_),
    .Q_N(_14658_),
    .Q(\cpu.dcache.r_tag[6][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1528),
    .D(_00709_),
    .Q_N(_14657_),
    .Q(\cpu.dcache.r_tag[6][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1529),
    .D(_00710_),
    .Q_N(_14656_),
    .Q(\cpu.dcache.r_tag[6][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1530),
    .D(_00711_),
    .Q_N(_14655_),
    .Q(\cpu.dcache.r_tag[6][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1531),
    .D(_00712_),
    .Q_N(_14654_),
    .Q(\cpu.dcache.r_tag[6][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1532),
    .D(_00713_),
    .Q_N(_14653_),
    .Q(\cpu.dcache.r_tag[6][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1533),
    .D(_00714_),
    .Q_N(_14652_),
    .Q(\cpu.dcache.r_tag[6][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1534),
    .D(_00715_),
    .Q_N(_14651_),
    .Q(\cpu.dcache.r_tag[6][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1535),
    .D(_00716_),
    .Q_N(_14650_),
    .Q(\cpu.dcache.r_tag[6][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1536),
    .D(_00717_),
    .Q_N(_14649_),
    .Q(\cpu.dcache.r_tag[6][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1537),
    .D(_00718_),
    .Q_N(_14648_),
    .Q(\cpu.dcache.r_tag[6][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1538),
    .D(_00719_),
    .Q_N(_14647_),
    .Q(\cpu.dcache.r_tag[6][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1539),
    .D(_00720_),
    .Q_N(_14646_),
    .Q(\cpu.dcache.r_tag[6][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1540),
    .D(_00721_),
    .Q_N(_14645_),
    .Q(\cpu.dcache.r_tag[6][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1541),
    .D(_00722_),
    .Q_N(_14644_),
    .Q(\cpu.dcache.r_tag[7][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1542),
    .D(_00723_),
    .Q_N(_14643_),
    .Q(\cpu.dcache.r_tag[7][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1543),
    .D(_00724_),
    .Q_N(_14642_),
    .Q(\cpu.dcache.r_tag[7][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1544),
    .D(_00725_),
    .Q_N(_14641_),
    .Q(\cpu.dcache.r_tag[7][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1545),
    .D(_00726_),
    .Q_N(_14640_),
    .Q(\cpu.dcache.r_tag[7][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1546),
    .D(_00727_),
    .Q_N(_14639_),
    .Q(\cpu.dcache.r_tag[7][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1547),
    .D(_00728_),
    .Q_N(_14638_),
    .Q(\cpu.dcache.r_tag[7][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1548),
    .D(_00729_),
    .Q_N(_14637_),
    .Q(\cpu.dcache.r_tag[7][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1549),
    .D(_00730_),
    .Q_N(_14636_),
    .Q(\cpu.dcache.r_tag[7][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1550),
    .D(_00731_),
    .Q_N(_14635_),
    .Q(\cpu.dcache.r_tag[7][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1551),
    .D(_00732_),
    .Q_N(_14634_),
    .Q(\cpu.dcache.r_tag[7][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1552),
    .D(_00733_),
    .Q_N(_14633_),
    .Q(\cpu.dcache.r_tag[7][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1553),
    .D(_00734_),
    .Q_N(_14632_),
    .Q(\cpu.dcache.r_tag[7][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1554),
    .D(_00735_),
    .Q_N(_14631_),
    .Q(\cpu.dcache.r_tag[7][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1555),
    .D(_00736_),
    .Q_N(_14630_),
    .Q(\cpu.dcache.r_tag[7][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1556),
    .D(_00737_),
    .Q_N(_14629_),
    .Q(\cpu.dcache.r_tag[7][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1557),
    .D(_00738_),
    .Q_N(_14628_),
    .Q(\cpu.dcache.r_tag[7][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1558),
    .D(_00739_),
    .Q_N(_14627_),
    .Q(\cpu.dcache.r_tag[7][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1559),
    .D(_00740_),
    .Q_N(_14626_),
    .Q(\cpu.dcache.r_tag[7][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1560),
    .D(_00741_),
    .Q_N(_14625_),
    .Q(\cpu.dcache.r_valid[0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1561),
    .D(_00742_),
    .Q_N(_14624_),
    .Q(\cpu.dcache.r_valid[1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1562),
    .D(_00743_),
    .Q_N(_14623_),
    .Q(\cpu.dcache.r_valid[2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1563),
    .D(_00744_),
    .Q_N(_14622_),
    .Q(\cpu.dcache.r_valid[3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1564),
    .D(_00745_),
    .Q_N(_14621_),
    .Q(\cpu.dcache.r_valid[4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1565),
    .D(_00746_),
    .Q_N(_14620_),
    .Q(\cpu.dcache.r_valid[5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1566),
    .D(_00747_),
    .Q_N(_14619_),
    .Q(\cpu.dcache.r_valid[6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1567),
    .D(_00748_),
    .Q_N(_14618_),
    .Q(\cpu.dcache.r_valid[7] ));
 sg13g2_dfrbp_1 \cpu.dec.r_br$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1568),
    .D(_00749_),
    .Q_N(_14617_),
    .Q(\cpu.br ));
 sg13g2_dfrbp_1 \cpu.dec.r_cond[0]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1569),
    .D(_00750_),
    .Q_N(_00298_),
    .Q(\cpu.cond[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_cond[1]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1570),
    .D(_00751_),
    .Q_N(_14616_),
    .Q(\cpu.cond[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_cond[2]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1571),
    .D(_00752_),
    .Q_N(_00273_),
    .Q(\cpu.cond[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_div$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1572),
    .D(_00753_),
    .Q_N(_14615_),
    .Q(\cpu.dec.div ));
 sg13g2_dfrbp_1 \cpu.dec.r_flush_all$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1573),
    .D(_00754_),
    .Q_N(_14614_),
    .Q(\cpu.dec.do_flush_all ));
 sg13g2_dfrbp_1 \cpu.dec.r_flush_write$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1574),
    .D(_00755_),
    .Q_N(_14613_),
    .Q(\cpu.dec.do_flush_write ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[0]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1575),
    .D(_00756_),
    .Q_N(_14612_),
    .Q(\cpu.dec.imm[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[10]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1576),
    .D(_00757_),
    .Q_N(_14611_),
    .Q(\cpu.dec.imm[10] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[11]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1577),
    .D(_00758_),
    .Q_N(_14610_),
    .Q(\cpu.dec.imm[11] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[12]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1578),
    .D(_00759_),
    .Q_N(_14609_),
    .Q(\cpu.dec.imm[12] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[13]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1579),
    .D(_00760_),
    .Q_N(_14608_),
    .Q(\cpu.dec.imm[13] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[14]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1580),
    .D(_00761_),
    .Q_N(_14607_),
    .Q(\cpu.dec.imm[14] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[15]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1581),
    .D(_00762_),
    .Q_N(_14606_),
    .Q(\cpu.dec.imm[15] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[1]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1582),
    .D(_00763_),
    .Q_N(_14605_),
    .Q(\cpu.dec.imm[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[2]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1583),
    .D(_00764_),
    .Q_N(_14604_),
    .Q(\cpu.dec.imm[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[3]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1584),
    .D(_00765_),
    .Q_N(_14603_),
    .Q(\cpu.dec.imm[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[4]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1585),
    .D(_00766_),
    .Q_N(_14602_),
    .Q(\cpu.dec.imm[4] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[5]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1586),
    .D(_00767_),
    .Q_N(_14601_),
    .Q(\cpu.dec.imm[5] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[6]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1587),
    .D(_00768_),
    .Q_N(_14600_),
    .Q(\cpu.dec.imm[6] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[7]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1588),
    .D(_00769_),
    .Q_N(_14599_),
    .Q(\cpu.dec.imm[7] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[8]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1589),
    .D(_00770_),
    .Q_N(_14598_),
    .Q(\cpu.dec.imm[8] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[9]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1590),
    .D(_00771_),
    .Q_N(_14597_),
    .Q(\cpu.dec.imm[9] ));
 sg13g2_dfrbp_1 \cpu.dec.r_inv_mmu$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1591),
    .D(_00772_),
    .Q_N(_14596_),
    .Q(\cpu.dec.do_inv_mmu ));
 sg13g2_dfrbp_1 \cpu.dec.r_io$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1592),
    .D(_00773_),
    .Q_N(_14595_),
    .Q(\cpu.dec.io ));
 sg13g2_dfrbp_1 \cpu.dec.r_jmp$_SDFFCE_PP0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1593),
    .D(_00774_),
    .Q_N(_00258_),
    .Q(\cpu.dec.jmp ));
 sg13g2_dfrbp_1 \cpu.dec.r_load$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1594),
    .D(_00775_),
    .Q_N(_14594_),
    .Q(\cpu.dec.load ));
 sg13g2_dfrbp_1 \cpu.dec.r_mult$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1595),
    .D(_00776_),
    .Q_N(_14593_),
    .Q(\cpu.dec.mult ));
 sg13g2_dfrbp_1 \cpu.dec.r_needs_rs2$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1596),
    .D(_00777_),
    .Q_N(_15005_),
    .Q(\cpu.dec.needs_rs2 ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[10]$_DFF_P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1597),
    .D(_00011_),
    .Q_N(_15006_),
    .Q(\cpu.dec.r_op[10] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[1]$_DFF_P_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1598),
    .D(_00012_),
    .Q_N(_15007_),
    .Q(\cpu.dec.r_op[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[2]$_DFF_P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1599),
    .D(_00013_),
    .Q_N(_15008_),
    .Q(\cpu.dec.r_op[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[3]$_DFF_P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1600),
    .D(_00014_),
    .Q_N(_15009_),
    .Q(\cpu.dec.r_op[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[4]$_DFF_P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1601),
    .D(_00015_),
    .Q_N(_15010_),
    .Q(\cpu.dec.r_op[4] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[5]$_DFF_P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1602),
    .D(_00016_),
    .Q_N(_15011_),
    .Q(\cpu.dec.r_op[5] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[6]$_DFF_P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1603),
    .D(_00017_),
    .Q_N(_15012_),
    .Q(\cpu.dec.r_op[6] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[7]$_DFF_P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1604),
    .D(_00018_),
    .Q_N(_15013_),
    .Q(\cpu.dec.r_op[7] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[8]$_DFF_P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1605),
    .D(_00019_),
    .Q_N(_15014_),
    .Q(\cpu.dec.r_op[8] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[9]$_DFF_P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1606),
    .D(_00020_),
    .Q_N(_14592_),
    .Q(\cpu.dec.r_op[9] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[0]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1607),
    .D(_00778_),
    .Q_N(_14591_),
    .Q(\cpu.dec.r_rd[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[1]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1608),
    .D(_00779_),
    .Q_N(_14590_),
    .Q(\cpu.dec.r_rd[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[2]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1609),
    .D(_00780_),
    .Q_N(_14589_),
    .Q(\cpu.dec.r_rd[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[3]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1610),
    .D(_00781_),
    .Q_N(_15015_),
    .Q(\cpu.dec.r_rd[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_ready$_DFF_P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1611),
    .D(_00052_),
    .Q_N(_14588_),
    .Q(\cpu.dec.iready ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[0]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1612),
    .D(_00782_),
    .Q_N(_14587_),
    .Q(\cpu.dec.r_rs1[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[1]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1613),
    .D(_00783_),
    .Q_N(_14586_),
    .Q(\cpu.dec.r_rs1[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[2]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1614),
    .D(_00784_),
    .Q_N(_14585_),
    .Q(\cpu.dec.r_rs1[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[3]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1615),
    .D(_00785_),
    .Q_N(_14584_),
    .Q(\cpu.dec.r_rs1[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[0]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1616),
    .D(_00786_),
    .Q_N(_14583_),
    .Q(\cpu.dec.r_rs2[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[1]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1617),
    .D(_00787_),
    .Q_N(_14582_),
    .Q(\cpu.dec.r_rs2[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[2]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1618),
    .D(_00788_),
    .Q_N(_14581_),
    .Q(\cpu.dec.r_rs2[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[3]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1619),
    .D(_00789_),
    .Q_N(_14580_),
    .Q(\cpu.dec.r_rs2[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2_inv$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1620),
    .D(_00790_),
    .Q_N(_14579_),
    .Q(\cpu.dec.r_rs2_inv ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2_pc$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1621),
    .D(_00791_),
    .Q_N(_14578_),
    .Q(\cpu.dec.r_rs2_pc ));
 sg13g2_dfrbp_1 \cpu.dec.r_set_cc$_SDFFCE_PP0P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1622),
    .D(_00792_),
    .Q_N(_14577_),
    .Q(\cpu.dec.r_set_cc ));
 sg13g2_dfrbp_1 \cpu.dec.r_store$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1623),
    .D(_00793_),
    .Q_N(_00310_),
    .Q(\cpu.dec.r_store ));
 sg13g2_dfrbp_1 \cpu.dec.r_swapsp$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1624),
    .D(_00794_),
    .Q_N(_14576_),
    .Q(\cpu.dec.r_swapsp ));
 sg13g2_dfrbp_1 \cpu.dec.r_sys_call$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1625),
    .D(_00795_),
    .Q_N(_00274_),
    .Q(\cpu.dec.r_sys_call ));
 sg13g2_dfrbp_1 \cpu.dec.r_trap$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1626),
    .D(_00796_),
    .Q_N(_14575_),
    .Q(\cpu.dec.r_trap ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_mmu_d_proxy$_SDFFE_PP0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1627),
    .D(_00797_),
    .Q_N(_14574_),
    .Q(\cpu.ex.genblk3.r_mmu_d_proxy ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_mmu_enable$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1628),
    .D(_00798_),
    .Q_N(_00192_),
    .Q(\cpu.ex.genblk3.r_mmu_enable ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_prev_supmode$_SDFFE_PN1P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1629),
    .D(_00799_),
    .Q_N(_15016_),
    .Q(\cpu.ex.genblk3.r_prev_supmode ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_supmode$_DFF_P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1630),
    .D(\cpu.ex.genblk3.c_supmode ),
    .Q_N(_00193_),
    .Q(\cpu.dec.supmode ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_user_io$_SDFFE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1631),
    .D(_00800_),
    .Q_N(_14573_),
    .Q(\cpu.dec.user_io ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[0]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1632),
    .D(_00801_),
    .Q_N(_14572_),
    .Q(\cpu.ex.r_10[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[10]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1633),
    .D(_00802_),
    .Q_N(_14571_),
    .Q(\cpu.ex.r_10[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[11]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1634),
    .D(_00803_),
    .Q_N(_14570_),
    .Q(\cpu.ex.r_10[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[12]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1635),
    .D(_00804_),
    .Q_N(_14569_),
    .Q(\cpu.ex.r_10[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[13]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1636),
    .D(_00805_),
    .Q_N(_14568_),
    .Q(\cpu.ex.r_10[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[14]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1637),
    .D(_00806_),
    .Q_N(_14567_),
    .Q(\cpu.ex.r_10[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[15]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1638),
    .D(_00807_),
    .Q_N(_14566_),
    .Q(\cpu.ex.r_10[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[1]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1639),
    .D(_00808_),
    .Q_N(_14565_),
    .Q(\cpu.ex.r_10[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[2]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1640),
    .D(_00809_),
    .Q_N(_14564_),
    .Q(\cpu.ex.r_10[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[3]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1641),
    .D(_00810_),
    .Q_N(_14563_),
    .Q(\cpu.ex.r_10[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[4]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1642),
    .D(_00811_),
    .Q_N(_14562_),
    .Q(\cpu.ex.r_10[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[5]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1643),
    .D(_00812_),
    .Q_N(_14561_),
    .Q(\cpu.ex.r_10[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[6]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1644),
    .D(_00813_),
    .Q_N(_14560_),
    .Q(\cpu.ex.r_10[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[7]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1645),
    .D(_00814_),
    .Q_N(_14559_),
    .Q(\cpu.ex.r_10[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[8]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1646),
    .D(_00815_),
    .Q_N(_14558_),
    .Q(\cpu.ex.r_10[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[9]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1647),
    .D(_00816_),
    .Q_N(_14557_),
    .Q(\cpu.ex.r_10[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[0]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1648),
    .D(_00817_),
    .Q_N(_14556_),
    .Q(\cpu.ex.r_11[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[10]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1649),
    .D(_00818_),
    .Q_N(_14555_),
    .Q(\cpu.ex.r_11[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[11]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1650),
    .D(_00819_),
    .Q_N(_14554_),
    .Q(\cpu.ex.r_11[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[12]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1651),
    .D(_00820_),
    .Q_N(_14553_),
    .Q(\cpu.ex.r_11[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[13]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1652),
    .D(_00821_),
    .Q_N(_14552_),
    .Q(\cpu.ex.r_11[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[14]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1653),
    .D(_00822_),
    .Q_N(_14551_),
    .Q(\cpu.ex.r_11[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[15]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1654),
    .D(_00823_),
    .Q_N(_14550_),
    .Q(\cpu.ex.r_11[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[1]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1655),
    .D(_00824_),
    .Q_N(_14549_),
    .Q(\cpu.ex.r_11[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[2]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1656),
    .D(_00825_),
    .Q_N(_14548_),
    .Q(\cpu.ex.r_11[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[3]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1657),
    .D(_00826_),
    .Q_N(_14547_),
    .Q(\cpu.ex.r_11[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[4]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1658),
    .D(_00827_),
    .Q_N(_14546_),
    .Q(\cpu.ex.r_11[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[5]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1659),
    .D(_00828_),
    .Q_N(_14545_),
    .Q(\cpu.ex.r_11[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[6]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1660),
    .D(_00829_),
    .Q_N(_14544_),
    .Q(\cpu.ex.r_11[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[7]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1661),
    .D(_00830_),
    .Q_N(_14543_),
    .Q(\cpu.ex.r_11[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[8]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1662),
    .D(_00831_),
    .Q_N(_14542_),
    .Q(\cpu.ex.r_11[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[9]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1663),
    .D(_00832_),
    .Q_N(_14541_),
    .Q(\cpu.ex.r_11[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[0]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1664),
    .D(_00833_),
    .Q_N(_14540_),
    .Q(\cpu.ex.r_12[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[10]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1665),
    .D(_00834_),
    .Q_N(_14539_),
    .Q(\cpu.ex.r_12[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[11]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1666),
    .D(_00835_),
    .Q_N(_14538_),
    .Q(\cpu.ex.r_12[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[12]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1667),
    .D(_00836_),
    .Q_N(_14537_),
    .Q(\cpu.ex.r_12[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[13]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1668),
    .D(_00837_),
    .Q_N(_14536_),
    .Q(\cpu.ex.r_12[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[14]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1669),
    .D(_00838_),
    .Q_N(_14535_),
    .Q(\cpu.ex.r_12[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[15]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1670),
    .D(_00839_),
    .Q_N(_14534_),
    .Q(\cpu.ex.r_12[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[1]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1671),
    .D(_00840_),
    .Q_N(_14533_),
    .Q(\cpu.ex.r_12[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[2]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1672),
    .D(_00841_),
    .Q_N(_14532_),
    .Q(\cpu.ex.r_12[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[3]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1673),
    .D(_00842_),
    .Q_N(_14531_),
    .Q(\cpu.ex.r_12[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[4]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1674),
    .D(_00843_),
    .Q_N(_14530_),
    .Q(\cpu.ex.r_12[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[5]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1675),
    .D(_00844_),
    .Q_N(_14529_),
    .Q(\cpu.ex.r_12[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[6]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1676),
    .D(_00845_),
    .Q_N(_14528_),
    .Q(\cpu.ex.r_12[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[7]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1677),
    .D(_00846_),
    .Q_N(_14527_),
    .Q(\cpu.ex.r_12[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[8]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1678),
    .D(_00847_),
    .Q_N(_14526_),
    .Q(\cpu.ex.r_12[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[9]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1679),
    .D(_00848_),
    .Q_N(_14525_),
    .Q(\cpu.ex.r_12[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[0]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1680),
    .D(_00849_),
    .Q_N(_14524_),
    .Q(\cpu.ex.r_13[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[10]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1681),
    .D(_00850_),
    .Q_N(_14523_),
    .Q(\cpu.ex.r_13[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[11]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1682),
    .D(_00851_),
    .Q_N(_14522_),
    .Q(\cpu.ex.r_13[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[12]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1683),
    .D(_00852_),
    .Q_N(_14521_),
    .Q(\cpu.ex.r_13[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[13]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1684),
    .D(_00853_),
    .Q_N(_14520_),
    .Q(\cpu.ex.r_13[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[14]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1685),
    .D(_00854_),
    .Q_N(_14519_),
    .Q(\cpu.ex.r_13[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[15]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1686),
    .D(_00855_),
    .Q_N(_14518_),
    .Q(\cpu.ex.r_13[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[1]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1687),
    .D(_00856_),
    .Q_N(_14517_),
    .Q(\cpu.ex.r_13[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[2]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1688),
    .D(_00857_),
    .Q_N(_14516_),
    .Q(\cpu.ex.r_13[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[3]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1689),
    .D(_00858_),
    .Q_N(_14515_),
    .Q(\cpu.ex.r_13[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[4]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1690),
    .D(_00859_),
    .Q_N(_14514_),
    .Q(\cpu.ex.r_13[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[5]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1691),
    .D(_00860_),
    .Q_N(_14513_),
    .Q(\cpu.ex.r_13[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[6]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1692),
    .D(_00861_),
    .Q_N(_14512_),
    .Q(\cpu.ex.r_13[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[7]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1693),
    .D(_00862_),
    .Q_N(_14511_),
    .Q(\cpu.ex.r_13[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[8]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1694),
    .D(_00863_),
    .Q_N(_14510_),
    .Q(\cpu.ex.r_13[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[9]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1695),
    .D(_00864_),
    .Q_N(_14509_),
    .Q(\cpu.ex.r_13[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[0]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1696),
    .D(_00865_),
    .Q_N(_14508_),
    .Q(\cpu.ex.r_14[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[10]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1697),
    .D(_00866_),
    .Q_N(_14507_),
    .Q(\cpu.ex.r_14[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[11]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1698),
    .D(_00867_),
    .Q_N(_14506_),
    .Q(\cpu.ex.r_14[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[12]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1699),
    .D(_00868_),
    .Q_N(_14505_),
    .Q(\cpu.ex.r_14[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[13]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1700),
    .D(_00869_),
    .Q_N(_14504_),
    .Q(\cpu.ex.r_14[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[14]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1701),
    .D(_00870_),
    .Q_N(_14503_),
    .Q(\cpu.ex.r_14[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[15]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1702),
    .D(_00871_),
    .Q_N(_14502_),
    .Q(\cpu.ex.r_14[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[1]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1703),
    .D(_00872_),
    .Q_N(_14501_),
    .Q(\cpu.ex.r_14[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[2]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1704),
    .D(_00873_),
    .Q_N(_14500_),
    .Q(\cpu.ex.r_14[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[3]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1705),
    .D(_00874_),
    .Q_N(_14499_),
    .Q(\cpu.ex.r_14[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[4]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1706),
    .D(_00875_),
    .Q_N(_14498_),
    .Q(\cpu.ex.r_14[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[5]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1707),
    .D(_00876_),
    .Q_N(_14497_),
    .Q(\cpu.ex.r_14[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[6]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1708),
    .D(_00877_),
    .Q_N(_14496_),
    .Q(\cpu.ex.r_14[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[7]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1709),
    .D(_00878_),
    .Q_N(_14495_),
    .Q(\cpu.ex.r_14[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[8]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1710),
    .D(_00879_),
    .Q_N(_14494_),
    .Q(\cpu.ex.r_14[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[9]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1711),
    .D(_00880_),
    .Q_N(_14493_),
    .Q(\cpu.ex.r_14[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[0]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1712),
    .D(_00881_),
    .Q_N(_14492_),
    .Q(\cpu.ex.r_15[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[10]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1713),
    .D(_00882_),
    .Q_N(_00268_),
    .Q(\cpu.ex.r_15[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[11]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1714),
    .D(_00883_),
    .Q_N(_00269_),
    .Q(\cpu.ex.r_15[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[12]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1715),
    .D(_00884_),
    .Q_N(_00270_),
    .Q(\cpu.ex.r_15[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[13]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1716),
    .D(_00885_),
    .Q_N(_00271_),
    .Q(\cpu.ex.r_15[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[14]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1717),
    .D(_00886_),
    .Q_N(_00272_),
    .Q(\cpu.ex.r_15[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[15]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1718),
    .D(_00887_),
    .Q_N(_14491_),
    .Q(\cpu.ex.r_15[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[1]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1719),
    .D(_00888_),
    .Q_N(_00259_),
    .Q(\cpu.ex.r_15[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[2]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1720),
    .D(_00889_),
    .Q_N(_00260_),
    .Q(\cpu.ex.r_15[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[3]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1721),
    .D(_00890_),
    .Q_N(_00261_),
    .Q(\cpu.ex.r_15[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[4]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1722),
    .D(_00891_),
    .Q_N(_00262_),
    .Q(\cpu.ex.r_15[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[5]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1723),
    .D(_00892_),
    .Q_N(_00263_),
    .Q(\cpu.ex.r_15[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[6]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1724),
    .D(_00893_),
    .Q_N(_00264_),
    .Q(\cpu.ex.r_15[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[7]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1725),
    .D(_00894_),
    .Q_N(_00265_),
    .Q(\cpu.ex.r_15[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[8]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1726),
    .D(_00895_),
    .Q_N(_00266_),
    .Q(\cpu.ex.r_15[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[9]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1727),
    .D(_00896_),
    .Q_N(_00267_),
    .Q(\cpu.ex.r_15[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[0]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1728),
    .D(_00897_),
    .Q_N(_14490_),
    .Q(\cpu.ex.r_8[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[10]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1729),
    .D(_00898_),
    .Q_N(_14489_),
    .Q(\cpu.ex.r_8[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[11]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1730),
    .D(_00899_),
    .Q_N(_14488_),
    .Q(\cpu.ex.r_8[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[12]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1731),
    .D(_00900_),
    .Q_N(_14487_),
    .Q(\cpu.ex.r_8[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[13]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1732),
    .D(_00901_),
    .Q_N(_14486_),
    .Q(\cpu.ex.r_8[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[14]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1733),
    .D(_00902_),
    .Q_N(_14485_),
    .Q(\cpu.ex.r_8[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[15]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1734),
    .D(_00903_),
    .Q_N(_14484_),
    .Q(\cpu.ex.r_8[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[1]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1735),
    .D(_00904_),
    .Q_N(_14483_),
    .Q(\cpu.ex.r_8[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[2]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1736),
    .D(_00905_),
    .Q_N(_14482_),
    .Q(\cpu.ex.r_8[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[3]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1737),
    .D(_00906_),
    .Q_N(_14481_),
    .Q(\cpu.ex.r_8[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[4]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1738),
    .D(_00907_),
    .Q_N(_14480_),
    .Q(\cpu.ex.r_8[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[5]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1739),
    .D(_00908_),
    .Q_N(_14479_),
    .Q(\cpu.ex.r_8[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[6]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1740),
    .D(_00909_),
    .Q_N(_14478_),
    .Q(\cpu.ex.r_8[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[7]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1741),
    .D(_00910_),
    .Q_N(_14477_),
    .Q(\cpu.ex.r_8[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[8]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1742),
    .D(_00911_),
    .Q_N(_14476_),
    .Q(\cpu.ex.r_8[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[9]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1743),
    .D(_00912_),
    .Q_N(_14475_),
    .Q(\cpu.ex.r_8[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[0]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1744),
    .D(_00913_),
    .Q_N(_14474_),
    .Q(\cpu.ex.r_9[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[10]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1745),
    .D(_00914_),
    .Q_N(_14473_),
    .Q(\cpu.ex.r_9[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[11]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1746),
    .D(_00915_),
    .Q_N(_14472_),
    .Q(\cpu.ex.r_9[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[12]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1747),
    .D(_00916_),
    .Q_N(_14471_),
    .Q(\cpu.ex.r_9[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[13]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1748),
    .D(_00917_),
    .Q_N(_14470_),
    .Q(\cpu.ex.r_9[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[14]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1749),
    .D(_00918_),
    .Q_N(_14469_),
    .Q(\cpu.ex.r_9[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[15]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1750),
    .D(_00919_),
    .Q_N(_14468_),
    .Q(\cpu.ex.r_9[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[1]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1751),
    .D(_00920_),
    .Q_N(_14467_),
    .Q(\cpu.ex.r_9[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[2]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1752),
    .D(_00921_),
    .Q_N(_14466_),
    .Q(\cpu.ex.r_9[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[3]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1753),
    .D(_00922_),
    .Q_N(_14465_),
    .Q(\cpu.ex.r_9[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[4]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1754),
    .D(_00923_),
    .Q_N(_14464_),
    .Q(\cpu.ex.r_9[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[5]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1755),
    .D(_00924_),
    .Q_N(_14463_),
    .Q(\cpu.ex.r_9[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[6]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1756),
    .D(_00925_),
    .Q_N(_14462_),
    .Q(\cpu.ex.r_9[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[7]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1757),
    .D(_00926_),
    .Q_N(_14461_),
    .Q(\cpu.ex.r_9[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[8]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1758),
    .D(_00927_),
    .Q_N(_14460_),
    .Q(\cpu.ex.r_9[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[9]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1759),
    .D(_00928_),
    .Q_N(_15017_),
    .Q(\cpu.ex.r_9[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_branch_stall$_DFF_P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1760),
    .D(_00053_),
    .Q_N(_14459_),
    .Q(\cpu.ex.r_branch_stall ));
 sg13g2_dfrbp_1 \cpu.ex.r_cc$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1761),
    .D(_00929_),
    .Q_N(_14458_),
    .Q(\cpu.ex.r_cc ));
 sg13g2_dfrbp_1 \cpu.ex.r_d_flush_all$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1762),
    .D(_00930_),
    .Q_N(_15018_),
    .Q(\cpu.d_flush_all ));
 sg13g2_dfrbp_1 \cpu.ex.r_div_running$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1763),
    .D(\cpu.ex.c_div_running ),
    .Q_N(_14457_),
    .Q(\cpu.ex.r_div_running ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[0]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1764),
    .D(_00931_),
    .Q_N(_14456_),
    .Q(\cpu.ex.r_epc[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[10]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1765),
    .D(_00932_),
    .Q_N(_14455_),
    .Q(\cpu.ex.r_epc[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[11]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1766),
    .D(_00933_),
    .Q_N(_14454_),
    .Q(\cpu.ex.r_epc[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[12]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1767),
    .D(_00934_),
    .Q_N(_14453_),
    .Q(\cpu.ex.r_epc[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[13]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1768),
    .D(_00935_),
    .Q_N(_14452_),
    .Q(\cpu.ex.r_epc[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[14]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1769),
    .D(_00936_),
    .Q_N(_14451_),
    .Q(\cpu.ex.r_epc[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[1]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1770),
    .D(_00937_),
    .Q_N(_14450_),
    .Q(\cpu.ex.r_epc[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[2]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1771),
    .D(_00938_),
    .Q_N(_14449_),
    .Q(\cpu.ex.r_epc[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[3]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1772),
    .D(_00939_),
    .Q_N(_14448_),
    .Q(\cpu.ex.r_epc[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[4]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1773),
    .D(_00940_),
    .Q_N(_14447_),
    .Q(\cpu.ex.r_epc[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[5]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1774),
    .D(_00941_),
    .Q_N(_14446_),
    .Q(\cpu.ex.r_epc[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[6]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1775),
    .D(_00942_),
    .Q_N(_14445_),
    .Q(\cpu.ex.r_epc[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[7]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1776),
    .D(_00943_),
    .Q_N(_14444_),
    .Q(\cpu.ex.r_epc[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[8]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1777),
    .D(_00944_),
    .Q_N(_14443_),
    .Q(\cpu.ex.r_epc[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[9]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1778),
    .D(_00945_),
    .Q_N(_14442_),
    .Q(\cpu.ex.r_epc[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_fetch$_SDFF_PN1_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1779),
    .D(_00946_),
    .Q_N(_00189_),
    .Q(\cpu.ex.ifetch ));
 sg13g2_dfrbp_1 \cpu.ex.r_flush_write$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1780),
    .D(_00947_),
    .Q_N(_14441_),
    .Q(\cpu.dcache.flush_write ));
 sg13g2_dfrbp_1 \cpu.ex.r_i_flush_all$_SDFF_PP0_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1781),
    .D(_00948_),
    .Q_N(_14440_),
    .Q(\cpu.ex.i_flush_all ));
 sg13g2_dfrbp_1 \cpu.ex.r_ie$_SDFFE_PP0P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1782),
    .D(_00949_),
    .Q_N(_14439_),
    .Q(\cpu.ex.r_ie ));
 sg13g2_dfrbp_1 \cpu.ex.r_io_access$_SDFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1783),
    .D(_00950_),
    .Q_N(_00197_),
    .Q(\cpu.ex.io_access ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[0]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1784),
    .D(_00951_),
    .Q_N(_14438_),
    .Q(\cpu.ex.r_lr[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[10]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1785),
    .D(_00952_),
    .Q_N(_14437_),
    .Q(\cpu.ex.r_lr[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[11]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1786),
    .D(_00953_),
    .Q_N(_14436_),
    .Q(\cpu.ex.r_lr[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[12]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1787),
    .D(_00954_),
    .Q_N(_14435_),
    .Q(\cpu.ex.r_lr[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[13]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1788),
    .D(_00955_),
    .Q_N(_14434_),
    .Q(\cpu.ex.r_lr[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[14]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1789),
    .D(_00956_),
    .Q_N(_14433_),
    .Q(\cpu.ex.r_lr[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[1]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1790),
    .D(_00957_),
    .Q_N(_14432_),
    .Q(\cpu.ex.r_lr[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[2]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1791),
    .D(_00958_),
    .Q_N(_14431_),
    .Q(\cpu.ex.r_lr[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[3]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1792),
    .D(_00959_),
    .Q_N(_14430_),
    .Q(\cpu.ex.r_lr[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[4]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1793),
    .D(_00960_),
    .Q_N(_14429_),
    .Q(\cpu.ex.r_lr[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[5]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1794),
    .D(_00961_),
    .Q_N(_14428_),
    .Q(\cpu.ex.r_lr[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[6]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1795),
    .D(_00962_),
    .Q_N(_14427_),
    .Q(\cpu.ex.r_lr[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[7]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1796),
    .D(_00963_),
    .Q_N(_14426_),
    .Q(\cpu.ex.r_lr[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[8]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1797),
    .D(_00964_),
    .Q_N(_14425_),
    .Q(\cpu.ex.r_lr[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[9]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1798),
    .D(_00965_),
    .Q_N(_15019_),
    .Q(\cpu.ex.r_lr[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[0]$_DFF_P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1799),
    .D(\cpu.ex.c_mult[0] ),
    .Q_N(_15020_),
    .Q(\cpu.ex.r_mult[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[10]$_DFF_P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1800),
    .D(\cpu.ex.c_mult[10] ),
    .Q_N(_00167_),
    .Q(\cpu.ex.r_mult[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[11]$_DFF_P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1801),
    .D(\cpu.ex.c_mult[11] ),
    .Q_N(_00168_),
    .Q(\cpu.ex.r_mult[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[12]$_DFF_P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1802),
    .D(\cpu.ex.c_mult[12] ),
    .Q_N(_00169_),
    .Q(\cpu.ex.r_mult[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[13]$_DFF_P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1803),
    .D(\cpu.ex.c_mult[13] ),
    .Q_N(_00170_),
    .Q(\cpu.ex.r_mult[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[14]$_DFF_P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1804),
    .D(\cpu.ex.c_mult[14] ),
    .Q_N(_00171_),
    .Q(\cpu.ex.r_mult[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[15]$_DFF_P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1805),
    .D(\cpu.ex.c_mult[15] ),
    .Q_N(_14424_),
    .Q(\cpu.ex.r_mult[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[16]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1806),
    .D(_00966_),
    .Q_N(_00309_),
    .Q(\cpu.ex.r_mult[16] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[17]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1807),
    .D(_00967_),
    .Q_N(_00308_),
    .Q(\cpu.ex.r_mult[17] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[18]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1808),
    .D(_00968_),
    .Q_N(_00307_),
    .Q(\cpu.ex.r_mult[18] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[19]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1809),
    .D(_00969_),
    .Q_N(_00306_),
    .Q(\cpu.ex.r_mult[19] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[1]$_DFF_P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1810),
    .D(\cpu.ex.c_mult[1] ),
    .Q_N(_14423_),
    .Q(\cpu.ex.r_mult[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[20]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1811),
    .D(_00970_),
    .Q_N(_00305_),
    .Q(\cpu.ex.r_mult[20] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[21]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1812),
    .D(_00971_),
    .Q_N(_00304_),
    .Q(\cpu.ex.r_mult[21] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[22]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1813),
    .D(_00972_),
    .Q_N(_14422_),
    .Q(\cpu.ex.r_mult[22] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[23]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1814),
    .D(_00973_),
    .Q_N(_00303_),
    .Q(\cpu.ex.r_mult[23] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[24]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1815),
    .D(_00974_),
    .Q_N(_00302_),
    .Q(\cpu.ex.r_mult[24] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[25]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1816),
    .D(_00975_),
    .Q_N(_00301_),
    .Q(\cpu.ex.r_mult[25] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[26]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1817),
    .D(_00976_),
    .Q_N(_14421_),
    .Q(\cpu.ex.r_mult[26] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[27]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1818),
    .D(_00977_),
    .Q_N(_00300_),
    .Q(\cpu.ex.r_mult[27] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[28]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1819),
    .D(_00978_),
    .Q_N(_14420_),
    .Q(\cpu.ex.r_mult[28] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[29]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1820),
    .D(_00979_),
    .Q_N(_15021_),
    .Q(\cpu.ex.r_mult[29] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[2]$_DFF_P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1821),
    .D(\cpu.ex.c_mult[2] ),
    .Q_N(_00120_),
    .Q(\cpu.ex.r_mult[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[30]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1822),
    .D(_00980_),
    .Q_N(_00299_),
    .Q(\cpu.ex.r_mult[30] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[31]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1823),
    .D(_00981_),
    .Q_N(_15022_),
    .Q(\cpu.ex.r_mult[31] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[3]$_DFF_P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1824),
    .D(\cpu.ex.c_mult[3] ),
    .Q_N(_00127_),
    .Q(\cpu.ex.r_mult[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[4]$_DFF_P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1825),
    .D(\cpu.ex.c_mult[4] ),
    .Q_N(_00139_),
    .Q(\cpu.ex.r_mult[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[5]$_DFF_P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1826),
    .D(\cpu.ex.c_mult[5] ),
    .Q_N(_00151_),
    .Q(\cpu.ex.r_mult[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[6]$_DFF_P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1827),
    .D(\cpu.ex.c_mult[6] ),
    .Q_N(_00163_),
    .Q(\cpu.ex.r_mult[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[7]$_DFF_P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1828),
    .D(\cpu.ex.c_mult[7] ),
    .Q_N(_00164_),
    .Q(\cpu.ex.r_mult[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[8]$_DFF_P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1829),
    .D(\cpu.ex.c_mult[8] ),
    .Q_N(_00165_),
    .Q(\cpu.ex.r_mult[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[9]$_DFF_P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1830),
    .D(\cpu.ex.c_mult[9] ),
    .Q_N(_00166_),
    .Q(\cpu.ex.r_mult[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[0]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1831),
    .D(\cpu.ex.c_mult_off[0] ),
    .Q_N(_15023_),
    .Q(\cpu.ex.r_mult_off[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[1]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1832),
    .D(\cpu.ex.c_mult_off[1] ),
    .Q_N(_15024_),
    .Q(\cpu.ex.r_mult_off[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[2]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1833),
    .D(\cpu.ex.c_mult_off[2] ),
    .Q_N(_15025_),
    .Q(\cpu.ex.r_mult_off[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[3]$_DFF_P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1834),
    .D(\cpu.ex.c_mult_off[3] ),
    .Q_N(_15026_),
    .Q(\cpu.ex.r_mult_off[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_running$_DFF_P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1835),
    .D(\cpu.ex.c_mult_running ),
    .Q_N(_00199_),
    .Q(\cpu.ex.r_mult_running ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[0]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1836),
    .D(_00982_),
    .Q_N(_00200_),
    .Q(\cpu.ex.pc[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[10]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1837),
    .D(_00983_),
    .Q_N(_00290_),
    .Q(\cpu.ex.pc[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[11]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1838),
    .D(_00984_),
    .Q_N(_00289_),
    .Q(\cpu.ex.pc[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[12]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1839),
    .D(_00985_),
    .Q_N(_00196_),
    .Q(\cpu.ex.pc[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[13]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1840),
    .D(_00986_),
    .Q_N(_00195_),
    .Q(\cpu.ex.pc[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[14]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1841),
    .D(_00987_),
    .Q_N(_00194_),
    .Q(\cpu.ex.pc[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[1]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1842),
    .D(_00988_),
    .Q_N(_00297_),
    .Q(\cpu.ex.pc[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[2]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1843),
    .D(_00989_),
    .Q_N(_00191_),
    .Q(\cpu.ex.pc[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[3]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1844),
    .D(_00990_),
    .Q_N(_00190_),
    .Q(\cpu.ex.pc[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[4]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1845),
    .D(_00991_),
    .Q_N(_00296_),
    .Q(\cpu.ex.pc[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[5]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1846),
    .D(_00992_),
    .Q_N(_00295_),
    .Q(\cpu.ex.pc[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[6]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1847),
    .D(_00993_),
    .Q_N(_00294_),
    .Q(\cpu.ex.pc[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[7]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1848),
    .D(_00994_),
    .Q_N(_00293_),
    .Q(\cpu.ex.pc[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[8]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1849),
    .D(_00995_),
    .Q_N(_00292_),
    .Q(\cpu.ex.pc[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[9]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1850),
    .D(_00996_),
    .Q_N(_00291_),
    .Q(\cpu.ex.pc[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_prev_ie$_SDFFE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1851),
    .D(_00997_),
    .Q_N(_14419_),
    .Q(\cpu.ex.r_prev_ie ));
 sg13g2_dfrbp_1 \cpu.ex.r_read_stall$_SDFFE_PN0P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1852),
    .D(_00998_),
    .Q_N(_00198_),
    .Q(\cpu.ex.r_read_stall ));
 sg13g2_dfrbp_1 \cpu.ex.r_set_cc$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1853),
    .D(_00999_),
    .Q_N(_14418_),
    .Q(\cpu.ex.r_set_cc ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[0]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1854),
    .D(_01000_),
    .Q_N(_14417_),
    .Q(\cpu.ex.r_sp[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[10]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1855),
    .D(_01001_),
    .Q_N(_14416_),
    .Q(\cpu.ex.r_sp[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[11]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1856),
    .D(_01002_),
    .Q_N(_14415_),
    .Q(\cpu.ex.r_sp[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[12]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1857),
    .D(_01003_),
    .Q_N(_14414_),
    .Q(\cpu.ex.r_sp[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[13]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1858),
    .D(_01004_),
    .Q_N(_14413_),
    .Q(\cpu.ex.r_sp[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[14]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1859),
    .D(_01005_),
    .Q_N(_14412_),
    .Q(\cpu.ex.r_sp[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[1]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1860),
    .D(_01006_),
    .Q_N(_14411_),
    .Q(\cpu.ex.r_sp[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[2]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1861),
    .D(_01007_),
    .Q_N(_14410_),
    .Q(\cpu.ex.r_sp[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[3]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1862),
    .D(_01008_),
    .Q_N(_14409_),
    .Q(\cpu.ex.r_sp[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[4]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1863),
    .D(_01009_),
    .Q_N(_14408_),
    .Q(\cpu.ex.r_sp[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[5]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1864),
    .D(_01010_),
    .Q_N(_14407_),
    .Q(\cpu.ex.r_sp[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[6]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1865),
    .D(_01011_),
    .Q_N(_14406_),
    .Q(\cpu.ex.r_sp[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[7]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1866),
    .D(_01012_),
    .Q_N(_14405_),
    .Q(\cpu.ex.r_sp[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[8]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1867),
    .D(_01013_),
    .Q_N(_14404_),
    .Q(\cpu.ex.r_sp[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[9]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1868),
    .D(_01014_),
    .Q_N(_14403_),
    .Q(\cpu.ex.r_sp[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1869),
    .D(_01015_),
    .Q_N(_14402_),
    .Q(\cpu.ex.r_stmp[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[10]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1870),
    .D(_01016_),
    .Q_N(_14401_),
    .Q(\cpu.ex.r_stmp[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[11]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1871),
    .D(_01017_),
    .Q_N(_14400_),
    .Q(\cpu.ex.r_stmp[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[12]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1872),
    .D(_01018_),
    .Q_N(_14399_),
    .Q(\cpu.ex.r_stmp[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[13]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1873),
    .D(_01019_),
    .Q_N(_14398_),
    .Q(\cpu.ex.r_stmp[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[14]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1874),
    .D(_01020_),
    .Q_N(_14397_),
    .Q(\cpu.ex.r_stmp[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[15]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1875),
    .D(_01021_),
    .Q_N(_14396_),
    .Q(\cpu.ex.r_stmp[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[1]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1876),
    .D(_01022_),
    .Q_N(_14395_),
    .Q(\cpu.ex.r_stmp[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[2]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1877),
    .D(_01023_),
    .Q_N(_14394_),
    .Q(\cpu.ex.r_stmp[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[3]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1878),
    .D(_01024_),
    .Q_N(_14393_),
    .Q(\cpu.ex.r_stmp[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[4]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1879),
    .D(_01025_),
    .Q_N(_14392_),
    .Q(\cpu.ex.r_stmp[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[5]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1880),
    .D(_01026_),
    .Q_N(_14391_),
    .Q(\cpu.ex.r_stmp[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[6]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1881),
    .D(_01027_),
    .Q_N(_14390_),
    .Q(\cpu.ex.r_stmp[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[7]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1882),
    .D(_01028_),
    .Q_N(_14389_),
    .Q(\cpu.ex.r_stmp[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[8]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1883),
    .D(_01029_),
    .Q_N(_14388_),
    .Q(\cpu.ex.r_stmp[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[9]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1884),
    .D(_01030_),
    .Q_N(_14387_),
    .Q(\cpu.ex.r_stmp[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[0]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1885),
    .D(_01031_),
    .Q_N(_00257_),
    .Q(\cpu.ex.mmu_reg_data[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[10]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1886),
    .D(_01032_),
    .Q_N(_00239_),
    .Q(\cpu.addr[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[11]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1887),
    .D(_01033_),
    .Q_N(_00241_),
    .Q(\cpu.addr[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[12]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1888),
    .D(_01034_),
    .Q_N(_14386_),
    .Q(\cpu.addr[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[13]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1889),
    .D(_01035_),
    .Q_N(_14385_),
    .Q(\cpu.addr[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[14]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1890),
    .D(_01036_),
    .Q_N(_14384_),
    .Q(\cpu.addr[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[15]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1891),
    .D(_01037_),
    .Q_N(_14383_),
    .Q(\cpu.addr[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[1]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1892),
    .D(_01038_),
    .Q_N(_00275_),
    .Q(\cpu.addr[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[2]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1893),
    .D(_01039_),
    .Q_N(_14382_),
    .Q(\cpu.addr[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[3]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1894),
    .D(_01040_),
    .Q_N(_00228_),
    .Q(\cpu.addr[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[4]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1895),
    .D(_01041_),
    .Q_N(_00227_),
    .Q(\cpu.addr[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[5]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1896),
    .D(_01042_),
    .Q_N(_00229_),
    .Q(\cpu.addr[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[6]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1897),
    .D(_01043_),
    .Q_N(_00231_),
    .Q(\cpu.addr[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[7]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1898),
    .D(_01044_),
    .Q_N(_00233_),
    .Q(\cpu.addr[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[8]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1899),
    .D(_01045_),
    .Q_N(_00235_),
    .Q(\cpu.addr[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[9]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1900),
    .D(_01046_),
    .Q_N(_00237_),
    .Q(\cpu.addr[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1901),
    .D(_01047_),
    .Q_N(_14381_),
    .Q(\cpu.ex.r_wb_addr[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1902),
    .D(_01048_),
    .Q_N(_14380_),
    .Q(\cpu.ex.r_wb_addr[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[2]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1903),
    .D(_01049_),
    .Q_N(_14379_),
    .Q(\cpu.ex.r_wb_addr[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[3]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1904),
    .D(_01050_),
    .Q_N(_14378_),
    .Q(\cpu.ex.r_wb_addr[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_swapsp$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1905),
    .D(_01051_),
    .Q_N(_15027_),
    .Q(\cpu.ex.r_wb_swapsp ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_valid$_DFF_P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1906),
    .D(_00054_),
    .Q_N(_00256_),
    .Q(\cpu.ex.r_wb_valid ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[0]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1907),
    .D(_01052_),
    .Q_N(_00223_),
    .Q(\cpu.dcache.wdata[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[10]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1908),
    .D(_01053_),
    .Q_N(_14377_),
    .Q(\cpu.dcache.wdata[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[11]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1909),
    .D(_01054_),
    .Q_N(_14376_),
    .Q(\cpu.dcache.wdata[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[12]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1910),
    .D(_01055_),
    .Q_N(_14375_),
    .Q(\cpu.dcache.wdata[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[13]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1911),
    .D(_01056_),
    .Q_N(_14374_),
    .Q(\cpu.dcache.wdata[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[14]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1912),
    .D(_01057_),
    .Q_N(_14373_),
    .Q(\cpu.dcache.wdata[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[15]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1913),
    .D(_01058_),
    .Q_N(_14372_),
    .Q(\cpu.dcache.wdata[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[1]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1914),
    .D(_01059_),
    .Q_N(_00178_),
    .Q(\cpu.dcache.wdata[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[2]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1915),
    .D(_01060_),
    .Q_N(_00179_),
    .Q(\cpu.dcache.wdata[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[3]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1916),
    .D(_01061_),
    .Q_N(_00287_),
    .Q(\cpu.dcache.wdata[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[4]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1917),
    .D(_01062_),
    .Q_N(_00180_),
    .Q(\cpu.dcache.wdata[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[5]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1918),
    .D(_01063_),
    .Q_N(_00181_),
    .Q(\cpu.dcache.wdata[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[6]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1919),
    .D(_01064_),
    .Q_N(_00182_),
    .Q(\cpu.dcache.wdata[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[7]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1920),
    .D(_01065_),
    .Q_N(_00281_),
    .Q(\cpu.dcache.wdata[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[8]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1921),
    .D(_01066_),
    .Q_N(_14371_),
    .Q(\cpu.dcache.wdata[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[9]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1922),
    .D(_01067_),
    .Q_N(_14370_),
    .Q(\cpu.dcache.wdata[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wmask[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1923),
    .D(_01068_),
    .Q_N(_14369_),
    .Q(\cpu.ex.r_wmask[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wmask[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1924),
    .D(_01069_),
    .Q_N(_14368_),
    .Q(\cpu.ex.r_wmask[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[0]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1925),
    .D(_01070_),
    .Q_N(_00288_),
    .Q(\cpu.ex.mmu_read[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[1]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1926),
    .D(_01071_),
    .Q_N(_14367_),
    .Q(\cpu.ex.mmu_read[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[2]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1927),
    .D(_01072_),
    .Q_N(_00188_),
    .Q(\cpu.ex.mmu_read[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[3]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1928),
    .D(_01073_),
    .Q_N(_14366_),
    .Q(\cpu.ex.mmu_read[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_ins$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1929),
    .D(_01074_),
    .Q_N(_00255_),
    .Q(\cpu.ex.mmu_read[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_sup$_SDFFE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1930),
    .D(_01075_),
    .Q_N(_14365_),
    .Q(\cpu.ex.mmu_read[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_type$_SDFFE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1931),
    .D(_01076_),
    .Q_N(_14364_),
    .Q(\cpu.ex.mmu_read[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1932),
    .D(_01077_),
    .Q_N(_14363_),
    .Q(\cpu.genblk1.mmu.r_valid_d[0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1933),
    .D(_01078_),
    .Q_N(_14362_),
    .Q(\cpu.genblk1.mmu.r_valid_d[10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1934),
    .D(_01079_),
    .Q_N(_14361_),
    .Q(\cpu.genblk1.mmu.r_valid_d[11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1935),
    .D(_01080_),
    .Q_N(_14360_),
    .Q(\cpu.genblk1.mmu.r_valid_d[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1936),
    .D(_01081_),
    .Q_N(_14359_),
    .Q(\cpu.genblk1.mmu.r_valid_d[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1937),
    .D(_01082_),
    .Q_N(_14358_),
    .Q(\cpu.genblk1.mmu.r_valid_d[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1938),
    .D(_01083_),
    .Q_N(_14357_),
    .Q(\cpu.genblk1.mmu.r_valid_d[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1939),
    .D(_01084_),
    .Q_N(_14356_),
    .Q(\cpu.genblk1.mmu.r_valid_d[16] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1940),
    .D(_01085_),
    .Q_N(_14355_),
    .Q(\cpu.genblk1.mmu.r_valid_d[17] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1941),
    .D(_01086_),
    .Q_N(_14354_),
    .Q(\cpu.genblk1.mmu.r_valid_d[18] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1942),
    .D(_01087_),
    .Q_N(_14353_),
    .Q(\cpu.genblk1.mmu.r_valid_d[19] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1943),
    .D(_01088_),
    .Q_N(_14352_),
    .Q(\cpu.genblk1.mmu.r_valid_d[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1944),
    .D(_01089_),
    .Q_N(_14351_),
    .Q(\cpu.genblk1.mmu.r_valid_d[20] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1945),
    .D(_01090_),
    .Q_N(_14350_),
    .Q(\cpu.genblk1.mmu.r_valid_d[21] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1946),
    .D(_01091_),
    .Q_N(_14349_),
    .Q(\cpu.genblk1.mmu.r_valid_d[22] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1947),
    .D(_01092_),
    .Q_N(_14348_),
    .Q(\cpu.genblk1.mmu.r_valid_d[23] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1948),
    .D(_01093_),
    .Q_N(_14347_),
    .Q(\cpu.genblk1.mmu.r_valid_d[24] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1949),
    .D(_01094_),
    .Q_N(_14346_),
    .Q(\cpu.genblk1.mmu.r_valid_d[25] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1950),
    .D(_01095_),
    .Q_N(_14345_),
    .Q(\cpu.genblk1.mmu.r_valid_d[26] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1951),
    .D(_01096_),
    .Q_N(_14344_),
    .Q(\cpu.genblk1.mmu.r_valid_d[27] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1952),
    .D(_01097_),
    .Q_N(_14343_),
    .Q(\cpu.genblk1.mmu.r_valid_d[28] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1953),
    .D(_01098_),
    .Q_N(_14342_),
    .Q(\cpu.genblk1.mmu.r_valid_d[29] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1954),
    .D(_01099_),
    .Q_N(_14341_),
    .Q(\cpu.genblk1.mmu.r_valid_d[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1955),
    .D(_01100_),
    .Q_N(_14340_),
    .Q(\cpu.genblk1.mmu.r_valid_d[30] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1956),
    .D(_01101_),
    .Q_N(_14339_),
    .Q(\cpu.genblk1.mmu.r_valid_d[31] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1957),
    .D(_01102_),
    .Q_N(_14338_),
    .Q(\cpu.genblk1.mmu.r_valid_d[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1958),
    .D(_01103_),
    .Q_N(_14337_),
    .Q(\cpu.genblk1.mmu.r_valid_d[4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1959),
    .D(_01104_),
    .Q_N(_14336_),
    .Q(\cpu.genblk1.mmu.r_valid_d[5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1960),
    .D(_01105_),
    .Q_N(_14335_),
    .Q(\cpu.genblk1.mmu.r_valid_d[6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1961),
    .D(_01106_),
    .Q_N(_14334_),
    .Q(\cpu.genblk1.mmu.r_valid_d[7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1962),
    .D(_01107_),
    .Q_N(_14333_),
    .Q(\cpu.genblk1.mmu.r_valid_d[8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1963),
    .D(_01108_),
    .Q_N(_14332_),
    .Q(\cpu.genblk1.mmu.r_valid_d[9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1964),
    .D(_01109_),
    .Q_N(_14331_),
    .Q(\cpu.genblk1.mmu.r_valid_i[0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1965),
    .D(_01110_),
    .Q_N(_14330_),
    .Q(\cpu.genblk1.mmu.r_valid_i[10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1966),
    .D(_01111_),
    .Q_N(_14329_),
    .Q(\cpu.genblk1.mmu.r_valid_i[11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1967),
    .D(_01112_),
    .Q_N(_14328_),
    .Q(\cpu.genblk1.mmu.r_valid_i[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1968),
    .D(_01113_),
    .Q_N(_14327_),
    .Q(\cpu.genblk1.mmu.r_valid_i[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1969),
    .D(_01114_),
    .Q_N(_14326_),
    .Q(\cpu.genblk1.mmu.r_valid_i[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1970),
    .D(_01115_),
    .Q_N(_14325_),
    .Q(\cpu.genblk1.mmu.r_valid_i[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1971),
    .D(_01116_),
    .Q_N(_14324_),
    .Q(\cpu.genblk1.mmu.r_valid_i[16] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1972),
    .D(_01117_),
    .Q_N(_14323_),
    .Q(\cpu.genblk1.mmu.r_valid_i[17] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1973),
    .D(_01118_),
    .Q_N(_14322_),
    .Q(\cpu.genblk1.mmu.r_valid_i[18] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1974),
    .D(_01119_),
    .Q_N(_14321_),
    .Q(\cpu.genblk1.mmu.r_valid_i[19] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1975),
    .D(_01120_),
    .Q_N(_14320_),
    .Q(\cpu.genblk1.mmu.r_valid_i[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1976),
    .D(_01121_),
    .Q_N(_14319_),
    .Q(\cpu.genblk1.mmu.r_valid_i[20] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1977),
    .D(_01122_),
    .Q_N(_14318_),
    .Q(\cpu.genblk1.mmu.r_valid_i[21] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1978),
    .D(_01123_),
    .Q_N(_14317_),
    .Q(\cpu.genblk1.mmu.r_valid_i[22] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1979),
    .D(_01124_),
    .Q_N(_14316_),
    .Q(\cpu.genblk1.mmu.r_valid_i[23] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1980),
    .D(_01125_),
    .Q_N(_14315_),
    .Q(\cpu.genblk1.mmu.r_valid_i[24] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1981),
    .D(_01126_),
    .Q_N(_14314_),
    .Q(\cpu.genblk1.mmu.r_valid_i[25] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1982),
    .D(_01127_),
    .Q_N(_14313_),
    .Q(\cpu.genblk1.mmu.r_valid_i[26] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1983),
    .D(_01128_),
    .Q_N(_14312_),
    .Q(\cpu.genblk1.mmu.r_valid_i[27] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1984),
    .D(_01129_),
    .Q_N(_14311_),
    .Q(\cpu.genblk1.mmu.r_valid_i[28] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1985),
    .D(_01130_),
    .Q_N(_14310_),
    .Q(\cpu.genblk1.mmu.r_valid_i[29] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1986),
    .D(_01131_),
    .Q_N(_14309_),
    .Q(\cpu.genblk1.mmu.r_valid_i[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1987),
    .D(_01132_),
    .Q_N(_14308_),
    .Q(\cpu.genblk1.mmu.r_valid_i[30] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1988),
    .D(_01133_),
    .Q_N(_14307_),
    .Q(\cpu.genblk1.mmu.r_valid_i[31] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1989),
    .D(_01134_),
    .Q_N(_14306_),
    .Q(\cpu.genblk1.mmu.r_valid_i[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1990),
    .D(_01135_),
    .Q_N(_14305_),
    .Q(\cpu.genblk1.mmu.r_valid_i[4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1991),
    .D(_01136_),
    .Q_N(_14304_),
    .Q(\cpu.genblk1.mmu.r_valid_i[5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1992),
    .D(_01137_),
    .Q_N(_14303_),
    .Q(\cpu.genblk1.mmu.r_valid_i[6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1993),
    .D(_01138_),
    .Q_N(_14302_),
    .Q(\cpu.genblk1.mmu.r_valid_i[7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1994),
    .D(_01139_),
    .Q_N(_14301_),
    .Q(\cpu.genblk1.mmu.r_valid_i[8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1995),
    .D(_01140_),
    .Q_N(_14300_),
    .Q(\cpu.genblk1.mmu.r_valid_i[9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1996),
    .D(_01141_),
    .Q_N(_14299_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1997),
    .D(_01142_),
    .Q_N(_14298_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1998),
    .D(_01143_),
    .Q_N(_14297_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1999),
    .D(_01144_),
    .Q_N(_14296_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2000),
    .D(_01145_),
    .Q_N(_14295_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2001),
    .D(_01146_),
    .Q_N(_14294_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2002),
    .D(_01147_),
    .Q_N(_14293_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2003),
    .D(_01148_),
    .Q_N(_14292_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2004),
    .D(_01149_),
    .Q_N(_14291_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2005),
    .D(_01150_),
    .Q_N(_14290_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2006),
    .D(_01151_),
    .Q_N(_14289_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2007),
    .D(_01152_),
    .Q_N(_14288_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][0]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2008),
    .D(_01153_),
    .Q_N(_14287_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][10]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2009),
    .D(_01154_),
    .Q_N(_14286_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][11]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2010),
    .D(_01155_),
    .Q_N(_14285_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][1]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2011),
    .D(_01156_),
    .Q_N(_14284_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][2]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2012),
    .D(_01157_),
    .Q_N(_14283_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][3]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2013),
    .D(_01158_),
    .Q_N(_14282_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][4]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2014),
    .D(_01159_),
    .Q_N(_14281_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][5]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2015),
    .D(_01160_),
    .Q_N(_14280_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][6]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2016),
    .D(_01161_),
    .Q_N(_14279_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][7]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2017),
    .D(_01162_),
    .Q_N(_14278_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][8]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2018),
    .D(_01163_),
    .Q_N(_14277_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][9]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2019),
    .D(_01164_),
    .Q_N(_14276_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][0]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2020),
    .D(_01165_),
    .Q_N(_14275_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][10]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2021),
    .D(_01166_),
    .Q_N(_14274_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][11]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2022),
    .D(_01167_),
    .Q_N(_14273_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][1]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2023),
    .D(_01168_),
    .Q_N(_14272_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][2]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2024),
    .D(_01169_),
    .Q_N(_14271_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][3]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2025),
    .D(_01170_),
    .Q_N(_14270_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][4]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2026),
    .D(_01171_),
    .Q_N(_14269_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][5]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2027),
    .D(_01172_),
    .Q_N(_14268_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][6]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2028),
    .D(_01173_),
    .Q_N(_14267_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][7]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2029),
    .D(_01174_),
    .Q_N(_14266_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][8]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2030),
    .D(_01175_),
    .Q_N(_14265_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][9]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2031),
    .D(_01176_),
    .Q_N(_14264_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][0]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2032),
    .D(_01177_),
    .Q_N(_14263_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][10]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2033),
    .D(_01178_),
    .Q_N(_14262_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][11]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2034),
    .D(_01179_),
    .Q_N(_14261_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][1]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2035),
    .D(_01180_),
    .Q_N(_14260_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][2]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2036),
    .D(_01181_),
    .Q_N(_14259_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][3]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2037),
    .D(_01182_),
    .Q_N(_14258_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][4]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2038),
    .D(_01183_),
    .Q_N(_14257_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][5]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2039),
    .D(_01184_),
    .Q_N(_14256_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][6]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2040),
    .D(_01185_),
    .Q_N(_14255_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][7]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2041),
    .D(_01186_),
    .Q_N(_14254_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][8]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2042),
    .D(_01187_),
    .Q_N(_14253_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][9]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2043),
    .D(_01188_),
    .Q_N(_14252_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][0]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2044),
    .D(_01189_),
    .Q_N(_14251_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][10]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2045),
    .D(_01190_),
    .Q_N(_14250_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][11]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2046),
    .D(_01191_),
    .Q_N(_14249_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][1]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2047),
    .D(_01192_),
    .Q_N(_14248_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][2]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2048),
    .D(_01193_),
    .Q_N(_14247_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][3]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2049),
    .D(_01194_),
    .Q_N(_14246_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][4]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2050),
    .D(_01195_),
    .Q_N(_14245_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][5]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2051),
    .D(_01196_),
    .Q_N(_14244_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][6]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2052),
    .D(_01197_),
    .Q_N(_14243_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][7]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2053),
    .D(_01198_),
    .Q_N(_14242_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][8]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2054),
    .D(_01199_),
    .Q_N(_14241_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][9]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2055),
    .D(_01200_),
    .Q_N(_14240_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][0]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2056),
    .D(_01201_),
    .Q_N(_14239_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][10]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2057),
    .D(_01202_),
    .Q_N(_14238_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][11]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2058),
    .D(_01203_),
    .Q_N(_14237_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][1]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2059),
    .D(_01204_),
    .Q_N(_14236_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][2]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2060),
    .D(_01205_),
    .Q_N(_14235_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][3]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2061),
    .D(_01206_),
    .Q_N(_14234_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][4]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2062),
    .D(_01207_),
    .Q_N(_14233_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][5]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2063),
    .D(_01208_),
    .Q_N(_14232_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][6]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2064),
    .D(_01209_),
    .Q_N(_14231_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][7]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2065),
    .D(_01210_),
    .Q_N(_14230_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][8]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2066),
    .D(_01211_),
    .Q_N(_14229_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][9]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2067),
    .D(_01212_),
    .Q_N(_14228_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][0]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2068),
    .D(_01213_),
    .Q_N(_14227_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][10]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2069),
    .D(_01214_),
    .Q_N(_14226_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][11]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2070),
    .D(_01215_),
    .Q_N(_14225_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][1]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2071),
    .D(_01216_),
    .Q_N(_14224_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][2]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2072),
    .D(_01217_),
    .Q_N(_14223_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][3]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2073),
    .D(_01218_),
    .Q_N(_14222_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][4]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2074),
    .D(_01219_),
    .Q_N(_14221_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][5]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2075),
    .D(_01220_),
    .Q_N(_14220_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][6]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2076),
    .D(_01221_),
    .Q_N(_14219_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][7]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2077),
    .D(_01222_),
    .Q_N(_14218_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][8]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2078),
    .D(_01223_),
    .Q_N(_14217_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][9]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2079),
    .D(_01224_),
    .Q_N(_14216_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][0]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2080),
    .D(_01225_),
    .Q_N(_14215_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][10]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2081),
    .D(_01226_),
    .Q_N(_14214_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][11]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2082),
    .D(_01227_),
    .Q_N(_14213_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][1]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2083),
    .D(_01228_),
    .Q_N(_14212_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][2]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2084),
    .D(_01229_),
    .Q_N(_14211_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][3]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2085),
    .D(_01230_),
    .Q_N(_14210_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][4]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2086),
    .D(_01231_),
    .Q_N(_14209_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][5]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2087),
    .D(_01232_),
    .Q_N(_14208_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][6]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2088),
    .D(_01233_),
    .Q_N(_14207_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][7]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2089),
    .D(_01234_),
    .Q_N(_14206_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][8]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2090),
    .D(_01235_),
    .Q_N(_14205_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][9]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2091),
    .D(_01236_),
    .Q_N(_14204_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][0]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2092),
    .D(_01237_),
    .Q_N(_14203_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][10]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2093),
    .D(_01238_),
    .Q_N(_14202_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][11]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2094),
    .D(_01239_),
    .Q_N(_14201_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][1]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2095),
    .D(_01240_),
    .Q_N(_14200_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][2]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2096),
    .D(_01241_),
    .Q_N(_14199_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][3]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2097),
    .D(_01242_),
    .Q_N(_14198_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][4]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2098),
    .D(_01243_),
    .Q_N(_14197_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][5]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2099),
    .D(_01244_),
    .Q_N(_14196_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][6]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2100),
    .D(_01245_),
    .Q_N(_14195_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][7]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2101),
    .D(_01246_),
    .Q_N(_14194_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][8]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2102),
    .D(_01247_),
    .Q_N(_14193_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][9]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2103),
    .D(_01248_),
    .Q_N(_14192_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][0]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2104),
    .D(_01249_),
    .Q_N(_14191_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][10]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2105),
    .D(_01250_),
    .Q_N(_14190_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][11]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2106),
    .D(_01251_),
    .Q_N(_14189_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][1]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2107),
    .D(_01252_),
    .Q_N(_14188_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][2]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2108),
    .D(_01253_),
    .Q_N(_14187_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][3]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2109),
    .D(_01254_),
    .Q_N(_14186_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][4]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2110),
    .D(_01255_),
    .Q_N(_14185_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][5]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2111),
    .D(_01256_),
    .Q_N(_14184_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][6]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2112),
    .D(_01257_),
    .Q_N(_14183_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][7]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2113),
    .D(_01258_),
    .Q_N(_14182_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][8]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2114),
    .D(_01259_),
    .Q_N(_14181_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][9]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2115),
    .D(_01260_),
    .Q_N(_14180_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][0]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2116),
    .D(_01261_),
    .Q_N(_14179_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][10]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2117),
    .D(_01262_),
    .Q_N(_14178_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][11]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2118),
    .D(_01263_),
    .Q_N(_14177_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][1]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2119),
    .D(_01264_),
    .Q_N(_14176_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][2]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2120),
    .D(_01265_),
    .Q_N(_14175_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][3]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2121),
    .D(_01266_),
    .Q_N(_14174_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][4]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2122),
    .D(_01267_),
    .Q_N(_14173_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][5]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2123),
    .D(_01268_),
    .Q_N(_14172_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][6]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2124),
    .D(_01269_),
    .Q_N(_14171_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][7]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2125),
    .D(_01270_),
    .Q_N(_14170_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][8]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2126),
    .D(_01271_),
    .Q_N(_14169_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][9]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2127),
    .D(_01272_),
    .Q_N(_14168_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2128),
    .D(_01273_),
    .Q_N(_14167_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2129),
    .D(_01274_),
    .Q_N(_14166_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2130),
    .D(_01275_),
    .Q_N(_14165_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2131),
    .D(_01276_),
    .Q_N(_14164_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2132),
    .D(_01277_),
    .Q_N(_14163_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2133),
    .D(_01278_),
    .Q_N(_14162_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2134),
    .D(_01279_),
    .Q_N(_14161_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2135),
    .D(_01280_),
    .Q_N(_14160_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2136),
    .D(_01281_),
    .Q_N(_14159_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2137),
    .D(_01282_),
    .Q_N(_14158_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2138),
    .D(_01283_),
    .Q_N(_14157_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2139),
    .D(_01284_),
    .Q_N(_14156_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][0]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2140),
    .D(_01285_),
    .Q_N(_14155_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][10]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2141),
    .D(_01286_),
    .Q_N(_14154_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][11]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2142),
    .D(_01287_),
    .Q_N(_14153_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][1]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2143),
    .D(_01288_),
    .Q_N(_14152_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][2]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2144),
    .D(_01289_),
    .Q_N(_14151_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][3]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2145),
    .D(_01290_),
    .Q_N(_14150_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][4]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2146),
    .D(_01291_),
    .Q_N(_14149_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][5]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2147),
    .D(_01292_),
    .Q_N(_14148_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][6]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2148),
    .D(_01293_),
    .Q_N(_14147_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][7]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2149),
    .D(_01294_),
    .Q_N(_14146_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][8]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2150),
    .D(_01295_),
    .Q_N(_14145_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][9]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2151),
    .D(_01296_),
    .Q_N(_14144_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][0]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2152),
    .D(_01297_),
    .Q_N(_14143_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][10]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2153),
    .D(_01298_),
    .Q_N(_14142_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][11]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2154),
    .D(_01299_),
    .Q_N(_14141_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][1]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2155),
    .D(_01300_),
    .Q_N(_14140_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][2]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2156),
    .D(_01301_),
    .Q_N(_14139_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][3]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2157),
    .D(_01302_),
    .Q_N(_14138_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][4]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2158),
    .D(_01303_),
    .Q_N(_14137_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][5]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2159),
    .D(_01304_),
    .Q_N(_14136_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][6]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2160),
    .D(_01305_),
    .Q_N(_14135_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][7]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2161),
    .D(_01306_),
    .Q_N(_14134_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][8]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2162),
    .D(_01307_),
    .Q_N(_14133_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][9]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2163),
    .D(_01308_),
    .Q_N(_14132_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][0]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2164),
    .D(_01309_),
    .Q_N(_14131_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][10]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2165),
    .D(_01310_),
    .Q_N(_14130_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][11]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2166),
    .D(_01311_),
    .Q_N(_14129_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][1]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2167),
    .D(_01312_),
    .Q_N(_14128_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][2]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2168),
    .D(_01313_),
    .Q_N(_14127_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][3]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2169),
    .D(_01314_),
    .Q_N(_14126_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][4]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2170),
    .D(_01315_),
    .Q_N(_14125_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][5]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2171),
    .D(_01316_),
    .Q_N(_14124_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][6]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2172),
    .D(_01317_),
    .Q_N(_14123_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][7]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2173),
    .D(_01318_),
    .Q_N(_14122_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][8]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2174),
    .D(_01319_),
    .Q_N(_14121_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][9]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2175),
    .D(_01320_),
    .Q_N(_14120_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][0]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2176),
    .D(_01321_),
    .Q_N(_14119_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][10]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2177),
    .D(_01322_),
    .Q_N(_14118_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][11]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2178),
    .D(_01323_),
    .Q_N(_14117_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][1]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2179),
    .D(_01324_),
    .Q_N(_14116_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][2]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2180),
    .D(_01325_),
    .Q_N(_14115_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][3]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2181),
    .D(_01326_),
    .Q_N(_14114_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][4]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2182),
    .D(_01327_),
    .Q_N(_14113_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][5]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2183),
    .D(_01328_),
    .Q_N(_14112_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][6]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2184),
    .D(_01329_),
    .Q_N(_14111_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][7]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2185),
    .D(_01330_),
    .Q_N(_14110_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][8]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2186),
    .D(_01331_),
    .Q_N(_14109_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][9]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2187),
    .D(_01332_),
    .Q_N(_14108_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][0]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2188),
    .D(_01333_),
    .Q_N(_14107_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][10]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2189),
    .D(_01334_),
    .Q_N(_14106_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][11]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2190),
    .D(_01335_),
    .Q_N(_14105_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][1]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2191),
    .D(_01336_),
    .Q_N(_14104_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][2]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2192),
    .D(_01337_),
    .Q_N(_14103_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][3]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2193),
    .D(_01338_),
    .Q_N(_14102_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][4]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2194),
    .D(_01339_),
    .Q_N(_14101_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][5]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2195),
    .D(_01340_),
    .Q_N(_14100_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][6]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2196),
    .D(_01341_),
    .Q_N(_14099_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][7]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2197),
    .D(_01342_),
    .Q_N(_14098_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][8]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2198),
    .D(_01343_),
    .Q_N(_14097_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][9]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2199),
    .D(_01344_),
    .Q_N(_14096_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][0]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2200),
    .D(_01345_),
    .Q_N(_14095_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][10]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2201),
    .D(_01346_),
    .Q_N(_14094_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][11]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2202),
    .D(_01347_),
    .Q_N(_14093_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][1]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2203),
    .D(_01348_),
    .Q_N(_14092_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][2]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2204),
    .D(_01349_),
    .Q_N(_14091_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][3]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2205),
    .D(_01350_),
    .Q_N(_14090_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][4]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2206),
    .D(_01351_),
    .Q_N(_14089_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][5]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2207),
    .D(_01352_),
    .Q_N(_14088_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][6]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2208),
    .D(_01353_),
    .Q_N(_14087_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][7]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2209),
    .D(_01354_),
    .Q_N(_14086_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][8]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2210),
    .D(_01355_),
    .Q_N(_14085_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][9]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2211),
    .D(_01356_),
    .Q_N(_14084_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][0]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2212),
    .D(_01357_),
    .Q_N(_14083_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][10]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2213),
    .D(_01358_),
    .Q_N(_14082_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][11]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2214),
    .D(_01359_),
    .Q_N(_14081_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][1]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2215),
    .D(_01360_),
    .Q_N(_14080_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][2]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2216),
    .D(_01361_),
    .Q_N(_14079_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][3]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2217),
    .D(_01362_),
    .Q_N(_14078_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][4]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2218),
    .D(_01363_),
    .Q_N(_14077_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][5]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2219),
    .D(_01364_),
    .Q_N(_14076_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][6]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2220),
    .D(_01365_),
    .Q_N(_14075_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][7]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2221),
    .D(_01366_),
    .Q_N(_14074_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][8]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2222),
    .D(_01367_),
    .Q_N(_14073_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][9]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2223),
    .D(_01368_),
    .Q_N(_14072_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][0]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2224),
    .D(_01369_),
    .Q_N(_14071_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][10]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2225),
    .D(_01370_),
    .Q_N(_14070_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][11]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2226),
    .D(_01371_),
    .Q_N(_14069_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][1]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2227),
    .D(_01372_),
    .Q_N(_14068_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][2]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2228),
    .D(_01373_),
    .Q_N(_14067_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][3]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2229),
    .D(_01374_),
    .Q_N(_14066_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][4]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2230),
    .D(_01375_),
    .Q_N(_14065_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][5]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2231),
    .D(_01376_),
    .Q_N(_14064_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][6]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2232),
    .D(_01377_),
    .Q_N(_14063_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][7]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2233),
    .D(_01378_),
    .Q_N(_14062_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][8]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2234),
    .D(_01379_),
    .Q_N(_14061_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][9]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2235),
    .D(_01380_),
    .Q_N(_14060_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][0]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2236),
    .D(_01381_),
    .Q_N(_14059_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][10]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2237),
    .D(_01382_),
    .Q_N(_14058_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][11]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2238),
    .D(_01383_),
    .Q_N(_14057_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][1]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2239),
    .D(_01384_),
    .Q_N(_14056_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][2]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2240),
    .D(_01385_),
    .Q_N(_14055_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][3]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2241),
    .D(_01386_),
    .Q_N(_14054_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][4]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2242),
    .D(_01387_),
    .Q_N(_14053_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][5]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2243),
    .D(_01388_),
    .Q_N(_14052_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][6]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2244),
    .D(_01389_),
    .Q_N(_14051_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][7]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2245),
    .D(_01390_),
    .Q_N(_14050_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][8]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2246),
    .D(_01391_),
    .Q_N(_14049_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][9]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2247),
    .D(_01392_),
    .Q_N(_14048_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][0]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2248),
    .D(_01393_),
    .Q_N(_14047_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][10]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2249),
    .D(_01394_),
    .Q_N(_14046_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][11]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2250),
    .D(_01395_),
    .Q_N(_14045_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][1]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2251),
    .D(_01396_),
    .Q_N(_14044_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][2]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2252),
    .D(_01397_),
    .Q_N(_14043_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][3]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2253),
    .D(_01398_),
    .Q_N(_14042_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][4]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2254),
    .D(_01399_),
    .Q_N(_14041_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][5]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2255),
    .D(_01400_),
    .Q_N(_14040_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][6]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2256),
    .D(_01401_),
    .Q_N(_14039_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][7]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2257),
    .D(_01402_),
    .Q_N(_14038_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][8]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2258),
    .D(_01403_),
    .Q_N(_14037_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][9]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2259),
    .D(_01404_),
    .Q_N(_14036_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2260),
    .D(_01405_),
    .Q_N(_14035_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2261),
    .D(_01406_),
    .Q_N(_14034_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2262),
    .D(_01407_),
    .Q_N(_14033_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2263),
    .D(_01408_),
    .Q_N(_14032_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2264),
    .D(_01409_),
    .Q_N(_14031_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2265),
    .D(_01410_),
    .Q_N(_14030_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2266),
    .D(_01411_),
    .Q_N(_14029_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2267),
    .D(_01412_),
    .Q_N(_14028_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2268),
    .D(_01413_),
    .Q_N(_14027_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2269),
    .D(_01414_),
    .Q_N(_14026_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2270),
    .D(_01415_),
    .Q_N(_14025_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2271),
    .D(_01416_),
    .Q_N(_14024_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][0]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2272),
    .D(_01417_),
    .Q_N(_14023_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][10]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2273),
    .D(_01418_),
    .Q_N(_14022_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][11]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2274),
    .D(_01419_),
    .Q_N(_14021_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][1]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2275),
    .D(_01420_),
    .Q_N(_14020_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][2]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2276),
    .D(_01421_),
    .Q_N(_14019_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][3]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2277),
    .D(_01422_),
    .Q_N(_14018_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][4]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2278),
    .D(_01423_),
    .Q_N(_14017_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][5]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2279),
    .D(_01424_),
    .Q_N(_14016_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][6]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2280),
    .D(_01425_),
    .Q_N(_14015_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][7]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2281),
    .D(_01426_),
    .Q_N(_14014_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][8]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2282),
    .D(_01427_),
    .Q_N(_14013_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][9]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2283),
    .D(_01428_),
    .Q_N(_14012_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][0]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2284),
    .D(_01429_),
    .Q_N(_14011_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][10]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2285),
    .D(_01430_),
    .Q_N(_14010_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][11]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2286),
    .D(_01431_),
    .Q_N(_14009_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][1]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2287),
    .D(_01432_),
    .Q_N(_14008_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][2]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2288),
    .D(_01433_),
    .Q_N(_14007_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][3]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2289),
    .D(_01434_),
    .Q_N(_14006_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][4]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2290),
    .D(_01435_),
    .Q_N(_14005_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][5]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2291),
    .D(_01436_),
    .Q_N(_14004_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][6]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2292),
    .D(_01437_),
    .Q_N(_14003_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][7]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2293),
    .D(_01438_),
    .Q_N(_14002_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][8]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2294),
    .D(_01439_),
    .Q_N(_14001_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][9]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2295),
    .D(_01440_),
    .Q_N(_14000_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2296),
    .D(_01441_),
    .Q_N(_13999_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2297),
    .D(_01442_),
    .Q_N(_13998_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2298),
    .D(_01443_),
    .Q_N(_13997_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2299),
    .D(_01444_),
    .Q_N(_13996_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2300),
    .D(_01445_),
    .Q_N(_13995_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2301),
    .D(_01446_),
    .Q_N(_13994_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2302),
    .D(_01447_),
    .Q_N(_13993_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2303),
    .D(_01448_),
    .Q_N(_13992_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2304),
    .D(_01449_),
    .Q_N(_13991_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2305),
    .D(_01450_),
    .Q_N(_13990_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2306),
    .D(_01451_),
    .Q_N(_13989_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2307),
    .D(_01452_),
    .Q_N(_13988_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2308),
    .D(_01453_),
    .Q_N(_13987_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2309),
    .D(_01454_),
    .Q_N(_13986_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2310),
    .D(_01455_),
    .Q_N(_13985_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2311),
    .D(_01456_),
    .Q_N(_13984_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2312),
    .D(_01457_),
    .Q_N(_13983_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2313),
    .D(_01458_),
    .Q_N(_13982_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2314),
    .D(_01459_),
    .Q_N(_13981_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2315),
    .D(_01460_),
    .Q_N(_13980_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2316),
    .D(_01461_),
    .Q_N(_13979_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2317),
    .D(_01462_),
    .Q_N(_13978_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2318),
    .D(_01463_),
    .Q_N(_13977_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2319),
    .D(_01464_),
    .Q_N(_13976_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2320),
    .D(_01465_),
    .Q_N(_13975_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2321),
    .D(_01466_),
    .Q_N(_13974_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2322),
    .D(_01467_),
    .Q_N(_13973_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2323),
    .D(_01468_),
    .Q_N(_13972_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2324),
    .D(_01469_),
    .Q_N(_13971_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2325),
    .D(_01470_),
    .Q_N(_13970_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2326),
    .D(_01471_),
    .Q_N(_13969_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2327),
    .D(_01472_),
    .Q_N(_13968_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2328),
    .D(_01473_),
    .Q_N(_13967_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2329),
    .D(_01474_),
    .Q_N(_13966_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2330),
    .D(_01475_),
    .Q_N(_13965_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2331),
    .D(_01476_),
    .Q_N(_13964_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2332),
    .D(_01477_),
    .Q_N(_13963_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2333),
    .D(_01478_),
    .Q_N(_13962_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2334),
    .D(_01479_),
    .Q_N(_13961_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2335),
    .D(_01480_),
    .Q_N(_13960_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2336),
    .D(_01481_),
    .Q_N(_13959_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2337),
    .D(_01482_),
    .Q_N(_13958_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2338),
    .D(_01483_),
    .Q_N(_13957_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2339),
    .D(_01484_),
    .Q_N(_13956_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2340),
    .D(_01485_),
    .Q_N(_13955_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2341),
    .D(_01486_),
    .Q_N(_13954_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2342),
    .D(_01487_),
    .Q_N(_13953_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2343),
    .D(_01488_),
    .Q_N(_13952_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2344),
    .D(_01489_),
    .Q_N(_13951_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2345),
    .D(_01490_),
    .Q_N(_13950_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2346),
    .D(_01491_),
    .Q_N(_13949_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2347),
    .D(_01492_),
    .Q_N(_13948_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2348),
    .D(_01493_),
    .Q_N(_13947_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2349),
    .D(_01494_),
    .Q_N(_13946_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2350),
    .D(_01495_),
    .Q_N(_13945_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2351),
    .D(_01496_),
    .Q_N(_13944_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2352),
    .D(_01497_),
    .Q_N(_13943_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2353),
    .D(_01498_),
    .Q_N(_13942_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2354),
    .D(_01499_),
    .Q_N(_13941_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2355),
    .D(_01500_),
    .Q_N(_13940_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][0]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2356),
    .D(_01501_),
    .Q_N(_13939_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][10]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2357),
    .D(_01502_),
    .Q_N(_13938_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][11]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2358),
    .D(_01503_),
    .Q_N(_13937_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][1]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2359),
    .D(_01504_),
    .Q_N(_13936_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][2]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2360),
    .D(_01505_),
    .Q_N(_13935_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][3]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2361),
    .D(_01506_),
    .Q_N(_13934_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][4]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net2362),
    .D(_01507_),
    .Q_N(_13933_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][5]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2363),
    .D(_01508_),
    .Q_N(_13932_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][6]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2364),
    .D(_01509_),
    .Q_N(_13931_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][7]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2365),
    .D(_01510_),
    .Q_N(_13930_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][8]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2366),
    .D(_01511_),
    .Q_N(_13929_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][9]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2367),
    .D(_01512_),
    .Q_N(_13928_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][0]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2368),
    .D(_01513_),
    .Q_N(_13927_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][10]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2369),
    .D(_01514_),
    .Q_N(_13926_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][11]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2370),
    .D(_01515_),
    .Q_N(_13925_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][1]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2371),
    .D(_01516_),
    .Q_N(_13924_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][2]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2372),
    .D(_01517_),
    .Q_N(_13923_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][3]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2373),
    .D(_01518_),
    .Q_N(_13922_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][4]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2374),
    .D(_01519_),
    .Q_N(_13921_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][5]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2375),
    .D(_01520_),
    .Q_N(_13920_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][6]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2376),
    .D(_01521_),
    .Q_N(_13919_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][7]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2377),
    .D(_01522_),
    .Q_N(_13918_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][8]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2378),
    .D(_01523_),
    .Q_N(_13917_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][9]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2379),
    .D(_01524_),
    .Q_N(_13916_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2380),
    .D(_01525_),
    .Q_N(_13915_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2381),
    .D(_01526_),
    .Q_N(_13914_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2382),
    .D(_01527_),
    .Q_N(_13913_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2383),
    .D(_01528_),
    .Q_N(_13912_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2384),
    .D(_01529_),
    .Q_N(_13911_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2385),
    .D(_01530_),
    .Q_N(_13910_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2386),
    .D(_01531_),
    .Q_N(_13909_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2387),
    .D(_01532_),
    .Q_N(_13908_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2388),
    .D(_01533_),
    .Q_N(_13907_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2389),
    .D(_01534_),
    .Q_N(_13906_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2390),
    .D(_01535_),
    .Q_N(_13905_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2391),
    .D(_01536_),
    .Q_N(_13904_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][0]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2392),
    .D(_01537_),
    .Q_N(_13903_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][10]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2393),
    .D(_01538_),
    .Q_N(_13902_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][11]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2394),
    .D(_01539_),
    .Q_N(_13901_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][1]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2395),
    .D(_01540_),
    .Q_N(_13900_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][2]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2396),
    .D(_01541_),
    .Q_N(_13899_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][3]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2397),
    .D(_01542_),
    .Q_N(_13898_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][4]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2398),
    .D(_01543_),
    .Q_N(_13897_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][5]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2399),
    .D(_01544_),
    .Q_N(_13896_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][6]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net2400),
    .D(_01545_),
    .Q_N(_13895_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][7]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2401),
    .D(_01546_),
    .Q_N(_13894_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][8]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2402),
    .D(_01547_),
    .Q_N(_13893_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][9]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2403),
    .D(_01548_),
    .Q_N(_13892_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][0]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2404),
    .D(_01549_),
    .Q_N(_13891_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][10]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2405),
    .D(_01550_),
    .Q_N(_13890_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][11]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2406),
    .D(_01551_),
    .Q_N(_13889_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][1]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2407),
    .D(_01552_),
    .Q_N(_13888_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][2]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2408),
    .D(_01553_),
    .Q_N(_13887_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][3]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2409),
    .D(_01554_),
    .Q_N(_13886_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][4]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2410),
    .D(_01555_),
    .Q_N(_13885_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][5]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2411),
    .D(_01556_),
    .Q_N(_13884_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][6]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2412),
    .D(_01557_),
    .Q_N(_13883_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][7]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2413),
    .D(_01558_),
    .Q_N(_13882_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][8]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2414),
    .D(_01559_),
    .Q_N(_13881_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][9]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2415),
    .D(_01560_),
    .Q_N(_13880_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][0]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2416),
    .D(_01561_),
    .Q_N(_13879_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][10]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2417),
    .D(_01562_),
    .Q_N(_13878_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][11]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2418),
    .D(_01563_),
    .Q_N(_13877_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][1]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2419),
    .D(_01564_),
    .Q_N(_13876_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][2]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2420),
    .D(_01565_),
    .Q_N(_13875_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][3]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2421),
    .D(_01566_),
    .Q_N(_13874_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][4]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2422),
    .D(_01567_),
    .Q_N(_13873_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][5]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2423),
    .D(_01568_),
    .Q_N(_13872_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][6]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2424),
    .D(_01569_),
    .Q_N(_13871_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][7]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2425),
    .D(_01570_),
    .Q_N(_13870_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][8]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2426),
    .D(_01571_),
    .Q_N(_13869_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][9]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2427),
    .D(_01572_),
    .Q_N(_13868_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][0]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2428),
    .D(_01573_),
    .Q_N(_13867_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][10]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2429),
    .D(_01574_),
    .Q_N(_13866_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][11]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2430),
    .D(_01575_),
    .Q_N(_13865_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][1]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2431),
    .D(_01576_),
    .Q_N(_13864_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][2]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2432),
    .D(_01577_),
    .Q_N(_13863_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][3]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2433),
    .D(_01578_),
    .Q_N(_13862_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][4]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2434),
    .D(_01579_),
    .Q_N(_13861_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][5]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2435),
    .D(_01580_),
    .Q_N(_13860_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][6]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2436),
    .D(_01581_),
    .Q_N(_13859_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][7]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2437),
    .D(_01582_),
    .Q_N(_13858_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][8]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2438),
    .D(_01583_),
    .Q_N(_13857_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][9]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2439),
    .D(_01584_),
    .Q_N(_13856_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][0]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2440),
    .D(_01585_),
    .Q_N(_13855_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][10]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2441),
    .D(_01586_),
    .Q_N(_13854_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][11]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2442),
    .D(_01587_),
    .Q_N(_13853_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][1]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2443),
    .D(_01588_),
    .Q_N(_13852_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][2]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2444),
    .D(_01589_),
    .Q_N(_13851_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][3]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2445),
    .D(_01590_),
    .Q_N(_13850_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][4]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net2446),
    .D(_01591_),
    .Q_N(_13849_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][5]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2447),
    .D(_01592_),
    .Q_N(_13848_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][6]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2448),
    .D(_01593_),
    .Q_N(_13847_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][7]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2449),
    .D(_01594_),
    .Q_N(_13846_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][8]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2450),
    .D(_01595_),
    .Q_N(_13845_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][9]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2451),
    .D(_01596_),
    .Q_N(_13844_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][0]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2452),
    .D(_01597_),
    .Q_N(_13843_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][10]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2453),
    .D(_01598_),
    .Q_N(_13842_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][11]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2454),
    .D(_01599_),
    .Q_N(_13841_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][1]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2455),
    .D(_01600_),
    .Q_N(_13840_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][2]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2456),
    .D(_01601_),
    .Q_N(_13839_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][3]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2457),
    .D(_01602_),
    .Q_N(_13838_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][4]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2458),
    .D(_01603_),
    .Q_N(_13837_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][5]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2459),
    .D(_01604_),
    .Q_N(_13836_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][6]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2460),
    .D(_01605_),
    .Q_N(_13835_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][7]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2461),
    .D(_01606_),
    .Q_N(_13834_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][8]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2462),
    .D(_01607_),
    .Q_N(_13833_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][9]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2463),
    .D(_01608_),
    .Q_N(_13832_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][0]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2464),
    .D(_01609_),
    .Q_N(_13831_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][10]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2465),
    .D(_01610_),
    .Q_N(_13830_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][11]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2466),
    .D(_01611_),
    .Q_N(_13829_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][1]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2467),
    .D(_01612_),
    .Q_N(_13828_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][2]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2468),
    .D(_01613_),
    .Q_N(_13827_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][3]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2469),
    .D(_01614_),
    .Q_N(_13826_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][4]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2470),
    .D(_01615_),
    .Q_N(_13825_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][5]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2471),
    .D(_01616_),
    .Q_N(_13824_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][6]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2472),
    .D(_01617_),
    .Q_N(_13823_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][7]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2473),
    .D(_01618_),
    .Q_N(_13822_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][8]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2474),
    .D(_01619_),
    .Q_N(_13821_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][9]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2475),
    .D(_01620_),
    .Q_N(_13820_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][0]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2476),
    .D(_01621_),
    .Q_N(_13819_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][10]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2477),
    .D(_01622_),
    .Q_N(_13818_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][11]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2478),
    .D(_01623_),
    .Q_N(_13817_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][1]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2479),
    .D(_01624_),
    .Q_N(_13816_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][2]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2480),
    .D(_01625_),
    .Q_N(_13815_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][3]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2481),
    .D(_01626_),
    .Q_N(_13814_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][4]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2482),
    .D(_01627_),
    .Q_N(_13813_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][5]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2483),
    .D(_01628_),
    .Q_N(_13812_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][6]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2484),
    .D(_01629_),
    .Q_N(_13811_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][7]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2485),
    .D(_01630_),
    .Q_N(_13810_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][8]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2486),
    .D(_01631_),
    .Q_N(_13809_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][9]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2487),
    .D(_01632_),
    .Q_N(_13808_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][0]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2488),
    .D(_01633_),
    .Q_N(_13807_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][10]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2489),
    .D(_01634_),
    .Q_N(_13806_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][11]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2490),
    .D(_01635_),
    .Q_N(_13805_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][1]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2491),
    .D(_01636_),
    .Q_N(_13804_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][2]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2492),
    .D(_01637_),
    .Q_N(_13803_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][3]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2493),
    .D(_01638_),
    .Q_N(_13802_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][4]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2494),
    .D(_01639_),
    .Q_N(_13801_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][5]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2495),
    .D(_01640_),
    .Q_N(_13800_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][6]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2496),
    .D(_01641_),
    .Q_N(_13799_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][7]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2497),
    .D(_01642_),
    .Q_N(_13798_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][8]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2498),
    .D(_01643_),
    .Q_N(_13797_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][9]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2499),
    .D(_01644_),
    .Q_N(_13796_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][0]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2500),
    .D(_01645_),
    .Q_N(_13795_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][10]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2501),
    .D(_01646_),
    .Q_N(_13794_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][11]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2502),
    .D(_01647_),
    .Q_N(_13793_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][1]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2503),
    .D(_01648_),
    .Q_N(_13792_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][2]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2504),
    .D(_01649_),
    .Q_N(_13791_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][3]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2505),
    .D(_01650_),
    .Q_N(_13790_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][4]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2506),
    .D(_01651_),
    .Q_N(_13789_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][5]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2507),
    .D(_01652_),
    .Q_N(_13788_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][6]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2508),
    .D(_01653_),
    .Q_N(_13787_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][7]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2509),
    .D(_01654_),
    .Q_N(_13786_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][8]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2510),
    .D(_01655_),
    .Q_N(_13785_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][9]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2511),
    .D(_01656_),
    .Q_N(_13784_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2512),
    .D(_01657_),
    .Q_N(_13783_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2513),
    .D(_01658_),
    .Q_N(_13782_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2514),
    .D(_01659_),
    .Q_N(_13781_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2515),
    .D(_01660_),
    .Q_N(_13780_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2516),
    .D(_01661_),
    .Q_N(_13779_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2517),
    .D(_01662_),
    .Q_N(_13778_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2518),
    .D(_01663_),
    .Q_N(_13777_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2519),
    .D(_01664_),
    .Q_N(_13776_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2520),
    .D(_01665_),
    .Q_N(_13775_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2521),
    .D(_01666_),
    .Q_N(_13774_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2522),
    .D(_01667_),
    .Q_N(_13773_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2523),
    .D(_01668_),
    .Q_N(_13772_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][0]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2524),
    .D(_01669_),
    .Q_N(_13771_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][10]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2525),
    .D(_01670_),
    .Q_N(_13770_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][11]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2526),
    .D(_01671_),
    .Q_N(_13769_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][1]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2527),
    .D(_01672_),
    .Q_N(_13768_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][2]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2528),
    .D(_01673_),
    .Q_N(_13767_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][3]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2529),
    .D(_01674_),
    .Q_N(_13766_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][4]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2530),
    .D(_01675_),
    .Q_N(_13765_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][5]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2531),
    .D(_01676_),
    .Q_N(_13764_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][6]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2532),
    .D(_01677_),
    .Q_N(_13763_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][7]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2533),
    .D(_01678_),
    .Q_N(_13762_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][8]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2534),
    .D(_01679_),
    .Q_N(_13761_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][9]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2535),
    .D(_01680_),
    .Q_N(_13760_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][0]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2536),
    .D(_01681_),
    .Q_N(_13759_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][10]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2537),
    .D(_01682_),
    .Q_N(_13758_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][11]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2538),
    .D(_01683_),
    .Q_N(_13757_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][1]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2539),
    .D(_01684_),
    .Q_N(_13756_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][2]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2540),
    .D(_01685_),
    .Q_N(_13755_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][3]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2541),
    .D(_01686_),
    .Q_N(_13754_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][4]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2542),
    .D(_01687_),
    .Q_N(_13753_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][5]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2543),
    .D(_01688_),
    .Q_N(_13752_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][6]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2544),
    .D(_01689_),
    .Q_N(_13751_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][7]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2545),
    .D(_01690_),
    .Q_N(_13750_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][8]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2546),
    .D(_01691_),
    .Q_N(_13749_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][9]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2547),
    .D(_01692_),
    .Q_N(_13748_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][0]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2548),
    .D(_01693_),
    .Q_N(_13747_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][10]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2549),
    .D(_01694_),
    .Q_N(_13746_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][11]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2550),
    .D(_01695_),
    .Q_N(_13745_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][1]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2551),
    .D(_01696_),
    .Q_N(_13744_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][2]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2552),
    .D(_01697_),
    .Q_N(_13743_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][3]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2553),
    .D(_01698_),
    .Q_N(_13742_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][4]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2554),
    .D(_01699_),
    .Q_N(_13741_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][5]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2555),
    .D(_01700_),
    .Q_N(_13740_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][6]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2556),
    .D(_01701_),
    .Q_N(_13739_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][7]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2557),
    .D(_01702_),
    .Q_N(_13738_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][8]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2558),
    .D(_01703_),
    .Q_N(_13737_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][9]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2559),
    .D(_01704_),
    .Q_N(_13736_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][0]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2560),
    .D(_01705_),
    .Q_N(_13735_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][10]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2561),
    .D(_01706_),
    .Q_N(_13734_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][11]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2562),
    .D(_01707_),
    .Q_N(_13733_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][1]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2563),
    .D(_01708_),
    .Q_N(_13732_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][2]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2564),
    .D(_01709_),
    .Q_N(_13731_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][3]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2565),
    .D(_01710_),
    .Q_N(_13730_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][4]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2566),
    .D(_01711_),
    .Q_N(_13729_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][5]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2567),
    .D(_01712_),
    .Q_N(_13728_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][6]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2568),
    .D(_01713_),
    .Q_N(_13727_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][7]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2569),
    .D(_01714_),
    .Q_N(_13726_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][8]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2570),
    .D(_01715_),
    .Q_N(_13725_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][9]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2571),
    .D(_01716_),
    .Q_N(_13724_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][0]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2572),
    .D(_01717_),
    .Q_N(_13723_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][10]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2573),
    .D(_01718_),
    .Q_N(_13722_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][11]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2574),
    .D(_01719_),
    .Q_N(_13721_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][1]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2575),
    .D(_01720_),
    .Q_N(_13720_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][2]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2576),
    .D(_01721_),
    .Q_N(_13719_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][3]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2577),
    .D(_01722_),
    .Q_N(_13718_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][4]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2578),
    .D(_01723_),
    .Q_N(_13717_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][5]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2579),
    .D(_01724_),
    .Q_N(_13716_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][6]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2580),
    .D(_01725_),
    .Q_N(_13715_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][7]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2581),
    .D(_01726_),
    .Q_N(_13714_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][8]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2582),
    .D(_01727_),
    .Q_N(_13713_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][9]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2583),
    .D(_01728_),
    .Q_N(_13712_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][0]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2584),
    .D(_01729_),
    .Q_N(_13711_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][10]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2585),
    .D(_01730_),
    .Q_N(_13710_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][11]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2586),
    .D(_01731_),
    .Q_N(_13709_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][1]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2587),
    .D(_01732_),
    .Q_N(_13708_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][2]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2588),
    .D(_01733_),
    .Q_N(_13707_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][3]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2589),
    .D(_01734_),
    .Q_N(_13706_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][4]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2590),
    .D(_01735_),
    .Q_N(_13705_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][5]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2591),
    .D(_01736_),
    .Q_N(_13704_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][6]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2592),
    .D(_01737_),
    .Q_N(_13703_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][7]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2593),
    .D(_01738_),
    .Q_N(_13702_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][8]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2594),
    .D(_01739_),
    .Q_N(_13701_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][9]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2595),
    .D(_01740_),
    .Q_N(_13700_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][0]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2596),
    .D(_01741_),
    .Q_N(_13699_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][10]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2597),
    .D(_01742_),
    .Q_N(_13698_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][11]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2598),
    .D(_01743_),
    .Q_N(_13697_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][1]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2599),
    .D(_01744_),
    .Q_N(_13696_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][2]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2600),
    .D(_01745_),
    .Q_N(_13695_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][3]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2601),
    .D(_01746_),
    .Q_N(_13694_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][4]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2602),
    .D(_01747_),
    .Q_N(_13693_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][5]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2603),
    .D(_01748_),
    .Q_N(_13692_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][6]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2604),
    .D(_01749_),
    .Q_N(_13691_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][7]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2605),
    .D(_01750_),
    .Q_N(_13690_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][8]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2606),
    .D(_01751_),
    .Q_N(_13689_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][9]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2607),
    .D(_01752_),
    .Q_N(_13688_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][0]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2608),
    .D(_01753_),
    .Q_N(_13687_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][10]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2609),
    .D(_01754_),
    .Q_N(_13686_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][11]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2610),
    .D(_01755_),
    .Q_N(_13685_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][1]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2611),
    .D(_01756_),
    .Q_N(_13684_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][2]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2612),
    .D(_01757_),
    .Q_N(_13683_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][3]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2613),
    .D(_01758_),
    .Q_N(_13682_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][4]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2614),
    .D(_01759_),
    .Q_N(_13681_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][5]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2615),
    .D(_01760_),
    .Q_N(_13680_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][6]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2616),
    .D(_01761_),
    .Q_N(_13679_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][7]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2617),
    .D(_01762_),
    .Q_N(_13678_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][8]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2618),
    .D(_01763_),
    .Q_N(_13677_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][9]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2619),
    .D(_01764_),
    .Q_N(_13676_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][0]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2620),
    .D(_01765_),
    .Q_N(_13675_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][10]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2621),
    .D(_01766_),
    .Q_N(_13674_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][11]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2622),
    .D(_01767_),
    .Q_N(_13673_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][1]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2623),
    .D(_01768_),
    .Q_N(_13672_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][2]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2624),
    .D(_01769_),
    .Q_N(_13671_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][3]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2625),
    .D(_01770_),
    .Q_N(_13670_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][4]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2626),
    .D(_01771_),
    .Q_N(_13669_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][5]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2627),
    .D(_01772_),
    .Q_N(_13668_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][6]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2628),
    .D(_01773_),
    .Q_N(_13667_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][7]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2629),
    .D(_01774_),
    .Q_N(_13666_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][8]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2630),
    .D(_01775_),
    .Q_N(_13665_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][9]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2631),
    .D(_01776_),
    .Q_N(_13664_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][0]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2632),
    .D(_01777_),
    .Q_N(_13663_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][10]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2633),
    .D(_01778_),
    .Q_N(_13662_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][11]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2634),
    .D(_01779_),
    .Q_N(_13661_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][1]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2635),
    .D(_01780_),
    .Q_N(_13660_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][2]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2636),
    .D(_01781_),
    .Q_N(_13659_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][3]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2637),
    .D(_01782_),
    .Q_N(_13658_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][4]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2638),
    .D(_01783_),
    .Q_N(_13657_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][5]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2639),
    .D(_01784_),
    .Q_N(_13656_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][6]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2640),
    .D(_01785_),
    .Q_N(_13655_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][7]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2641),
    .D(_01786_),
    .Q_N(_13654_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][8]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2642),
    .D(_01787_),
    .Q_N(_13653_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][9]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2643),
    .D(_01788_),
    .Q_N(_13652_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2644),
    .D(_01789_),
    .Q_N(_13651_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2645),
    .D(_01790_),
    .Q_N(_13650_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2646),
    .D(_01791_),
    .Q_N(_13649_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2647),
    .D(_01792_),
    .Q_N(_13648_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2648),
    .D(_01793_),
    .Q_N(_13647_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2649),
    .D(_01794_),
    .Q_N(_13646_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2650),
    .D(_01795_),
    .Q_N(_13645_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2651),
    .D(_01796_),
    .Q_N(_13644_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2652),
    .D(_01797_),
    .Q_N(_13643_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2653),
    .D(_01798_),
    .Q_N(_13642_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2654),
    .D(_01799_),
    .Q_N(_13641_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2655),
    .D(_01800_),
    .Q_N(_13640_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][0]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2656),
    .D(_01801_),
    .Q_N(_13639_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][10]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2657),
    .D(_01802_),
    .Q_N(_13638_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][11]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2658),
    .D(_01803_),
    .Q_N(_13637_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][1]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2659),
    .D(_01804_),
    .Q_N(_13636_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][2]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2660),
    .D(_01805_),
    .Q_N(_13635_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][3]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2661),
    .D(_01806_),
    .Q_N(_13634_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][4]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2662),
    .D(_01807_),
    .Q_N(_13633_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][5]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2663),
    .D(_01808_),
    .Q_N(_13632_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][6]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2664),
    .D(_01809_),
    .Q_N(_13631_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][7]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2665),
    .D(_01810_),
    .Q_N(_13630_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][8]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2666),
    .D(_01811_),
    .Q_N(_13629_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][9]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2667),
    .D(_01812_),
    .Q_N(_13628_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][0]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2668),
    .D(_01813_),
    .Q_N(_13627_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][10]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2669),
    .D(_01814_),
    .Q_N(_13626_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][11]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2670),
    .D(_01815_),
    .Q_N(_13625_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][1]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2671),
    .D(_01816_),
    .Q_N(_13624_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][2]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2672),
    .D(_01817_),
    .Q_N(_13623_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][3]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2673),
    .D(_01818_),
    .Q_N(_13622_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][4]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2674),
    .D(_01819_),
    .Q_N(_13621_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][5]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2675),
    .D(_01820_),
    .Q_N(_13620_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][6]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2676),
    .D(_01821_),
    .Q_N(_13619_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][7]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2677),
    .D(_01822_),
    .Q_N(_13618_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][8]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2678),
    .D(_01823_),
    .Q_N(_13617_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][9]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2679),
    .D(_01824_),
    .Q_N(_13616_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2680),
    .D(_01825_),
    .Q_N(_13615_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2681),
    .D(_01826_),
    .Q_N(_13614_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2682),
    .D(_01827_),
    .Q_N(_13613_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2683),
    .D(_01828_),
    .Q_N(_13612_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2684),
    .D(_01829_),
    .Q_N(_13611_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2685),
    .D(_01830_),
    .Q_N(_13610_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2686),
    .D(_01831_),
    .Q_N(_13609_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2687),
    .D(_01832_),
    .Q_N(_13608_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2688),
    .D(_01833_),
    .Q_N(_13607_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2689),
    .D(_01834_),
    .Q_N(_13606_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2690),
    .D(_01835_),
    .Q_N(_13605_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2691),
    .D(_01836_),
    .Q_N(_13604_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2692),
    .D(_01837_),
    .Q_N(_13603_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2693),
    .D(_01838_),
    .Q_N(_13602_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2694),
    .D(_01839_),
    .Q_N(_13601_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2695),
    .D(_01840_),
    .Q_N(_13600_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2696),
    .D(_01841_),
    .Q_N(_13599_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2697),
    .D(_01842_),
    .Q_N(_13598_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2698),
    .D(_01843_),
    .Q_N(_13597_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2699),
    .D(_01844_),
    .Q_N(_13596_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2700),
    .D(_01845_),
    .Q_N(_13595_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net2701),
    .D(_01846_),
    .Q_N(_13594_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2702),
    .D(_01847_),
    .Q_N(_13593_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2703),
    .D(_01848_),
    .Q_N(_13592_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2704),
    .D(_01849_),
    .Q_N(_13591_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2705),
    .D(_01850_),
    .Q_N(_13590_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2706),
    .D(_01851_),
    .Q_N(_13589_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2707),
    .D(_01852_),
    .Q_N(_13588_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2708),
    .D(_01853_),
    .Q_N(_13587_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2709),
    .D(_01854_),
    .Q_N(_13586_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2710),
    .D(_01855_),
    .Q_N(_13585_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2711),
    .D(_01856_),
    .Q_N(_13584_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2712),
    .D(_01857_),
    .Q_N(_13583_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2713),
    .D(_01858_),
    .Q_N(_13582_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2714),
    .D(_01859_),
    .Q_N(_13581_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2715),
    .D(_01860_),
    .Q_N(_13580_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2716),
    .D(_01861_),
    .Q_N(_13579_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2717),
    .D(_01862_),
    .Q_N(_13578_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2718),
    .D(_01863_),
    .Q_N(_13577_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2719),
    .D(_01864_),
    .Q_N(_13576_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2720),
    .D(_01865_),
    .Q_N(_13575_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2721),
    .D(_01866_),
    .Q_N(_13574_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2722),
    .D(_01867_),
    .Q_N(_13573_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2723),
    .D(_01868_),
    .Q_N(_13572_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2724),
    .D(_01869_),
    .Q_N(_13571_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2725),
    .D(_01870_),
    .Q_N(_13570_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2726),
    .D(_01871_),
    .Q_N(_13569_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2727),
    .D(_01872_),
    .Q_N(_13568_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2728),
    .D(_01873_),
    .Q_N(_13567_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2729),
    .D(_01874_),
    .Q_N(_13566_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2730),
    .D(_01875_),
    .Q_N(_13565_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2731),
    .D(_01876_),
    .Q_N(_13564_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2732),
    .D(_01877_),
    .Q_N(_13563_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2733),
    .D(_01878_),
    .Q_N(_13562_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2734),
    .D(_01879_),
    .Q_N(_13561_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2735),
    .D(_01880_),
    .Q_N(_13560_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2736),
    .D(_01881_),
    .Q_N(_13559_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2737),
    .D(_01882_),
    .Q_N(_13558_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2738),
    .D(_01883_),
    .Q_N(_13557_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2739),
    .D(_01884_),
    .Q_N(_13556_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][0]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2740),
    .D(_01885_),
    .Q_N(_13555_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][10]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2741),
    .D(_01886_),
    .Q_N(_13554_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][11]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2742),
    .D(_01887_),
    .Q_N(_13553_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][1]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2743),
    .D(_01888_),
    .Q_N(_13552_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][2]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2744),
    .D(_01889_),
    .Q_N(_13551_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][3]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2745),
    .D(_01890_),
    .Q_N(_13550_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][4]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net2746),
    .D(_01891_),
    .Q_N(_13549_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][5]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2747),
    .D(_01892_),
    .Q_N(_13548_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][6]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2748),
    .D(_01893_),
    .Q_N(_13547_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][7]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net2749),
    .D(_01894_),
    .Q_N(_13546_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][8]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2750),
    .D(_01895_),
    .Q_N(_13545_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][9]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2751),
    .D(_01896_),
    .Q_N(_13544_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][0]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2752),
    .D(_01897_),
    .Q_N(_13543_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][10]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2753),
    .D(_01898_),
    .Q_N(_13542_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][11]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2754),
    .D(_01899_),
    .Q_N(_13541_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][1]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2755),
    .D(_01900_),
    .Q_N(_13540_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][2]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2756),
    .D(_01901_),
    .Q_N(_13539_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][3]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2757),
    .D(_01902_),
    .Q_N(_13538_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][4]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net2758),
    .D(_01903_),
    .Q_N(_13537_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][5]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2759),
    .D(_01904_),
    .Q_N(_13536_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][6]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2760),
    .D(_01905_),
    .Q_N(_13535_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][7]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net2761),
    .D(_01906_),
    .Q_N(_13534_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][8]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2762),
    .D(_01907_),
    .Q_N(_13533_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][9]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2763),
    .D(_01908_),
    .Q_N(_13532_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[0]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2764),
    .D(_01909_),
    .Q_N(_13531_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[10]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2765),
    .D(_01910_),
    .Q_N(_13530_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[11]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2766),
    .D(_01911_),
    .Q_N(_13529_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[12]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2767),
    .D(_01912_),
    .Q_N(_13528_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[13]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2768),
    .D(_01913_),
    .Q_N(_13527_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[14]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2769),
    .D(_01914_),
    .Q_N(_13526_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[15]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2770),
    .D(_01915_),
    .Q_N(_13525_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[16]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2771),
    .D(_01916_),
    .Q_N(_13524_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[16] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[17]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2772),
    .D(_01917_),
    .Q_N(_13523_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[17] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[18]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2773),
    .D(_01918_),
    .Q_N(_13522_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[18] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[19]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2774),
    .D(_01919_),
    .Q_N(_13521_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[19] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[1]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2775),
    .D(_01920_),
    .Q_N(_13520_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[20]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2776),
    .D(_01921_),
    .Q_N(_13519_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[20] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[21]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2777),
    .D(_01922_),
    .Q_N(_13518_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[21] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[22]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2778),
    .D(_01923_),
    .Q_N(_13517_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[22] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[23]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2779),
    .D(_01924_),
    .Q_N(_13516_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[23] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[24]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2780),
    .D(_01925_),
    .Q_N(_13515_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[24] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[25]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2781),
    .D(_01926_),
    .Q_N(_13514_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[25] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[26]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2782),
    .D(_01927_),
    .Q_N(_13513_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[26] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[27]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2783),
    .D(_01928_),
    .Q_N(_13512_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[27] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[28]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2784),
    .D(_01929_),
    .Q_N(_13511_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[28] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[29]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2785),
    .D(_01930_),
    .Q_N(_13510_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[29] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[2]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2786),
    .D(_01931_),
    .Q_N(_13509_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[30]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2787),
    .D(_01932_),
    .Q_N(_13508_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[30] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[31]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2788),
    .D(_01933_),
    .Q_N(_13507_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[31] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[3]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2789),
    .D(_01934_),
    .Q_N(_13506_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[4]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2790),
    .D(_01935_),
    .Q_N(_13505_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[5]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2791),
    .D(_01936_),
    .Q_N(_13504_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[6]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2792),
    .D(_01937_),
    .Q_N(_13503_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[7]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2793),
    .D(_01938_),
    .Q_N(_13502_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[8]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2794),
    .D(_01939_),
    .Q_N(_13501_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[9]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2795),
    .D(_01940_),
    .Q_N(_13500_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[9] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2796),
    .D(_01941_),
    .Q_N(_13499_),
    .Q(\cpu.gpio.r_enable_in[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2797),
    .D(_01942_),
    .Q_N(_13498_),
    .Q(\cpu.gpio.r_enable_in[1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2798),
    .D(_01943_),
    .Q_N(_13497_),
    .Q(\cpu.gpio.r_enable_in[2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net2799),
    .D(_01944_),
    .Q_N(_13496_),
    .Q(\cpu.gpio.r_enable_in[3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2800),
    .D(_01945_),
    .Q_N(_13495_),
    .Q(\cpu.gpio.r_enable_in[4] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2801),
    .D(_01946_),
    .Q_N(_13494_),
    .Q(\cpu.gpio.r_enable_in[5] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net2802),
    .D(_01947_),
    .Q_N(_13493_),
    .Q(\cpu.gpio.r_enable_in[6] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net2803),
    .D(_01948_),
    .Q_N(_13492_),
    .Q(\cpu.gpio.r_enable_in[7] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2804),
    .D(_01949_),
    .Q_N(_13491_),
    .Q(\cpu.gpio.r_enable_io[4] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2805),
    .D(_01950_),
    .Q_N(_13490_),
    .Q(\cpu.gpio.r_enable_io[5] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2806),
    .D(_01951_),
    .Q_N(_13489_),
    .Q(\cpu.gpio.r_enable_io[6] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2807),
    .D(_01952_),
    .Q_N(_13488_),
    .Q(\cpu.gpio.r_enable_io[7] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2808),
    .D(_01953_),
    .Q_N(_13487_),
    .Q(net7));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2809),
    .D(_01954_),
    .Q_N(_13486_),
    .Q(net8));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2810),
    .D(_01955_),
    .Q_N(_13485_),
    .Q(net9));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2811),
    .D(_01956_),
    .Q_N(_13484_),
    .Q(net10));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[0]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2812),
    .D(_01957_),
    .Q_N(_13483_),
    .Q(\cpu.gpio.genblk2[4].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[1]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2813),
    .D(_01958_),
    .Q_N(_13482_),
    .Q(\cpu.gpio.genblk2[5].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[2]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2814),
    .D(_01959_),
    .Q_N(_13481_),
    .Q(\cpu.gpio.genblk2[6].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[3]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2815),
    .D(_01960_),
    .Q_N(_13480_),
    .Q(\cpu.gpio.genblk2[7].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[0]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2816),
    .D(_01961_),
    .Q_N(_13479_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[1]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2817),
    .D(_01962_),
    .Q_N(_13478_),
    .Q(\cpu.gpio.genblk1[4].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[2]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2818),
    .D(_01963_),
    .Q_N(_13477_),
    .Q(\cpu.gpio.genblk1[5].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[3]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2819),
    .D(_01964_),
    .Q_N(_13476_),
    .Q(\cpu.gpio.genblk1[6].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[4]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2820),
    .D(_01965_),
    .Q_N(_13475_),
    .Q(\cpu.gpio.genblk1[7].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2821),
    .D(_01966_),
    .Q_N(_13474_),
    .Q(\cpu.gpio.r_spi_miso_src[0][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2822),
    .D(_01967_),
    .Q_N(_00100_),
    .Q(\cpu.gpio.r_spi_miso_src[0][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2823),
    .D(_01968_),
    .Q_N(_00110_),
    .Q(\cpu.gpio.r_spi_miso_src[0][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2824),
    .D(_01969_),
    .Q_N(_00119_),
    .Q(\cpu.gpio.r_spi_miso_src[0][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2825),
    .D(_01970_),
    .Q_N(_13473_),
    .Q(\cpu.gpio.r_spi_miso_src[1][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2826),
    .D(_01971_),
    .Q_N(_00138_),
    .Q(\cpu.gpio.r_spi_miso_src[1][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2827),
    .D(_01972_),
    .Q_N(_00150_),
    .Q(\cpu.gpio.r_spi_miso_src[1][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2828),
    .D(_01973_),
    .Q_N(_00162_),
    .Q(\cpu.gpio.r_spi_miso_src[1][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2829),
    .D(_01974_),
    .Q_N(_13472_),
    .Q(\cpu.gpio.r_src_io[4][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2830),
    .D(_01975_),
    .Q_N(_13471_),
    .Q(\cpu.gpio.r_src_io[4][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2831),
    .D(_01976_),
    .Q_N(_00187_),
    .Q(\cpu.gpio.r_src_io[4][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2832),
    .D(_01977_),
    .Q_N(_13470_),
    .Q(\cpu.gpio.r_src_io[4][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2833),
    .D(_01978_),
    .Q_N(_13469_),
    .Q(\cpu.gpio.r_src_io[5][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2834),
    .D(_01979_),
    .Q_N(_13468_),
    .Q(\cpu.gpio.r_src_io[5][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2835),
    .D(_01980_),
    .Q_N(_00186_),
    .Q(\cpu.gpio.r_src_io[5][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2836),
    .D(_01981_),
    .Q_N(_13467_),
    .Q(\cpu.gpio.r_src_io[5][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2837),
    .D(_01982_),
    .Q_N(_13466_),
    .Q(\cpu.gpio.r_src_io[6][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2838),
    .D(_01983_),
    .Q_N(_00096_),
    .Q(\cpu.gpio.r_src_io[6][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2839),
    .D(_01984_),
    .Q_N(_00106_),
    .Q(\cpu.gpio.r_src_io[6][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2840),
    .D(_01985_),
    .Q_N(_00116_),
    .Q(\cpu.gpio.r_src_io[6][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2841),
    .D(_01986_),
    .Q_N(_13465_),
    .Q(\cpu.gpio.r_src_io[7][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2842),
    .D(_01987_),
    .Q_N(_00134_),
    .Q(\cpu.gpio.r_src_io[7][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2843),
    .D(_01988_),
    .Q_N(_00146_),
    .Q(\cpu.gpio.r_src_io[7][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2844),
    .D(_01989_),
    .Q_N(_00158_),
    .Q(\cpu.gpio.r_src_io[7][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2845),
    .D(_01990_),
    .Q_N(_13464_),
    .Q(\cpu.gpio.r_src_o[3][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2846),
    .D(_01991_),
    .Q_N(_00137_),
    .Q(\cpu.gpio.r_src_o[3][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2847),
    .D(_01992_),
    .Q_N(_00149_),
    .Q(\cpu.gpio.r_src_o[3][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2848),
    .D(_01993_),
    .Q_N(_00161_),
    .Q(\cpu.gpio.r_src_o[3][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2849),
    .D(_01994_),
    .Q_N(_13463_),
    .Q(\cpu.gpio.r_src_o[4][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2850),
    .D(_01995_),
    .Q_N(_00098_),
    .Q(\cpu.gpio.r_src_o[4][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2851),
    .D(_01996_),
    .Q_N(_00108_),
    .Q(\cpu.gpio.r_src_o[4][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2852),
    .D(_01997_),
    .Q_N(_00118_),
    .Q(\cpu.gpio.r_src_o[4][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2853),
    .D(_01998_),
    .Q_N(_13462_),
    .Q(\cpu.gpio.r_src_o[5][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2854),
    .D(_01999_),
    .Q_N(_00136_),
    .Q(\cpu.gpio.r_src_o[5][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2855),
    .D(_02000_),
    .Q_N(_00148_),
    .Q(\cpu.gpio.r_src_o[5][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2856),
    .D(_02001_),
    .Q_N(_00160_),
    .Q(\cpu.gpio.r_src_o[5][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2857),
    .D(_02002_),
    .Q_N(_13461_),
    .Q(\cpu.gpio.r_src_o[6][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2858),
    .D(_02003_),
    .Q_N(_00097_),
    .Q(\cpu.gpio.r_src_o[6][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2859),
    .D(_02004_),
    .Q_N(_00107_),
    .Q(\cpu.gpio.r_src_o[6][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2860),
    .D(_02005_),
    .Q_N(_00117_),
    .Q(\cpu.gpio.r_src_o[6][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2861),
    .D(_02006_),
    .Q_N(_13460_),
    .Q(\cpu.gpio.r_src_o[7][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2862),
    .D(_02007_),
    .Q_N(_00135_),
    .Q(\cpu.gpio.r_src_o[7][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2863),
    .D(_02008_),
    .Q_N(_00147_),
    .Q(\cpu.gpio.r_src_o[7][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2864),
    .D(_02009_),
    .Q_N(_00159_),
    .Q(\cpu.gpio.r_src_o[7][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_uart_rx_src[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2865),
    .D(_02010_),
    .Q_N(_13459_),
    .Q(\cpu.gpio.r_uart_rx_src[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_uart_rx_src[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2866),
    .D(_02011_),
    .Q_N(_00099_),
    .Q(\cpu.gpio.r_uart_rx_src[1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_uart_rx_src[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2867),
    .D(_02012_),
    .Q_N(_00109_),
    .Q(\cpu.gpio.r_uart_rx_src[2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2868),
    .D(_02013_),
    .Q_N(_13458_),
    .Q(\cpu.icache.r_data[0][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2869),
    .D(_02014_),
    .Q_N(_00205_),
    .Q(\cpu.icache.r_data[0][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2870),
    .D(_02015_),
    .Q_N(_00207_),
    .Q(\cpu.icache.r_data[0][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2871),
    .D(_02016_),
    .Q_N(_00213_),
    .Q(\cpu.icache.r_data[0][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2872),
    .D(_02017_),
    .Q_N(_13457_),
    .Q(\cpu.icache.r_data[0][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2873),
    .D(_02018_),
    .Q_N(_00201_),
    .Q(\cpu.icache.r_data[0][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2874),
    .D(_02019_),
    .Q_N(_00203_),
    .Q(\cpu.icache.r_data[0][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2875),
    .D(_02020_),
    .Q_N(_13456_),
    .Q(\cpu.icache.r_data[0][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2876),
    .D(_02021_),
    .Q_N(_13455_),
    .Q(\cpu.icache.r_data[0][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2877),
    .D(_02022_),
    .Q_N(_00216_),
    .Q(\cpu.icache.r_data[0][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][19]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2878),
    .D(_02023_),
    .Q_N(_00218_),
    .Q(\cpu.icache.r_data[0][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2879),
    .D(_02024_),
    .Q_N(_13454_),
    .Q(\cpu.icache.r_data[0][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][20]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2880),
    .D(_02025_),
    .Q_N(_00220_),
    .Q(\cpu.icache.r_data[0][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][21]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2881),
    .D(_02026_),
    .Q_N(_00210_),
    .Q(\cpu.icache.r_data[0][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][22]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2882),
    .D(_02027_),
    .Q_N(_00212_),
    .Q(\cpu.icache.r_data[0][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][23]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2883),
    .D(_02028_),
    .Q_N(_00173_),
    .Q(\cpu.icache.r_data[0][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][24]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2884),
    .D(_02029_),
    .Q_N(_00175_),
    .Q(\cpu.icache.r_data[0][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][25]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2885),
    .D(_02030_),
    .Q_N(_00177_),
    .Q(\cpu.icache.r_data[0][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][26]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2886),
    .D(_02031_),
    .Q_N(_00206_),
    .Q(\cpu.icache.r_data[0][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][27]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2887),
    .D(_02032_),
    .Q_N(_00208_),
    .Q(\cpu.icache.r_data[0][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][28]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2888),
    .D(_02033_),
    .Q_N(_00214_),
    .Q(\cpu.icache.r_data[0][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][29]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2889),
    .D(_02034_),
    .Q_N(_13453_),
    .Q(\cpu.icache.r_data[0][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2890),
    .D(_02035_),
    .Q_N(_00215_),
    .Q(\cpu.icache.r_data[0][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][30]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2891),
    .D(_02036_),
    .Q_N(_00202_),
    .Q(\cpu.icache.r_data[0][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][31]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2892),
    .D(_02037_),
    .Q_N(_00204_),
    .Q(\cpu.icache.r_data[0][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2893),
    .D(_02038_),
    .Q_N(_00217_),
    .Q(\cpu.icache.r_data[0][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2894),
    .D(_02039_),
    .Q_N(_00219_),
    .Q(\cpu.icache.r_data[0][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2895),
    .D(_02040_),
    .Q_N(_00209_),
    .Q(\cpu.icache.r_data[0][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2896),
    .D(_02041_),
    .Q_N(_00211_),
    .Q(\cpu.icache.r_data[0][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2897),
    .D(_02042_),
    .Q_N(_00172_),
    .Q(\cpu.icache.r_data[0][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2898),
    .D(_02043_),
    .Q_N(_00174_),
    .Q(\cpu.icache.r_data[0][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2899),
    .D(_02044_),
    .Q_N(_00176_),
    .Q(\cpu.icache.r_data[0][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2900),
    .D(_02045_),
    .Q_N(_13452_),
    .Q(\cpu.icache.r_data[1][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2901),
    .D(_02046_),
    .Q_N(_13451_),
    .Q(\cpu.icache.r_data[1][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2902),
    .D(_02047_),
    .Q_N(_13450_),
    .Q(\cpu.icache.r_data[1][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2903),
    .D(_02048_),
    .Q_N(_13449_),
    .Q(\cpu.icache.r_data[1][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2904),
    .D(_02049_),
    .Q_N(_13448_),
    .Q(\cpu.icache.r_data[1][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2905),
    .D(_02050_),
    .Q_N(_13447_),
    .Q(\cpu.icache.r_data[1][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net2906),
    .D(_02051_),
    .Q_N(_13446_),
    .Q(\cpu.icache.r_data[1][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2907),
    .D(_02052_),
    .Q_N(_13445_),
    .Q(\cpu.icache.r_data[1][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2908),
    .D(_02053_),
    .Q_N(_13444_),
    .Q(\cpu.icache.r_data[1][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2909),
    .D(_02054_),
    .Q_N(_13443_),
    .Q(\cpu.icache.r_data[1][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][19]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2910),
    .D(_02055_),
    .Q_N(_13442_),
    .Q(\cpu.icache.r_data[1][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2911),
    .D(_02056_),
    .Q_N(_13441_),
    .Q(\cpu.icache.r_data[1][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][20]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2912),
    .D(_02057_),
    .Q_N(_13440_),
    .Q(\cpu.icache.r_data[1][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][21]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2913),
    .D(_02058_),
    .Q_N(_13439_),
    .Q(\cpu.icache.r_data[1][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][22]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2914),
    .D(_02059_),
    .Q_N(_13438_),
    .Q(\cpu.icache.r_data[1][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][23]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2915),
    .D(_02060_),
    .Q_N(_13437_),
    .Q(\cpu.icache.r_data[1][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][24]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2916),
    .D(_02061_),
    .Q_N(_13436_),
    .Q(\cpu.icache.r_data[1][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][25]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2917),
    .D(_02062_),
    .Q_N(_13435_),
    .Q(\cpu.icache.r_data[1][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][26]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2918),
    .D(_02063_),
    .Q_N(_13434_),
    .Q(\cpu.icache.r_data[1][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][27]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2919),
    .D(_02064_),
    .Q_N(_13433_),
    .Q(\cpu.icache.r_data[1][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][28]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2920),
    .D(_02065_),
    .Q_N(_13432_),
    .Q(\cpu.icache.r_data[1][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][29]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2921),
    .D(_02066_),
    .Q_N(_13431_),
    .Q(\cpu.icache.r_data[1][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2922),
    .D(_02067_),
    .Q_N(_13430_),
    .Q(\cpu.icache.r_data[1][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][30]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2923),
    .D(_02068_),
    .Q_N(_13429_),
    .Q(\cpu.icache.r_data[1][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][31]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2924),
    .D(_02069_),
    .Q_N(_13428_),
    .Q(\cpu.icache.r_data[1][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2925),
    .D(_02070_),
    .Q_N(_13427_),
    .Q(\cpu.icache.r_data[1][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2926),
    .D(_02071_),
    .Q_N(_13426_),
    .Q(\cpu.icache.r_data[1][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2927),
    .D(_02072_),
    .Q_N(_13425_),
    .Q(\cpu.icache.r_data[1][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2928),
    .D(_02073_),
    .Q_N(_13424_),
    .Q(\cpu.icache.r_data[1][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2929),
    .D(_02074_),
    .Q_N(_13423_),
    .Q(\cpu.icache.r_data[1][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2930),
    .D(_02075_),
    .Q_N(_13422_),
    .Q(\cpu.icache.r_data[1][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2931),
    .D(_02076_),
    .Q_N(_13421_),
    .Q(\cpu.icache.r_data[1][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2932),
    .D(_02077_),
    .Q_N(_13420_),
    .Q(\cpu.icache.r_data[2][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2933),
    .D(_02078_),
    .Q_N(_13419_),
    .Q(\cpu.icache.r_data[2][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2934),
    .D(_02079_),
    .Q_N(_13418_),
    .Q(\cpu.icache.r_data[2][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2935),
    .D(_02080_),
    .Q_N(_13417_),
    .Q(\cpu.icache.r_data[2][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2936),
    .D(_02081_),
    .Q_N(_13416_),
    .Q(\cpu.icache.r_data[2][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2937),
    .D(_02082_),
    .Q_N(_13415_),
    .Q(\cpu.icache.r_data[2][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2938),
    .D(_02083_),
    .Q_N(_13414_),
    .Q(\cpu.icache.r_data[2][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2939),
    .D(_02084_),
    .Q_N(_13413_),
    .Q(\cpu.icache.r_data[2][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2940),
    .D(_02085_),
    .Q_N(_13412_),
    .Q(\cpu.icache.r_data[2][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2941),
    .D(_02086_),
    .Q_N(_13411_),
    .Q(\cpu.icache.r_data[2][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][19]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2942),
    .D(_02087_),
    .Q_N(_13410_),
    .Q(\cpu.icache.r_data[2][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2943),
    .D(_02088_),
    .Q_N(_13409_),
    .Q(\cpu.icache.r_data[2][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][20]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2944),
    .D(_02089_),
    .Q_N(_13408_),
    .Q(\cpu.icache.r_data[2][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][21]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2945),
    .D(_02090_),
    .Q_N(_13407_),
    .Q(\cpu.icache.r_data[2][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][22]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2946),
    .D(_02091_),
    .Q_N(_13406_),
    .Q(\cpu.icache.r_data[2][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][23]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2947),
    .D(_02092_),
    .Q_N(_13405_),
    .Q(\cpu.icache.r_data[2][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][24]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2948),
    .D(_02093_),
    .Q_N(_13404_),
    .Q(\cpu.icache.r_data[2][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][25]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2949),
    .D(_02094_),
    .Q_N(_13403_),
    .Q(\cpu.icache.r_data[2][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][26]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2950),
    .D(_02095_),
    .Q_N(_13402_),
    .Q(\cpu.icache.r_data[2][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][27]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2951),
    .D(_02096_),
    .Q_N(_13401_),
    .Q(\cpu.icache.r_data[2][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][28]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2952),
    .D(_02097_),
    .Q_N(_13400_),
    .Q(\cpu.icache.r_data[2][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][29]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2953),
    .D(_02098_),
    .Q_N(_13399_),
    .Q(\cpu.icache.r_data[2][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2954),
    .D(_02099_),
    .Q_N(_13398_),
    .Q(\cpu.icache.r_data[2][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][30]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2955),
    .D(_02100_),
    .Q_N(_13397_),
    .Q(\cpu.icache.r_data[2][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][31]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2956),
    .D(_02101_),
    .Q_N(_13396_),
    .Q(\cpu.icache.r_data[2][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2957),
    .D(_02102_),
    .Q_N(_13395_),
    .Q(\cpu.icache.r_data[2][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2958),
    .D(_02103_),
    .Q_N(_13394_),
    .Q(\cpu.icache.r_data[2][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2959),
    .D(_02104_),
    .Q_N(_13393_),
    .Q(\cpu.icache.r_data[2][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2960),
    .D(_02105_),
    .Q_N(_13392_),
    .Q(\cpu.icache.r_data[2][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2961),
    .D(_02106_),
    .Q_N(_13391_),
    .Q(\cpu.icache.r_data[2][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2962),
    .D(_02107_),
    .Q_N(_13390_),
    .Q(\cpu.icache.r_data[2][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2963),
    .D(_02108_),
    .Q_N(_13389_),
    .Q(\cpu.icache.r_data[2][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2964),
    .D(_02109_),
    .Q_N(_13388_),
    .Q(\cpu.icache.r_data[3][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2965),
    .D(_02110_),
    .Q_N(_13387_),
    .Q(\cpu.icache.r_data[3][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2966),
    .D(_02111_),
    .Q_N(_13386_),
    .Q(\cpu.icache.r_data[3][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2967),
    .D(_02112_),
    .Q_N(_13385_),
    .Q(\cpu.icache.r_data[3][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2968),
    .D(_02113_),
    .Q_N(_13384_),
    .Q(\cpu.icache.r_data[3][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2969),
    .D(_02114_),
    .Q_N(_13383_),
    .Q(\cpu.icache.r_data[3][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2970),
    .D(_02115_),
    .Q_N(_13382_),
    .Q(\cpu.icache.r_data[3][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2971),
    .D(_02116_),
    .Q_N(_13381_),
    .Q(\cpu.icache.r_data[3][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2972),
    .D(_02117_),
    .Q_N(_13380_),
    .Q(\cpu.icache.r_data[3][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2973),
    .D(_02118_),
    .Q_N(_13379_),
    .Q(\cpu.icache.r_data[3][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][19]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2974),
    .D(_02119_),
    .Q_N(_13378_),
    .Q(\cpu.icache.r_data[3][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2975),
    .D(_02120_),
    .Q_N(_13377_),
    .Q(\cpu.icache.r_data[3][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][20]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2976),
    .D(_02121_),
    .Q_N(_13376_),
    .Q(\cpu.icache.r_data[3][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][21]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2977),
    .D(_02122_),
    .Q_N(_13375_),
    .Q(\cpu.icache.r_data[3][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][22]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2978),
    .D(_02123_),
    .Q_N(_13374_),
    .Q(\cpu.icache.r_data[3][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][23]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2979),
    .D(_02124_),
    .Q_N(_13373_),
    .Q(\cpu.icache.r_data[3][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][24]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2980),
    .D(_02125_),
    .Q_N(_13372_),
    .Q(\cpu.icache.r_data[3][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][25]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2981),
    .D(_02126_),
    .Q_N(_13371_),
    .Q(\cpu.icache.r_data[3][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][26]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2982),
    .D(_02127_),
    .Q_N(_13370_),
    .Q(\cpu.icache.r_data[3][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][27]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2983),
    .D(_02128_),
    .Q_N(_13369_),
    .Q(\cpu.icache.r_data[3][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][28]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2984),
    .D(_02129_),
    .Q_N(_13368_),
    .Q(\cpu.icache.r_data[3][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][29]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2985),
    .D(_02130_),
    .Q_N(_13367_),
    .Q(\cpu.icache.r_data[3][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2986),
    .D(_02131_),
    .Q_N(_13366_),
    .Q(\cpu.icache.r_data[3][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][30]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2987),
    .D(_02132_),
    .Q_N(_13365_),
    .Q(\cpu.icache.r_data[3][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][31]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2988),
    .D(_02133_),
    .Q_N(_13364_),
    .Q(\cpu.icache.r_data[3][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2989),
    .D(_02134_),
    .Q_N(_13363_),
    .Q(\cpu.icache.r_data[3][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2990),
    .D(_02135_),
    .Q_N(_13362_),
    .Q(\cpu.icache.r_data[3][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2991),
    .D(_02136_),
    .Q_N(_13361_),
    .Q(\cpu.icache.r_data[3][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2992),
    .D(_02137_),
    .Q_N(_13360_),
    .Q(\cpu.icache.r_data[3][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2993),
    .D(_02138_),
    .Q_N(_13359_),
    .Q(\cpu.icache.r_data[3][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2994),
    .D(_02139_),
    .Q_N(_13358_),
    .Q(\cpu.icache.r_data[3][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2995),
    .D(_02140_),
    .Q_N(_13357_),
    .Q(\cpu.icache.r_data[3][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2996),
    .D(_02141_),
    .Q_N(_13356_),
    .Q(\cpu.icache.r_data[4][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2997),
    .D(_02142_),
    .Q_N(_13355_),
    .Q(\cpu.icache.r_data[4][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2998),
    .D(_02143_),
    .Q_N(_13354_),
    .Q(\cpu.icache.r_data[4][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2999),
    .D(_02144_),
    .Q_N(_13353_),
    .Q(\cpu.icache.r_data[4][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3000),
    .D(_02145_),
    .Q_N(_13352_),
    .Q(\cpu.icache.r_data[4][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3001),
    .D(_02146_),
    .Q_N(_13351_),
    .Q(\cpu.icache.r_data[4][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3002),
    .D(_02147_),
    .Q_N(_13350_),
    .Q(\cpu.icache.r_data[4][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net3003),
    .D(_02148_),
    .Q_N(_13349_),
    .Q(\cpu.icache.r_data[4][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net3004),
    .D(_02149_),
    .Q_N(_13348_),
    .Q(\cpu.icache.r_data[4][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net3005),
    .D(_02150_),
    .Q_N(_13347_),
    .Q(\cpu.icache.r_data[4][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][19]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net3006),
    .D(_02151_),
    .Q_N(_13346_),
    .Q(\cpu.icache.r_data[4][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net3007),
    .D(_02152_),
    .Q_N(_13345_),
    .Q(\cpu.icache.r_data[4][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][20]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net3008),
    .D(_02153_),
    .Q_N(_13344_),
    .Q(\cpu.icache.r_data[4][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][21]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net3009),
    .D(_02154_),
    .Q_N(_13343_),
    .Q(\cpu.icache.r_data[4][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][22]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net3010),
    .D(_02155_),
    .Q_N(_13342_),
    .Q(\cpu.icache.r_data[4][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][23]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3011),
    .D(_02156_),
    .Q_N(_13341_),
    .Q(\cpu.icache.r_data[4][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][24]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3012),
    .D(_02157_),
    .Q_N(_13340_),
    .Q(\cpu.icache.r_data[4][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][25]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3013),
    .D(_02158_),
    .Q_N(_13339_),
    .Q(\cpu.icache.r_data[4][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][26]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3014),
    .D(_02159_),
    .Q_N(_13338_),
    .Q(\cpu.icache.r_data[4][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][27]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3015),
    .D(_02160_),
    .Q_N(_13337_),
    .Q(\cpu.icache.r_data[4][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][28]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3016),
    .D(_02161_),
    .Q_N(_13336_),
    .Q(\cpu.icache.r_data[4][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][29]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3017),
    .D(_02162_),
    .Q_N(_13335_),
    .Q(\cpu.icache.r_data[4][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net3018),
    .D(_02163_),
    .Q_N(_13334_),
    .Q(\cpu.icache.r_data[4][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][30]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net3019),
    .D(_02164_),
    .Q_N(_13333_),
    .Q(\cpu.icache.r_data[4][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][31]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3020),
    .D(_02165_),
    .Q_N(_13332_),
    .Q(\cpu.icache.r_data[4][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3021),
    .D(_02166_),
    .Q_N(_13331_),
    .Q(\cpu.icache.r_data[4][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net3022),
    .D(_02167_),
    .Q_N(_13330_),
    .Q(\cpu.icache.r_data[4][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net3023),
    .D(_02168_),
    .Q_N(_13329_),
    .Q(\cpu.icache.r_data[4][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net3024),
    .D(_02169_),
    .Q_N(_13328_),
    .Q(\cpu.icache.r_data[4][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net3025),
    .D(_02170_),
    .Q_N(_13327_),
    .Q(\cpu.icache.r_data[4][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3026),
    .D(_02171_),
    .Q_N(_13326_),
    .Q(\cpu.icache.r_data[4][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3027),
    .D(_02172_),
    .Q_N(_13325_),
    .Q(\cpu.icache.r_data[4][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net3028),
    .D(_02173_),
    .Q_N(_13324_),
    .Q(\cpu.icache.r_data[5][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3029),
    .D(_02174_),
    .Q_N(_13323_),
    .Q(\cpu.icache.r_data[5][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3030),
    .D(_02175_),
    .Q_N(_13322_),
    .Q(\cpu.icache.r_data[5][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3031),
    .D(_02176_),
    .Q_N(_13321_),
    .Q(\cpu.icache.r_data[5][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3032),
    .D(_02177_),
    .Q_N(_13320_),
    .Q(\cpu.icache.r_data[5][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net3033),
    .D(_02178_),
    .Q_N(_13319_),
    .Q(\cpu.icache.r_data[5][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3034),
    .D(_02179_),
    .Q_N(_13318_),
    .Q(\cpu.icache.r_data[5][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net3035),
    .D(_02180_),
    .Q_N(_13317_),
    .Q(\cpu.icache.r_data[5][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net3036),
    .D(_02181_),
    .Q_N(_13316_),
    .Q(\cpu.icache.r_data[5][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net3037),
    .D(_02182_),
    .Q_N(_13315_),
    .Q(\cpu.icache.r_data[5][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][19]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net3038),
    .D(_02183_),
    .Q_N(_13314_),
    .Q(\cpu.icache.r_data[5][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3039),
    .D(_02184_),
    .Q_N(_13313_),
    .Q(\cpu.icache.r_data[5][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][20]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net3040),
    .D(_02185_),
    .Q_N(_13312_),
    .Q(\cpu.icache.r_data[5][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][21]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net3041),
    .D(_02186_),
    .Q_N(_13311_),
    .Q(\cpu.icache.r_data[5][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][22]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net3042),
    .D(_02187_),
    .Q_N(_13310_),
    .Q(\cpu.icache.r_data[5][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][23]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3043),
    .D(_02188_),
    .Q_N(_13309_),
    .Q(\cpu.icache.r_data[5][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][24]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3044),
    .D(_02189_),
    .Q_N(_13308_),
    .Q(\cpu.icache.r_data[5][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][25]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3045),
    .D(_02190_),
    .Q_N(_13307_),
    .Q(\cpu.icache.r_data[5][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][26]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3046),
    .D(_02191_),
    .Q_N(_13306_),
    .Q(\cpu.icache.r_data[5][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][27]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3047),
    .D(_02192_),
    .Q_N(_13305_),
    .Q(\cpu.icache.r_data[5][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][28]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net3048),
    .D(_02193_),
    .Q_N(_13304_),
    .Q(\cpu.icache.r_data[5][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][29]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net3049),
    .D(_02194_),
    .Q_N(_13303_),
    .Q(\cpu.icache.r_data[5][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net3050),
    .D(_02195_),
    .Q_N(_13302_),
    .Q(\cpu.icache.r_data[5][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][30]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3051),
    .D(_02196_),
    .Q_N(_13301_),
    .Q(\cpu.icache.r_data[5][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][31]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net3052),
    .D(_02197_),
    .Q_N(_13300_),
    .Q(\cpu.icache.r_data[5][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net3053),
    .D(_02198_),
    .Q_N(_13299_),
    .Q(\cpu.icache.r_data[5][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net3054),
    .D(_02199_),
    .Q_N(_13298_),
    .Q(\cpu.icache.r_data[5][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3055),
    .D(_02200_),
    .Q_N(_13297_),
    .Q(\cpu.icache.r_data[5][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net3056),
    .D(_02201_),
    .Q_N(_13296_),
    .Q(\cpu.icache.r_data[5][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net3057),
    .D(_02202_),
    .Q_N(_13295_),
    .Q(\cpu.icache.r_data[5][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3058),
    .D(_02203_),
    .Q_N(_13294_),
    .Q(\cpu.icache.r_data[5][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3059),
    .D(_02204_),
    .Q_N(_13293_),
    .Q(\cpu.icache.r_data[5][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3060),
    .D(_02205_),
    .Q_N(_13292_),
    .Q(\cpu.icache.r_data[6][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3061),
    .D(_02206_),
    .Q_N(_13291_),
    .Q(\cpu.icache.r_data[6][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3062),
    .D(_02207_),
    .Q_N(_13290_),
    .Q(\cpu.icache.r_data[6][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3063),
    .D(_02208_),
    .Q_N(_13289_),
    .Q(\cpu.icache.r_data[6][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3064),
    .D(_02209_),
    .Q_N(_13288_),
    .Q(\cpu.icache.r_data[6][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3065),
    .D(_02210_),
    .Q_N(_13287_),
    .Q(\cpu.icache.r_data[6][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3066),
    .D(_02211_),
    .Q_N(_13286_),
    .Q(\cpu.icache.r_data[6][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net3067),
    .D(_02212_),
    .Q_N(_13285_),
    .Q(\cpu.icache.r_data[6][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net3068),
    .D(_02213_),
    .Q_N(_13284_),
    .Q(\cpu.icache.r_data[6][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net3069),
    .D(_02214_),
    .Q_N(_13283_),
    .Q(\cpu.icache.r_data[6][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][19]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net3070),
    .D(_02215_),
    .Q_N(_13282_),
    .Q(\cpu.icache.r_data[6][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net3071),
    .D(_02216_),
    .Q_N(_13281_),
    .Q(\cpu.icache.r_data[6][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][20]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net3072),
    .D(_02217_),
    .Q_N(_13280_),
    .Q(\cpu.icache.r_data[6][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][21]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net3073),
    .D(_02218_),
    .Q_N(_13279_),
    .Q(\cpu.icache.r_data[6][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][22]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net3074),
    .D(_02219_),
    .Q_N(_13278_),
    .Q(\cpu.icache.r_data[6][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][23]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3075),
    .D(_02220_),
    .Q_N(_13277_),
    .Q(\cpu.icache.r_data[6][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][24]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3076),
    .D(_02221_),
    .Q_N(_13276_),
    .Q(\cpu.icache.r_data[6][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][25]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3077),
    .D(_02222_),
    .Q_N(_13275_),
    .Q(\cpu.icache.r_data[6][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][26]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3078),
    .D(_02223_),
    .Q_N(_13274_),
    .Q(\cpu.icache.r_data[6][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][27]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3079),
    .D(_02224_),
    .Q_N(_13273_),
    .Q(\cpu.icache.r_data[6][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][28]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net3080),
    .D(_02225_),
    .Q_N(_13272_),
    .Q(\cpu.icache.r_data[6][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][29]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net3081),
    .D(_02226_),
    .Q_N(_13271_),
    .Q(\cpu.icache.r_data[6][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net3082),
    .D(_02227_),
    .Q_N(_13270_),
    .Q(\cpu.icache.r_data[6][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][30]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net3083),
    .D(_02228_),
    .Q_N(_13269_),
    .Q(\cpu.icache.r_data[6][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][31]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3084),
    .D(_02229_),
    .Q_N(_13268_),
    .Q(\cpu.icache.r_data[6][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3085),
    .D(_02230_),
    .Q_N(_13267_),
    .Q(\cpu.icache.r_data[6][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net3086),
    .D(_02231_),
    .Q_N(_13266_),
    .Q(\cpu.icache.r_data[6][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net3087),
    .D(_02232_),
    .Q_N(_13265_),
    .Q(\cpu.icache.r_data[6][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net3088),
    .D(_02233_),
    .Q_N(_13264_),
    .Q(\cpu.icache.r_data[6][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3089),
    .D(_02234_),
    .Q_N(_13263_),
    .Q(\cpu.icache.r_data[6][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3090),
    .D(_02235_),
    .Q_N(_13262_),
    .Q(\cpu.icache.r_data[6][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3091),
    .D(_02236_),
    .Q_N(_13261_),
    .Q(\cpu.icache.r_data[6][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net3092),
    .D(_02237_),
    .Q_N(_13260_),
    .Q(\cpu.icache.r_data[7][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3093),
    .D(_02238_),
    .Q_N(_13259_),
    .Q(\cpu.icache.r_data[7][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3094),
    .D(_02239_),
    .Q_N(_13258_),
    .Q(\cpu.icache.r_data[7][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3095),
    .D(_02240_),
    .Q_N(_13257_),
    .Q(\cpu.icache.r_data[7][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3096),
    .D(_02241_),
    .Q_N(_13256_),
    .Q(\cpu.icache.r_data[7][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3097),
    .D(_02242_),
    .Q_N(_13255_),
    .Q(\cpu.icache.r_data[7][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3098),
    .D(_02243_),
    .Q_N(_13254_),
    .Q(\cpu.icache.r_data[7][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net3099),
    .D(_02244_),
    .Q_N(_13253_),
    .Q(\cpu.icache.r_data[7][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net3100),
    .D(_02245_),
    .Q_N(_13252_),
    .Q(\cpu.icache.r_data[7][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net3101),
    .D(_02246_),
    .Q_N(_13251_),
    .Q(\cpu.icache.r_data[7][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][19]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net3102),
    .D(_02247_),
    .Q_N(_13250_),
    .Q(\cpu.icache.r_data[7][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net3103),
    .D(_02248_),
    .Q_N(_13249_),
    .Q(\cpu.icache.r_data[7][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][20]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net3104),
    .D(_02249_),
    .Q_N(_13248_),
    .Q(\cpu.icache.r_data[7][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][21]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net3105),
    .D(_02250_),
    .Q_N(_13247_),
    .Q(\cpu.icache.r_data[7][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][22]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net3106),
    .D(_02251_),
    .Q_N(_13246_),
    .Q(\cpu.icache.r_data[7][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][23]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3107),
    .D(_02252_),
    .Q_N(_13245_),
    .Q(\cpu.icache.r_data[7][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][24]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3108),
    .D(_02253_),
    .Q_N(_13244_),
    .Q(\cpu.icache.r_data[7][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][25]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3109),
    .D(_02254_),
    .Q_N(_13243_),
    .Q(\cpu.icache.r_data[7][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][26]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3110),
    .D(_02255_),
    .Q_N(_13242_),
    .Q(\cpu.icache.r_data[7][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][27]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3111),
    .D(_02256_),
    .Q_N(_13241_),
    .Q(\cpu.icache.r_data[7][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][28]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net3112),
    .D(_02257_),
    .Q_N(_13240_),
    .Q(\cpu.icache.r_data[7][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][29]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3113),
    .D(_02258_),
    .Q_N(_13239_),
    .Q(\cpu.icache.r_data[7][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net3114),
    .D(_02259_),
    .Q_N(_13238_),
    .Q(\cpu.icache.r_data[7][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][30]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net3115),
    .D(_02260_),
    .Q_N(_13237_),
    .Q(\cpu.icache.r_data[7][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][31]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3116),
    .D(_02261_),
    .Q_N(_13236_),
    .Q(\cpu.icache.r_data[7][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net3117),
    .D(_02262_),
    .Q_N(_13235_),
    .Q(\cpu.icache.r_data[7][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net3118),
    .D(_02263_),
    .Q_N(_13234_),
    .Q(\cpu.icache.r_data[7][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net3119),
    .D(_02264_),
    .Q_N(_13233_),
    .Q(\cpu.icache.r_data[7][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net3120),
    .D(_02265_),
    .Q_N(_13232_),
    .Q(\cpu.icache.r_data[7][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net3121),
    .D(_02266_),
    .Q_N(_13231_),
    .Q(\cpu.icache.r_data[7][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3122),
    .D(_02267_),
    .Q_N(_13230_),
    .Q(\cpu.icache.r_data[7][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3123),
    .D(_02268_),
    .Q_N(_13229_),
    .Q(\cpu.icache.r_data[7][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_offset[0]$_SDFF_PN0_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net3124),
    .D(_02269_),
    .Q_N(_00316_),
    .Q(\cpu.icache.r_offset[0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_offset[1]$_SDFF_PN0_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net3125),
    .D(_02270_),
    .Q_N(_13228_),
    .Q(\cpu.icache.r_offset[1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_offset[2]$_SDFF_PN0_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3126),
    .D(_02271_),
    .Q_N(_00254_),
    .Q(\cpu.icache.r_offset[2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3127),
    .D(_02272_),
    .Q_N(_13227_),
    .Q(\cpu.icache.r_tag[0][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3128),
    .D(_02273_),
    .Q_N(_13226_),
    .Q(\cpu.icache.r_tag[0][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3129),
    .D(_02274_),
    .Q_N(_13225_),
    .Q(\cpu.icache.r_tag[0][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3130),
    .D(_02275_),
    .Q_N(_13224_),
    .Q(\cpu.icache.r_tag[0][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3131),
    .D(_02276_),
    .Q_N(_13223_),
    .Q(\cpu.icache.r_tag[0][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3132),
    .D(_02277_),
    .Q_N(_13222_),
    .Q(\cpu.icache.r_tag[0][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3133),
    .D(_02278_),
    .Q_N(_13221_),
    .Q(\cpu.icache.r_tag[0][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3134),
    .D(_02279_),
    .Q_N(_13220_),
    .Q(\cpu.icache.r_tag[0][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3135),
    .D(_02280_),
    .Q_N(_13219_),
    .Q(\cpu.icache.r_tag[0][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3136),
    .D(_02281_),
    .Q_N(_13218_),
    .Q(\cpu.icache.r_tag[0][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3137),
    .D(_02282_),
    .Q_N(_13217_),
    .Q(\cpu.icache.r_tag[0][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3138),
    .D(_02283_),
    .Q_N(_13216_),
    .Q(\cpu.icache.r_tag[0][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3139),
    .D(_02284_),
    .Q_N(_13215_),
    .Q(\cpu.icache.r_tag[0][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3140),
    .D(_02285_),
    .Q_N(_13214_),
    .Q(\cpu.icache.r_tag[0][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3141),
    .D(_02286_),
    .Q_N(_13213_),
    .Q(\cpu.icache.r_tag[0][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3142),
    .D(_02287_),
    .Q_N(_13212_),
    .Q(\cpu.icache.r_tag[0][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3143),
    .D(_02288_),
    .Q_N(_13211_),
    .Q(\cpu.icache.r_tag[0][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3144),
    .D(_02289_),
    .Q_N(_13210_),
    .Q(\cpu.icache.r_tag[0][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3145),
    .D(_02290_),
    .Q_N(_13209_),
    .Q(\cpu.icache.r_tag[0][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3146),
    .D(_02291_),
    .Q_N(_13208_),
    .Q(\cpu.icache.r_tag[1][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3147),
    .D(_02292_),
    .Q_N(_13207_),
    .Q(\cpu.icache.r_tag[1][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3148),
    .D(_02293_),
    .Q_N(_13206_),
    .Q(\cpu.icache.r_tag[1][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3149),
    .D(_02294_),
    .Q_N(_13205_),
    .Q(\cpu.icache.r_tag[1][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3150),
    .D(_02295_),
    .Q_N(_13204_),
    .Q(\cpu.icache.r_tag[1][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3151),
    .D(_02296_),
    .Q_N(_13203_),
    .Q(\cpu.icache.r_tag[1][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3152),
    .D(_02297_),
    .Q_N(_13202_),
    .Q(\cpu.icache.r_tag[1][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3153),
    .D(_02298_),
    .Q_N(_13201_),
    .Q(\cpu.icache.r_tag[1][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3154),
    .D(_02299_),
    .Q_N(_13200_),
    .Q(\cpu.icache.r_tag[1][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3155),
    .D(_02300_),
    .Q_N(_13199_),
    .Q(\cpu.icache.r_tag[1][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3156),
    .D(_02301_),
    .Q_N(_13198_),
    .Q(\cpu.icache.r_tag[1][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3157),
    .D(_02302_),
    .Q_N(_13197_),
    .Q(\cpu.icache.r_tag[1][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3158),
    .D(_02303_),
    .Q_N(_13196_),
    .Q(\cpu.icache.r_tag[1][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3159),
    .D(_02304_),
    .Q_N(_13195_),
    .Q(\cpu.icache.r_tag[1][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3160),
    .D(_02305_),
    .Q_N(_13194_),
    .Q(\cpu.icache.r_tag[1][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3161),
    .D(_02306_),
    .Q_N(_13193_),
    .Q(\cpu.icache.r_tag[1][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3162),
    .D(_02307_),
    .Q_N(_13192_),
    .Q(\cpu.icache.r_tag[1][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3163),
    .D(_02308_),
    .Q_N(_13191_),
    .Q(\cpu.icache.r_tag[1][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3164),
    .D(_02309_),
    .Q_N(_13190_),
    .Q(\cpu.icache.r_tag[1][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3165),
    .D(_02310_),
    .Q_N(_13189_),
    .Q(\cpu.icache.r_tag[2][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3166),
    .D(_02311_),
    .Q_N(_13188_),
    .Q(\cpu.icache.r_tag[2][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3167),
    .D(_02312_),
    .Q_N(_13187_),
    .Q(\cpu.icache.r_tag[2][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3168),
    .D(_02313_),
    .Q_N(_13186_),
    .Q(\cpu.icache.r_tag[2][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3169),
    .D(_02314_),
    .Q_N(_13185_),
    .Q(\cpu.icache.r_tag[2][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3170),
    .D(_02315_),
    .Q_N(_13184_),
    .Q(\cpu.icache.r_tag[2][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3171),
    .D(_02316_),
    .Q_N(_13183_),
    .Q(\cpu.icache.r_tag[2][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3172),
    .D(_02317_),
    .Q_N(_13182_),
    .Q(\cpu.icache.r_tag[2][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3173),
    .D(_02318_),
    .Q_N(_13181_),
    .Q(\cpu.icache.r_tag[2][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3174),
    .D(_02319_),
    .Q_N(_13180_),
    .Q(\cpu.icache.r_tag[2][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3175),
    .D(_02320_),
    .Q_N(_13179_),
    .Q(\cpu.icache.r_tag[2][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3176),
    .D(_02321_),
    .Q_N(_13178_),
    .Q(\cpu.icache.r_tag[2][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3177),
    .D(_02322_),
    .Q_N(_13177_),
    .Q(\cpu.icache.r_tag[2][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3178),
    .D(_02323_),
    .Q_N(_13176_),
    .Q(\cpu.icache.r_tag[2][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3179),
    .D(_02324_),
    .Q_N(_13175_),
    .Q(\cpu.icache.r_tag[2][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3180),
    .D(_02325_),
    .Q_N(_13174_),
    .Q(\cpu.icache.r_tag[2][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3181),
    .D(_02326_),
    .Q_N(_13173_),
    .Q(\cpu.icache.r_tag[2][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3182),
    .D(_02327_),
    .Q_N(_13172_),
    .Q(\cpu.icache.r_tag[2][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3183),
    .D(_02328_),
    .Q_N(_13171_),
    .Q(\cpu.icache.r_tag[2][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3184),
    .D(_02329_),
    .Q_N(_13170_),
    .Q(\cpu.icache.r_tag[3][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3185),
    .D(_02330_),
    .Q_N(_13169_),
    .Q(\cpu.icache.r_tag[3][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3186),
    .D(_02331_),
    .Q_N(_13168_),
    .Q(\cpu.icache.r_tag[3][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3187),
    .D(_02332_),
    .Q_N(_13167_),
    .Q(\cpu.icache.r_tag[3][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3188),
    .D(_02333_),
    .Q_N(_13166_),
    .Q(\cpu.icache.r_tag[3][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3189),
    .D(_02334_),
    .Q_N(_13165_),
    .Q(\cpu.icache.r_tag[3][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3190),
    .D(_02335_),
    .Q_N(_13164_),
    .Q(\cpu.icache.r_tag[3][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3191),
    .D(_02336_),
    .Q_N(_13163_),
    .Q(\cpu.icache.r_tag[3][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3192),
    .D(_02337_),
    .Q_N(_13162_),
    .Q(\cpu.icache.r_tag[3][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3193),
    .D(_02338_),
    .Q_N(_13161_),
    .Q(\cpu.icache.r_tag[3][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3194),
    .D(_02339_),
    .Q_N(_13160_),
    .Q(\cpu.icache.r_tag[3][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3195),
    .D(_02340_),
    .Q_N(_13159_),
    .Q(\cpu.icache.r_tag[3][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3196),
    .D(_02341_),
    .Q_N(_13158_),
    .Q(\cpu.icache.r_tag[3][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3197),
    .D(_02342_),
    .Q_N(_13157_),
    .Q(\cpu.icache.r_tag[3][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3198),
    .D(_02343_),
    .Q_N(_13156_),
    .Q(\cpu.icache.r_tag[3][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3199),
    .D(_02344_),
    .Q_N(_13155_),
    .Q(\cpu.icache.r_tag[3][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3200),
    .D(_02345_),
    .Q_N(_13154_),
    .Q(\cpu.icache.r_tag[3][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3201),
    .D(_02346_),
    .Q_N(_13153_),
    .Q(\cpu.icache.r_tag[3][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3202),
    .D(_02347_),
    .Q_N(_13152_),
    .Q(\cpu.icache.r_tag[3][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3203),
    .D(_02348_),
    .Q_N(_13151_),
    .Q(\cpu.icache.r_tag[4][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3204),
    .D(_02349_),
    .Q_N(_13150_),
    .Q(\cpu.icache.r_tag[4][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3205),
    .D(_02350_),
    .Q_N(_13149_),
    .Q(\cpu.icache.r_tag[4][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3206),
    .D(_02351_),
    .Q_N(_13148_),
    .Q(\cpu.icache.r_tag[4][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3207),
    .D(_02352_),
    .Q_N(_13147_),
    .Q(\cpu.icache.r_tag[4][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3208),
    .D(_02353_),
    .Q_N(_13146_),
    .Q(\cpu.icache.r_tag[4][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3209),
    .D(_02354_),
    .Q_N(_13145_),
    .Q(\cpu.icache.r_tag[4][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3210),
    .D(_02355_),
    .Q_N(_13144_),
    .Q(\cpu.icache.r_tag[4][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3211),
    .D(_02356_),
    .Q_N(_13143_),
    .Q(\cpu.icache.r_tag[4][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3212),
    .D(_02357_),
    .Q_N(_13142_),
    .Q(\cpu.icache.r_tag[4][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3213),
    .D(_02358_),
    .Q_N(_13141_),
    .Q(\cpu.icache.r_tag[4][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3214),
    .D(_02359_),
    .Q_N(_13140_),
    .Q(\cpu.icache.r_tag[4][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3215),
    .D(_02360_),
    .Q_N(_13139_),
    .Q(\cpu.icache.r_tag[4][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3216),
    .D(_02361_),
    .Q_N(_13138_),
    .Q(\cpu.icache.r_tag[4][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3217),
    .D(_02362_),
    .Q_N(_13137_),
    .Q(\cpu.icache.r_tag[4][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3218),
    .D(_02363_),
    .Q_N(_13136_),
    .Q(\cpu.icache.r_tag[4][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3219),
    .D(_02364_),
    .Q_N(_13135_),
    .Q(\cpu.icache.r_tag[4][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3220),
    .D(_02365_),
    .Q_N(_13134_),
    .Q(\cpu.icache.r_tag[4][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3221),
    .D(_02366_),
    .Q_N(_13133_),
    .Q(\cpu.icache.r_tag[4][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3222),
    .D(_02367_),
    .Q_N(_13132_),
    .Q(\cpu.icache.r_tag[5][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3223),
    .D(_02368_),
    .Q_N(_13131_),
    .Q(\cpu.icache.r_tag[5][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3224),
    .D(_02369_),
    .Q_N(_13130_),
    .Q(\cpu.icache.r_tag[5][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3225),
    .D(_02370_),
    .Q_N(_13129_),
    .Q(\cpu.icache.r_tag[5][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3226),
    .D(_02371_),
    .Q_N(_13128_),
    .Q(\cpu.icache.r_tag[5][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3227),
    .D(_02372_),
    .Q_N(_13127_),
    .Q(\cpu.icache.r_tag[5][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3228),
    .D(_02373_),
    .Q_N(_13126_),
    .Q(\cpu.icache.r_tag[5][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3229),
    .D(_02374_),
    .Q_N(_13125_),
    .Q(\cpu.icache.r_tag[5][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3230),
    .D(_02375_),
    .Q_N(_13124_),
    .Q(\cpu.icache.r_tag[5][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3231),
    .D(_02376_),
    .Q_N(_13123_),
    .Q(\cpu.icache.r_tag[5][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3232),
    .D(_02377_),
    .Q_N(_13122_),
    .Q(\cpu.icache.r_tag[5][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3233),
    .D(_02378_),
    .Q_N(_13121_),
    .Q(\cpu.icache.r_tag[5][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3234),
    .D(_02379_),
    .Q_N(_13120_),
    .Q(\cpu.icache.r_tag[5][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3235),
    .D(_02380_),
    .Q_N(_13119_),
    .Q(\cpu.icache.r_tag[5][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3236),
    .D(_02381_),
    .Q_N(_13118_),
    .Q(\cpu.icache.r_tag[5][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3237),
    .D(_02382_),
    .Q_N(_13117_),
    .Q(\cpu.icache.r_tag[5][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3238),
    .D(_02383_),
    .Q_N(_13116_),
    .Q(\cpu.icache.r_tag[5][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3239),
    .D(_02384_),
    .Q_N(_13115_),
    .Q(\cpu.icache.r_tag[5][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3240),
    .D(_02385_),
    .Q_N(_13114_),
    .Q(\cpu.icache.r_tag[5][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3241),
    .D(_02386_),
    .Q_N(_13113_),
    .Q(\cpu.icache.r_tag[6][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3242),
    .D(_02387_),
    .Q_N(_13112_),
    .Q(\cpu.icache.r_tag[6][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3243),
    .D(_02388_),
    .Q_N(_13111_),
    .Q(\cpu.icache.r_tag[6][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3244),
    .D(_02389_),
    .Q_N(_13110_),
    .Q(\cpu.icache.r_tag[6][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3245),
    .D(_02390_),
    .Q_N(_13109_),
    .Q(\cpu.icache.r_tag[6][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3246),
    .D(_02391_),
    .Q_N(_13108_),
    .Q(\cpu.icache.r_tag[6][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3247),
    .D(_02392_),
    .Q_N(_13107_),
    .Q(\cpu.icache.r_tag[6][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3248),
    .D(_02393_),
    .Q_N(_13106_),
    .Q(\cpu.icache.r_tag[6][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3249),
    .D(_02394_),
    .Q_N(_13105_),
    .Q(\cpu.icache.r_tag[6][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3250),
    .D(_02395_),
    .Q_N(_13104_),
    .Q(\cpu.icache.r_tag[6][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3251),
    .D(_02396_),
    .Q_N(_13103_),
    .Q(\cpu.icache.r_tag[6][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3252),
    .D(_02397_),
    .Q_N(_13102_),
    .Q(\cpu.icache.r_tag[6][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3253),
    .D(_02398_),
    .Q_N(_13101_),
    .Q(\cpu.icache.r_tag[6][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3254),
    .D(_02399_),
    .Q_N(_13100_),
    .Q(\cpu.icache.r_tag[6][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3255),
    .D(_02400_),
    .Q_N(_13099_),
    .Q(\cpu.icache.r_tag[6][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3256),
    .D(_02401_),
    .Q_N(_13098_),
    .Q(\cpu.icache.r_tag[6][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3257),
    .D(_02402_),
    .Q_N(_13097_),
    .Q(\cpu.icache.r_tag[6][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3258),
    .D(_02403_),
    .Q_N(_13096_),
    .Q(\cpu.icache.r_tag[6][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3259),
    .D(_02404_),
    .Q_N(_13095_),
    .Q(\cpu.icache.r_tag[6][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3260),
    .D(_02405_),
    .Q_N(_13094_),
    .Q(\cpu.icache.r_tag[7][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3261),
    .D(_02406_),
    .Q_N(_13093_),
    .Q(\cpu.icache.r_tag[7][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3262),
    .D(_02407_),
    .Q_N(_13092_),
    .Q(\cpu.icache.r_tag[7][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3263),
    .D(_02408_),
    .Q_N(_13091_),
    .Q(\cpu.icache.r_tag[7][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3264),
    .D(_02409_),
    .Q_N(_13090_),
    .Q(\cpu.icache.r_tag[7][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3265),
    .D(_02410_),
    .Q_N(_13089_),
    .Q(\cpu.icache.r_tag[7][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3266),
    .D(_02411_),
    .Q_N(_13088_),
    .Q(\cpu.icache.r_tag[7][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3267),
    .D(_02412_),
    .Q_N(_13087_),
    .Q(\cpu.icache.r_tag[7][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3268),
    .D(_02413_),
    .Q_N(_13086_),
    .Q(\cpu.icache.r_tag[7][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3269),
    .D(_02414_),
    .Q_N(_13085_),
    .Q(\cpu.icache.r_tag[7][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3270),
    .D(_02415_),
    .Q_N(_13084_),
    .Q(\cpu.icache.r_tag[7][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3271),
    .D(_02416_),
    .Q_N(_13083_),
    .Q(\cpu.icache.r_tag[7][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3272),
    .D(_02417_),
    .Q_N(_13082_),
    .Q(\cpu.icache.r_tag[7][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3273),
    .D(_02418_),
    .Q_N(_13081_),
    .Q(\cpu.icache.r_tag[7][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3274),
    .D(_02419_),
    .Q_N(_13080_),
    .Q(\cpu.icache.r_tag[7][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3275),
    .D(_02420_),
    .Q_N(_13079_),
    .Q(\cpu.icache.r_tag[7][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3276),
    .D(_02421_),
    .Q_N(_13078_),
    .Q(\cpu.icache.r_tag[7][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3277),
    .D(_02422_),
    .Q_N(_13077_),
    .Q(\cpu.icache.r_tag[7][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3278),
    .D(_02423_),
    .Q_N(_13076_),
    .Q(\cpu.icache.r_tag[7][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3279),
    .D(_02424_),
    .Q_N(_13075_),
    .Q(\cpu.icache.r_valid[0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net3280),
    .D(_02425_),
    .Q_N(_13074_),
    .Q(\cpu.icache.r_valid[1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net3281),
    .D(_02426_),
    .Q_N(_13073_),
    .Q(\cpu.icache.r_valid[2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3282),
    .D(_02427_),
    .Q_N(_13072_),
    .Q(\cpu.icache.r_valid[3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3283),
    .D(_02428_),
    .Q_N(_13071_),
    .Q(\cpu.icache.r_valid[4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3284),
    .D(_02429_),
    .Q_N(_13070_),
    .Q(\cpu.icache.r_valid[5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3285),
    .D(_02430_),
    .Q_N(_13069_),
    .Q(\cpu.icache.r_valid[6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3286),
    .D(_02431_),
    .Q_N(_13068_),
    .Q(\cpu.icache.r_valid[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3287),
    .D(_02432_),
    .Q_N(_13067_),
    .Q(\cpu.intr.r_clock ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[0]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3288),
    .D(_02433_),
    .Q_N(_13066_),
    .Q(\cpu.intr.r_clock_cmp[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[10]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net3289),
    .D(_02434_),
    .Q_N(_13065_),
    .Q(\cpu.intr.r_clock_cmp[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[11]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3290),
    .D(_02435_),
    .Q_N(_13064_),
    .Q(\cpu.intr.r_clock_cmp[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[12]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3291),
    .D(_02436_),
    .Q_N(_13063_),
    .Q(\cpu.intr.r_clock_cmp[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[13]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3292),
    .D(_02437_),
    .Q_N(_13062_),
    .Q(\cpu.intr.r_clock_cmp[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[14]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3293),
    .D(_02438_),
    .Q_N(_13061_),
    .Q(\cpu.intr.r_clock_cmp[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[15]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net3294),
    .D(_02439_),
    .Q_N(_13060_),
    .Q(\cpu.intr.r_clock_cmp[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[16]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3295),
    .D(_02440_),
    .Q_N(_13059_),
    .Q(\cpu.intr.r_clock_cmp[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[17]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3296),
    .D(_02441_),
    .Q_N(_13058_),
    .Q(\cpu.intr.r_clock_cmp[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[18]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3297),
    .D(_02442_),
    .Q_N(_13057_),
    .Q(\cpu.intr.r_clock_cmp[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[19]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3298),
    .D(_02443_),
    .Q_N(_13056_),
    .Q(\cpu.intr.r_clock_cmp[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[1]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3299),
    .D(_02444_),
    .Q_N(_13055_),
    .Q(\cpu.intr.r_clock_cmp[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[20]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3300),
    .D(_02445_),
    .Q_N(_13054_),
    .Q(\cpu.intr.r_clock_cmp[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[21]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3301),
    .D(_02446_),
    .Q_N(_13053_),
    .Q(\cpu.intr.r_clock_cmp[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[22]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3302),
    .D(_02447_),
    .Q_N(_13052_),
    .Q(\cpu.intr.r_clock_cmp[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[23]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3303),
    .D(_02448_),
    .Q_N(_13051_),
    .Q(\cpu.intr.r_clock_cmp[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[24]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3304),
    .D(_02449_),
    .Q_N(_13050_),
    .Q(\cpu.intr.r_clock_cmp[24] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[25]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3305),
    .D(_02450_),
    .Q_N(_13049_),
    .Q(\cpu.intr.r_clock_cmp[25] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[26]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net3306),
    .D(_02451_),
    .Q_N(_13048_),
    .Q(\cpu.intr.r_clock_cmp[26] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[27]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3307),
    .D(_02452_),
    .Q_N(_13047_),
    .Q(\cpu.intr.r_clock_cmp[27] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[28]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3308),
    .D(_02453_),
    .Q_N(_13046_),
    .Q(\cpu.intr.r_clock_cmp[28] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[29]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3309),
    .D(_02454_),
    .Q_N(_13045_),
    .Q(\cpu.intr.r_clock_cmp[29] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[2]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3310),
    .D(_02455_),
    .Q_N(_13044_),
    .Q(\cpu.intr.r_clock_cmp[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[30]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3311),
    .D(_02456_),
    .Q_N(_13043_),
    .Q(\cpu.intr.r_clock_cmp[30] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[31]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net3312),
    .D(_02457_),
    .Q_N(_13042_),
    .Q(\cpu.intr.r_clock_cmp[31] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[3]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3313),
    .D(_02458_),
    .Q_N(_13041_),
    .Q(\cpu.intr.r_clock_cmp[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[4]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3314),
    .D(_02459_),
    .Q_N(_13040_),
    .Q(\cpu.intr.r_clock_cmp[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[5]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3315),
    .D(_02460_),
    .Q_N(_13039_),
    .Q(\cpu.intr.r_clock_cmp[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[6]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3316),
    .D(_02461_),
    .Q_N(_13038_),
    .Q(\cpu.intr.r_clock_cmp[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[7]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3317),
    .D(_02462_),
    .Q_N(_13037_),
    .Q(\cpu.intr.r_clock_cmp[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[8]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3318),
    .D(_02463_),
    .Q_N(_13036_),
    .Q(\cpu.intr.r_clock_cmp[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[9]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3319),
    .D(_02464_),
    .Q_N(_15028_),
    .Q(\cpu.intr.r_clock_cmp[9] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[0]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3320),
    .D(_00036_),
    .Q_N(_00286_),
    .Q(\cpu.intr.r_clock_count[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[10]$_DFF_P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3321),
    .D(_00037_),
    .Q_N(_15029_),
    .Q(\cpu.intr.r_clock_count[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[11]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3322),
    .D(_00038_),
    .Q_N(_15030_),
    .Q(\cpu.intr.r_clock_count[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[12]$_DFF_P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3323),
    .D(_00039_),
    .Q_N(_15031_),
    .Q(\cpu.intr.r_clock_count[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[13]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3324),
    .D(_00040_),
    .Q_N(_15032_),
    .Q(\cpu.intr.r_clock_count[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[14]$_DFF_P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3325),
    .D(_00041_),
    .Q_N(_15033_),
    .Q(\cpu.intr.r_clock_count[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[15]$_DFF_P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3326),
    .D(_00042_),
    .Q_N(_13035_),
    .Q(\cpu.intr.r_clock_count[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[16]$_DFFE_PN_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net3327),
    .D(_02465_),
    .Q_N(_13034_),
    .Q(\cpu.intr.r_clock_count[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[17]$_DFFE_PN_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3328),
    .D(_02466_),
    .Q_N(_13033_),
    .Q(\cpu.intr.r_clock_count[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[18]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3329),
    .D(_02467_),
    .Q_N(_13032_),
    .Q(\cpu.intr.r_clock_count[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[19]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3330),
    .D(_02468_),
    .Q_N(_15034_),
    .Q(\cpu.intr.r_clock_count[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[1]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3331),
    .D(_00043_),
    .Q_N(_13031_),
    .Q(\cpu.intr.r_clock_count[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[20]$_DFFE_PN_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3332),
    .D(_02469_),
    .Q_N(_13030_),
    .Q(\cpu.intr.r_clock_count[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[21]$_DFFE_PN_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3333),
    .D(_02470_),
    .Q_N(_13029_),
    .Q(\cpu.intr.r_clock_count[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[22]$_DFFE_PN_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3334),
    .D(_02471_),
    .Q_N(_13028_),
    .Q(\cpu.intr.r_clock_count[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[23]$_DFFE_PN_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3335),
    .D(_02472_),
    .Q_N(_13027_),
    .Q(\cpu.intr.r_clock_count[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[24]$_DFFE_PN_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3336),
    .D(_02473_),
    .Q_N(_13026_),
    .Q(\cpu.intr.r_clock_count[24] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[25]$_DFFE_PN_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3337),
    .D(_02474_),
    .Q_N(_13025_),
    .Q(\cpu.intr.r_clock_count[25] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[26]$_DFFE_PN_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3338),
    .D(_02475_),
    .Q_N(_13024_),
    .Q(\cpu.intr.r_clock_count[26] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[27]$_DFFE_PN_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3339),
    .D(_02476_),
    .Q_N(_13023_),
    .Q(\cpu.intr.r_clock_count[27] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[28]$_DFFE_PN_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3340),
    .D(_02477_),
    .Q_N(_13022_),
    .Q(\cpu.intr.r_clock_count[28] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[29]$_DFFE_PN_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3341),
    .D(_02478_),
    .Q_N(_15035_),
    .Q(\cpu.intr.r_clock_count[29] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[2]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3342),
    .D(_00044_),
    .Q_N(_13021_),
    .Q(\cpu.intr.r_clock_count[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[30]$_DFFE_PN_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3343),
    .D(_02479_),
    .Q_N(_13020_),
    .Q(\cpu.intr.r_clock_count[30] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[31]$_DFFE_PN_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3344),
    .D(_02480_),
    .Q_N(_15036_),
    .Q(\cpu.intr.r_clock_count[31] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[3]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3345),
    .D(_00045_),
    .Q_N(_15037_),
    .Q(\cpu.intr.r_clock_count[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[4]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3346),
    .D(_00046_),
    .Q_N(_15038_),
    .Q(\cpu.intr.r_clock_count[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[5]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3347),
    .D(_00047_),
    .Q_N(_15039_),
    .Q(\cpu.intr.r_clock_count[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[6]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3348),
    .D(_00048_),
    .Q_N(_15040_),
    .Q(\cpu.intr.r_clock_count[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[7]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3349),
    .D(_00049_),
    .Q_N(_15041_),
    .Q(\cpu.intr.r_clock_count[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[8]$_DFF_P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3350),
    .D(_00050_),
    .Q_N(_15042_),
    .Q(\cpu.intr.r_clock_count[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[9]$_DFF_P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3351),
    .D(_00051_),
    .Q_N(_13019_),
    .Q(\cpu.intr.r_clock_count[9] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3352),
    .D(_02481_),
    .Q_N(_13018_),
    .Q(\cpu.intr.r_enable[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3353),
    .D(_02482_),
    .Q_N(_13017_),
    .Q(\cpu.intr.r_enable[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3354),
    .D(_02483_),
    .Q_N(_13016_),
    .Q(\cpu.intr.r_enable[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3355),
    .D(_02484_),
    .Q_N(_13015_),
    .Q(\cpu.intr.r_enable[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3356),
    .D(_02485_),
    .Q_N(_13014_),
    .Q(\cpu.intr.r_enable[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3357),
    .D(_02486_),
    .Q_N(_13013_),
    .Q(\cpu.intr.r_enable[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3358),
    .D(_02487_),
    .Q_N(_15043_),
    .Q(\cpu.intr.r_timer ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[0]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3359),
    .D(_00055_),
    .Q_N(_00285_),
    .Q(\cpu.intr.r_timer_count[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[10]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3360),
    .D(_00056_),
    .Q_N(_15044_),
    .Q(\cpu.intr.r_timer_count[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[11]$_DFF_P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net3361),
    .D(_00057_),
    .Q_N(_15045_),
    .Q(\cpu.intr.r_timer_count[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[12]$_DFF_P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net3362),
    .D(_00058_),
    .Q_N(_15046_),
    .Q(\cpu.intr.r_timer_count[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[13]$_DFF_P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net3363),
    .D(_00059_),
    .Q_N(_15047_),
    .Q(\cpu.intr.r_timer_count[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[14]$_DFF_P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net3364),
    .D(_00060_),
    .Q_N(_15048_),
    .Q(\cpu.intr.r_timer_count[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[15]$_DFF_P_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net3365),
    .D(_00061_),
    .Q_N(_15049_),
    .Q(\cpu.intr.r_timer_count[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[16]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net3366),
    .D(_00062_),
    .Q_N(_15050_),
    .Q(\cpu.intr.r_timer_count[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[17]$_DFF_P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3367),
    .D(_00063_),
    .Q_N(_15051_),
    .Q(\cpu.intr.r_timer_count[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[18]$_DFF_P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3368),
    .D(_00064_),
    .Q_N(_15052_),
    .Q(\cpu.intr.r_timer_count[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[19]$_DFF_P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3369),
    .D(_00065_),
    .Q_N(_15053_),
    .Q(\cpu.intr.r_timer_count[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[1]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net3370),
    .D(_00066_),
    .Q_N(_15054_),
    .Q(\cpu.intr.r_timer_count[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[20]$_DFF_P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3371),
    .D(_00067_),
    .Q_N(_15055_),
    .Q(\cpu.intr.r_timer_count[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[21]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net3372),
    .D(_00068_),
    .Q_N(_15056_),
    .Q(\cpu.intr.r_timer_count[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[22]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net3373),
    .D(_00069_),
    .Q_N(_15057_),
    .Q(\cpu.intr.r_timer_count[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[23]$_DFF_P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3374),
    .D(_00070_),
    .Q_N(_15058_),
    .Q(\cpu.intr.r_timer_count[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[2]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net3375),
    .D(_00071_),
    .Q_N(_15059_),
    .Q(\cpu.intr.r_timer_count[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[3]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net3376),
    .D(_00072_),
    .Q_N(_15060_),
    .Q(\cpu.intr.r_timer_count[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[4]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net3377),
    .D(_00073_),
    .Q_N(_15061_),
    .Q(\cpu.intr.r_timer_count[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[5]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3378),
    .D(_00074_),
    .Q_N(_15062_),
    .Q(\cpu.intr.r_timer_count[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[6]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3379),
    .D(_00075_),
    .Q_N(_15063_),
    .Q(\cpu.intr.r_timer_count[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[7]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3380),
    .D(_00076_),
    .Q_N(_15064_),
    .Q(\cpu.intr.r_timer_count[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[8]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3381),
    .D(_00077_),
    .Q_N(_15065_),
    .Q(\cpu.intr.r_timer_count[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[9]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3382),
    .D(_00078_),
    .Q_N(_13012_),
    .Q(\cpu.intr.r_timer_count[9] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[0]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3383),
    .D(_02488_),
    .Q_N(_13011_),
    .Q(\cpu.intr.r_timer_reload[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[10]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net3384),
    .D(_02489_),
    .Q_N(_13010_),
    .Q(\cpu.intr.r_timer_reload[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[11]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net3385),
    .D(_02490_),
    .Q_N(_13009_),
    .Q(\cpu.intr.r_timer_reload[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[12]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net3386),
    .D(_02491_),
    .Q_N(_13008_),
    .Q(\cpu.intr.r_timer_reload[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[13]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net3387),
    .D(_02492_),
    .Q_N(_13007_),
    .Q(\cpu.intr.r_timer_reload[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[14]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net3388),
    .D(_02493_),
    .Q_N(_13006_),
    .Q(\cpu.intr.r_timer_reload[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[15]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net3389),
    .D(_02494_),
    .Q_N(_13005_),
    .Q(\cpu.intr.r_timer_reload[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[16]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net3390),
    .D(_02495_),
    .Q_N(_13004_),
    .Q(\cpu.intr.r_timer_reload[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[17]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3391),
    .D(_02496_),
    .Q_N(_13003_),
    .Q(\cpu.intr.r_timer_reload[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[18]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3392),
    .D(_02497_),
    .Q_N(_13002_),
    .Q(\cpu.intr.r_timer_reload[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[19]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3393),
    .D(_02498_),
    .Q_N(_13001_),
    .Q(\cpu.intr.r_timer_reload[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[1]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3394),
    .D(_02499_),
    .Q_N(_13000_),
    .Q(\cpu.intr.r_timer_reload[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[20]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3395),
    .D(_02500_),
    .Q_N(_12999_),
    .Q(\cpu.intr.r_timer_reload[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[21]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3396),
    .D(_02501_),
    .Q_N(_12998_),
    .Q(\cpu.intr.r_timer_reload[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[22]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net3397),
    .D(_02502_),
    .Q_N(_12997_),
    .Q(\cpu.intr.r_timer_reload[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[23]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3398),
    .D(_02503_),
    .Q_N(_12996_),
    .Q(\cpu.intr.r_timer_reload[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[2]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3399),
    .D(_02504_),
    .Q_N(_12995_),
    .Q(\cpu.intr.r_timer_reload[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[3]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3400),
    .D(_02505_),
    .Q_N(_12994_),
    .Q(\cpu.intr.r_timer_reload[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[4]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3401),
    .D(_02506_),
    .Q_N(_12993_),
    .Q(\cpu.intr.r_timer_reload[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[5]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3402),
    .D(_02507_),
    .Q_N(_12992_),
    .Q(\cpu.intr.r_timer_reload[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[6]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3403),
    .D(_02508_),
    .Q_N(_12991_),
    .Q(\cpu.intr.r_timer_reload[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[7]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3404),
    .D(_02509_),
    .Q_N(_12990_),
    .Q(\cpu.intr.r_timer_reload[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[8]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3405),
    .D(_02510_),
    .Q_N(_12989_),
    .Q(\cpu.intr.r_timer_reload[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[9]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3406),
    .D(_02511_),
    .Q_N(_12988_),
    .Q(\cpu.intr.r_timer_reload[9] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[0]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3407),
    .D(_02512_),
    .Q_N(_00183_),
    .Q(\cpu.qspi.r_count[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[1]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3408),
    .D(_02513_),
    .Q_N(_12987_),
    .Q(\cpu.qspi.r_count[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[2]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3409),
    .D(_02514_),
    .Q_N(_00184_),
    .Q(\cpu.qspi.r_count[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[3]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3410),
    .D(_02515_),
    .Q_N(_12986_),
    .Q(\cpu.qspi.r_count[3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[4]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3411),
    .D(_02516_),
    .Q_N(_00252_),
    .Q(\cpu.qspi.r_count[4] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_cs[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3412),
    .D(_02517_),
    .Q_N(_12985_),
    .Q(net19));
 sg13g2_dfrbp_1 \cpu.qspi.r_cs[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3413),
    .D(_02518_),
    .Q_N(_12984_),
    .Q(net20));
 sg13g2_dfrbp_1 \cpu.qspi.r_cs[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net3414),
    .D(_02519_),
    .Q_N(_12983_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[11] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_ind$_SDFFE_PN0N_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3415),
    .D(_02520_),
    .Q_N(_12982_),
    .Q(\cpu.qspi.r_ind ));
 sg13g2_dfrbp_1 \cpu.qspi.r_mask[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3416),
    .D(_02521_),
    .Q_N(_12981_),
    .Q(\cpu.qspi.r_mask[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_mask[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3417),
    .D(_02522_),
    .Q_N(_12980_),
    .Q(\cpu.qspi.r_mask[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_mask[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3418),
    .D(_02523_),
    .Q_N(_12979_),
    .Q(\cpu.qspi.r_mask[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_quad[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3419),
    .D(_02524_),
    .Q_N(_12978_),
    .Q(\cpu.qspi.r_quad[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_quad[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3420),
    .D(_02525_),
    .Q_N(_12977_),
    .Q(\cpu.qspi.r_quad[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_quad[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3421),
    .D(_02526_),
    .Q_N(_12976_),
    .Q(\cpu.qspi.r_quad[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3422),
    .D(_02527_),
    .Q_N(_12975_),
    .Q(\cpu.qspi.r_read_delay[0][0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3423),
    .D(_02528_),
    .Q_N(_12974_),
    .Q(\cpu.qspi.r_read_delay[0][1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][2]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3424),
    .D(_02529_),
    .Q_N(_12973_),
    .Q(\cpu.qspi.r_read_delay[0][2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3425),
    .D(_02530_),
    .Q_N(_12972_),
    .Q(\cpu.qspi.r_read_delay[0][3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3426),
    .D(_02531_),
    .Q_N(_12971_),
    .Q(\cpu.qspi.r_read_delay[1][0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3427),
    .D(_02532_),
    .Q_N(_12970_),
    .Q(\cpu.qspi.r_read_delay[1][1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][2]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3428),
    .D(_02533_),
    .Q_N(_12969_),
    .Q(\cpu.qspi.r_read_delay[1][2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3429),
    .D(_02534_),
    .Q_N(_12968_),
    .Q(\cpu.qspi.r_read_delay[1][3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3430),
    .D(_02535_),
    .Q_N(_12967_),
    .Q(\cpu.qspi.r_read_delay[2][0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3431),
    .D(_02536_),
    .Q_N(_12966_),
    .Q(\cpu.qspi.r_read_delay[2][1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][2]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3432),
    .D(_02537_),
    .Q_N(_12965_),
    .Q(\cpu.qspi.r_read_delay[2][2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3433),
    .D(_02538_),
    .Q_N(_12964_),
    .Q(\cpu.qspi.r_read_delay[2][3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_rom_mode[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3434),
    .D(_02539_),
    .Q_N(_12963_),
    .Q(\cpu.qspi.r_rom_mode[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_rom_mode[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3435),
    .D(_02540_),
    .Q_N(_15066_),
    .Q(\cpu.qspi.r_rom_mode[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_rstrobe_d$_DFF_P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net3436),
    .D(\cpu.qspi.c_rstrobe_d ),
    .Q_N(_15067_),
    .Q(\cpu.d_rstrobe_d ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[0]$_DFF_P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3437),
    .D(_00021_),
    .Q_N(_00277_),
    .Q(\cpu.qspi.r_state[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[10]$_DFF_P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3438),
    .D(_00008_),
    .Q_N(_15068_),
    .Q(\cpu.qspi.r_state[10] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[11]$_DFF_P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3439),
    .D(_00022_),
    .Q_N(_15069_),
    .Q(\cpu.qspi.r_state[11] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[12]$_DFF_P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3440),
    .D(_00023_),
    .Q_N(_15070_),
    .Q(\cpu.qspi.r_state[12] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[13]$_DFF_P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net3441),
    .D(_00009_),
    .Q_N(_15071_),
    .Q(\cpu.qspi.r_state[13] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[14]$_DFF_P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3442),
    .D(_00024_),
    .Q_N(_15072_),
    .Q(\cpu.qspi.r_state[14] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[15]$_DFF_P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net3443),
    .D(_00010_),
    .Q_N(_15073_),
    .Q(\cpu.qspi.r_state[15] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[16]$_DFF_P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3444),
    .D(_00025_),
    .Q_N(_15074_),
    .Q(\cpu.qspi.r_state[16] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[17]$_DFF_P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3445),
    .D(_00026_),
    .Q_N(_15075_),
    .Q(\cpu.qspi.r_state[17] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[1]$_DFF_P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net3446),
    .D(_00001_),
    .Q_N(_15076_),
    .Q(\cpu.qspi.r_state[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[2]$_DFF_P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3447),
    .D(_00027_),
    .Q_N(_15077_),
    .Q(\cpu.qspi.r_state[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[3]$_DFF_P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net3448),
    .D(_00002_),
    .Q_N(_15078_),
    .Q(\cpu.qspi.r_state[3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[4]$_DFF_P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3449),
    .D(_00028_),
    .Q_N(_15079_),
    .Q(\cpu.qspi.r_state[4] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[5]$_DFF_P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3450),
    .D(_00003_),
    .Q_N(_15080_),
    .Q(\cpu.qspi.r_state[5] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[6]$_DFF_P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3451),
    .D(_00004_),
    .Q_N(_15081_),
    .Q(\cpu.qspi.r_state[6] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[7]$_DFF_P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3452),
    .D(_00005_),
    .Q_N(_15082_),
    .Q(\cpu.qspi.r_state[7] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[8]$_DFF_P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net3453),
    .D(_00006_),
    .Q_N(_00185_),
    .Q(\cpu.qspi.r_state[8] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[9]$_DFF_P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3454),
    .D(_00007_),
    .Q_N(_12962_),
    .Q(\cpu.qspi.r_state[9] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_oe[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3455),
    .D(_02541_),
    .Q_N(_12961_),
    .Q(net3));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_oe[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3456),
    .D(_02542_),
    .Q_N(_12960_),
    .Q(net6));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3457),
    .D(_02543_),
    .Q_N(_12959_),
    .Q(net11));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3458),
    .D(_02544_),
    .Q_N(_12958_),
    .Q(net12));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3459),
    .D(_02545_),
    .Q_N(_12957_),
    .Q(net13));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3460),
    .D(_02546_),
    .Q_N(_15083_),
    .Q(net14));
 sg13g2_dfrbp_1 \cpu.qspi.r_wstrobe_d$_DFF_P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net3461),
    .D(\cpu.qspi.c_wstrobe_d ),
    .Q_N(_15084_),
    .Q(\cpu.d_wstrobe_d ));
 sg13g2_dfrbp_1 \cpu.qspi.r_wstrobe_i$_DFF_P_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net3462),
    .D(\cpu.qspi.c_wstrobe_i ),
    .Q_N(_00253_),
    .Q(\cpu.i_wstrobe_d ));
 sg13g2_dfrbp_1 \cpu.r_clk_invert$_DFFE_PN_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net3463),
    .D(_02547_),
    .Q_N(_12956_),
    .Q(\cpu.r_clk_invert ));
 sg13g2_dfrbp_1 \cpu.spi.r_bits[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3464),
    .D(_02548_),
    .Q_N(_12955_),
    .Q(\cpu.spi.r_bits[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_bits[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3465),
    .D(_02549_),
    .Q_N(_12954_),
    .Q(\cpu.spi.r_bits[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_bits[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3466),
    .D(_02550_),
    .Q_N(_12953_),
    .Q(\cpu.spi.r_bits[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3467),
    .D(_02551_),
    .Q_N(_00314_),
    .Q(\cpu.spi.r_clk_count[0][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3468),
    .D(_02552_),
    .Q_N(_00095_),
    .Q(\cpu.spi.r_clk_count[0][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3469),
    .D(_02553_),
    .Q_N(_00105_),
    .Q(\cpu.spi.r_clk_count[0][2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3470),
    .D(_02554_),
    .Q_N(_00115_),
    .Q(\cpu.spi.r_clk_count[0][3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3471),
    .D(_02555_),
    .Q_N(_00126_),
    .Q(\cpu.spi.r_clk_count[0][4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3472),
    .D(_02556_),
    .Q_N(_00133_),
    .Q(\cpu.spi.r_clk_count[0][5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3473),
    .D(_02557_),
    .Q_N(_00145_),
    .Q(\cpu.spi.r_clk_count[0][6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3474),
    .D(_02558_),
    .Q_N(_00157_),
    .Q(\cpu.spi.r_clk_count[0][7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3475),
    .D(_02559_),
    .Q_N(_00313_),
    .Q(\cpu.spi.r_clk_count[1][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3476),
    .D(_02560_),
    .Q_N(_00094_),
    .Q(\cpu.spi.r_clk_count[1][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3477),
    .D(_02561_),
    .Q_N(_00104_),
    .Q(\cpu.spi.r_clk_count[1][2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3478),
    .D(_02562_),
    .Q_N(_00114_),
    .Q(\cpu.spi.r_clk_count[1][3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3479),
    .D(_02563_),
    .Q_N(_00125_),
    .Q(\cpu.spi.r_clk_count[1][4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3480),
    .D(_02564_),
    .Q_N(_00132_),
    .Q(\cpu.spi.r_clk_count[1][5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3481),
    .D(_02565_),
    .Q_N(_00144_),
    .Q(\cpu.spi.r_clk_count[1][6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3482),
    .D(_02566_),
    .Q_N(_00156_),
    .Q(\cpu.spi.r_clk_count[1][7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3483),
    .D(_02567_),
    .Q_N(_12952_),
    .Q(\cpu.spi.r_clk_count[2][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3484),
    .D(_02568_),
    .Q_N(_12951_),
    .Q(\cpu.spi.r_clk_count[2][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3485),
    .D(_02569_),
    .Q_N(_12950_),
    .Q(\cpu.spi.r_clk_count[2][2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3486),
    .D(_02570_),
    .Q_N(_12949_),
    .Q(\cpu.spi.r_clk_count[2][3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3487),
    .D(_02571_),
    .Q_N(_12948_),
    .Q(\cpu.spi.r_clk_count[2][4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3488),
    .D(_02572_),
    .Q_N(_12947_),
    .Q(\cpu.spi.r_clk_count[2][5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3489),
    .D(_02573_),
    .Q_N(_12946_),
    .Q(\cpu.spi.r_clk_count[2][6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3490),
    .D(_02574_),
    .Q_N(_12945_),
    .Q(\cpu.spi.r_clk_count[2][7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3491),
    .D(_02575_),
    .Q_N(_12944_),
    .Q(\cpu.spi.r_count[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3492),
    .D(_02576_),
    .Q_N(_12943_),
    .Q(\cpu.spi.r_count[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3493),
    .D(_02577_),
    .Q_N(_12942_),
    .Q(\cpu.spi.r_count[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3494),
    .D(_02578_),
    .Q_N(_12941_),
    .Q(\cpu.spi.r_count[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3495),
    .D(_02579_),
    .Q_N(_12940_),
    .Q(\cpu.spi.r_count[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3496),
    .D(_02580_),
    .Q_N(_12939_),
    .Q(\cpu.spi.r_count[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3497),
    .D(_02581_),
    .Q_N(_12938_),
    .Q(\cpu.spi.r_count[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3498),
    .D(_02582_),
    .Q_N(_12937_),
    .Q(\cpu.spi.r_count[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_cs[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3499),
    .D(_02583_),
    .Q_N(_12936_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_cs[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3500),
    .D(_02584_),
    .Q_N(_12935_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_cs[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3501),
    .D(_02585_),
    .Q_N(_12934_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[8] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[0]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3502),
    .D(_02586_),
    .Q_N(_12933_),
    .Q(\cpu.spi.r_in[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[1]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3503),
    .D(_02587_),
    .Q_N(_12932_),
    .Q(\cpu.spi.r_in[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[2]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3504),
    .D(_02588_),
    .Q_N(_12931_),
    .Q(\cpu.spi.r_in[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[3]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3505),
    .D(_02589_),
    .Q_N(_12930_),
    .Q(\cpu.spi.r_in[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[4]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3506),
    .D(_02590_),
    .Q_N(_12929_),
    .Q(\cpu.spi.r_in[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[5]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3507),
    .D(_02591_),
    .Q_N(_12928_),
    .Q(\cpu.spi.r_in[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[6]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3508),
    .D(_02592_),
    .Q_N(_12927_),
    .Q(\cpu.spi.r_in[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[7]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3509),
    .D(_02593_),
    .Q_N(_00222_),
    .Q(\cpu.spi.r_in[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_interrupt$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3510),
    .D(_02594_),
    .Q_N(_12926_),
    .Q(\cpu.intr.spi_intr ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[0][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3511),
    .D(_02595_),
    .Q_N(_00224_),
    .Q(\cpu.spi.r_mode[0][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[0][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3512),
    .D(_02596_),
    .Q_N(_12925_),
    .Q(\cpu.spi.r_mode[0][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[1][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3513),
    .D(_02597_),
    .Q_N(_12924_),
    .Q(\cpu.spi.r_mode[1][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[1][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3514),
    .D(_02598_),
    .Q_N(_12923_),
    .Q(\cpu.spi.r_mode[1][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[2][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3515),
    .D(_02599_),
    .Q_N(_12922_),
    .Q(\cpu.spi.r_mode[2][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[2][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3516),
    .D(_02600_),
    .Q_N(_12921_),
    .Q(\cpu.spi.r_mode[2][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3517),
    .D(_02601_),
    .Q_N(_12920_),
    .Q(\cpu.spi.r_out[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3518),
    .D(_02602_),
    .Q_N(_12919_),
    .Q(\cpu.spi.r_out[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3519),
    .D(_02603_),
    .Q_N(_12918_),
    .Q(\cpu.spi.r_out[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3520),
    .D(_02604_),
    .Q_N(_12917_),
    .Q(\cpu.spi.r_out[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[4]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3521),
    .D(_02605_),
    .Q_N(_12916_),
    .Q(\cpu.spi.r_out[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[5]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3522),
    .D(_02606_),
    .Q_N(_12915_),
    .Q(\cpu.spi.r_out[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[6]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3523),
    .D(_02607_),
    .Q_N(_12914_),
    .Q(\cpu.spi.r_out[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[7]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3524),
    .D(_02608_),
    .Q_N(_12913_),
    .Q(\cpu.spi.r_out[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_ready$_SDFFE_PN1P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3525),
    .D(_02609_),
    .Q_N(_12912_),
    .Q(\cpu.spi.r_ready ));
 sg13g2_dfrbp_1 \cpu.spi.r_searching$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3526),
    .D(_02610_),
    .Q_N(_00221_),
    .Q(\cpu.spi.r_searching ));
 sg13g2_dfrbp_1 \cpu.spi.r_sel[0]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3527),
    .D(_02611_),
    .Q_N(_12911_),
    .Q(\cpu.spi.r_sel[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_sel[1]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3528),
    .D(_02612_),
    .Q_N(_12910_),
    .Q(\cpu.spi.r_sel[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_src[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3529),
    .D(_02613_),
    .Q_N(_00282_),
    .Q(\cpu.spi.r_src[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_src[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3530),
    .D(_02614_),
    .Q_N(_00283_),
    .Q(\cpu.spi.r_src[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_src[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3531),
    .D(_02615_),
    .Q_N(_15085_),
    .Q(\cpu.spi.r_src[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[0]$_DFF_P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3532),
    .D(_00029_),
    .Q_N(_15086_),
    .Q(\cpu.spi.r_state[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[1]$_DFF_P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3533),
    .D(_00030_),
    .Q_N(_00225_),
    .Q(\cpu.spi.r_state[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[2]$_DFF_P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3534),
    .D(_00031_),
    .Q_N(_15087_),
    .Q(\cpu.spi.r_state[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[3]$_DFF_P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3535),
    .D(_00032_),
    .Q_N(_15088_),
    .Q(\cpu.spi.r_state[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[4]$_DFF_P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3536),
    .D(_00033_),
    .Q_N(_00278_),
    .Q(\cpu.spi.r_state[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[5]$_DFF_P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3537),
    .D(_00034_),
    .Q_N(_15089_),
    .Q(\cpu.spi.r_state[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[6]$_DFF_P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3538),
    .D(_00035_),
    .Q_N(_00226_),
    .Q(\cpu.spi.r_state[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[0]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3539),
    .D(_02616_),
    .Q_N(_12909_),
    .Q(\cpu.spi.r_timeout[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[1]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3540),
    .D(_02617_),
    .Q_N(_12908_),
    .Q(\cpu.spi.r_timeout[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[2]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3541),
    .D(_02618_),
    .Q_N(_12907_),
    .Q(\cpu.spi.r_timeout[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[3]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3542),
    .D(_02619_),
    .Q_N(_12906_),
    .Q(\cpu.spi.r_timeout[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[4]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3543),
    .D(_02620_),
    .Q_N(_12905_),
    .Q(\cpu.spi.r_timeout[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[5]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3544),
    .D(_02621_),
    .Q_N(_12904_),
    .Q(\cpu.spi.r_timeout[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[6]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3545),
    .D(_02622_),
    .Q_N(_12903_),
    .Q(\cpu.spi.r_timeout[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[7]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3546),
    .D(_02623_),
    .Q_N(_12902_),
    .Q(\cpu.spi.r_timeout[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[0]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3547),
    .D(_02624_),
    .Q_N(_00284_),
    .Q(\cpu.spi.r_timeout_count[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[1]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3548),
    .D(_02625_),
    .Q_N(_12901_),
    .Q(\cpu.spi.r_timeout_count[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[2]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3549),
    .D(_02626_),
    .Q_N(_12900_),
    .Q(\cpu.spi.r_timeout_count[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[3]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3550),
    .D(_02627_),
    .Q_N(_12899_),
    .Q(\cpu.spi.r_timeout_count[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[4]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3551),
    .D(_02628_),
    .Q_N(_12898_),
    .Q(\cpu.spi.r_timeout_count[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[5]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net3552),
    .D(_02629_),
    .Q_N(_12897_),
    .Q(\cpu.spi.r_timeout_count[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[6]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3553),
    .D(_02630_),
    .Q_N(_12896_),
    .Q(\cpu.spi.r_timeout_count[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[7]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3554),
    .D(_02631_),
    .Q_N(_15090_),
    .Q(\cpu.spi.r_timeout_count[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[0]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3555),
    .D(_00079_),
    .Q_N(_00279_),
    .Q(\cpu.uart.r_div[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[10]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3556),
    .D(_00080_),
    .Q_N(_15091_),
    .Q(\cpu.uart.r_div[10] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[11]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3557),
    .D(_00081_),
    .Q_N(_15092_),
    .Q(\cpu.uart.r_div[11] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[1]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3558),
    .D(_00082_),
    .Q_N(_15093_),
    .Q(\cpu.uart.r_div[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[2]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3559),
    .D(_00083_),
    .Q_N(_15094_),
    .Q(\cpu.uart.r_div[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[3]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3560),
    .D(_00084_),
    .Q_N(_15095_),
    .Q(\cpu.uart.r_div[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[4]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3561),
    .D(_00085_),
    .Q_N(_15096_),
    .Q(\cpu.uart.r_div[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[5]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3562),
    .D(_00086_),
    .Q_N(_15097_),
    .Q(\cpu.uart.r_div[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[6]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3563),
    .D(_00087_),
    .Q_N(_15098_),
    .Q(\cpu.uart.r_div[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[7]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3564),
    .D(_00088_),
    .Q_N(_15099_),
    .Q(\cpu.uart.r_div[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[8]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3565),
    .D(_00089_),
    .Q_N(_15100_),
    .Q(\cpu.uart.r_div[8] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[9]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3566),
    .D(_00090_),
    .Q_N(_12895_),
    .Q(\cpu.uart.r_div[9] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3567),
    .D(_02632_),
    .Q_N(_12894_),
    .Q(\cpu.uart.r_div_value[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3568),
    .D(_02633_),
    .Q_N(_12893_),
    .Q(\cpu.uart.r_div_value[10] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3569),
    .D(_02634_),
    .Q_N(_12892_),
    .Q(\cpu.uart.r_div_value[11] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3570),
    .D(_02635_),
    .Q_N(_12891_),
    .Q(\cpu.uart.r_div_value[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3571),
    .D(_02636_),
    .Q_N(_12890_),
    .Q(\cpu.uart.r_div_value[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3572),
    .D(_02637_),
    .Q_N(_12889_),
    .Q(\cpu.uart.r_div_value[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3573),
    .D(_02638_),
    .Q_N(_12888_),
    .Q(\cpu.uart.r_div_value[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3574),
    .D(_02639_),
    .Q_N(_12887_),
    .Q(\cpu.uart.r_div_value[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3575),
    .D(_02640_),
    .Q_N(_12886_),
    .Q(\cpu.uart.r_div_value[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3576),
    .D(_02641_),
    .Q_N(_12885_),
    .Q(\cpu.uart.r_div_value[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3577),
    .D(_02642_),
    .Q_N(_12884_),
    .Q(\cpu.uart.r_div_value[8] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3578),
    .D(_02643_),
    .Q_N(_12883_),
    .Q(\cpu.uart.r_div_value[9] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[0]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3579),
    .D(_02644_),
    .Q_N(_12882_),
    .Q(\cpu.uart.r_ib[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[1]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3580),
    .D(_02645_),
    .Q_N(_12881_),
    .Q(\cpu.uart.r_ib[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[2]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3581),
    .D(_02646_),
    .Q_N(_12880_),
    .Q(\cpu.uart.r_ib[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[3]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3582),
    .D(_02647_),
    .Q_N(_12879_),
    .Q(\cpu.uart.r_ib[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[4]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3583),
    .D(_02648_),
    .Q_N(_12878_),
    .Q(\cpu.uart.r_ib[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[5]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3584),
    .D(_02649_),
    .Q_N(_12877_),
    .Q(\cpu.uart.r_ib[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[6]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3585),
    .D(_02650_),
    .Q_N(_12876_),
    .Q(\cpu.uart.r_ib[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[0]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3586),
    .D(_02651_),
    .Q_N(_12875_),
    .Q(\cpu.uart.r_in[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[1]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3587),
    .D(_02652_),
    .Q_N(_12874_),
    .Q(\cpu.uart.r_in[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[2]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3588),
    .D(_02653_),
    .Q_N(_12873_),
    .Q(\cpu.uart.r_in[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[3]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3589),
    .D(_02654_),
    .Q_N(_12872_),
    .Q(\cpu.uart.r_in[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[4]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3590),
    .D(_02655_),
    .Q_N(_12871_),
    .Q(\cpu.uart.r_in[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[5]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3591),
    .D(_02656_),
    .Q_N(_12870_),
    .Q(\cpu.uart.r_in[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[6]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3592),
    .D(_02657_),
    .Q_N(_12869_),
    .Q(\cpu.uart.r_in[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[7]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3593),
    .D(_02658_),
    .Q_N(_12868_),
    .Q(\cpu.uart.r_in[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3594),
    .D(_02659_),
    .Q_N(_12867_),
    .Q(\cpu.uart.r_out[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3595),
    .D(_02660_),
    .Q_N(_12866_),
    .Q(\cpu.uart.r_out[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3596),
    .D(_02661_),
    .Q_N(_12865_),
    .Q(\cpu.uart.r_out[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3597),
    .D(_02662_),
    .Q_N(_12864_),
    .Q(\cpu.uart.r_out[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[4]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3598),
    .D(_02663_),
    .Q_N(_12863_),
    .Q(\cpu.uart.r_out[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[5]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3599),
    .D(_02664_),
    .Q_N(_12862_),
    .Q(\cpu.uart.r_out[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[6]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3600),
    .D(_02665_),
    .Q_N(_12861_),
    .Q(\cpu.uart.r_out[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[7]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3601),
    .D(_02666_),
    .Q_N(_15101_),
    .Q(\cpu.uart.r_out[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_r$_DFF_P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3602),
    .D(\cpu.gpio.uart_rx ),
    .Q_N(_12860_),
    .Q(\cpu.uart.r_r ));
 sg13g2_dfrbp_1 \cpu.uart.r_r_int$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3603),
    .D(_02667_),
    .Q_N(_12859_),
    .Q(\cpu.uart.r_r_int ));
 sg13g2_dfrbp_1 \cpu.uart.r_r_invert$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3604),
    .D(_02668_),
    .Q_N(_12858_),
    .Q(\cpu.uart.r_r_invert ));
 sg13g2_dfrbp_1 \cpu.uart.r_rcnt[0]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3605),
    .D(_02669_),
    .Q_N(_12857_),
    .Q(\cpu.uart.r_rcnt[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rcnt[1]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3606),
    .D(_02670_),
    .Q_N(_12856_),
    .Q(\cpu.uart.r_rcnt[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3607),
    .D(_02671_),
    .Q_N(_12855_),
    .Q(\cpu.uart.r_rstate[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3608),
    .D(_02672_),
    .Q_N(_12854_),
    .Q(\cpu.uart.r_rstate[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3609),
    .D(_02673_),
    .Q_N(_12853_),
    .Q(\cpu.uart.r_rstate[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3610),
    .D(_02674_),
    .Q_N(_12852_),
    .Q(\cpu.uart.r_rstate[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_x$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3611),
    .D(_02675_),
    .Q_N(_12851_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_x_int$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3612),
    .D(_02676_),
    .Q_N(_12850_),
    .Q(\cpu.uart.r_x_int ));
 sg13g2_dfrbp_1 \cpu.uart.r_x_invert$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3613),
    .D(_02677_),
    .Q_N(_00280_),
    .Q(\cpu.uart.r_x_invert ));
 sg13g2_dfrbp_1 \cpu.uart.r_xcnt[0]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3614),
    .D(_02678_),
    .Q_N(_12849_),
    .Q(\cpu.uart.r_xcnt[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xcnt[1]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3615),
    .D(_02679_),
    .Q_N(_12848_),
    .Q(\cpu.uart.r_xcnt[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3616),
    .D(_02680_),
    .Q_N(_12847_),
    .Q(\cpu.uart.r_xstate[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3617),
    .D(_02681_),
    .Q_N(_12846_),
    .Q(\cpu.uart.r_xstate[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3618),
    .D(_02682_),
    .Q_N(_12845_),
    .Q(\cpu.uart.r_xstate[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3619),
    .D(_02683_),
    .Q_N(_15102_),
    .Q(\cpu.uart.r_xstate[3] ));
 sg13g2_dfrbp_1 \r_reset$_DFF_P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3620),
    .D(_00000_),
    .Q_N(_12844_),
    .Q(r_reset));
 sg13g2_buf_1 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_1 input2 (.A(rst_n),
    .X(net2));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uio_oe[0]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uio_oe[1]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uio_oe[2]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_oe[3]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_oe[4]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_oe[5]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_oe[6]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_oe[7]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[0]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[1]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[2]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[3]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_out[4]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_out[5]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_out[6]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_out[7]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[0]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[1]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[2]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[3]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[4]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[5]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[6]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout27 (.A(_03801_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_06766_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_03729_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_07161_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_07995_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_04147_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_07084_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_02889_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_02844_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_02789_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_02754_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_02737_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_02725_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_12838_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_12802_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_12785_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_12774_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_12723_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_12686_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_12669_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_12661_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_12616_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_12573_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_12513_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_12479_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_12462_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_12452_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_12399_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_12358_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_12337_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_12324_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_12266_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_12207_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_12156_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_12124_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_11801_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_04828_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_04223_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_04031_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_02860_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_02835_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_12589_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_12563_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_11663_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_11658_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_10250_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_10249_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_10145_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_10134_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_10133_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_07270_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_07253_),
    .X(net78));
 sg13g2_buf_4 fanout79 (.X(net79),
    .A(_06751_));
 sg13g2_buf_4 fanout80 (.X(net80),
    .A(_06748_));
 sg13g2_buf_4 fanout81 (.X(net81),
    .A(_05777_));
 sg13g2_buf_2 fanout82 (.A(_05239_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_04829_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_04827_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_04824_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_04135_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_03028_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_11662_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_10021_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_09434_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_09264_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_09171_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_08208_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_07257_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_07256_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_06404_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_05143_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_05021_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_04097_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_11740_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_11689_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_11661_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_10276_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_10259_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_10239_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_09998_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_09433_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_09170_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_07255_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_06804_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_04096_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_03123_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_03114_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_03032_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_03012_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_11954_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_10238_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_09994_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_08974_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_08973_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_06879_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_06845_),
    .X(net122));
 sg13g2_buf_4 fanout123 (.X(net123),
    .A(_06754_));
 sg13g2_buf_2 fanout124 (.A(_06745_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_04256_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_04192_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_04095_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_03592_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_03492_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_03485_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_03479_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_11634_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_10181_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_04194_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_04180_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_04178_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_04167_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_04067_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_04062_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_04036_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_03566_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_03491_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_03487_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_03133_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_11914_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_11650_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_11594_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_10180_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_10030_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_10005_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_09201_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_09083_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_07639_),
    .X(net153));
 sg13g2_buf_4 fanout154 (.X(net154),
    .A(_07130_));
 sg13g2_buf_2 fanout155 (.A(_04274_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_04259_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_04149_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_04107_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_04093_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_04076_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_04032_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_03789_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_03558_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_03473_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_03262_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_03120_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_03018_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_03016_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_11926_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_11892_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_11886_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_11829_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_11644_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_11638_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_10567_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_10532_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_10015_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_10012_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_09198_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_09194_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_07699_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_07665_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_07646_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_07645_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_07521_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_07482_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_07481_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_07470_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_05173_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_04106_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_04070_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_03569_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_03537_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_03529_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_03510_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_03472_),
    .X(net196));
 sg13g2_buf_4 fanout197 (.X(net197),
    .A(_02981_));
 sg13g2_buf_4 fanout198 (.X(net198),
    .A(_02980_));
 sg13g2_buf_2 fanout199 (.A(_11925_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_11840_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_11806_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_11584_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_10753_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_10653_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_10061_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_10028_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_10014_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_10013_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_09239_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_09193_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_09151_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_08998_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_07464_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_05790_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_04822_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_04176_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_04043_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_03595_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_03507_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_03503_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_03474_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_03095_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_03023_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_03021_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_03014_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_03002_),
    .X(net226));
 sg13g2_buf_4 fanout227 (.X(net227),
    .A(_03000_));
 sg13g2_buf_4 fanout228 (.X(net228),
    .A(_02999_));
 sg13g2_buf_2 fanout229 (.A(_11735_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_11731_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_11700_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_11653_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_11290_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_11011_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_10908_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_10877_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_10060_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_09102_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_09040_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_09018_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_06373_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_06323_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_06273_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_06262_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_06226_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_06179_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_06169_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_06158_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_06123_),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(_06073_),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(_06061_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(_06028_),
    .X(net252));
 sg13g2_buf_4 fanout253 (.X(net253),
    .A(_06019_));
 sg13g2_buf_4 fanout254 (.X(net254),
    .A(_05986_));
 sg13g2_buf_4 fanout255 (.X(net255),
    .A(_05982_));
 sg13g2_buf_4 fanout256 (.X(net256),
    .A(_05976_));
 sg13g2_buf_4 fanout257 (.X(net257),
    .A(_05954_));
 sg13g2_buf_4 fanout258 (.X(net258),
    .A(_05942_));
 sg13g2_buf_4 fanout259 (.X(net259),
    .A(_05938_));
 sg13g2_buf_4 fanout260 (.X(net260),
    .A(_05925_));
 sg13g2_buf_4 fanout261 (.X(net261),
    .A(_05909_));
 sg13g2_buf_4 fanout262 (.X(net262),
    .A(_05893_));
 sg13g2_buf_4 fanout263 (.X(net263),
    .A(_05889_));
 sg13g2_buf_2 fanout264 (.A(_04963_),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(_03849_),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(_03520_),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(_03214_),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(_03117_),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(_03091_),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(_03015_),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(_12561_),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(_11714_),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(_11587_),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(_11382_),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(_11267_),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(_11038_),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(_10948_),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_10367_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(_10025_),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_09195_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_09173_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_08527_),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(_06640_),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(_06633_),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(_06592_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(_06590_),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(_06589_),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(_06517_),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(_06516_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(_06372_),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(_06363_),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(_06353_),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(_06343_),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(_06333_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(_06322_),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(_06313_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_06303_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(_06293_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(_06283_),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(_06272_),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(_06261_),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(_06251_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(_06237_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_06225_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(_06210_),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(_06199_),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_06189_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(_06178_),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(_06168_),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_06157_),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(_06147_),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(_06137_),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(_06122_),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(_06112_),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(_06094_),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(_06083_),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(_06072_),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(_06060_),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(_06050_),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(_06040_),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(_06027_),
    .X(net321));
 sg13g2_buf_4 fanout322 (.X(net322),
    .A(_06016_));
 sg13g2_buf_4 fanout323 (.X(net323),
    .A(_06013_));
 sg13g2_buf_4 fanout324 (.X(net324),
    .A(_06008_));
 sg13g2_buf_4 fanout325 (.X(net325),
    .A(_06002_));
 sg13g2_buf_4 fanout326 (.X(net326),
    .A(_05997_));
 sg13g2_buf_4 fanout327 (.X(net327),
    .A(_05993_));
 sg13g2_buf_4 fanout328 (.X(net328),
    .A(_05990_));
 sg13g2_buf_4 fanout329 (.X(net329),
    .A(_05972_));
 sg13g2_buf_4 fanout330 (.X(net330),
    .A(_05964_));
 sg13g2_buf_4 fanout331 (.X(net331),
    .A(_05959_));
 sg13g2_buf_4 fanout332 (.X(net332),
    .A(_05951_));
 sg13g2_buf_4 fanout333 (.X(net333),
    .A(_05945_));
 sg13g2_buf_4 fanout334 (.X(net334),
    .A(_05933_));
 sg13g2_buf_4 fanout335 (.X(net335),
    .A(_05921_));
 sg13g2_buf_4 fanout336 (.X(net336),
    .A(_05913_));
 sg13g2_buf_4 fanout337 (.X(net337),
    .A(_05905_));
 sg13g2_buf_4 fanout338 (.X(net338),
    .A(_05899_));
 sg13g2_buf_4 fanout339 (.X(net339),
    .A(_05882_));
 sg13g2_buf_4 fanout340 (.X(net340),
    .A(_05874_));
 sg13g2_buf_4 fanout341 (.X(net341),
    .A(_05865_));
 sg13g2_buf_4 fanout342 (.X(net342),
    .A(_05854_));
 sg13g2_buf_2 fanout343 (.A(_05002_),
    .X(net343));
 sg13g2_buf_2 fanout344 (.A(_03064_),
    .X(net344));
 sg13g2_buf_2 fanout345 (.A(_02833_),
    .X(net345));
 sg13g2_buf_2 fanout346 (.A(_11660_),
    .X(net346));
 sg13g2_buf_4 fanout347 (.X(net347),
    .A(_11192_));
 sg13g2_buf_2 fanout348 (.A(_10058_),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(_08558_),
    .X(net349));
 sg13g2_buf_2 fanout350 (.A(_06704_),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(_06702_),
    .X(net351));
 sg13g2_buf_2 fanout352 (.A(_06701_),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(_06681_),
    .X(net353));
 sg13g2_buf_2 fanout354 (.A(_06679_),
    .X(net354));
 sg13g2_buf_2 fanout355 (.A(_06678_),
    .X(net355));
 sg13g2_buf_2 fanout356 (.A(_06615_),
    .X(net356));
 sg13g2_buf_2 fanout357 (.A(_06613_),
    .X(net357));
 sg13g2_buf_2 fanout358 (.A(_06612_),
    .X(net358));
 sg13g2_buf_2 fanout359 (.A(_06588_),
    .X(net359));
 sg13g2_buf_2 fanout360 (.A(_06362_),
    .X(net360));
 sg13g2_buf_2 fanout361 (.A(_06352_),
    .X(net361));
 sg13g2_buf_2 fanout362 (.A(_06342_),
    .X(net362));
 sg13g2_buf_2 fanout363 (.A(_06332_),
    .X(net363));
 sg13g2_buf_2 fanout364 (.A(_06312_),
    .X(net364));
 sg13g2_buf_2 fanout365 (.A(_06302_),
    .X(net365));
 sg13g2_buf_2 fanout366 (.A(_06292_),
    .X(net366));
 sg13g2_buf_2 fanout367 (.A(_06282_),
    .X(net367));
 sg13g2_buf_2 fanout368 (.A(_06250_),
    .X(net368));
 sg13g2_buf_2 fanout369 (.A(_06236_),
    .X(net369));
 sg13g2_buf_2 fanout370 (.A(_06209_),
    .X(net370));
 sg13g2_buf_2 fanout371 (.A(_06198_),
    .X(net371));
 sg13g2_buf_2 fanout372 (.A(_06188_),
    .X(net372));
 sg13g2_buf_2 fanout373 (.A(_06146_),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(_06136_),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(_06111_),
    .X(net375));
 sg13g2_buf_2 fanout376 (.A(_06093_),
    .X(net376));
 sg13g2_buf_2 fanout377 (.A(_06082_),
    .X(net377));
 sg13g2_buf_2 fanout378 (.A(_06049_),
    .X(net378));
 sg13g2_buf_2 fanout379 (.A(_06039_),
    .X(net379));
 sg13g2_buf_2 fanout380 (.A(_04996_),
    .X(net380));
 sg13g2_buf_2 fanout381 (.A(_04952_),
    .X(net381));
 sg13g2_buf_2 fanout382 (.A(_04939_),
    .X(net382));
 sg13g2_buf_2 fanout383 (.A(_04912_),
    .X(net383));
 sg13g2_buf_2 fanout384 (.A(_03434_),
    .X(net384));
 sg13g2_buf_4 fanout385 (.X(net385),
    .A(_02985_));
 sg13g2_buf_2 fanout386 (.A(_02982_),
    .X(net386));
 sg13g2_buf_4 fanout387 (.X(net387),
    .A(_02946_));
 sg13g2_buf_2 fanout388 (.A(_02945_),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(_12332_),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(_12275_),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(_12261_),
    .X(net391));
 sg13g2_buf_2 fanout392 (.A(_12201_),
    .X(net392));
 sg13g2_buf_2 fanout393 (.A(_12195_),
    .X(net393));
 sg13g2_buf_2 fanout394 (.A(_12187_),
    .X(net394));
 sg13g2_buf_2 fanout395 (.A(_12175_),
    .X(net395));
 sg13g2_buf_2 fanout396 (.A(_12167_),
    .X(net396));
 sg13g2_buf_2 fanout397 (.A(_12150_),
    .X(net397));
 sg13g2_buf_2 fanout398 (.A(_11540_),
    .X(net398));
 sg13g2_buf_2 fanout399 (.A(_10256_),
    .X(net399));
 sg13g2_buf_2 fanout400 (.A(_09913_),
    .X(net400));
 sg13g2_buf_2 fanout401 (.A(_09890_),
    .X(net401));
 sg13g2_buf_2 fanout402 (.A(_09797_),
    .X(net402));
 sg13g2_buf_2 fanout403 (.A(_09768_),
    .X(net403));
 sg13g2_buf_2 fanout404 (.A(_09743_),
    .X(net404));
 sg13g2_buf_2 fanout405 (.A(_09722_),
    .X(net405));
 sg13g2_buf_2 fanout406 (.A(_09696_),
    .X(net406));
 sg13g2_buf_2 fanout407 (.A(_09649_),
    .X(net407));
 sg13g2_buf_2 fanout408 (.A(_09588_),
    .X(net408));
 sg13g2_buf_2 fanout409 (.A(_09565_),
    .X(net409));
 sg13g2_buf_2 fanout410 (.A(_09158_),
    .X(net410));
 sg13g2_buf_2 fanout411 (.A(_08960_),
    .X(net411));
 sg13g2_buf_2 fanout412 (.A(_08939_),
    .X(net412));
 sg13g2_buf_2 fanout413 (.A(_08918_),
    .X(net413));
 sg13g2_buf_2 fanout414 (.A(_08728_),
    .X(net414));
 sg13g2_buf_2 fanout415 (.A(_08634_),
    .X(net415));
 sg13g2_buf_2 fanout416 (.A(_08573_),
    .X(net416));
 sg13g2_buf_2 fanout417 (.A(_06700_),
    .X(net417));
 sg13g2_buf_2 fanout418 (.A(_06677_),
    .X(net418));
 sg13g2_buf_2 fanout419 (.A(_06611_),
    .X(net419));
 sg13g2_buf_2 fanout420 (.A(_06572_),
    .X(net420));
 sg13g2_buf_2 fanout421 (.A(_06565_),
    .X(net421));
 sg13g2_buf_2 fanout422 (.A(_06453_),
    .X(net422));
 sg13g2_buf_2 fanout423 (.A(_06452_),
    .X(net423));
 sg13g2_buf_2 fanout424 (.A(_06383_),
    .X(net424));
 sg13g2_buf_2 fanout425 (.A(_06382_),
    .X(net425));
 sg13g2_buf_2 fanout426 (.A(_06381_),
    .X(net426));
 sg13g2_buf_2 fanout427 (.A(_05005_),
    .X(net427));
 sg13g2_buf_2 fanout428 (.A(_04988_),
    .X(net428));
 sg13g2_buf_2 fanout429 (.A(_04934_),
    .X(net429));
 sg13g2_buf_2 fanout430 (.A(_04905_),
    .X(net430));
 sg13g2_buf_2 fanout431 (.A(_04844_),
    .X(net431));
 sg13g2_buf_2 fanout432 (.A(_04835_),
    .X(net432));
 sg13g2_buf_2 fanout433 (.A(_04831_),
    .X(net433));
 sg13g2_buf_2 fanout434 (.A(_03433_),
    .X(net434));
 sg13g2_buf_2 fanout435 (.A(_02734_),
    .X(net435));
 sg13g2_buf_2 fanout436 (.A(_12726_),
    .X(net436));
 sg13g2_buf_4 fanout437 (.X(net437),
    .A(_12558_));
 sg13g2_buf_2 fanout438 (.A(_12459_),
    .X(net438));
 sg13g2_buf_2 fanout439 (.A(_12331_),
    .X(net439));
 sg13g2_buf_2 fanout440 (.A(_12269_),
    .X(net440));
 sg13g2_buf_2 fanout441 (.A(_11707_),
    .X(net441));
 sg13g2_buf_2 fanout442 (.A(_11667_),
    .X(net442));
 sg13g2_buf_2 fanout443 (.A(_10255_),
    .X(net443));
 sg13g2_buf_2 fanout444 (.A(_10236_),
    .X(net444));
 sg13g2_buf_2 fanout445 (.A(_10121_),
    .X(net445));
 sg13g2_buf_2 fanout446 (.A(_09394_),
    .X(net446));
 sg13g2_buf_2 fanout447 (.A(_09276_),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(_08896_),
    .X(net448));
 sg13g2_buf_2 fanout449 (.A(_08854_),
    .X(net449));
 sg13g2_buf_2 fanout450 (.A(_08698_),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(_08660_),
    .X(net451));
 sg13g2_buf_2 fanout452 (.A(_08575_),
    .X(net452));
 sg13g2_buf_2 fanout453 (.A(_08572_),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(_07575_),
    .X(net454));
 sg13g2_buf_2 fanout455 (.A(_07478_),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(_06727_),
    .X(net456));
 sg13g2_buf_2 fanout457 (.A(_06725_),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(_06724_),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(_06658_),
    .X(net459));
 sg13g2_buf_2 fanout460 (.A(_06656_),
    .X(net460));
 sg13g2_buf_2 fanout461 (.A(_06655_),
    .X(net461));
 sg13g2_buf_2 fanout462 (.A(_06091_),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(_06037_),
    .X(net463));
 sg13g2_buf_2 fanout464 (.A(_05935_),
    .X(net464));
 sg13g2_buf_2 fanout465 (.A(_05876_),
    .X(net465));
 sg13g2_buf_2 fanout466 (.A(_05856_),
    .X(net466));
 sg13g2_buf_2 fanout467 (.A(_05132_),
    .X(net467));
 sg13g2_buf_2 fanout468 (.A(_04837_),
    .X(net468));
 sg13g2_buf_2 fanout469 (.A(_04830_),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(_04756_),
    .X(net470));
 sg13g2_buf_2 fanout471 (.A(_04752_),
    .X(net471));
 sg13g2_buf_2 fanout472 (.A(_03733_),
    .X(net472));
 sg13g2_buf_2 fanout473 (.A(_03463_),
    .X(net473));
 sg13g2_buf_2 fanout474 (.A(_03436_),
    .X(net474));
 sg13g2_buf_4 fanout475 (.X(net475),
    .A(_03432_));
 sg13g2_buf_2 fanout476 (.A(_03431_),
    .X(net476));
 sg13g2_buf_4 fanout477 (.X(net477),
    .A(_02993_));
 sg13g2_buf_4 fanout478 (.X(net478),
    .A(_02992_));
 sg13g2_buf_4 fanout479 (.X(net479),
    .A(_02990_));
 sg13g2_buf_4 fanout480 (.X(net480),
    .A(_02989_));
 sg13g2_buf_4 fanout481 (.X(net481),
    .A(_02979_));
 sg13g2_buf_4 fanout482 (.X(net482),
    .A(_02978_));
 sg13g2_buf_4 fanout483 (.X(net483),
    .A(_02970_));
 sg13g2_buf_4 fanout484 (.X(net484),
    .A(_02968_));
 sg13g2_buf_2 fanout485 (.A(_02733_),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(_12782_),
    .X(net486));
 sg13g2_buf_2 fanout487 (.A(_12570_),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(_12458_),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(_12330_),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(_11706_),
    .X(net490));
 sg13g2_buf_2 fanout491 (.A(_10463_),
    .X(net491));
 sg13g2_buf_2 fanout492 (.A(_10362_),
    .X(net492));
 sg13g2_buf_2 fanout493 (.A(_10235_),
    .X(net493));
 sg13g2_buf_2 fanout494 (.A(_10120_),
    .X(net494));
 sg13g2_buf_2 fanout495 (.A(_09465_),
    .X(net495));
 sg13g2_buf_2 fanout496 (.A(_09345_),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(_09275_),
    .X(net497));
 sg13g2_buf_4 fanout498 (.X(net498),
    .A(_09000_));
 sg13g2_buf_2 fanout499 (.A(_08981_),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(_08874_),
    .X(net500));
 sg13g2_buf_2 fanout501 (.A(_08661_),
    .X(net501));
 sg13g2_buf_2 fanout502 (.A(_08591_),
    .X(net502));
 sg13g2_buf_2 fanout503 (.A(_08574_),
    .X(net503));
 sg13g2_buf_2 fanout504 (.A(_08571_),
    .X(net504));
 sg13g2_buf_2 fanout505 (.A(_08523_),
    .X(net505));
 sg13g2_buf_2 fanout506 (.A(_07540_),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(_07537_),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(_06723_),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(_06654_),
    .X(net509));
 sg13g2_buf_2 fanout510 (.A(_05977_),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(_05926_),
    .X(net511));
 sg13g2_buf_2 fanout512 (.A(_05906_),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(_05866_),
    .X(net513));
 sg13g2_buf_2 fanout514 (.A(_05111_),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(_04949_),
    .X(net515));
 sg13g2_buf_2 fanout516 (.A(_04754_),
    .X(net516));
 sg13g2_buf_2 fanout517 (.A(_04751_),
    .X(net517));
 sg13g2_buf_2 fanout518 (.A(_04745_),
    .X(net518));
 sg13g2_buf_2 fanout519 (.A(_03732_),
    .X(net519));
 sg13g2_buf_4 fanout520 (.X(net520),
    .A(_03470_));
 sg13g2_buf_2 fanout521 (.A(_03465_),
    .X(net521));
 sg13g2_buf_4 fanout522 (.X(net522),
    .A(_03462_));
 sg13g2_buf_4 fanout523 (.X(net523),
    .A(_03439_));
 sg13g2_buf_4 fanout524 (.X(net524),
    .A(_03435_));
 sg13g2_buf_2 fanout525 (.A(_03429_),
    .X(net525));
 sg13g2_buf_4 fanout526 (.X(net526),
    .A(_03426_));
 sg13g2_buf_2 fanout527 (.A(_02967_),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(_02732_),
    .X(net528));
 sg13g2_buf_2 fanout529 (.A(_12781_),
    .X(net529));
 sg13g2_buf_2 fanout530 (.A(_12569_),
    .X(net530));
 sg13g2_buf_2 fanout531 (.A(_12557_),
    .X(net531));
 sg13g2_buf_2 fanout532 (.A(_11705_),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(_11698_),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(_11150_),
    .X(net534));
 sg13g2_buf_2 fanout535 (.A(_11120_),
    .X(net535));
 sg13g2_buf_2 fanout536 (.A(_10522_),
    .X(net536));
 sg13g2_buf_2 fanout537 (.A(_10470_),
    .X(net537));
 sg13g2_buf_2 fanout538 (.A(_10445_),
    .X(net538));
 sg13g2_buf_2 fanout539 (.A(_10420_),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(_10399_),
    .X(net540));
 sg13g2_buf_2 fanout541 (.A(_10389_),
    .X(net541));
 sg13g2_buf_4 fanout542 (.X(net542),
    .A(_10246_));
 sg13g2_buf_2 fanout543 (.A(_10240_),
    .X(net543));
 sg13g2_buf_2 fanout544 (.A(_10234_),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(_10119_),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(_09769_),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(_09697_),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(_09623_),
    .X(net548));
 sg13g2_buf_2 fanout549 (.A(_09518_),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(_09474_),
    .X(net550));
 sg13g2_buf_4 fanout551 (.X(net551),
    .A(_09344_));
 sg13g2_buf_4 fanout552 (.X(net552),
    .A(_08992_));
 sg13g2_buf_2 fanout553 (.A(_08747_),
    .X(net553));
 sg13g2_buf_2 fanout554 (.A(_08708_),
    .X(net554));
 sg13g2_buf_2 fanout555 (.A(_08703_),
    .X(net555));
 sg13g2_buf_2 fanout556 (.A(_08667_),
    .X(net556));
 sg13g2_buf_2 fanout557 (.A(_08597_),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(_08590_),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(_08580_),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(_08570_),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(_08227_),
    .X(net561));
 sg13g2_buf_2 fanout562 (.A(_08060_),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(_07957_),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(_07932_),
    .X(net564));
 sg13g2_buf_2 fanout565 (.A(_07841_),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(_07787_),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(_07763_),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(_07738_),
    .X(net568));
 sg13g2_buf_2 fanout569 (.A(_07696_),
    .X(net569));
 sg13g2_buf_2 fanout570 (.A(_07673_),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(_07624_),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(_07589_),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(_07545_),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(_07452_),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(_07436_),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(_07376_),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(_06814_),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(_06241_),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(_06234_),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(_06127_),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(_06120_),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(_05978_),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(_05955_),
    .X(net583));
 sg13g2_buf_2 fanout584 (.A(_05927_),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(_05867_),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(_04868_),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(_04744_),
    .X(net587));
 sg13g2_buf_4 fanout588 (.X(net588),
    .A(_04739_));
 sg13g2_buf_2 fanout589 (.A(_04225_),
    .X(net589));
 sg13g2_buf_2 fanout590 (.A(_03715_),
    .X(net590));
 sg13g2_buf_2 fanout591 (.A(_03714_),
    .X(net591));
 sg13g2_buf_2 fanout592 (.A(_03708_),
    .X(net592));
 sg13g2_buf_2 fanout593 (.A(_03703_),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(_03691_),
    .X(net594));
 sg13g2_buf_2 fanout595 (.A(_03690_),
    .X(net595));
 sg13g2_buf_4 fanout596 (.X(net596),
    .A(_03461_));
 sg13g2_buf_4 fanout597 (.X(net597),
    .A(_03459_));
 sg13g2_buf_4 fanout598 (.X(net598),
    .A(_03454_));
 sg13g2_buf_4 fanout599 (.X(net599),
    .A(_03451_));
 sg13g2_buf_4 fanout600 (.X(net600),
    .A(_03444_));
 sg13g2_buf_2 fanout601 (.A(_03427_),
    .X(net601));
 sg13g2_buf_2 fanout602 (.A(_02966_),
    .X(net602));
 sg13g2_buf_2 fanout603 (.A(_02731_),
    .X(net603));
 sg13g2_buf_2 fanout604 (.A(_12780_),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(_12658_),
    .X(net605));
 sg13g2_buf_2 fanout606 (.A(_12449_),
    .X(net606));
 sg13g2_buf_2 fanout607 (.A(_12128_),
    .X(net607));
 sg13g2_buf_2 fanout608 (.A(_12096_),
    .X(net608));
 sg13g2_buf_2 fanout609 (.A(_12068_),
    .X(net609));
 sg13g2_buf_2 fanout610 (.A(_12067_),
    .X(net610));
 sg13g2_buf_2 fanout611 (.A(_11222_),
    .X(net611));
 sg13g2_buf_2 fanout612 (.A(_11149_),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(_10482_),
    .X(net613));
 sg13g2_buf_4 fanout614 (.X(net614),
    .A(_10479_));
 sg13g2_buf_2 fanout615 (.A(_10469_),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(_10444_),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(_10419_),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(_10245_),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(_10174_),
    .X(net619));
 sg13g2_buf_2 fanout620 (.A(_10172_),
    .X(net620));
 sg13g2_buf_2 fanout621 (.A(_10118_),
    .X(net621));
 sg13g2_buf_2 fanout622 (.A(_09541_),
    .X(net622));
 sg13g2_buf_2 fanout623 (.A(_09535_),
    .X(net623));
 sg13g2_buf_2 fanout624 (.A(_09526_),
    .X(net624));
 sg13g2_buf_2 fanout625 (.A(_09517_),
    .X(net625));
 sg13g2_buf_2 fanout626 (.A(_09508_),
    .X(net626));
 sg13g2_buf_2 fanout627 (.A(_09504_),
    .X(net627));
 sg13g2_buf_2 fanout628 (.A(_09479_),
    .X(net628));
 sg13g2_buf_2 fanout629 (.A(_09461_),
    .X(net629));
 sg13g2_buf_2 fanout630 (.A(_09453_),
    .X(net630));
 sg13g2_buf_4 fanout631 (.X(net631),
    .A(_09390_));
 sg13g2_buf_2 fanout632 (.A(_09382_),
    .X(net632));
 sg13g2_buf_2 fanout633 (.A(_09343_),
    .X(net633));
 sg13g2_buf_2 fanout634 (.A(_08780_),
    .X(net634));
 sg13g2_buf_2 fanout635 (.A(_08666_),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(_08662_),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(_08604_),
    .X(net637));
 sg13g2_buf_2 fanout638 (.A(_08596_),
    .X(net638));
 sg13g2_buf_2 fanout639 (.A(_08589_),
    .X(net639));
 sg13g2_buf_2 fanout640 (.A(_08585_),
    .X(net640));
 sg13g2_buf_2 fanout641 (.A(_08579_),
    .X(net641));
 sg13g2_buf_2 fanout642 (.A(_08002_),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(_07165_),
    .X(net643));
 sg13g2_buf_2 fanout644 (.A(_06843_),
    .X(net644));
 sg13g2_buf_2 fanout645 (.A(_06239_),
    .X(net645));
 sg13g2_buf_2 fanout646 (.A(_06125_),
    .X(net646));
 sg13g2_buf_2 fanout647 (.A(_05979_),
    .X(net647));
 sg13g2_buf_2 fanout648 (.A(_05928_),
    .X(net648));
 sg13g2_buf_2 fanout649 (.A(_05868_),
    .X(net649));
 sg13g2_buf_2 fanout650 (.A(_05835_),
    .X(net650));
 sg13g2_buf_2 fanout651 (.A(_05434_),
    .X(net651));
 sg13g2_buf_2 fanout652 (.A(_05162_),
    .X(net652));
 sg13g2_buf_2 fanout653 (.A(_05131_),
    .X(net653));
 sg13g2_buf_2 fanout654 (.A(_04852_),
    .X(net654));
 sg13g2_buf_2 fanout655 (.A(_04818_),
    .X(net655));
 sg13g2_buf_2 fanout656 (.A(_03707_),
    .X(net656));
 sg13g2_buf_2 fanout657 (.A(_03701_),
    .X(net657));
 sg13g2_buf_2 fanout658 (.A(_03428_),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(_02965_),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(_02722_),
    .X(net660));
 sg13g2_buf_2 fanout661 (.A(_12319_),
    .X(net661));
 sg13g2_buf_2 fanout662 (.A(_12151_),
    .X(net662));
 sg13g2_buf_2 fanout663 (.A(_12110_),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(_12066_),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(_12059_),
    .X(net665));
 sg13g2_buf_2 fanout666 (.A(_12022_),
    .X(net666));
 sg13g2_buf_2 fanout667 (.A(_12004_),
    .X(net667));
 sg13g2_buf_2 fanout668 (.A(_11200_),
    .X(net668));
 sg13g2_buf_2 fanout669 (.A(_11174_),
    .X(net669));
 sg13g2_buf_2 fanout670 (.A(_11147_),
    .X(net670));
 sg13g2_buf_2 fanout671 (.A(_11085_),
    .X(net671));
 sg13g2_buf_2 fanout672 (.A(_11078_),
    .X(net672));
 sg13g2_buf_2 fanout673 (.A(_11052_),
    .X(net673));
 sg13g2_buf_2 fanout674 (.A(_10509_),
    .X(net674));
 sg13g2_buf_2 fanout675 (.A(_10486_),
    .X(net675));
 sg13g2_buf_2 fanout676 (.A(_10478_),
    .X(net676));
 sg13g2_buf_2 fanout677 (.A(_10443_),
    .X(net677));
 sg13g2_buf_4 fanout678 (.X(net678),
    .A(_10418_));
 sg13g2_buf_2 fanout679 (.A(_10412_),
    .X(net679));
 sg13g2_buf_2 fanout680 (.A(_10408_),
    .X(net680));
 sg13g2_buf_2 fanout681 (.A(_10173_),
    .X(net681));
 sg13g2_buf_2 fanout682 (.A(_10171_),
    .X(net682));
 sg13g2_buf_2 fanout683 (.A(_10126_),
    .X(net683));
 sg13g2_buf_2 fanout684 (.A(_10117_),
    .X(net684));
 sg13g2_buf_2 fanout685 (.A(_09990_),
    .X(net685));
 sg13g2_buf_2 fanout686 (.A(_09698_),
    .X(net686));
 sg13g2_buf_2 fanout687 (.A(_09682_),
    .X(net687));
 sg13g2_buf_8 fanout688 (.A(_09679_),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(_09671_),
    .X(net689));
 sg13g2_buf_8 fanout690 (.A(_09633_),
    .X(net690));
 sg13g2_buf_2 fanout691 (.A(_09580_),
    .X(net691));
 sg13g2_buf_8 fanout692 (.A(_09577_),
    .X(net692));
 sg13g2_buf_8 fanout693 (.A(_09573_),
    .X(net693));
 sg13g2_buf_8 fanout694 (.A(_09569_),
    .X(net694));
 sg13g2_buf_8 fanout695 (.A(_09556_),
    .X(net695));
 sg13g2_buf_8 fanout696 (.A(_09549_),
    .X(net696));
 sg13g2_buf_8 fanout697 (.A(_09544_),
    .X(net697));
 sg13g2_buf_4 fanout698 (.X(net698),
    .A(_09540_));
 sg13g2_buf_2 fanout699 (.A(_09529_),
    .X(net699));
 sg13g2_buf_2 fanout700 (.A(_09525_),
    .X(net700));
 sg13g2_buf_2 fanout701 (.A(_09521_),
    .X(net701));
 sg13g2_buf_2 fanout702 (.A(_09511_),
    .X(net702));
 sg13g2_buf_2 fanout703 (.A(_09507_),
    .X(net703));
 sg13g2_buf_2 fanout704 (.A(_09503_),
    .X(net704));
 sg13g2_buf_2 fanout705 (.A(_09447_),
    .X(net705));
 sg13g2_buf_2 fanout706 (.A(_09445_),
    .X(net706));
 sg13g2_buf_4 fanout707 (.X(net707),
    .A(_09389_));
 sg13g2_buf_2 fanout708 (.A(_09342_),
    .X(net708));
 sg13g2_buf_2 fanout709 (.A(_09283_),
    .X(net709));
 sg13g2_buf_4 fanout710 (.X(net710),
    .A(_09007_));
 sg13g2_buf_4 fanout711 (.X(net711),
    .A(_08802_));
 sg13g2_buf_4 fanout712 (.X(net712),
    .A(_08800_));
 sg13g2_buf_8 fanout713 (.A(_08714_),
    .X(net713));
 sg13g2_buf_8 fanout714 (.A(_08686_),
    .X(net714));
 sg13g2_buf_8 fanout715 (.A(_08619_),
    .X(net715));
 sg13g2_buf_8 fanout716 (.A(_08615_),
    .X(net716));
 sg13g2_buf_2 fanout717 (.A(_08578_),
    .X(net717));
 sg13g2_buf_8 fanout718 (.A(_08535_),
    .X(net718));
 sg13g2_buf_4 fanout719 (.X(net719),
    .A(_08530_));
 sg13g2_buf_2 fanout720 (.A(_06247_),
    .X(net720));
 sg13g2_buf_2 fanout721 (.A(_06245_),
    .X(net721));
 sg13g2_buf_2 fanout722 (.A(_06220_),
    .X(net722));
 sg13g2_buf_2 fanout723 (.A(_06218_),
    .X(net723));
 sg13g2_buf_2 fanout724 (.A(_06217_),
    .X(net724));
 sg13g2_buf_2 fanout725 (.A(_06216_),
    .X(net725));
 sg13g2_buf_2 fanout726 (.A(_06214_),
    .X(net726));
 sg13g2_buf_2 fanout727 (.A(_06133_),
    .X(net727));
 sg13g2_buf_2 fanout728 (.A(_06131_),
    .X(net728));
 sg13g2_buf_2 fanout729 (.A(_06104_),
    .X(net729));
 sg13g2_buf_2 fanout730 (.A(_06102_),
    .X(net730));
 sg13g2_buf_2 fanout731 (.A(_06101_),
    .X(net731));
 sg13g2_buf_2 fanout732 (.A(_06100_),
    .X(net732));
 sg13g2_buf_2 fanout733 (.A(_06098_),
    .X(net733));
 sg13g2_buf_2 fanout734 (.A(_06033_),
    .X(net734));
 sg13g2_buf_2 fanout735 (.A(_05983_),
    .X(net735));
 sg13g2_buf_2 fanout736 (.A(_05934_),
    .X(net736));
 sg13g2_buf_2 fanout737 (.A(_05875_),
    .X(net737));
 sg13g2_buf_2 fanout738 (.A(_05855_),
    .X(net738));
 sg13g2_buf_2 fanout739 (.A(_04741_),
    .X(net739));
 sg13g2_buf_2 fanout740 (.A(_03700_),
    .X(net740));
 sg13g2_buf_2 fanout741 (.A(_03698_),
    .X(net741));
 sg13g2_buf_2 fanout742 (.A(_03695_),
    .X(net742));
 sg13g2_buf_2 fanout743 (.A(_03430_),
    .X(net743));
 sg13g2_buf_2 fanout744 (.A(_03419_),
    .X(net744));
 sg13g2_buf_2 fanout745 (.A(_03247_),
    .X(net745));
 sg13g2_buf_2 fanout746 (.A(_02997_),
    .X(net746));
 sg13g2_buf_2 fanout747 (.A(_02996_),
    .X(net747));
 sg13g2_buf_2 fanout748 (.A(_02995_),
    .X(net748));
 sg13g2_buf_2 fanout749 (.A(_02972_),
    .X(net749));
 sg13g2_buf_2 fanout750 (.A(_02971_),
    .X(net750));
 sg13g2_buf_2 fanout751 (.A(_02969_),
    .X(net751));
 sg13g2_buf_2 fanout752 (.A(_02963_),
    .X(net752));
 sg13g2_buf_2 fanout753 (.A(_02957_),
    .X(net753));
 sg13g2_buf_2 fanout754 (.A(_02955_),
    .X(net754));
 sg13g2_buf_2 fanout755 (.A(_02952_),
    .X(net755));
 sg13g2_buf_2 fanout756 (.A(_02944_),
    .X(net756));
 sg13g2_buf_2 fanout757 (.A(_12771_),
    .X(net757));
 sg13g2_buf_2 fanout758 (.A(_12656_),
    .X(net758));
 sg13g2_buf_2 fanout759 (.A(_12447_),
    .X(net759));
 sg13g2_buf_2 fanout760 (.A(_12062_),
    .X(net760));
 sg13g2_buf_2 fanout761 (.A(_12058_),
    .X(net761));
 sg13g2_buf_2 fanout762 (.A(_11682_),
    .X(net762));
 sg13g2_buf_2 fanout763 (.A(_11215_),
    .X(net763));
 sg13g2_buf_2 fanout764 (.A(_11152_),
    .X(net764));
 sg13g2_buf_2 fanout765 (.A(_11104_),
    .X(net765));
 sg13g2_buf_2 fanout766 (.A(_11100_),
    .X(net766));
 sg13g2_buf_2 fanout767 (.A(_11094_),
    .X(net767));
 sg13g2_buf_2 fanout768 (.A(_11092_),
    .X(net768));
 sg13g2_buf_2 fanout769 (.A(_11080_),
    .X(net769));
 sg13g2_buf_2 fanout770 (.A(_11077_),
    .X(net770));
 sg13g2_buf_2 fanout771 (.A(_11073_),
    .X(net771));
 sg13g2_buf_2 fanout772 (.A(_11063_),
    .X(net772));
 sg13g2_buf_2 fanout773 (.A(_11059_),
    .X(net773));
 sg13g2_buf_2 fanout774 (.A(_10598_),
    .X(net774));
 sg13g2_buf_2 fanout775 (.A(_10594_),
    .X(net775));
 sg13g2_buf_2 fanout776 (.A(_10508_),
    .X(net776));
 sg13g2_buf_2 fanout777 (.A(_10492_),
    .X(net777));
 sg13g2_buf_2 fanout778 (.A(_10477_),
    .X(net778));
 sg13g2_buf_2 fanout779 (.A(_10475_),
    .X(net779));
 sg13g2_buf_2 fanout780 (.A(_10442_),
    .X(net780));
 sg13g2_buf_2 fanout781 (.A(_10430_),
    .X(net781));
 sg13g2_buf_2 fanout782 (.A(_10417_),
    .X(net782));
 sg13g2_buf_2 fanout783 (.A(_10411_),
    .X(net783));
 sg13g2_buf_2 fanout784 (.A(_10407_),
    .X(net784));
 sg13g2_buf_2 fanout785 (.A(_10176_),
    .X(net785));
 sg13g2_buf_2 fanout786 (.A(_10170_),
    .X(net786));
 sg13g2_buf_2 fanout787 (.A(_10116_),
    .X(net787));
 sg13g2_buf_2 fanout788 (.A(_09952_),
    .X(net788));
 sg13g2_buf_8 fanout789 (.A(_09753_),
    .X(net789));
 sg13g2_buf_4 fanout790 (.X(net790),
    .A(_09684_));
 sg13g2_buf_2 fanout791 (.A(_09680_),
    .X(net791));
 sg13g2_buf_8 fanout792 (.A(_09637_),
    .X(net792));
 sg13g2_buf_4 fanout793 (.X(net793),
    .A(_09634_));
 sg13g2_buf_4 fanout794 (.X(net794),
    .A(_09576_));
 sg13g2_buf_4 fanout795 (.X(net795),
    .A(_09570_));
 sg13g2_buf_2 fanout796 (.A(_09568_),
    .X(net796));
 sg13g2_buf_4 fanout797 (.X(net797),
    .A(_09557_));
 sg13g2_buf_4 fanout798 (.X(net798),
    .A(_09552_));
 sg13g2_buf_4 fanout799 (.X(net799),
    .A(_09550_));
 sg13g2_buf_4 fanout800 (.X(net800),
    .A(_09546_));
 sg13g2_buf_4 fanout801 (.X(net801),
    .A(_09539_));
 sg13g2_buf_2 fanout802 (.A(_09485_),
    .X(net802));
 sg13g2_buf_4 fanout803 (.X(net803),
    .A(_09444_));
 sg13g2_buf_2 fanout804 (.A(_09388_),
    .X(net804));
 sg13g2_buf_4 fanout805 (.X(net805),
    .A(_09379_));
 sg13g2_buf_2 fanout806 (.A(_09349_),
    .X(net806));
 sg13g2_buf_2 fanout807 (.A(_09341_),
    .X(net807));
 sg13g2_buf_2 fanout808 (.A(_09065_),
    .X(net808));
 sg13g2_buf_2 fanout809 (.A(_08978_),
    .X(net809));
 sg13g2_buf_2 fanout810 (.A(_08801_),
    .X(net810));
 sg13g2_buf_2 fanout811 (.A(_08762_),
    .X(net811));
 sg13g2_buf_4 fanout812 (.X(net812),
    .A(_08732_));
 sg13g2_buf_4 fanout813 (.X(net813),
    .A(_08715_));
 sg13g2_buf_2 fanout814 (.A(_08706_),
    .X(net814));
 sg13g2_buf_4 fanout815 (.X(net815),
    .A(_08693_));
 sg13g2_buf_4 fanout816 (.X(net816),
    .A(_08689_));
 sg13g2_buf_4 fanout817 (.X(net817),
    .A(_08687_));
 sg13g2_buf_8 fanout818 (.A(_08648_),
    .X(net818));
 sg13g2_buf_4 fanout819 (.X(net819),
    .A(_08622_));
 sg13g2_buf_4 fanout820 (.X(net820),
    .A(_08617_));
 sg13g2_buf_4 fanout821 (.X(net821),
    .A(_08614_));
 sg13g2_buf_4 fanout822 (.X(net822),
    .A(_08608_));
 sg13g2_buf_2 fanout823 (.A(_08601_),
    .X(net823));
 sg13g2_buf_8 fanout824 (.A(_08544_),
    .X(net824));
 sg13g2_buf_4 fanout825 (.X(net825),
    .A(_08538_));
 sg13g2_buf_4 fanout826 (.X(net826),
    .A(_08534_));
 sg13g2_buf_4 fanout827 (.X(net827),
    .A(_08529_));
 sg13g2_buf_2 fanout828 (.A(_08003_),
    .X(net828));
 sg13g2_buf_2 fanout829 (.A(_07044_),
    .X(net829));
 sg13g2_buf_2 fanout830 (.A(_06913_),
    .X(net830));
 sg13g2_buf_2 fanout831 (.A(_06849_),
    .X(net831));
 sg13g2_buf_2 fanout832 (.A(_06548_),
    .X(net832));
 sg13g2_buf_2 fanout833 (.A(_06547_),
    .X(net833));
 sg13g2_buf_2 fanout834 (.A(_06546_),
    .X(net834));
 sg13g2_buf_2 fanout835 (.A(_06544_),
    .X(net835));
 sg13g2_buf_2 fanout836 (.A(_06513_),
    .X(net836));
 sg13g2_buf_2 fanout837 (.A(_06512_),
    .X(net837));
 sg13g2_buf_2 fanout838 (.A(_06510_),
    .X(net838));
 sg13g2_buf_2 fanout839 (.A(_06508_),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(_06499_),
    .X(net840));
 sg13g2_buf_2 fanout841 (.A(_06498_),
    .X(net841));
 sg13g2_buf_2 fanout842 (.A(_06497_),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(_06495_),
    .X(net843));
 sg13g2_buf_2 fanout844 (.A(_06478_),
    .X(net844));
 sg13g2_buf_2 fanout845 (.A(_06475_),
    .X(net845));
 sg13g2_buf_2 fanout846 (.A(_06474_),
    .X(net846));
 sg13g2_buf_2 fanout847 (.A(_06473_),
    .X(net847));
 sg13g2_buf_2 fanout848 (.A(_06470_),
    .X(net848));
 sg13g2_buf_2 fanout849 (.A(_06469_),
    .X(net849));
 sg13g2_buf_2 fanout850 (.A(_06465_),
    .X(net850));
 sg13g2_buf_2 fanout851 (.A(_06460_),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(_06438_),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(_06432_),
    .X(net853));
 sg13g2_buf_2 fanout854 (.A(_06426_),
    .X(net854));
 sg13g2_buf_2 fanout855 (.A(_06413_),
    .X(net855));
 sg13g2_buf_2 fanout856 (.A(_06267_),
    .X(net856));
 sg13g2_buf_2 fanout857 (.A(_06219_),
    .X(net857));
 sg13g2_buf_2 fanout858 (.A(_06152_),
    .X(net858));
 sg13g2_buf_2 fanout859 (.A(_06103_),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(_05987_),
    .X(net860));
 sg13g2_buf_2 fanout861 (.A(_05973_),
    .X(net861));
 sg13g2_buf_2 fanout862 (.A(_05966_),
    .X(net862));
 sg13g2_buf_2 fanout863 (.A(_05965_),
    .X(net863));
 sg13g2_buf_2 fanout864 (.A(_05939_),
    .X(net864));
 sg13g2_buf_2 fanout865 (.A(_05922_),
    .X(net865));
 sg13g2_buf_2 fanout866 (.A(_05915_),
    .X(net866));
 sg13g2_buf_2 fanout867 (.A(_05914_),
    .X(net867));
 sg13g2_buf_2 fanout868 (.A(_05894_),
    .X(net868));
 sg13g2_buf_2 fanout869 (.A(_05883_),
    .X(net869));
 sg13g2_buf_2 fanout870 (.A(_05823_),
    .X(net870));
 sg13g2_buf_2 fanout871 (.A(_05761_),
    .X(net871));
 sg13g2_buf_2 fanout872 (.A(_04887_),
    .X(net872));
 sg13g2_buf_2 fanout873 (.A(_04742_),
    .X(net873));
 sg13g2_buf_2 fanout874 (.A(_04740_),
    .X(net874));
 sg13g2_buf_2 fanout875 (.A(_03697_),
    .X(net875));
 sg13g2_buf_2 fanout876 (.A(_03694_),
    .X(net876));
 sg13g2_buf_2 fanout877 (.A(_03586_),
    .X(net877));
 sg13g2_buf_2 fanout878 (.A(_03455_),
    .X(net878));
 sg13g2_buf_2 fanout879 (.A(_03446_),
    .X(net879));
 sg13g2_buf_2 fanout880 (.A(_03418_),
    .X(net880));
 sg13g2_buf_2 fanout881 (.A(_02998_),
    .X(net881));
 sg13g2_buf_2 fanout882 (.A(_02977_),
    .X(net882));
 sg13g2_buf_2 fanout883 (.A(_02975_),
    .X(net883));
 sg13g2_buf_2 fanout884 (.A(_02974_),
    .X(net884));
 sg13g2_buf_2 fanout885 (.A(_02962_),
    .X(net885));
 sg13g2_buf_2 fanout886 (.A(_02961_),
    .X(net886));
 sg13g2_buf_2 fanout887 (.A(_02956_),
    .X(net887));
 sg13g2_buf_2 fanout888 (.A(_02954_),
    .X(net888));
 sg13g2_buf_2 fanout889 (.A(_02951_),
    .X(net889));
 sg13g2_buf_2 fanout890 (.A(_02943_),
    .X(net890));
 sg13g2_buf_2 fanout891 (.A(_02925_),
    .X(net891));
 sg13g2_buf_2 fanout892 (.A(_12814_),
    .X(net892));
 sg13g2_buf_2 fanout893 (.A(_12807_),
    .X(net893));
 sg13g2_buf_2 fanout894 (.A(_12694_),
    .X(net894));
 sg13g2_buf_2 fanout895 (.A(_12226_),
    .X(net895));
 sg13g2_buf_2 fanout896 (.A(_12215_),
    .X(net896));
 sg13g2_buf_2 fanout897 (.A(_12141_),
    .X(net897));
 sg13g2_buf_2 fanout898 (.A(_12080_),
    .X(net898));
 sg13g2_buf_2 fanout899 (.A(_12057_),
    .X(net899));
 sg13g2_buf_2 fanout900 (.A(_12051_),
    .X(net900));
 sg13g2_buf_2 fanout901 (.A(_11087_),
    .X(net901));
 sg13g2_buf_2 fanout902 (.A(_11069_),
    .X(net902));
 sg13g2_buf_2 fanout903 (.A(_11058_),
    .X(net903));
 sg13g2_buf_2 fanout904 (.A(_11055_),
    .X(net904));
 sg13g2_buf_2 fanout905 (.A(_11050_),
    .X(net905));
 sg13g2_buf_2 fanout906 (.A(_10528_),
    .X(net906));
 sg13g2_buf_2 fanout907 (.A(_10504_),
    .X(net907));
 sg13g2_buf_2 fanout908 (.A(_10438_),
    .X(net908));
 sg13g2_buf_2 fanout909 (.A(_10426_),
    .X(net909));
 sg13g2_buf_2 fanout910 (.A(_10424_),
    .X(net910));
 sg13g2_buf_2 fanout911 (.A(_10422_),
    .X(net911));
 sg13g2_buf_2 fanout912 (.A(_10416_),
    .X(net912));
 sg13g2_buf_2 fanout913 (.A(_10410_),
    .X(net913));
 sg13g2_buf_2 fanout914 (.A(_10406_),
    .X(net914));
 sg13g2_buf_2 fanout915 (.A(_10374_),
    .X(net915));
 sg13g2_buf_2 fanout916 (.A(_10282_),
    .X(net916));
 sg13g2_buf_2 fanout917 (.A(_10264_),
    .X(net917));
 sg13g2_buf_2 fanout918 (.A(_10244_),
    .X(net918));
 sg13g2_buf_2 fanout919 (.A(_10241_),
    .X(net919));
 sg13g2_buf_2 fanout920 (.A(_10202_),
    .X(net920));
 sg13g2_buf_2 fanout921 (.A(_10196_),
    .X(net921));
 sg13g2_buf_2 fanout922 (.A(_10175_),
    .X(net922));
 sg13g2_buf_2 fanout923 (.A(_10115_),
    .X(net923));
 sg13g2_buf_4 fanout924 (.X(net924),
    .A(_09754_));
 sg13g2_buf_4 fanout925 (.X(net925),
    .A(_09652_));
 sg13g2_buf_2 fanout926 (.A(_09632_),
    .X(net926));
 sg13g2_buf_4 fanout927 (.X(net927),
    .A(_09542_));
 sg13g2_buf_2 fanout928 (.A(_09514_),
    .X(net928));
 sg13g2_buf_2 fanout929 (.A(_09495_),
    .X(net929));
 sg13g2_buf_4 fanout930 (.X(net930),
    .A(_09443_));
 sg13g2_buf_2 fanout931 (.A(_09386_),
    .X(net931));
 sg13g2_buf_2 fanout932 (.A(_09378_),
    .X(net932));
 sg13g2_buf_2 fanout933 (.A(_09352_),
    .X(net933));
 sg13g2_buf_2 fanout934 (.A(_09340_),
    .X(net934));
 sg13g2_buf_2 fanout935 (.A(_09064_),
    .X(net935));
 sg13g2_buf_2 fanout936 (.A(_09013_),
    .X(net936));
 sg13g2_buf_2 fanout937 (.A(_08977_),
    .X(net937));
 sg13g2_buf_2 fanout938 (.A(_08808_),
    .X(net938));
 sg13g2_buf_2 fanout939 (.A(_08779_),
    .X(net939));
 sg13g2_buf_2 fanout940 (.A(_08759_),
    .X(net940));
 sg13g2_buf_2 fanout941 (.A(_08679_),
    .X(net941));
 sg13g2_buf_4 fanout942 (.X(net942),
    .A(_08671_));
 sg13g2_buf_4 fanout943 (.X(net943),
    .A(_08670_));
 sg13g2_buf_2 fanout944 (.A(_08649_),
    .X(net944));
 sg13g2_buf_2 fanout945 (.A(_08616_),
    .X(net945));
 sg13g2_buf_4 fanout946 (.X(net946),
    .A(_08606_));
 sg13g2_buf_2 fanout947 (.A(_08600_),
    .X(net947));
 sg13g2_buf_2 fanout948 (.A(_08592_),
    .X(net948));
 sg13g2_buf_2 fanout949 (.A(_08582_),
    .X(net949));
 sg13g2_buf_2 fanout950 (.A(_08566_),
    .X(net950));
 sg13g2_buf_4 fanout951 (.X(net951),
    .A(_08551_));
 sg13g2_buf_4 fanout952 (.X(net952),
    .A(_08546_));
 sg13g2_buf_4 fanout953 (.X(net953),
    .A(_08543_));
 sg13g2_buf_4 fanout954 (.X(net954),
    .A(_08537_));
 sg13g2_buf_2 fanout955 (.A(_08533_),
    .X(net955));
 sg13g2_buf_4 fanout956 (.X(net956),
    .A(_08405_));
 sg13g2_buf_2 fanout957 (.A(_08392_),
    .X(net957));
 sg13g2_buf_2 fanout958 (.A(_07143_),
    .X(net958));
 sg13g2_buf_2 fanout959 (.A(_07134_),
    .X(net959));
 sg13g2_buf_2 fanout960 (.A(_07132_),
    .X(net960));
 sg13g2_buf_2 fanout961 (.A(_07120_),
    .X(net961));
 sg13g2_buf_2 fanout962 (.A(_07117_),
    .X(net962));
 sg13g2_buf_2 fanout963 (.A(_07033_),
    .X(net963));
 sg13g2_buf_2 fanout964 (.A(_07031_),
    .X(net964));
 sg13g2_buf_2 fanout965 (.A(_06854_),
    .X(net965));
 sg13g2_buf_2 fanout966 (.A(_06824_),
    .X(net966));
 sg13g2_buf_2 fanout967 (.A(_05967_),
    .X(net967));
 sg13g2_buf_2 fanout968 (.A(_05946_),
    .X(net968));
 sg13g2_buf_2 fanout969 (.A(_05916_),
    .X(net969));
 sg13g2_buf_2 fanout970 (.A(_05846_),
    .X(net970));
 sg13g2_buf_2 fanout971 (.A(_05836_),
    .X(net971));
 sg13g2_buf_2 fanout972 (.A(_05829_),
    .X(net972));
 sg13g2_buf_2 fanout973 (.A(_05815_),
    .X(net973));
 sg13g2_buf_2 fanout974 (.A(_05748_),
    .X(net974));
 sg13g2_buf_2 fanout975 (.A(_05311_),
    .X(net975));
 sg13g2_buf_2 fanout976 (.A(_05137_),
    .X(net976));
 sg13g2_buf_2 fanout977 (.A(_04913_),
    .X(net977));
 sg13g2_buf_2 fanout978 (.A(_04732_),
    .X(net978));
 sg13g2_buf_2 fanout979 (.A(_04278_),
    .X(net979));
 sg13g2_buf_2 fanout980 (.A(_04211_),
    .X(net980));
 sg13g2_buf_2 fanout981 (.A(_02976_),
    .X(net981));
 sg13g2_buf_2 fanout982 (.A(_02960_),
    .X(net982));
 sg13g2_buf_2 fanout983 (.A(_02953_),
    .X(net983));
 sg13g2_buf_4 fanout984 (.X(net984),
    .A(_02950_));
 sg13g2_buf_2 fanout985 (.A(_02785_),
    .X(net985));
 sg13g2_buf_2 fanout986 (.A(_12751_),
    .X(net986));
 sg13g2_buf_2 fanout987 (.A(_12748_),
    .X(net987));
 sg13g2_buf_2 fanout988 (.A(_12740_),
    .X(net988));
 sg13g2_buf_2 fanout989 (.A(_12711_),
    .X(net989));
 sg13g2_buf_2 fanout990 (.A(_12705_),
    .X(net990));
 sg13g2_buf_2 fanout991 (.A(_12613_),
    .X(net991));
 sg13g2_buf_2 fanout992 (.A(_12425_),
    .X(net992));
 sg13g2_buf_2 fanout993 (.A(_12417_),
    .X(net993));
 sg13g2_buf_2 fanout994 (.A(_12390_),
    .X(net994));
 sg13g2_buf_2 fanout995 (.A(_12386_),
    .X(net995));
 sg13g2_buf_2 fanout996 (.A(_12383_),
    .X(net996));
 sg13g2_buf_2 fanout997 (.A(_12381_),
    .X(net997));
 sg13g2_buf_2 fanout998 (.A(_12376_),
    .X(net998));
 sg13g2_buf_2 fanout999 (.A(_12256_),
    .X(net999));
 sg13g2_buf_2 fanout1000 (.A(_12252_),
    .X(net1000));
 sg13g2_buf_2 fanout1001 (.A(_12248_),
    .X(net1001));
 sg13g2_buf_2 fanout1002 (.A(_12244_),
    .X(net1002));
 sg13g2_buf_2 fanout1003 (.A(_12232_),
    .X(net1003));
 sg13g2_buf_4 fanout1004 (.X(net1004),
    .A(_12229_));
 sg13g2_buf_4 fanout1005 (.X(net1005),
    .A(_12223_));
 sg13g2_buf_4 fanout1006 (.X(net1006),
    .A(_12218_));
 sg13g2_buf_2 fanout1007 (.A(_12208_),
    .X(net1007));
 sg13g2_buf_2 fanout1008 (.A(_12177_),
    .X(net1008));
 sg13g2_buf_2 fanout1009 (.A(_12131_),
    .X(net1009));
 sg13g2_buf_4 fanout1010 (.X(net1010),
    .A(_12127_));
 sg13g2_buf_2 fanout1011 (.A(_12117_),
    .X(net1011));
 sg13g2_buf_2 fanout1012 (.A(_12041_),
    .X(net1012));
 sg13g2_buf_2 fanout1013 (.A(_12040_),
    .X(net1013));
 sg13g2_buf_2 fanout1014 (.A(_12038_),
    .X(net1014));
 sg13g2_buf_2 fanout1015 (.A(_12034_),
    .X(net1015));
 sg13g2_buf_2 fanout1016 (.A(_11469_),
    .X(net1016));
 sg13g2_buf_2 fanout1017 (.A(_11098_),
    .X(net1017));
 sg13g2_buf_2 fanout1018 (.A(_11068_),
    .X(net1018));
 sg13g2_buf_2 fanout1019 (.A(_11057_),
    .X(net1019));
 sg13g2_buf_2 fanout1020 (.A(_11054_),
    .X(net1020));
 sg13g2_buf_2 fanout1021 (.A(_11049_),
    .X(net1021));
 sg13g2_buf_2 fanout1022 (.A(_10572_),
    .X(net1022));
 sg13g2_buf_2 fanout1023 (.A(_10569_),
    .X(net1023));
 sg13g2_buf_2 fanout1024 (.A(_10542_),
    .X(net1024));
 sg13g2_buf_2 fanout1025 (.A(_10409_),
    .X(net1025));
 sg13g2_buf_2 fanout1026 (.A(_10401_),
    .X(net1026));
 sg13g2_buf_2 fanout1027 (.A(_10400_),
    .X(net1027));
 sg13g2_buf_2 fanout1028 (.A(_10395_),
    .X(net1028));
 sg13g2_buf_2 fanout1029 (.A(_10373_),
    .X(net1029));
 sg13g2_buf_2 fanout1030 (.A(_10370_),
    .X(net1030));
 sg13g2_buf_2 fanout1031 (.A(_10288_),
    .X(net1031));
 sg13g2_buf_2 fanout1032 (.A(_10275_),
    .X(net1032));
 sg13g2_buf_2 fanout1033 (.A(_10269_),
    .X(net1033));
 sg13g2_buf_2 fanout1034 (.A(_10230_),
    .X(net1034));
 sg13g2_buf_2 fanout1035 (.A(_10227_),
    .X(net1035));
 sg13g2_buf_2 fanout1036 (.A(_10221_),
    .X(net1036));
 sg13g2_buf_2 fanout1037 (.A(_10215_),
    .X(net1037));
 sg13g2_buf_2 fanout1038 (.A(_10209_),
    .X(net1038));
 sg13g2_buf_2 fanout1039 (.A(_10201_),
    .X(net1039));
 sg13g2_buf_2 fanout1040 (.A(_10195_),
    .X(net1040));
 sg13g2_buf_2 fanout1041 (.A(_10187_),
    .X(net1041));
 sg13g2_buf_2 fanout1042 (.A(_10123_),
    .X(net1042));
 sg13g2_buf_2 fanout1043 (.A(_10037_),
    .X(net1043));
 sg13g2_buf_2 fanout1044 (.A(_10024_),
    .X(net1044));
 sg13g2_buf_2 fanout1045 (.A(_10020_),
    .X(net1045));
 sg13g2_buf_2 fanout1046 (.A(_09992_),
    .X(net1046));
 sg13g2_buf_2 fanout1047 (.A(_09963_),
    .X(net1047));
 sg13g2_buf_2 fanout1048 (.A(_09613_),
    .X(net1048));
 sg13g2_buf_2 fanout1049 (.A(_09432_),
    .X(net1049));
 sg13g2_buf_2 fanout1050 (.A(_09430_),
    .X(net1050));
 sg13g2_buf_2 fanout1051 (.A(_09380_),
    .X(net1051));
 sg13g2_buf_2 fanout1052 (.A(_09358_),
    .X(net1052));
 sg13g2_buf_2 fanout1053 (.A(_09357_),
    .X(net1053));
 sg13g2_buf_2 fanout1054 (.A(_09347_),
    .X(net1054));
 sg13g2_buf_2 fanout1055 (.A(_09339_),
    .X(net1055));
 sg13g2_buf_4 fanout1056 (.X(net1056),
    .A(_09279_));
 sg13g2_buf_2 fanout1057 (.A(_09263_),
    .X(net1057));
 sg13g2_buf_2 fanout1058 (.A(_09157_),
    .X(net1058));
 sg13g2_buf_2 fanout1059 (.A(_09120_),
    .X(net1059));
 sg13g2_buf_2 fanout1060 (.A(_08976_),
    .X(net1060));
 sg13g2_buf_4 fanout1061 (.X(net1061),
    .A(_08669_));
 sg13g2_buf_2 fanout1062 (.A(_08645_),
    .X(net1062));
 sg13g2_buf_2 fanout1063 (.A(_08605_),
    .X(net1063));
 sg13g2_buf_4 fanout1064 (.X(net1064),
    .A(_08599_));
 sg13g2_buf_4 fanout1065 (.X(net1065),
    .A(_08545_));
 sg13g2_buf_2 fanout1066 (.A(_08536_),
    .X(net1066));
 sg13g2_buf_2 fanout1067 (.A(_08532_),
    .X(net1067));
 sg13g2_buf_2 fanout1068 (.A(_08531_),
    .X(net1068));
 sg13g2_buf_2 fanout1069 (.A(_08457_),
    .X(net1069));
 sg13g2_buf_4 fanout1070 (.X(net1070),
    .A(_08449_));
 sg13g2_buf_4 fanout1071 (.X(net1071),
    .A(_08439_));
 sg13g2_buf_4 fanout1072 (.X(net1072),
    .A(_08422_));
 sg13g2_buf_4 fanout1073 (.X(net1073),
    .A(_08384_));
 sg13g2_buf_2 fanout1074 (.A(_08381_),
    .X(net1074));
 sg13g2_buf_4 fanout1075 (.X(net1075),
    .A(_08377_));
 sg13g2_buf_2 fanout1076 (.A(_08175_),
    .X(net1076));
 sg13g2_buf_2 fanout1077 (.A(_08172_),
    .X(net1077));
 sg13g2_buf_2 fanout1078 (.A(_08158_),
    .X(net1078));
 sg13g2_buf_2 fanout1079 (.A(_07867_),
    .X(net1079));
 sg13g2_buf_2 fanout1080 (.A(_07224_),
    .X(net1080));
 sg13g2_buf_2 fanout1081 (.A(_07118_),
    .X(net1081));
 sg13g2_buf_2 fanout1082 (.A(_07116_),
    .X(net1082));
 sg13g2_buf_2 fanout1083 (.A(_05803_),
    .X(net1083));
 sg13g2_buf_2 fanout1084 (.A(_12653_),
    .X(net1084));
 sg13g2_buf_2 fanout1085 (.A(_12650_),
    .X(net1085));
 sg13g2_buf_2 fanout1086 (.A(_12638_),
    .X(net1086));
 sg13g2_buf_2 fanout1087 (.A(_12635_),
    .X(net1087));
 sg13g2_buf_2 fanout1088 (.A(_12405_),
    .X(net1088));
 sg13g2_buf_2 fanout1089 (.A(_12400_),
    .X(net1089));
 sg13g2_buf_2 fanout1090 (.A(_12351_),
    .X(net1090));
 sg13g2_buf_2 fanout1091 (.A(_12348_),
    .X(net1091));
 sg13g2_buf_2 fanout1092 (.A(_12228_),
    .X(net1092));
 sg13g2_buf_2 fanout1093 (.A(_12222_),
    .X(net1093));
 sg13g2_buf_2 fanout1094 (.A(_12217_),
    .X(net1094));
 sg13g2_buf_1 fanout1095 (.A(_12189_),
    .X(net1095));
 sg13g2_buf_1 fanout1096 (.A(_12176_),
    .X(net1096));
 sg13g2_buf_1 fanout1097 (.A(_12169_),
    .X(net1097));
 sg13g2_buf_1 fanout1098 (.A(_12158_),
    .X(net1098));
 sg13g2_buf_2 fanout1099 (.A(_12132_),
    .X(net1099));
 sg13g2_buf_2 fanout1100 (.A(_12129_),
    .X(net1100));
 sg13g2_buf_2 fanout1101 (.A(_12126_),
    .X(net1101));
 sg13g2_buf_2 fanout1102 (.A(_12101_),
    .X(net1102));
 sg13g2_buf_2 fanout1103 (.A(_12085_),
    .X(net1103));
 sg13g2_buf_2 fanout1104 (.A(_12083_),
    .X(net1104));
 sg13g2_buf_2 fanout1105 (.A(_12076_),
    .X(net1105));
 sg13g2_buf_2 fanout1106 (.A(_10754_),
    .X(net1106));
 sg13g2_buf_2 fanout1107 (.A(_10645_),
    .X(net1107));
 sg13g2_buf_2 fanout1108 (.A(_10637_),
    .X(net1108));
 sg13g2_buf_2 fanout1109 (.A(_10584_),
    .X(net1109));
 sg13g2_buf_2 fanout1110 (.A(_10379_),
    .X(net1110));
 sg13g2_buf_2 fanout1111 (.A(_10353_),
    .X(net1111));
 sg13g2_buf_2 fanout1112 (.A(_10352_),
    .X(net1112));
 sg13g2_buf_2 fanout1113 (.A(_10350_),
    .X(net1113));
 sg13g2_buf_2 fanout1114 (.A(_10349_),
    .X(net1114));
 sg13g2_buf_2 fanout1115 (.A(_10347_),
    .X(net1115));
 sg13g2_buf_2 fanout1116 (.A(_10208_),
    .X(net1116));
 sg13g2_buf_2 fanout1117 (.A(_10036_),
    .X(net1117));
 sg13g2_buf_2 fanout1118 (.A(_10023_),
    .X(net1118));
 sg13g2_buf_2 fanout1119 (.A(_09987_),
    .X(net1119));
 sg13g2_buf_2 fanout1120 (.A(_09828_),
    .X(net1120));
 sg13g2_buf_2 fanout1121 (.A(_09490_),
    .X(net1121));
 sg13g2_buf_2 fanout1122 (.A(_09476_),
    .X(net1122));
 sg13g2_buf_2 fanout1123 (.A(_09440_),
    .X(net1123));
 sg13g2_buf_2 fanout1124 (.A(_09365_),
    .X(net1124));
 sg13g2_buf_2 fanout1125 (.A(_09262_),
    .X(net1125));
 sg13g2_buf_2 fanout1126 (.A(_08564_),
    .X(net1126));
 sg13g2_buf_4 fanout1127 (.X(net1127),
    .A(_08561_));
 sg13g2_buf_2 fanout1128 (.A(_08559_),
    .X(net1128));
 sg13g2_buf_2 fanout1129 (.A(_08452_),
    .X(net1129));
 sg13g2_buf_2 fanout1130 (.A(_08441_),
    .X(net1130));
 sg13g2_buf_4 fanout1131 (.X(net1131),
    .A(_08438_));
 sg13g2_buf_2 fanout1132 (.A(_08394_),
    .X(net1132));
 sg13g2_buf_4 fanout1133 (.X(net1133),
    .A(_08379_));
 sg13g2_buf_2 fanout1134 (.A(_08375_),
    .X(net1134));
 sg13g2_buf_2 fanout1135 (.A(_08372_),
    .X(net1135));
 sg13g2_tiehi _27759__1136 (.L_HI(net1136));
 sg13g2_tiehi _27760__1137 (.L_HI(net1137));
 sg13g2_tiehi _27761__1138 (.L_HI(net1138));
 sg13g2_tiehi _27762__1139 (.L_HI(net1139));
 sg13g2_tiehi _27763__1140 (.L_HI(net1140));
 sg13g2_tiehi \cpu.dcache.r_data[0][0]$_DFFE_PP__1141  (.L_HI(net1141));
 sg13g2_tiehi \cpu.dcache.r_data[0][10]$_DFFE_PP__1142  (.L_HI(net1142));
 sg13g2_tiehi \cpu.dcache.r_data[0][11]$_DFFE_PP__1143  (.L_HI(net1143));
 sg13g2_tiehi \cpu.dcache.r_data[0][12]$_DFFE_PP__1144  (.L_HI(net1144));
 sg13g2_tiehi \cpu.dcache.r_data[0][13]$_DFFE_PP__1145  (.L_HI(net1145));
 sg13g2_tiehi \cpu.dcache.r_data[0][14]$_DFFE_PP__1146  (.L_HI(net1146));
 sg13g2_tiehi \cpu.dcache.r_data[0][15]$_DFFE_PP__1147  (.L_HI(net1147));
 sg13g2_tiehi \cpu.dcache.r_data[0][16]$_DFFE_PP__1148  (.L_HI(net1148));
 sg13g2_tiehi \cpu.dcache.r_data[0][17]$_DFFE_PP__1149  (.L_HI(net1149));
 sg13g2_tiehi \cpu.dcache.r_data[0][18]$_DFFE_PP__1150  (.L_HI(net1150));
 sg13g2_tiehi \cpu.dcache.r_data[0][19]$_DFFE_PP__1151  (.L_HI(net1151));
 sg13g2_tiehi \cpu.dcache.r_data[0][1]$_DFFE_PP__1152  (.L_HI(net1152));
 sg13g2_tiehi \cpu.dcache.r_data[0][20]$_DFFE_PP__1153  (.L_HI(net1153));
 sg13g2_tiehi \cpu.dcache.r_data[0][21]$_DFFE_PP__1154  (.L_HI(net1154));
 sg13g2_tiehi \cpu.dcache.r_data[0][22]$_DFFE_PP__1155  (.L_HI(net1155));
 sg13g2_tiehi \cpu.dcache.r_data[0][23]$_DFFE_PP__1156  (.L_HI(net1156));
 sg13g2_tiehi \cpu.dcache.r_data[0][24]$_DFFE_PP__1157  (.L_HI(net1157));
 sg13g2_tiehi \cpu.dcache.r_data[0][25]$_DFFE_PP__1158  (.L_HI(net1158));
 sg13g2_tiehi \cpu.dcache.r_data[0][26]$_DFFE_PP__1159  (.L_HI(net1159));
 sg13g2_tiehi \cpu.dcache.r_data[0][27]$_DFFE_PP__1160  (.L_HI(net1160));
 sg13g2_tiehi \cpu.dcache.r_data[0][28]$_DFFE_PP__1161  (.L_HI(net1161));
 sg13g2_tiehi \cpu.dcache.r_data[0][29]$_DFFE_PP__1162  (.L_HI(net1162));
 sg13g2_tiehi \cpu.dcache.r_data[0][2]$_DFFE_PP__1163  (.L_HI(net1163));
 sg13g2_tiehi \cpu.dcache.r_data[0][30]$_DFFE_PP__1164  (.L_HI(net1164));
 sg13g2_tiehi \cpu.dcache.r_data[0][31]$_DFFE_PP__1165  (.L_HI(net1165));
 sg13g2_tiehi \cpu.dcache.r_data[0][3]$_DFFE_PP__1166  (.L_HI(net1166));
 sg13g2_tiehi \cpu.dcache.r_data[0][4]$_DFFE_PP__1167  (.L_HI(net1167));
 sg13g2_tiehi \cpu.dcache.r_data[0][5]$_DFFE_PP__1168  (.L_HI(net1168));
 sg13g2_tiehi \cpu.dcache.r_data[0][6]$_DFFE_PP__1169  (.L_HI(net1169));
 sg13g2_tiehi \cpu.dcache.r_data[0][7]$_DFFE_PP__1170  (.L_HI(net1170));
 sg13g2_tiehi \cpu.dcache.r_data[0][8]$_DFFE_PP__1171  (.L_HI(net1171));
 sg13g2_tiehi \cpu.dcache.r_data[0][9]$_DFFE_PP__1172  (.L_HI(net1172));
 sg13g2_tiehi \cpu.dcache.r_data[1][0]$_DFFE_PP__1173  (.L_HI(net1173));
 sg13g2_tiehi \cpu.dcache.r_data[1][10]$_DFFE_PP__1174  (.L_HI(net1174));
 sg13g2_tiehi \cpu.dcache.r_data[1][11]$_DFFE_PP__1175  (.L_HI(net1175));
 sg13g2_tiehi \cpu.dcache.r_data[1][12]$_DFFE_PP__1176  (.L_HI(net1176));
 sg13g2_tiehi \cpu.dcache.r_data[1][13]$_DFFE_PP__1177  (.L_HI(net1177));
 sg13g2_tiehi \cpu.dcache.r_data[1][14]$_DFFE_PP__1178  (.L_HI(net1178));
 sg13g2_tiehi \cpu.dcache.r_data[1][15]$_DFFE_PP__1179  (.L_HI(net1179));
 sg13g2_tiehi \cpu.dcache.r_data[1][16]$_DFFE_PP__1180  (.L_HI(net1180));
 sg13g2_tiehi \cpu.dcache.r_data[1][17]$_DFFE_PP__1181  (.L_HI(net1181));
 sg13g2_tiehi \cpu.dcache.r_data[1][18]$_DFFE_PP__1182  (.L_HI(net1182));
 sg13g2_tiehi \cpu.dcache.r_data[1][19]$_DFFE_PP__1183  (.L_HI(net1183));
 sg13g2_tiehi \cpu.dcache.r_data[1][1]$_DFFE_PP__1184  (.L_HI(net1184));
 sg13g2_tiehi \cpu.dcache.r_data[1][20]$_DFFE_PP__1185  (.L_HI(net1185));
 sg13g2_tiehi \cpu.dcache.r_data[1][21]$_DFFE_PP__1186  (.L_HI(net1186));
 sg13g2_tiehi \cpu.dcache.r_data[1][22]$_DFFE_PP__1187  (.L_HI(net1187));
 sg13g2_tiehi \cpu.dcache.r_data[1][23]$_DFFE_PP__1188  (.L_HI(net1188));
 sg13g2_tiehi \cpu.dcache.r_data[1][24]$_DFFE_PP__1189  (.L_HI(net1189));
 sg13g2_tiehi \cpu.dcache.r_data[1][25]$_DFFE_PP__1190  (.L_HI(net1190));
 sg13g2_tiehi \cpu.dcache.r_data[1][26]$_DFFE_PP__1191  (.L_HI(net1191));
 sg13g2_tiehi \cpu.dcache.r_data[1][27]$_DFFE_PP__1192  (.L_HI(net1192));
 sg13g2_tiehi \cpu.dcache.r_data[1][28]$_DFFE_PP__1193  (.L_HI(net1193));
 sg13g2_tiehi \cpu.dcache.r_data[1][29]$_DFFE_PP__1194  (.L_HI(net1194));
 sg13g2_tiehi \cpu.dcache.r_data[1][2]$_DFFE_PP__1195  (.L_HI(net1195));
 sg13g2_tiehi \cpu.dcache.r_data[1][30]$_DFFE_PP__1196  (.L_HI(net1196));
 sg13g2_tiehi \cpu.dcache.r_data[1][31]$_DFFE_PP__1197  (.L_HI(net1197));
 sg13g2_tiehi \cpu.dcache.r_data[1][3]$_DFFE_PP__1198  (.L_HI(net1198));
 sg13g2_tiehi \cpu.dcache.r_data[1][4]$_DFFE_PP__1199  (.L_HI(net1199));
 sg13g2_tiehi \cpu.dcache.r_data[1][5]$_DFFE_PP__1200  (.L_HI(net1200));
 sg13g2_tiehi \cpu.dcache.r_data[1][6]$_DFFE_PP__1201  (.L_HI(net1201));
 sg13g2_tiehi \cpu.dcache.r_data[1][7]$_DFFE_PP__1202  (.L_HI(net1202));
 sg13g2_tiehi \cpu.dcache.r_data[1][8]$_DFFE_PP__1203  (.L_HI(net1203));
 sg13g2_tiehi \cpu.dcache.r_data[1][9]$_DFFE_PP__1204  (.L_HI(net1204));
 sg13g2_tiehi \cpu.dcache.r_data[2][0]$_DFFE_PP__1205  (.L_HI(net1205));
 sg13g2_tiehi \cpu.dcache.r_data[2][10]$_DFFE_PP__1206  (.L_HI(net1206));
 sg13g2_tiehi \cpu.dcache.r_data[2][11]$_DFFE_PP__1207  (.L_HI(net1207));
 sg13g2_tiehi \cpu.dcache.r_data[2][12]$_DFFE_PP__1208  (.L_HI(net1208));
 sg13g2_tiehi \cpu.dcache.r_data[2][13]$_DFFE_PP__1209  (.L_HI(net1209));
 sg13g2_tiehi \cpu.dcache.r_data[2][14]$_DFFE_PP__1210  (.L_HI(net1210));
 sg13g2_tiehi \cpu.dcache.r_data[2][15]$_DFFE_PP__1211  (.L_HI(net1211));
 sg13g2_tiehi \cpu.dcache.r_data[2][16]$_DFFE_PP__1212  (.L_HI(net1212));
 sg13g2_tiehi \cpu.dcache.r_data[2][17]$_DFFE_PP__1213  (.L_HI(net1213));
 sg13g2_tiehi \cpu.dcache.r_data[2][18]$_DFFE_PP__1214  (.L_HI(net1214));
 sg13g2_tiehi \cpu.dcache.r_data[2][19]$_DFFE_PP__1215  (.L_HI(net1215));
 sg13g2_tiehi \cpu.dcache.r_data[2][1]$_DFFE_PP__1216  (.L_HI(net1216));
 sg13g2_tiehi \cpu.dcache.r_data[2][20]$_DFFE_PP__1217  (.L_HI(net1217));
 sg13g2_tiehi \cpu.dcache.r_data[2][21]$_DFFE_PP__1218  (.L_HI(net1218));
 sg13g2_tiehi \cpu.dcache.r_data[2][22]$_DFFE_PP__1219  (.L_HI(net1219));
 sg13g2_tiehi \cpu.dcache.r_data[2][23]$_DFFE_PP__1220  (.L_HI(net1220));
 sg13g2_tiehi \cpu.dcache.r_data[2][24]$_DFFE_PP__1221  (.L_HI(net1221));
 sg13g2_tiehi \cpu.dcache.r_data[2][25]$_DFFE_PP__1222  (.L_HI(net1222));
 sg13g2_tiehi \cpu.dcache.r_data[2][26]$_DFFE_PP__1223  (.L_HI(net1223));
 sg13g2_tiehi \cpu.dcache.r_data[2][27]$_DFFE_PP__1224  (.L_HI(net1224));
 sg13g2_tiehi \cpu.dcache.r_data[2][28]$_DFFE_PP__1225  (.L_HI(net1225));
 sg13g2_tiehi \cpu.dcache.r_data[2][29]$_DFFE_PP__1226  (.L_HI(net1226));
 sg13g2_tiehi \cpu.dcache.r_data[2][2]$_DFFE_PP__1227  (.L_HI(net1227));
 sg13g2_tiehi \cpu.dcache.r_data[2][30]$_DFFE_PP__1228  (.L_HI(net1228));
 sg13g2_tiehi \cpu.dcache.r_data[2][31]$_DFFE_PP__1229  (.L_HI(net1229));
 sg13g2_tiehi \cpu.dcache.r_data[2][3]$_DFFE_PP__1230  (.L_HI(net1230));
 sg13g2_tiehi \cpu.dcache.r_data[2][4]$_DFFE_PP__1231  (.L_HI(net1231));
 sg13g2_tiehi \cpu.dcache.r_data[2][5]$_DFFE_PP__1232  (.L_HI(net1232));
 sg13g2_tiehi \cpu.dcache.r_data[2][6]$_DFFE_PP__1233  (.L_HI(net1233));
 sg13g2_tiehi \cpu.dcache.r_data[2][7]$_DFFE_PP__1234  (.L_HI(net1234));
 sg13g2_tiehi \cpu.dcache.r_data[2][8]$_DFFE_PP__1235  (.L_HI(net1235));
 sg13g2_tiehi \cpu.dcache.r_data[2][9]$_DFFE_PP__1236  (.L_HI(net1236));
 sg13g2_tiehi \cpu.dcache.r_data[3][0]$_DFFE_PP__1237  (.L_HI(net1237));
 sg13g2_tiehi \cpu.dcache.r_data[3][10]$_DFFE_PP__1238  (.L_HI(net1238));
 sg13g2_tiehi \cpu.dcache.r_data[3][11]$_DFFE_PP__1239  (.L_HI(net1239));
 sg13g2_tiehi \cpu.dcache.r_data[3][12]$_DFFE_PP__1240  (.L_HI(net1240));
 sg13g2_tiehi \cpu.dcache.r_data[3][13]$_DFFE_PP__1241  (.L_HI(net1241));
 sg13g2_tiehi \cpu.dcache.r_data[3][14]$_DFFE_PP__1242  (.L_HI(net1242));
 sg13g2_tiehi \cpu.dcache.r_data[3][15]$_DFFE_PP__1243  (.L_HI(net1243));
 sg13g2_tiehi \cpu.dcache.r_data[3][16]$_DFFE_PP__1244  (.L_HI(net1244));
 sg13g2_tiehi \cpu.dcache.r_data[3][17]$_DFFE_PP__1245  (.L_HI(net1245));
 sg13g2_tiehi \cpu.dcache.r_data[3][18]$_DFFE_PP__1246  (.L_HI(net1246));
 sg13g2_tiehi \cpu.dcache.r_data[3][19]$_DFFE_PP__1247  (.L_HI(net1247));
 sg13g2_tiehi \cpu.dcache.r_data[3][1]$_DFFE_PP__1248  (.L_HI(net1248));
 sg13g2_tiehi \cpu.dcache.r_data[3][20]$_DFFE_PP__1249  (.L_HI(net1249));
 sg13g2_tiehi \cpu.dcache.r_data[3][21]$_DFFE_PP__1250  (.L_HI(net1250));
 sg13g2_tiehi \cpu.dcache.r_data[3][22]$_DFFE_PP__1251  (.L_HI(net1251));
 sg13g2_tiehi \cpu.dcache.r_data[3][23]$_DFFE_PP__1252  (.L_HI(net1252));
 sg13g2_tiehi \cpu.dcache.r_data[3][24]$_DFFE_PP__1253  (.L_HI(net1253));
 sg13g2_tiehi \cpu.dcache.r_data[3][25]$_DFFE_PP__1254  (.L_HI(net1254));
 sg13g2_tiehi \cpu.dcache.r_data[3][26]$_DFFE_PP__1255  (.L_HI(net1255));
 sg13g2_tiehi \cpu.dcache.r_data[3][27]$_DFFE_PP__1256  (.L_HI(net1256));
 sg13g2_tiehi \cpu.dcache.r_data[3][28]$_DFFE_PP__1257  (.L_HI(net1257));
 sg13g2_tiehi \cpu.dcache.r_data[3][29]$_DFFE_PP__1258  (.L_HI(net1258));
 sg13g2_tiehi \cpu.dcache.r_data[3][2]$_DFFE_PP__1259  (.L_HI(net1259));
 sg13g2_tiehi \cpu.dcache.r_data[3][30]$_DFFE_PP__1260  (.L_HI(net1260));
 sg13g2_tiehi \cpu.dcache.r_data[3][31]$_DFFE_PP__1261  (.L_HI(net1261));
 sg13g2_tiehi \cpu.dcache.r_data[3][3]$_DFFE_PP__1262  (.L_HI(net1262));
 sg13g2_tiehi \cpu.dcache.r_data[3][4]$_DFFE_PP__1263  (.L_HI(net1263));
 sg13g2_tiehi \cpu.dcache.r_data[3][5]$_DFFE_PP__1264  (.L_HI(net1264));
 sg13g2_tiehi \cpu.dcache.r_data[3][6]$_DFFE_PP__1265  (.L_HI(net1265));
 sg13g2_tiehi \cpu.dcache.r_data[3][7]$_DFFE_PP__1266  (.L_HI(net1266));
 sg13g2_tiehi \cpu.dcache.r_data[3][8]$_DFFE_PP__1267  (.L_HI(net1267));
 sg13g2_tiehi \cpu.dcache.r_data[3][9]$_DFFE_PP__1268  (.L_HI(net1268));
 sg13g2_tiehi \cpu.dcache.r_data[4][0]$_DFFE_PP__1269  (.L_HI(net1269));
 sg13g2_tiehi \cpu.dcache.r_data[4][10]$_DFFE_PP__1270  (.L_HI(net1270));
 sg13g2_tiehi \cpu.dcache.r_data[4][11]$_DFFE_PP__1271  (.L_HI(net1271));
 sg13g2_tiehi \cpu.dcache.r_data[4][12]$_DFFE_PP__1272  (.L_HI(net1272));
 sg13g2_tiehi \cpu.dcache.r_data[4][13]$_DFFE_PP__1273  (.L_HI(net1273));
 sg13g2_tiehi \cpu.dcache.r_data[4][14]$_DFFE_PP__1274  (.L_HI(net1274));
 sg13g2_tiehi \cpu.dcache.r_data[4][15]$_DFFE_PP__1275  (.L_HI(net1275));
 sg13g2_tiehi \cpu.dcache.r_data[4][16]$_DFFE_PP__1276  (.L_HI(net1276));
 sg13g2_tiehi \cpu.dcache.r_data[4][17]$_DFFE_PP__1277  (.L_HI(net1277));
 sg13g2_tiehi \cpu.dcache.r_data[4][18]$_DFFE_PP__1278  (.L_HI(net1278));
 sg13g2_tiehi \cpu.dcache.r_data[4][19]$_DFFE_PP__1279  (.L_HI(net1279));
 sg13g2_tiehi \cpu.dcache.r_data[4][1]$_DFFE_PP__1280  (.L_HI(net1280));
 sg13g2_tiehi \cpu.dcache.r_data[4][20]$_DFFE_PP__1281  (.L_HI(net1281));
 sg13g2_tiehi \cpu.dcache.r_data[4][21]$_DFFE_PP__1282  (.L_HI(net1282));
 sg13g2_tiehi \cpu.dcache.r_data[4][22]$_DFFE_PP__1283  (.L_HI(net1283));
 sg13g2_tiehi \cpu.dcache.r_data[4][23]$_DFFE_PP__1284  (.L_HI(net1284));
 sg13g2_tiehi \cpu.dcache.r_data[4][24]$_DFFE_PP__1285  (.L_HI(net1285));
 sg13g2_tiehi \cpu.dcache.r_data[4][25]$_DFFE_PP__1286  (.L_HI(net1286));
 sg13g2_tiehi \cpu.dcache.r_data[4][26]$_DFFE_PP__1287  (.L_HI(net1287));
 sg13g2_tiehi \cpu.dcache.r_data[4][27]$_DFFE_PP__1288  (.L_HI(net1288));
 sg13g2_tiehi \cpu.dcache.r_data[4][28]$_DFFE_PP__1289  (.L_HI(net1289));
 sg13g2_tiehi \cpu.dcache.r_data[4][29]$_DFFE_PP__1290  (.L_HI(net1290));
 sg13g2_tiehi \cpu.dcache.r_data[4][2]$_DFFE_PP__1291  (.L_HI(net1291));
 sg13g2_tiehi \cpu.dcache.r_data[4][30]$_DFFE_PP__1292  (.L_HI(net1292));
 sg13g2_tiehi \cpu.dcache.r_data[4][31]$_DFFE_PP__1293  (.L_HI(net1293));
 sg13g2_tiehi \cpu.dcache.r_data[4][3]$_DFFE_PP__1294  (.L_HI(net1294));
 sg13g2_tiehi \cpu.dcache.r_data[4][4]$_DFFE_PP__1295  (.L_HI(net1295));
 sg13g2_tiehi \cpu.dcache.r_data[4][5]$_DFFE_PP__1296  (.L_HI(net1296));
 sg13g2_tiehi \cpu.dcache.r_data[4][6]$_DFFE_PP__1297  (.L_HI(net1297));
 sg13g2_tiehi \cpu.dcache.r_data[4][7]$_DFFE_PP__1298  (.L_HI(net1298));
 sg13g2_tiehi \cpu.dcache.r_data[4][8]$_DFFE_PP__1299  (.L_HI(net1299));
 sg13g2_tiehi \cpu.dcache.r_data[4][9]$_DFFE_PP__1300  (.L_HI(net1300));
 sg13g2_tiehi \cpu.dcache.r_data[5][0]$_DFFE_PP__1301  (.L_HI(net1301));
 sg13g2_tiehi \cpu.dcache.r_data[5][10]$_DFFE_PP__1302  (.L_HI(net1302));
 sg13g2_tiehi \cpu.dcache.r_data[5][11]$_DFFE_PP__1303  (.L_HI(net1303));
 sg13g2_tiehi \cpu.dcache.r_data[5][12]$_DFFE_PP__1304  (.L_HI(net1304));
 sg13g2_tiehi \cpu.dcache.r_data[5][13]$_DFFE_PP__1305  (.L_HI(net1305));
 sg13g2_tiehi \cpu.dcache.r_data[5][14]$_DFFE_PP__1306  (.L_HI(net1306));
 sg13g2_tiehi \cpu.dcache.r_data[5][15]$_DFFE_PP__1307  (.L_HI(net1307));
 sg13g2_tiehi \cpu.dcache.r_data[5][16]$_DFFE_PP__1308  (.L_HI(net1308));
 sg13g2_tiehi \cpu.dcache.r_data[5][17]$_DFFE_PP__1309  (.L_HI(net1309));
 sg13g2_tiehi \cpu.dcache.r_data[5][18]$_DFFE_PP__1310  (.L_HI(net1310));
 sg13g2_tiehi \cpu.dcache.r_data[5][19]$_DFFE_PP__1311  (.L_HI(net1311));
 sg13g2_tiehi \cpu.dcache.r_data[5][1]$_DFFE_PP__1312  (.L_HI(net1312));
 sg13g2_tiehi \cpu.dcache.r_data[5][20]$_DFFE_PP__1313  (.L_HI(net1313));
 sg13g2_tiehi \cpu.dcache.r_data[5][21]$_DFFE_PP__1314  (.L_HI(net1314));
 sg13g2_tiehi \cpu.dcache.r_data[5][22]$_DFFE_PP__1315  (.L_HI(net1315));
 sg13g2_tiehi \cpu.dcache.r_data[5][23]$_DFFE_PP__1316  (.L_HI(net1316));
 sg13g2_tiehi \cpu.dcache.r_data[5][24]$_DFFE_PP__1317  (.L_HI(net1317));
 sg13g2_tiehi \cpu.dcache.r_data[5][25]$_DFFE_PP__1318  (.L_HI(net1318));
 sg13g2_tiehi \cpu.dcache.r_data[5][26]$_DFFE_PP__1319  (.L_HI(net1319));
 sg13g2_tiehi \cpu.dcache.r_data[5][27]$_DFFE_PP__1320  (.L_HI(net1320));
 sg13g2_tiehi \cpu.dcache.r_data[5][28]$_DFFE_PP__1321  (.L_HI(net1321));
 sg13g2_tiehi \cpu.dcache.r_data[5][29]$_DFFE_PP__1322  (.L_HI(net1322));
 sg13g2_tiehi \cpu.dcache.r_data[5][2]$_DFFE_PP__1323  (.L_HI(net1323));
 sg13g2_tiehi \cpu.dcache.r_data[5][30]$_DFFE_PP__1324  (.L_HI(net1324));
 sg13g2_tiehi \cpu.dcache.r_data[5][31]$_DFFE_PP__1325  (.L_HI(net1325));
 sg13g2_tiehi \cpu.dcache.r_data[5][3]$_DFFE_PP__1326  (.L_HI(net1326));
 sg13g2_tiehi \cpu.dcache.r_data[5][4]$_DFFE_PP__1327  (.L_HI(net1327));
 sg13g2_tiehi \cpu.dcache.r_data[5][5]$_DFFE_PP__1328  (.L_HI(net1328));
 sg13g2_tiehi \cpu.dcache.r_data[5][6]$_DFFE_PP__1329  (.L_HI(net1329));
 sg13g2_tiehi \cpu.dcache.r_data[5][7]$_DFFE_PP__1330  (.L_HI(net1330));
 sg13g2_tiehi \cpu.dcache.r_data[5][8]$_DFFE_PP__1331  (.L_HI(net1331));
 sg13g2_tiehi \cpu.dcache.r_data[5][9]$_DFFE_PP__1332  (.L_HI(net1332));
 sg13g2_tiehi \cpu.dcache.r_data[6][0]$_DFFE_PP__1333  (.L_HI(net1333));
 sg13g2_tiehi \cpu.dcache.r_data[6][10]$_DFFE_PP__1334  (.L_HI(net1334));
 sg13g2_tiehi \cpu.dcache.r_data[6][11]$_DFFE_PP__1335  (.L_HI(net1335));
 sg13g2_tiehi \cpu.dcache.r_data[6][12]$_DFFE_PP__1336  (.L_HI(net1336));
 sg13g2_tiehi \cpu.dcache.r_data[6][13]$_DFFE_PP__1337  (.L_HI(net1337));
 sg13g2_tiehi \cpu.dcache.r_data[6][14]$_DFFE_PP__1338  (.L_HI(net1338));
 sg13g2_tiehi \cpu.dcache.r_data[6][15]$_DFFE_PP__1339  (.L_HI(net1339));
 sg13g2_tiehi \cpu.dcache.r_data[6][16]$_DFFE_PP__1340  (.L_HI(net1340));
 sg13g2_tiehi \cpu.dcache.r_data[6][17]$_DFFE_PP__1341  (.L_HI(net1341));
 sg13g2_tiehi \cpu.dcache.r_data[6][18]$_DFFE_PP__1342  (.L_HI(net1342));
 sg13g2_tiehi \cpu.dcache.r_data[6][19]$_DFFE_PP__1343  (.L_HI(net1343));
 sg13g2_tiehi \cpu.dcache.r_data[6][1]$_DFFE_PP__1344  (.L_HI(net1344));
 sg13g2_tiehi \cpu.dcache.r_data[6][20]$_DFFE_PP__1345  (.L_HI(net1345));
 sg13g2_tiehi \cpu.dcache.r_data[6][21]$_DFFE_PP__1346  (.L_HI(net1346));
 sg13g2_tiehi \cpu.dcache.r_data[6][22]$_DFFE_PP__1347  (.L_HI(net1347));
 sg13g2_tiehi \cpu.dcache.r_data[6][23]$_DFFE_PP__1348  (.L_HI(net1348));
 sg13g2_tiehi \cpu.dcache.r_data[6][24]$_DFFE_PP__1349  (.L_HI(net1349));
 sg13g2_tiehi \cpu.dcache.r_data[6][25]$_DFFE_PP__1350  (.L_HI(net1350));
 sg13g2_tiehi \cpu.dcache.r_data[6][26]$_DFFE_PP__1351  (.L_HI(net1351));
 sg13g2_tiehi \cpu.dcache.r_data[6][27]$_DFFE_PP__1352  (.L_HI(net1352));
 sg13g2_tiehi \cpu.dcache.r_data[6][28]$_DFFE_PP__1353  (.L_HI(net1353));
 sg13g2_tiehi \cpu.dcache.r_data[6][29]$_DFFE_PP__1354  (.L_HI(net1354));
 sg13g2_tiehi \cpu.dcache.r_data[6][2]$_DFFE_PP__1355  (.L_HI(net1355));
 sg13g2_tiehi \cpu.dcache.r_data[6][30]$_DFFE_PP__1356  (.L_HI(net1356));
 sg13g2_tiehi \cpu.dcache.r_data[6][31]$_DFFE_PP__1357  (.L_HI(net1357));
 sg13g2_tiehi \cpu.dcache.r_data[6][3]$_DFFE_PP__1358  (.L_HI(net1358));
 sg13g2_tiehi \cpu.dcache.r_data[6][4]$_DFFE_PP__1359  (.L_HI(net1359));
 sg13g2_tiehi \cpu.dcache.r_data[6][5]$_DFFE_PP__1360  (.L_HI(net1360));
 sg13g2_tiehi \cpu.dcache.r_data[6][6]$_DFFE_PP__1361  (.L_HI(net1361));
 sg13g2_tiehi \cpu.dcache.r_data[6][7]$_DFFE_PP__1362  (.L_HI(net1362));
 sg13g2_tiehi \cpu.dcache.r_data[6][8]$_DFFE_PP__1363  (.L_HI(net1363));
 sg13g2_tiehi \cpu.dcache.r_data[6][9]$_DFFE_PP__1364  (.L_HI(net1364));
 sg13g2_tiehi \cpu.dcache.r_data[7][0]$_DFFE_PP__1365  (.L_HI(net1365));
 sg13g2_tiehi \cpu.dcache.r_data[7][10]$_DFFE_PP__1366  (.L_HI(net1366));
 sg13g2_tiehi \cpu.dcache.r_data[7][11]$_DFFE_PP__1367  (.L_HI(net1367));
 sg13g2_tiehi \cpu.dcache.r_data[7][12]$_DFFE_PP__1368  (.L_HI(net1368));
 sg13g2_tiehi \cpu.dcache.r_data[7][13]$_DFFE_PP__1369  (.L_HI(net1369));
 sg13g2_tiehi \cpu.dcache.r_data[7][14]$_DFFE_PP__1370  (.L_HI(net1370));
 sg13g2_tiehi \cpu.dcache.r_data[7][15]$_DFFE_PP__1371  (.L_HI(net1371));
 sg13g2_tiehi \cpu.dcache.r_data[7][16]$_DFFE_PP__1372  (.L_HI(net1372));
 sg13g2_tiehi \cpu.dcache.r_data[7][17]$_DFFE_PP__1373  (.L_HI(net1373));
 sg13g2_tiehi \cpu.dcache.r_data[7][18]$_DFFE_PP__1374  (.L_HI(net1374));
 sg13g2_tiehi \cpu.dcache.r_data[7][19]$_DFFE_PP__1375  (.L_HI(net1375));
 sg13g2_tiehi \cpu.dcache.r_data[7][1]$_DFFE_PP__1376  (.L_HI(net1376));
 sg13g2_tiehi \cpu.dcache.r_data[7][20]$_DFFE_PP__1377  (.L_HI(net1377));
 sg13g2_tiehi \cpu.dcache.r_data[7][21]$_DFFE_PP__1378  (.L_HI(net1378));
 sg13g2_tiehi \cpu.dcache.r_data[7][22]$_DFFE_PP__1379  (.L_HI(net1379));
 sg13g2_tiehi \cpu.dcache.r_data[7][23]$_DFFE_PP__1380  (.L_HI(net1380));
 sg13g2_tiehi \cpu.dcache.r_data[7][24]$_DFFE_PP__1381  (.L_HI(net1381));
 sg13g2_tiehi \cpu.dcache.r_data[7][25]$_DFFE_PP__1382  (.L_HI(net1382));
 sg13g2_tiehi \cpu.dcache.r_data[7][26]$_DFFE_PP__1383  (.L_HI(net1383));
 sg13g2_tiehi \cpu.dcache.r_data[7][27]$_DFFE_PP__1384  (.L_HI(net1384));
 sg13g2_tiehi \cpu.dcache.r_data[7][28]$_DFFE_PP__1385  (.L_HI(net1385));
 sg13g2_tiehi \cpu.dcache.r_data[7][29]$_DFFE_PP__1386  (.L_HI(net1386));
 sg13g2_tiehi \cpu.dcache.r_data[7][2]$_DFFE_PP__1387  (.L_HI(net1387));
 sg13g2_tiehi \cpu.dcache.r_data[7][30]$_DFFE_PP__1388  (.L_HI(net1388));
 sg13g2_tiehi \cpu.dcache.r_data[7][31]$_DFFE_PP__1389  (.L_HI(net1389));
 sg13g2_tiehi \cpu.dcache.r_data[7][3]$_DFFE_PP__1390  (.L_HI(net1390));
 sg13g2_tiehi \cpu.dcache.r_data[7][4]$_DFFE_PP__1391  (.L_HI(net1391));
 sg13g2_tiehi \cpu.dcache.r_data[7][5]$_DFFE_PP__1392  (.L_HI(net1392));
 sg13g2_tiehi \cpu.dcache.r_data[7][6]$_DFFE_PP__1393  (.L_HI(net1393));
 sg13g2_tiehi \cpu.dcache.r_data[7][7]$_DFFE_PP__1394  (.L_HI(net1394));
 sg13g2_tiehi \cpu.dcache.r_data[7][8]$_DFFE_PP__1395  (.L_HI(net1395));
 sg13g2_tiehi \cpu.dcache.r_data[7][9]$_DFFE_PP__1396  (.L_HI(net1396));
 sg13g2_tiehi \cpu.dcache.r_dirty[0]$_SDFFCE_PP1P__1397  (.L_HI(net1397));
 sg13g2_tiehi \cpu.dcache.r_dirty[1]$_SDFFCE_PP1P__1398  (.L_HI(net1398));
 sg13g2_tiehi \cpu.dcache.r_dirty[2]$_SDFFCE_PP1P__1399  (.L_HI(net1399));
 sg13g2_tiehi \cpu.dcache.r_dirty[3]$_SDFFCE_PP1P__1400  (.L_HI(net1400));
 sg13g2_tiehi \cpu.dcache.r_dirty[4]$_SDFFCE_PP1P__1401  (.L_HI(net1401));
 sg13g2_tiehi \cpu.dcache.r_dirty[5]$_SDFFCE_PP1P__1402  (.L_HI(net1402));
 sg13g2_tiehi \cpu.dcache.r_dirty[6]$_SDFFCE_PP1P__1403  (.L_HI(net1403));
 sg13g2_tiehi \cpu.dcache.r_dirty[7]$_SDFFCE_PP1P__1404  (.L_HI(net1404));
 sg13g2_tiehi \cpu.dcache.r_offset[0]$_SDFF_PN0__1405  (.L_HI(net1405));
 sg13g2_tiehi \cpu.dcache.r_offset[1]$_SDFF_PN0__1406  (.L_HI(net1406));
 sg13g2_tiehi \cpu.dcache.r_offset[2]$_SDFF_PN0__1407  (.L_HI(net1407));
 sg13g2_tiehi \cpu.dcache.r_tag[0][0]$_DFFE_PP__1408  (.L_HI(net1408));
 sg13g2_tiehi \cpu.dcache.r_tag[0][10]$_DFFE_PP__1409  (.L_HI(net1409));
 sg13g2_tiehi \cpu.dcache.r_tag[0][11]$_DFFE_PP__1410  (.L_HI(net1410));
 sg13g2_tiehi \cpu.dcache.r_tag[0][12]$_DFFE_PP__1411  (.L_HI(net1411));
 sg13g2_tiehi \cpu.dcache.r_tag[0][13]$_DFFE_PP__1412  (.L_HI(net1412));
 sg13g2_tiehi \cpu.dcache.r_tag[0][14]$_DFFE_PP__1413  (.L_HI(net1413));
 sg13g2_tiehi \cpu.dcache.r_tag[0][15]$_DFFE_PP__1414  (.L_HI(net1414));
 sg13g2_tiehi \cpu.dcache.r_tag[0][16]$_DFFE_PP__1415  (.L_HI(net1415));
 sg13g2_tiehi \cpu.dcache.r_tag[0][17]$_DFFE_PP__1416  (.L_HI(net1416));
 sg13g2_tiehi \cpu.dcache.r_tag[0][18]$_DFFE_PP__1417  (.L_HI(net1417));
 sg13g2_tiehi \cpu.dcache.r_tag[0][1]$_DFFE_PP__1418  (.L_HI(net1418));
 sg13g2_tiehi \cpu.dcache.r_tag[0][2]$_DFFE_PP__1419  (.L_HI(net1419));
 sg13g2_tiehi \cpu.dcache.r_tag[0][3]$_DFFE_PP__1420  (.L_HI(net1420));
 sg13g2_tiehi \cpu.dcache.r_tag[0][4]$_DFFE_PP__1421  (.L_HI(net1421));
 sg13g2_tiehi \cpu.dcache.r_tag[0][5]$_DFFE_PP__1422  (.L_HI(net1422));
 sg13g2_tiehi \cpu.dcache.r_tag[0][6]$_DFFE_PP__1423  (.L_HI(net1423));
 sg13g2_tiehi \cpu.dcache.r_tag[0][7]$_DFFE_PP__1424  (.L_HI(net1424));
 sg13g2_tiehi \cpu.dcache.r_tag[0][8]$_DFFE_PP__1425  (.L_HI(net1425));
 sg13g2_tiehi \cpu.dcache.r_tag[0][9]$_DFFE_PP__1426  (.L_HI(net1426));
 sg13g2_tiehi \cpu.dcache.r_tag[1][0]$_DFFE_PP__1427  (.L_HI(net1427));
 sg13g2_tiehi \cpu.dcache.r_tag[1][10]$_DFFE_PP__1428  (.L_HI(net1428));
 sg13g2_tiehi \cpu.dcache.r_tag[1][11]$_DFFE_PP__1429  (.L_HI(net1429));
 sg13g2_tiehi \cpu.dcache.r_tag[1][12]$_DFFE_PP__1430  (.L_HI(net1430));
 sg13g2_tiehi \cpu.dcache.r_tag[1][13]$_DFFE_PP__1431  (.L_HI(net1431));
 sg13g2_tiehi \cpu.dcache.r_tag[1][14]$_DFFE_PP__1432  (.L_HI(net1432));
 sg13g2_tiehi \cpu.dcache.r_tag[1][15]$_DFFE_PP__1433  (.L_HI(net1433));
 sg13g2_tiehi \cpu.dcache.r_tag[1][16]$_DFFE_PP__1434  (.L_HI(net1434));
 sg13g2_tiehi \cpu.dcache.r_tag[1][17]$_DFFE_PP__1435  (.L_HI(net1435));
 sg13g2_tiehi \cpu.dcache.r_tag[1][18]$_DFFE_PP__1436  (.L_HI(net1436));
 sg13g2_tiehi \cpu.dcache.r_tag[1][1]$_DFFE_PP__1437  (.L_HI(net1437));
 sg13g2_tiehi \cpu.dcache.r_tag[1][2]$_DFFE_PP__1438  (.L_HI(net1438));
 sg13g2_tiehi \cpu.dcache.r_tag[1][3]$_DFFE_PP__1439  (.L_HI(net1439));
 sg13g2_tiehi \cpu.dcache.r_tag[1][4]$_DFFE_PP__1440  (.L_HI(net1440));
 sg13g2_tiehi \cpu.dcache.r_tag[1][5]$_DFFE_PP__1441  (.L_HI(net1441));
 sg13g2_tiehi \cpu.dcache.r_tag[1][6]$_DFFE_PP__1442  (.L_HI(net1442));
 sg13g2_tiehi \cpu.dcache.r_tag[1][7]$_DFFE_PP__1443  (.L_HI(net1443));
 sg13g2_tiehi \cpu.dcache.r_tag[1][8]$_DFFE_PP__1444  (.L_HI(net1444));
 sg13g2_tiehi \cpu.dcache.r_tag[1][9]$_DFFE_PP__1445  (.L_HI(net1445));
 sg13g2_tiehi \cpu.dcache.r_tag[2][0]$_DFFE_PP__1446  (.L_HI(net1446));
 sg13g2_tiehi \cpu.dcache.r_tag[2][10]$_DFFE_PP__1447  (.L_HI(net1447));
 sg13g2_tiehi \cpu.dcache.r_tag[2][11]$_DFFE_PP__1448  (.L_HI(net1448));
 sg13g2_tiehi \cpu.dcache.r_tag[2][12]$_DFFE_PP__1449  (.L_HI(net1449));
 sg13g2_tiehi \cpu.dcache.r_tag[2][13]$_DFFE_PP__1450  (.L_HI(net1450));
 sg13g2_tiehi \cpu.dcache.r_tag[2][14]$_DFFE_PP__1451  (.L_HI(net1451));
 sg13g2_tiehi \cpu.dcache.r_tag[2][15]$_DFFE_PP__1452  (.L_HI(net1452));
 sg13g2_tiehi \cpu.dcache.r_tag[2][16]$_DFFE_PP__1453  (.L_HI(net1453));
 sg13g2_tiehi \cpu.dcache.r_tag[2][17]$_DFFE_PP__1454  (.L_HI(net1454));
 sg13g2_tiehi \cpu.dcache.r_tag[2][18]$_DFFE_PP__1455  (.L_HI(net1455));
 sg13g2_tiehi \cpu.dcache.r_tag[2][1]$_DFFE_PP__1456  (.L_HI(net1456));
 sg13g2_tiehi \cpu.dcache.r_tag[2][2]$_DFFE_PP__1457  (.L_HI(net1457));
 sg13g2_tiehi \cpu.dcache.r_tag[2][3]$_DFFE_PP__1458  (.L_HI(net1458));
 sg13g2_tiehi \cpu.dcache.r_tag[2][4]$_DFFE_PP__1459  (.L_HI(net1459));
 sg13g2_tiehi \cpu.dcache.r_tag[2][5]$_DFFE_PP__1460  (.L_HI(net1460));
 sg13g2_tiehi \cpu.dcache.r_tag[2][6]$_DFFE_PP__1461  (.L_HI(net1461));
 sg13g2_tiehi \cpu.dcache.r_tag[2][7]$_DFFE_PP__1462  (.L_HI(net1462));
 sg13g2_tiehi \cpu.dcache.r_tag[2][8]$_DFFE_PP__1463  (.L_HI(net1463));
 sg13g2_tiehi \cpu.dcache.r_tag[2][9]$_DFFE_PP__1464  (.L_HI(net1464));
 sg13g2_tiehi \cpu.dcache.r_tag[3][0]$_DFFE_PP__1465  (.L_HI(net1465));
 sg13g2_tiehi \cpu.dcache.r_tag[3][10]$_DFFE_PP__1466  (.L_HI(net1466));
 sg13g2_tiehi \cpu.dcache.r_tag[3][11]$_DFFE_PP__1467  (.L_HI(net1467));
 sg13g2_tiehi \cpu.dcache.r_tag[3][12]$_DFFE_PP__1468  (.L_HI(net1468));
 sg13g2_tiehi \cpu.dcache.r_tag[3][13]$_DFFE_PP__1469  (.L_HI(net1469));
 sg13g2_tiehi \cpu.dcache.r_tag[3][14]$_DFFE_PP__1470  (.L_HI(net1470));
 sg13g2_tiehi \cpu.dcache.r_tag[3][15]$_DFFE_PP__1471  (.L_HI(net1471));
 sg13g2_tiehi \cpu.dcache.r_tag[3][16]$_DFFE_PP__1472  (.L_HI(net1472));
 sg13g2_tiehi \cpu.dcache.r_tag[3][17]$_DFFE_PP__1473  (.L_HI(net1473));
 sg13g2_tiehi \cpu.dcache.r_tag[3][18]$_DFFE_PP__1474  (.L_HI(net1474));
 sg13g2_tiehi \cpu.dcache.r_tag[3][1]$_DFFE_PP__1475  (.L_HI(net1475));
 sg13g2_tiehi \cpu.dcache.r_tag[3][2]$_DFFE_PP__1476  (.L_HI(net1476));
 sg13g2_tiehi \cpu.dcache.r_tag[3][3]$_DFFE_PP__1477  (.L_HI(net1477));
 sg13g2_tiehi \cpu.dcache.r_tag[3][4]$_DFFE_PP__1478  (.L_HI(net1478));
 sg13g2_tiehi \cpu.dcache.r_tag[3][5]$_DFFE_PP__1479  (.L_HI(net1479));
 sg13g2_tiehi \cpu.dcache.r_tag[3][6]$_DFFE_PP__1480  (.L_HI(net1480));
 sg13g2_tiehi \cpu.dcache.r_tag[3][7]$_DFFE_PP__1481  (.L_HI(net1481));
 sg13g2_tiehi \cpu.dcache.r_tag[3][8]$_DFFE_PP__1482  (.L_HI(net1482));
 sg13g2_tiehi \cpu.dcache.r_tag[3][9]$_DFFE_PP__1483  (.L_HI(net1483));
 sg13g2_tiehi \cpu.dcache.r_tag[4][0]$_DFFE_PP__1484  (.L_HI(net1484));
 sg13g2_tiehi \cpu.dcache.r_tag[4][10]$_DFFE_PP__1485  (.L_HI(net1485));
 sg13g2_tiehi \cpu.dcache.r_tag[4][11]$_DFFE_PP__1486  (.L_HI(net1486));
 sg13g2_tiehi \cpu.dcache.r_tag[4][12]$_DFFE_PP__1487  (.L_HI(net1487));
 sg13g2_tiehi \cpu.dcache.r_tag[4][13]$_DFFE_PP__1488  (.L_HI(net1488));
 sg13g2_tiehi \cpu.dcache.r_tag[4][14]$_DFFE_PP__1489  (.L_HI(net1489));
 sg13g2_tiehi \cpu.dcache.r_tag[4][15]$_DFFE_PP__1490  (.L_HI(net1490));
 sg13g2_tiehi \cpu.dcache.r_tag[4][16]$_DFFE_PP__1491  (.L_HI(net1491));
 sg13g2_tiehi \cpu.dcache.r_tag[4][17]$_DFFE_PP__1492  (.L_HI(net1492));
 sg13g2_tiehi \cpu.dcache.r_tag[4][18]$_DFFE_PP__1493  (.L_HI(net1493));
 sg13g2_tiehi \cpu.dcache.r_tag[4][1]$_DFFE_PP__1494  (.L_HI(net1494));
 sg13g2_tiehi \cpu.dcache.r_tag[4][2]$_DFFE_PP__1495  (.L_HI(net1495));
 sg13g2_tiehi \cpu.dcache.r_tag[4][3]$_DFFE_PP__1496  (.L_HI(net1496));
 sg13g2_tiehi \cpu.dcache.r_tag[4][4]$_DFFE_PP__1497  (.L_HI(net1497));
 sg13g2_tiehi \cpu.dcache.r_tag[4][5]$_DFFE_PP__1498  (.L_HI(net1498));
 sg13g2_tiehi \cpu.dcache.r_tag[4][6]$_DFFE_PP__1499  (.L_HI(net1499));
 sg13g2_tiehi \cpu.dcache.r_tag[4][7]$_DFFE_PP__1500  (.L_HI(net1500));
 sg13g2_tiehi \cpu.dcache.r_tag[4][8]$_DFFE_PP__1501  (.L_HI(net1501));
 sg13g2_tiehi \cpu.dcache.r_tag[4][9]$_DFFE_PP__1502  (.L_HI(net1502));
 sg13g2_tiehi \cpu.dcache.r_tag[5][0]$_DFFE_PP__1503  (.L_HI(net1503));
 sg13g2_tiehi \cpu.dcache.r_tag[5][10]$_DFFE_PP__1504  (.L_HI(net1504));
 sg13g2_tiehi \cpu.dcache.r_tag[5][11]$_DFFE_PP__1505  (.L_HI(net1505));
 sg13g2_tiehi \cpu.dcache.r_tag[5][12]$_DFFE_PP__1506  (.L_HI(net1506));
 sg13g2_tiehi \cpu.dcache.r_tag[5][13]$_DFFE_PP__1507  (.L_HI(net1507));
 sg13g2_tiehi \cpu.dcache.r_tag[5][14]$_DFFE_PP__1508  (.L_HI(net1508));
 sg13g2_tiehi \cpu.dcache.r_tag[5][15]$_DFFE_PP__1509  (.L_HI(net1509));
 sg13g2_tiehi \cpu.dcache.r_tag[5][16]$_DFFE_PP__1510  (.L_HI(net1510));
 sg13g2_tiehi \cpu.dcache.r_tag[5][17]$_DFFE_PP__1511  (.L_HI(net1511));
 sg13g2_tiehi \cpu.dcache.r_tag[5][18]$_DFFE_PP__1512  (.L_HI(net1512));
 sg13g2_tiehi \cpu.dcache.r_tag[5][1]$_DFFE_PP__1513  (.L_HI(net1513));
 sg13g2_tiehi \cpu.dcache.r_tag[5][2]$_DFFE_PP__1514  (.L_HI(net1514));
 sg13g2_tiehi \cpu.dcache.r_tag[5][3]$_DFFE_PP__1515  (.L_HI(net1515));
 sg13g2_tiehi \cpu.dcache.r_tag[5][4]$_DFFE_PP__1516  (.L_HI(net1516));
 sg13g2_tiehi \cpu.dcache.r_tag[5][5]$_DFFE_PP__1517  (.L_HI(net1517));
 sg13g2_tiehi \cpu.dcache.r_tag[5][6]$_DFFE_PP__1518  (.L_HI(net1518));
 sg13g2_tiehi \cpu.dcache.r_tag[5][7]$_DFFE_PP__1519  (.L_HI(net1519));
 sg13g2_tiehi \cpu.dcache.r_tag[5][8]$_DFFE_PP__1520  (.L_HI(net1520));
 sg13g2_tiehi \cpu.dcache.r_tag[5][9]$_DFFE_PP__1521  (.L_HI(net1521));
 sg13g2_tiehi \cpu.dcache.r_tag[6][0]$_DFFE_PP__1522  (.L_HI(net1522));
 sg13g2_tiehi \cpu.dcache.r_tag[6][10]$_DFFE_PP__1523  (.L_HI(net1523));
 sg13g2_tiehi \cpu.dcache.r_tag[6][11]$_DFFE_PP__1524  (.L_HI(net1524));
 sg13g2_tiehi \cpu.dcache.r_tag[6][12]$_DFFE_PP__1525  (.L_HI(net1525));
 sg13g2_tiehi \cpu.dcache.r_tag[6][13]$_DFFE_PP__1526  (.L_HI(net1526));
 sg13g2_tiehi \cpu.dcache.r_tag[6][14]$_DFFE_PP__1527  (.L_HI(net1527));
 sg13g2_tiehi \cpu.dcache.r_tag[6][15]$_DFFE_PP__1528  (.L_HI(net1528));
 sg13g2_tiehi \cpu.dcache.r_tag[6][16]$_DFFE_PP__1529  (.L_HI(net1529));
 sg13g2_tiehi \cpu.dcache.r_tag[6][17]$_DFFE_PP__1530  (.L_HI(net1530));
 sg13g2_tiehi \cpu.dcache.r_tag[6][18]$_DFFE_PP__1531  (.L_HI(net1531));
 sg13g2_tiehi \cpu.dcache.r_tag[6][1]$_DFFE_PP__1532  (.L_HI(net1532));
 sg13g2_tiehi \cpu.dcache.r_tag[6][2]$_DFFE_PP__1533  (.L_HI(net1533));
 sg13g2_tiehi \cpu.dcache.r_tag[6][3]$_DFFE_PP__1534  (.L_HI(net1534));
 sg13g2_tiehi \cpu.dcache.r_tag[6][4]$_DFFE_PP__1535  (.L_HI(net1535));
 sg13g2_tiehi \cpu.dcache.r_tag[6][5]$_DFFE_PP__1536  (.L_HI(net1536));
 sg13g2_tiehi \cpu.dcache.r_tag[6][6]$_DFFE_PP__1537  (.L_HI(net1537));
 sg13g2_tiehi \cpu.dcache.r_tag[6][7]$_DFFE_PP__1538  (.L_HI(net1538));
 sg13g2_tiehi \cpu.dcache.r_tag[6][8]$_DFFE_PP__1539  (.L_HI(net1539));
 sg13g2_tiehi \cpu.dcache.r_tag[6][9]$_DFFE_PP__1540  (.L_HI(net1540));
 sg13g2_tiehi \cpu.dcache.r_tag[7][0]$_DFFE_PP__1541  (.L_HI(net1541));
 sg13g2_tiehi \cpu.dcache.r_tag[7][10]$_DFFE_PP__1542  (.L_HI(net1542));
 sg13g2_tiehi \cpu.dcache.r_tag[7][11]$_DFFE_PP__1543  (.L_HI(net1543));
 sg13g2_tiehi \cpu.dcache.r_tag[7][12]$_DFFE_PP__1544  (.L_HI(net1544));
 sg13g2_tiehi \cpu.dcache.r_tag[7][13]$_DFFE_PP__1545  (.L_HI(net1545));
 sg13g2_tiehi \cpu.dcache.r_tag[7][14]$_DFFE_PP__1546  (.L_HI(net1546));
 sg13g2_tiehi \cpu.dcache.r_tag[7][15]$_DFFE_PP__1547  (.L_HI(net1547));
 sg13g2_tiehi \cpu.dcache.r_tag[7][16]$_DFFE_PP__1548  (.L_HI(net1548));
 sg13g2_tiehi \cpu.dcache.r_tag[7][17]$_DFFE_PP__1549  (.L_HI(net1549));
 sg13g2_tiehi \cpu.dcache.r_tag[7][18]$_DFFE_PP__1550  (.L_HI(net1550));
 sg13g2_tiehi \cpu.dcache.r_tag[7][1]$_DFFE_PP__1551  (.L_HI(net1551));
 sg13g2_tiehi \cpu.dcache.r_tag[7][2]$_DFFE_PP__1552  (.L_HI(net1552));
 sg13g2_tiehi \cpu.dcache.r_tag[7][3]$_DFFE_PP__1553  (.L_HI(net1553));
 sg13g2_tiehi \cpu.dcache.r_tag[7][4]$_DFFE_PP__1554  (.L_HI(net1554));
 sg13g2_tiehi \cpu.dcache.r_tag[7][5]$_DFFE_PP__1555  (.L_HI(net1555));
 sg13g2_tiehi \cpu.dcache.r_tag[7][6]$_DFFE_PP__1556  (.L_HI(net1556));
 sg13g2_tiehi \cpu.dcache.r_tag[7][7]$_DFFE_PP__1557  (.L_HI(net1557));
 sg13g2_tiehi \cpu.dcache.r_tag[7][8]$_DFFE_PP__1558  (.L_HI(net1558));
 sg13g2_tiehi \cpu.dcache.r_tag[7][9]$_DFFE_PP__1559  (.L_HI(net1559));
 sg13g2_tiehi \cpu.dcache.r_valid[0]$_SDFFE_PP0P__1560  (.L_HI(net1560));
 sg13g2_tiehi \cpu.dcache.r_valid[1]$_SDFFE_PP0P__1561  (.L_HI(net1561));
 sg13g2_tiehi \cpu.dcache.r_valid[2]$_SDFFE_PP0P__1562  (.L_HI(net1562));
 sg13g2_tiehi \cpu.dcache.r_valid[3]$_SDFFE_PP0P__1563  (.L_HI(net1563));
 sg13g2_tiehi \cpu.dcache.r_valid[4]$_SDFFE_PP0P__1564  (.L_HI(net1564));
 sg13g2_tiehi \cpu.dcache.r_valid[5]$_SDFFE_PP0P__1565  (.L_HI(net1565));
 sg13g2_tiehi \cpu.dcache.r_valid[6]$_SDFFE_PP0P__1566  (.L_HI(net1566));
 sg13g2_tiehi \cpu.dcache.r_valid[7]$_SDFFE_PP0P__1567  (.L_HI(net1567));
 sg13g2_tiehi \cpu.dec.r_br$_DFFE_PP__1568  (.L_HI(net1568));
 sg13g2_tiehi \cpu.dec.r_cond[0]$_DFFE_PP__1569  (.L_HI(net1569));
 sg13g2_tiehi \cpu.dec.r_cond[1]$_DFFE_PP__1570  (.L_HI(net1570));
 sg13g2_tiehi \cpu.dec.r_cond[2]$_DFFE_PP__1571  (.L_HI(net1571));
 sg13g2_tiehi \cpu.dec.r_div$_DFFE_PP__1572  (.L_HI(net1572));
 sg13g2_tiehi \cpu.dec.r_flush_all$_DFFE_PP__1573  (.L_HI(net1573));
 sg13g2_tiehi \cpu.dec.r_flush_write$_DFFE_PP__1574  (.L_HI(net1574));
 sg13g2_tiehi \cpu.dec.r_imm[0]$_DFFE_PP__1575  (.L_HI(net1575));
 sg13g2_tiehi \cpu.dec.r_imm[10]$_DFFE_PP__1576  (.L_HI(net1576));
 sg13g2_tiehi \cpu.dec.r_imm[11]$_DFFE_PP__1577  (.L_HI(net1577));
 sg13g2_tiehi \cpu.dec.r_imm[12]$_DFFE_PP__1578  (.L_HI(net1578));
 sg13g2_tiehi \cpu.dec.r_imm[13]$_DFFE_PP__1579  (.L_HI(net1579));
 sg13g2_tiehi \cpu.dec.r_imm[14]$_DFFE_PP__1580  (.L_HI(net1580));
 sg13g2_tiehi \cpu.dec.r_imm[15]$_DFFE_PP__1581  (.L_HI(net1581));
 sg13g2_tiehi \cpu.dec.r_imm[1]$_DFFE_PP__1582  (.L_HI(net1582));
 sg13g2_tiehi \cpu.dec.r_imm[2]$_DFFE_PP__1583  (.L_HI(net1583));
 sg13g2_tiehi \cpu.dec.r_imm[3]$_DFFE_PP__1584  (.L_HI(net1584));
 sg13g2_tiehi \cpu.dec.r_imm[4]$_DFFE_PP__1585  (.L_HI(net1585));
 sg13g2_tiehi \cpu.dec.r_imm[5]$_DFFE_PP__1586  (.L_HI(net1586));
 sg13g2_tiehi \cpu.dec.r_imm[6]$_DFFE_PP__1587  (.L_HI(net1587));
 sg13g2_tiehi \cpu.dec.r_imm[7]$_DFFE_PP__1588  (.L_HI(net1588));
 sg13g2_tiehi \cpu.dec.r_imm[8]$_DFFE_PP__1589  (.L_HI(net1589));
 sg13g2_tiehi \cpu.dec.r_imm[9]$_DFFE_PP__1590  (.L_HI(net1590));
 sg13g2_tiehi \cpu.dec.r_inv_mmu$_DFFE_PP__1591  (.L_HI(net1591));
 sg13g2_tiehi \cpu.dec.r_io$_DFFE_PP__1592  (.L_HI(net1592));
 sg13g2_tiehi \cpu.dec.r_jmp$_SDFFCE_PP0P__1593  (.L_HI(net1593));
 sg13g2_tiehi \cpu.dec.r_load$_DFFE_PP__1594  (.L_HI(net1594));
 sg13g2_tiehi \cpu.dec.r_mult$_DFFE_PP__1595  (.L_HI(net1595));
 sg13g2_tiehi \cpu.dec.r_needs_rs2$_DFFE_PP__1596  (.L_HI(net1596));
 sg13g2_tiehi \cpu.dec.r_op[10]$_DFF_P__1597  (.L_HI(net1597));
 sg13g2_tiehi \cpu.dec.r_op[1]$_DFF_P__1598  (.L_HI(net1598));
 sg13g2_tiehi \cpu.dec.r_op[2]$_DFF_P__1599  (.L_HI(net1599));
 sg13g2_tiehi \cpu.dec.r_op[3]$_DFF_P__1600  (.L_HI(net1600));
 sg13g2_tiehi \cpu.dec.r_op[4]$_DFF_P__1601  (.L_HI(net1601));
 sg13g2_tiehi \cpu.dec.r_op[5]$_DFF_P__1602  (.L_HI(net1602));
 sg13g2_tiehi \cpu.dec.r_op[6]$_DFF_P__1603  (.L_HI(net1603));
 sg13g2_tiehi \cpu.dec.r_op[7]$_DFF_P__1604  (.L_HI(net1604));
 sg13g2_tiehi \cpu.dec.r_op[8]$_DFF_P__1605  (.L_HI(net1605));
 sg13g2_tiehi \cpu.dec.r_op[9]$_DFF_P__1606  (.L_HI(net1606));
 sg13g2_tiehi \cpu.dec.r_rd[0]$_DFFE_PP__1607  (.L_HI(net1607));
 sg13g2_tiehi \cpu.dec.r_rd[1]$_DFFE_PP__1608  (.L_HI(net1608));
 sg13g2_tiehi \cpu.dec.r_rd[2]$_DFFE_PP__1609  (.L_HI(net1609));
 sg13g2_tiehi \cpu.dec.r_rd[3]$_DFFE_PP__1610  (.L_HI(net1610));
 sg13g2_tiehi \cpu.dec.r_ready$_DFF_P__1611  (.L_HI(net1611));
 sg13g2_tiehi \cpu.dec.r_rs1[0]$_DFFE_PP__1612  (.L_HI(net1612));
 sg13g2_tiehi \cpu.dec.r_rs1[1]$_DFFE_PP__1613  (.L_HI(net1613));
 sg13g2_tiehi \cpu.dec.r_rs1[2]$_DFFE_PP__1614  (.L_HI(net1614));
 sg13g2_tiehi \cpu.dec.r_rs1[3]$_DFFE_PP__1615  (.L_HI(net1615));
 sg13g2_tiehi \cpu.dec.r_rs2[0]$_DFFE_PP__1616  (.L_HI(net1616));
 sg13g2_tiehi \cpu.dec.r_rs2[1]$_DFFE_PP__1617  (.L_HI(net1617));
 sg13g2_tiehi \cpu.dec.r_rs2[2]$_DFFE_PP__1618  (.L_HI(net1618));
 sg13g2_tiehi \cpu.dec.r_rs2[3]$_DFFE_PP__1619  (.L_HI(net1619));
 sg13g2_tiehi \cpu.dec.r_rs2_inv$_DFFE_PP__1620  (.L_HI(net1620));
 sg13g2_tiehi \cpu.dec.r_rs2_pc$_DFFE_PP__1621  (.L_HI(net1621));
 sg13g2_tiehi \cpu.dec.r_set_cc$_SDFFCE_PP0P__1622  (.L_HI(net1622));
 sg13g2_tiehi \cpu.dec.r_store$_DFFE_PP__1623  (.L_HI(net1623));
 sg13g2_tiehi \cpu.dec.r_swapsp$_DFFE_PP__1624  (.L_HI(net1624));
 sg13g2_tiehi \cpu.dec.r_sys_call$_DFFE_PP__1625  (.L_HI(net1625));
 sg13g2_tiehi \cpu.dec.r_trap$_DFFE_PP__1626  (.L_HI(net1626));
 sg13g2_tiehi \cpu.ex.genblk3.r_mmu_d_proxy$_SDFFE_PP0P__1627  (.L_HI(net1627));
 sg13g2_tiehi \cpu.ex.genblk3.r_mmu_enable$_SDFFE_PN0P__1628  (.L_HI(net1628));
 sg13g2_tiehi \cpu.ex.genblk3.r_prev_supmode$_SDFFE_PN1P__1629  (.L_HI(net1629));
 sg13g2_tiehi \cpu.ex.genblk3.r_supmode$_DFF_P__1630  (.L_HI(net1630));
 sg13g2_tiehi \cpu.ex.genblk3.r_user_io$_SDFFE_PN0P__1631  (.L_HI(net1631));
 sg13g2_tiehi \cpu.ex.r_10[0]$_DFFE_PP__1632  (.L_HI(net1632));
 sg13g2_tiehi \cpu.ex.r_10[10]$_DFFE_PP__1633  (.L_HI(net1633));
 sg13g2_tiehi \cpu.ex.r_10[11]$_DFFE_PP__1634  (.L_HI(net1634));
 sg13g2_tiehi \cpu.ex.r_10[12]$_DFFE_PP__1635  (.L_HI(net1635));
 sg13g2_tiehi \cpu.ex.r_10[13]$_DFFE_PP__1636  (.L_HI(net1636));
 sg13g2_tiehi \cpu.ex.r_10[14]$_DFFE_PP__1637  (.L_HI(net1637));
 sg13g2_tiehi \cpu.ex.r_10[15]$_DFFE_PP__1638  (.L_HI(net1638));
 sg13g2_tiehi \cpu.ex.r_10[1]$_DFFE_PP__1639  (.L_HI(net1639));
 sg13g2_tiehi \cpu.ex.r_10[2]$_DFFE_PP__1640  (.L_HI(net1640));
 sg13g2_tiehi \cpu.ex.r_10[3]$_DFFE_PP__1641  (.L_HI(net1641));
 sg13g2_tiehi \cpu.ex.r_10[4]$_DFFE_PP__1642  (.L_HI(net1642));
 sg13g2_tiehi \cpu.ex.r_10[5]$_DFFE_PP__1643  (.L_HI(net1643));
 sg13g2_tiehi \cpu.ex.r_10[6]$_DFFE_PP__1644  (.L_HI(net1644));
 sg13g2_tiehi \cpu.ex.r_10[7]$_DFFE_PP__1645  (.L_HI(net1645));
 sg13g2_tiehi \cpu.ex.r_10[8]$_DFFE_PP__1646  (.L_HI(net1646));
 sg13g2_tiehi \cpu.ex.r_10[9]$_DFFE_PP__1647  (.L_HI(net1647));
 sg13g2_tiehi \cpu.ex.r_11[0]$_DFFE_PP__1648  (.L_HI(net1648));
 sg13g2_tiehi \cpu.ex.r_11[10]$_DFFE_PP__1649  (.L_HI(net1649));
 sg13g2_tiehi \cpu.ex.r_11[11]$_DFFE_PP__1650  (.L_HI(net1650));
 sg13g2_tiehi \cpu.ex.r_11[12]$_DFFE_PP__1651  (.L_HI(net1651));
 sg13g2_tiehi \cpu.ex.r_11[13]$_DFFE_PP__1652  (.L_HI(net1652));
 sg13g2_tiehi \cpu.ex.r_11[14]$_DFFE_PP__1653  (.L_HI(net1653));
 sg13g2_tiehi \cpu.ex.r_11[15]$_DFFE_PP__1654  (.L_HI(net1654));
 sg13g2_tiehi \cpu.ex.r_11[1]$_DFFE_PP__1655  (.L_HI(net1655));
 sg13g2_tiehi \cpu.ex.r_11[2]$_DFFE_PP__1656  (.L_HI(net1656));
 sg13g2_tiehi \cpu.ex.r_11[3]$_DFFE_PP__1657  (.L_HI(net1657));
 sg13g2_tiehi \cpu.ex.r_11[4]$_DFFE_PP__1658  (.L_HI(net1658));
 sg13g2_tiehi \cpu.ex.r_11[5]$_DFFE_PP__1659  (.L_HI(net1659));
 sg13g2_tiehi \cpu.ex.r_11[6]$_DFFE_PP__1660  (.L_HI(net1660));
 sg13g2_tiehi \cpu.ex.r_11[7]$_DFFE_PP__1661  (.L_HI(net1661));
 sg13g2_tiehi \cpu.ex.r_11[8]$_DFFE_PP__1662  (.L_HI(net1662));
 sg13g2_tiehi \cpu.ex.r_11[9]$_DFFE_PP__1663  (.L_HI(net1663));
 sg13g2_tiehi \cpu.ex.r_12[0]$_DFFE_PP__1664  (.L_HI(net1664));
 sg13g2_tiehi \cpu.ex.r_12[10]$_DFFE_PP__1665  (.L_HI(net1665));
 sg13g2_tiehi \cpu.ex.r_12[11]$_DFFE_PP__1666  (.L_HI(net1666));
 sg13g2_tiehi \cpu.ex.r_12[12]$_DFFE_PP__1667  (.L_HI(net1667));
 sg13g2_tiehi \cpu.ex.r_12[13]$_DFFE_PP__1668  (.L_HI(net1668));
 sg13g2_tiehi \cpu.ex.r_12[14]$_DFFE_PP__1669  (.L_HI(net1669));
 sg13g2_tiehi \cpu.ex.r_12[15]$_DFFE_PP__1670  (.L_HI(net1670));
 sg13g2_tiehi \cpu.ex.r_12[1]$_DFFE_PP__1671  (.L_HI(net1671));
 sg13g2_tiehi \cpu.ex.r_12[2]$_DFFE_PP__1672  (.L_HI(net1672));
 sg13g2_tiehi \cpu.ex.r_12[3]$_DFFE_PP__1673  (.L_HI(net1673));
 sg13g2_tiehi \cpu.ex.r_12[4]$_DFFE_PP__1674  (.L_HI(net1674));
 sg13g2_tiehi \cpu.ex.r_12[5]$_DFFE_PP__1675  (.L_HI(net1675));
 sg13g2_tiehi \cpu.ex.r_12[6]$_DFFE_PP__1676  (.L_HI(net1676));
 sg13g2_tiehi \cpu.ex.r_12[7]$_DFFE_PP__1677  (.L_HI(net1677));
 sg13g2_tiehi \cpu.ex.r_12[8]$_DFFE_PP__1678  (.L_HI(net1678));
 sg13g2_tiehi \cpu.ex.r_12[9]$_DFFE_PP__1679  (.L_HI(net1679));
 sg13g2_tiehi \cpu.ex.r_13[0]$_DFFE_PP__1680  (.L_HI(net1680));
 sg13g2_tiehi \cpu.ex.r_13[10]$_DFFE_PP__1681  (.L_HI(net1681));
 sg13g2_tiehi \cpu.ex.r_13[11]$_DFFE_PP__1682  (.L_HI(net1682));
 sg13g2_tiehi \cpu.ex.r_13[12]$_DFFE_PP__1683  (.L_HI(net1683));
 sg13g2_tiehi \cpu.ex.r_13[13]$_DFFE_PP__1684  (.L_HI(net1684));
 sg13g2_tiehi \cpu.ex.r_13[14]$_DFFE_PP__1685  (.L_HI(net1685));
 sg13g2_tiehi \cpu.ex.r_13[15]$_DFFE_PP__1686  (.L_HI(net1686));
 sg13g2_tiehi \cpu.ex.r_13[1]$_DFFE_PP__1687  (.L_HI(net1687));
 sg13g2_tiehi \cpu.ex.r_13[2]$_DFFE_PP__1688  (.L_HI(net1688));
 sg13g2_tiehi \cpu.ex.r_13[3]$_DFFE_PP__1689  (.L_HI(net1689));
 sg13g2_tiehi \cpu.ex.r_13[4]$_DFFE_PP__1690  (.L_HI(net1690));
 sg13g2_tiehi \cpu.ex.r_13[5]$_DFFE_PP__1691  (.L_HI(net1691));
 sg13g2_tiehi \cpu.ex.r_13[6]$_DFFE_PP__1692  (.L_HI(net1692));
 sg13g2_tiehi \cpu.ex.r_13[7]$_DFFE_PP__1693  (.L_HI(net1693));
 sg13g2_tiehi \cpu.ex.r_13[8]$_DFFE_PP__1694  (.L_HI(net1694));
 sg13g2_tiehi \cpu.ex.r_13[9]$_DFFE_PP__1695  (.L_HI(net1695));
 sg13g2_tiehi \cpu.ex.r_14[0]$_DFFE_PP__1696  (.L_HI(net1696));
 sg13g2_tiehi \cpu.ex.r_14[10]$_DFFE_PP__1697  (.L_HI(net1697));
 sg13g2_tiehi \cpu.ex.r_14[11]$_DFFE_PP__1698  (.L_HI(net1698));
 sg13g2_tiehi \cpu.ex.r_14[12]$_DFFE_PP__1699  (.L_HI(net1699));
 sg13g2_tiehi \cpu.ex.r_14[13]$_DFFE_PP__1700  (.L_HI(net1700));
 sg13g2_tiehi \cpu.ex.r_14[14]$_DFFE_PP__1701  (.L_HI(net1701));
 sg13g2_tiehi \cpu.ex.r_14[15]$_DFFE_PP__1702  (.L_HI(net1702));
 sg13g2_tiehi \cpu.ex.r_14[1]$_DFFE_PP__1703  (.L_HI(net1703));
 sg13g2_tiehi \cpu.ex.r_14[2]$_DFFE_PP__1704  (.L_HI(net1704));
 sg13g2_tiehi \cpu.ex.r_14[3]$_DFFE_PP__1705  (.L_HI(net1705));
 sg13g2_tiehi \cpu.ex.r_14[4]$_DFFE_PP__1706  (.L_HI(net1706));
 sg13g2_tiehi \cpu.ex.r_14[5]$_DFFE_PP__1707  (.L_HI(net1707));
 sg13g2_tiehi \cpu.ex.r_14[6]$_DFFE_PP__1708  (.L_HI(net1708));
 sg13g2_tiehi \cpu.ex.r_14[7]$_DFFE_PP__1709  (.L_HI(net1709));
 sg13g2_tiehi \cpu.ex.r_14[8]$_DFFE_PP__1710  (.L_HI(net1710));
 sg13g2_tiehi \cpu.ex.r_14[9]$_DFFE_PP__1711  (.L_HI(net1711));
 sg13g2_tiehi \cpu.ex.r_15[0]$_DFFE_PP__1712  (.L_HI(net1712));
 sg13g2_tiehi \cpu.ex.r_15[10]$_DFFE_PP__1713  (.L_HI(net1713));
 sg13g2_tiehi \cpu.ex.r_15[11]$_DFFE_PP__1714  (.L_HI(net1714));
 sg13g2_tiehi \cpu.ex.r_15[12]$_DFFE_PP__1715  (.L_HI(net1715));
 sg13g2_tiehi \cpu.ex.r_15[13]$_DFFE_PP__1716  (.L_HI(net1716));
 sg13g2_tiehi \cpu.ex.r_15[14]$_DFFE_PP__1717  (.L_HI(net1717));
 sg13g2_tiehi \cpu.ex.r_15[15]$_DFFE_PP__1718  (.L_HI(net1718));
 sg13g2_tiehi \cpu.ex.r_15[1]$_DFFE_PP__1719  (.L_HI(net1719));
 sg13g2_tiehi \cpu.ex.r_15[2]$_DFFE_PP__1720  (.L_HI(net1720));
 sg13g2_tiehi \cpu.ex.r_15[3]$_DFFE_PP__1721  (.L_HI(net1721));
 sg13g2_tiehi \cpu.ex.r_15[4]$_DFFE_PP__1722  (.L_HI(net1722));
 sg13g2_tiehi \cpu.ex.r_15[5]$_DFFE_PP__1723  (.L_HI(net1723));
 sg13g2_tiehi \cpu.ex.r_15[6]$_DFFE_PP__1724  (.L_HI(net1724));
 sg13g2_tiehi \cpu.ex.r_15[7]$_DFFE_PP__1725  (.L_HI(net1725));
 sg13g2_tiehi \cpu.ex.r_15[8]$_DFFE_PP__1726  (.L_HI(net1726));
 sg13g2_tiehi \cpu.ex.r_15[9]$_DFFE_PP__1727  (.L_HI(net1727));
 sg13g2_tiehi \cpu.ex.r_8[0]$_DFFE_PP__1728  (.L_HI(net1728));
 sg13g2_tiehi \cpu.ex.r_8[10]$_DFFE_PP__1729  (.L_HI(net1729));
 sg13g2_tiehi \cpu.ex.r_8[11]$_DFFE_PP__1730  (.L_HI(net1730));
 sg13g2_tiehi \cpu.ex.r_8[12]$_DFFE_PP__1731  (.L_HI(net1731));
 sg13g2_tiehi \cpu.ex.r_8[13]$_DFFE_PP__1732  (.L_HI(net1732));
 sg13g2_tiehi \cpu.ex.r_8[14]$_DFFE_PP__1733  (.L_HI(net1733));
 sg13g2_tiehi \cpu.ex.r_8[15]$_DFFE_PP__1734  (.L_HI(net1734));
 sg13g2_tiehi \cpu.ex.r_8[1]$_DFFE_PP__1735  (.L_HI(net1735));
 sg13g2_tiehi \cpu.ex.r_8[2]$_DFFE_PP__1736  (.L_HI(net1736));
 sg13g2_tiehi \cpu.ex.r_8[3]$_DFFE_PP__1737  (.L_HI(net1737));
 sg13g2_tiehi \cpu.ex.r_8[4]$_DFFE_PP__1738  (.L_HI(net1738));
 sg13g2_tiehi \cpu.ex.r_8[5]$_DFFE_PP__1739  (.L_HI(net1739));
 sg13g2_tiehi \cpu.ex.r_8[6]$_DFFE_PP__1740  (.L_HI(net1740));
 sg13g2_tiehi \cpu.ex.r_8[7]$_DFFE_PP__1741  (.L_HI(net1741));
 sg13g2_tiehi \cpu.ex.r_8[8]$_DFFE_PP__1742  (.L_HI(net1742));
 sg13g2_tiehi \cpu.ex.r_8[9]$_DFFE_PP__1743  (.L_HI(net1743));
 sg13g2_tiehi \cpu.ex.r_9[0]$_DFFE_PP__1744  (.L_HI(net1744));
 sg13g2_tiehi \cpu.ex.r_9[10]$_DFFE_PP__1745  (.L_HI(net1745));
 sg13g2_tiehi \cpu.ex.r_9[11]$_DFFE_PP__1746  (.L_HI(net1746));
 sg13g2_tiehi \cpu.ex.r_9[12]$_DFFE_PP__1747  (.L_HI(net1747));
 sg13g2_tiehi \cpu.ex.r_9[13]$_DFFE_PP__1748  (.L_HI(net1748));
 sg13g2_tiehi \cpu.ex.r_9[14]$_DFFE_PP__1749  (.L_HI(net1749));
 sg13g2_tiehi \cpu.ex.r_9[15]$_DFFE_PP__1750  (.L_HI(net1750));
 sg13g2_tiehi \cpu.ex.r_9[1]$_DFFE_PP__1751  (.L_HI(net1751));
 sg13g2_tiehi \cpu.ex.r_9[2]$_DFFE_PP__1752  (.L_HI(net1752));
 sg13g2_tiehi \cpu.ex.r_9[3]$_DFFE_PP__1753  (.L_HI(net1753));
 sg13g2_tiehi \cpu.ex.r_9[4]$_DFFE_PP__1754  (.L_HI(net1754));
 sg13g2_tiehi \cpu.ex.r_9[5]$_DFFE_PP__1755  (.L_HI(net1755));
 sg13g2_tiehi \cpu.ex.r_9[6]$_DFFE_PP__1756  (.L_HI(net1756));
 sg13g2_tiehi \cpu.ex.r_9[7]$_DFFE_PP__1757  (.L_HI(net1757));
 sg13g2_tiehi \cpu.ex.r_9[8]$_DFFE_PP__1758  (.L_HI(net1758));
 sg13g2_tiehi \cpu.ex.r_9[9]$_DFFE_PP__1759  (.L_HI(net1759));
 sg13g2_tiehi \cpu.ex.r_branch_stall$_DFF_P__1760  (.L_HI(net1760));
 sg13g2_tiehi \cpu.ex.r_cc$_DFFE_PP__1761  (.L_HI(net1761));
 sg13g2_tiehi \cpu.ex.r_d_flush_all$_SDFF_PP0__1762  (.L_HI(net1762));
 sg13g2_tiehi \cpu.ex.r_div_running$_DFF_P__1763  (.L_HI(net1763));
 sg13g2_tiehi \cpu.ex.r_epc[0]$_DFFE_PP__1764  (.L_HI(net1764));
 sg13g2_tiehi \cpu.ex.r_epc[10]$_DFFE_PP__1765  (.L_HI(net1765));
 sg13g2_tiehi \cpu.ex.r_epc[11]$_DFFE_PP__1766  (.L_HI(net1766));
 sg13g2_tiehi \cpu.ex.r_epc[12]$_DFFE_PP__1767  (.L_HI(net1767));
 sg13g2_tiehi \cpu.ex.r_epc[13]$_DFFE_PP__1768  (.L_HI(net1768));
 sg13g2_tiehi \cpu.ex.r_epc[14]$_DFFE_PP__1769  (.L_HI(net1769));
 sg13g2_tiehi \cpu.ex.r_epc[1]$_DFFE_PP__1770  (.L_HI(net1770));
 sg13g2_tiehi \cpu.ex.r_epc[2]$_DFFE_PP__1771  (.L_HI(net1771));
 sg13g2_tiehi \cpu.ex.r_epc[3]$_DFFE_PP__1772  (.L_HI(net1772));
 sg13g2_tiehi \cpu.ex.r_epc[4]$_DFFE_PP__1773  (.L_HI(net1773));
 sg13g2_tiehi \cpu.ex.r_epc[5]$_DFFE_PP__1774  (.L_HI(net1774));
 sg13g2_tiehi \cpu.ex.r_epc[6]$_DFFE_PP__1775  (.L_HI(net1775));
 sg13g2_tiehi \cpu.ex.r_epc[7]$_DFFE_PP__1776  (.L_HI(net1776));
 sg13g2_tiehi \cpu.ex.r_epc[8]$_DFFE_PP__1777  (.L_HI(net1777));
 sg13g2_tiehi \cpu.ex.r_epc[9]$_DFFE_PP__1778  (.L_HI(net1778));
 sg13g2_tiehi \cpu.ex.r_fetch$_SDFF_PN1__1779  (.L_HI(net1779));
 sg13g2_tiehi \cpu.ex.r_flush_write$_SDFFE_PN0P__1780  (.L_HI(net1780));
 sg13g2_tiehi \cpu.ex.r_i_flush_all$_SDFF_PP0__1781  (.L_HI(net1781));
 sg13g2_tiehi \cpu.ex.r_ie$_SDFFE_PP0P__1782  (.L_HI(net1782));
 sg13g2_tiehi \cpu.ex.r_io_access$_SDFFE_PN0P__1783  (.L_HI(net1783));
 sg13g2_tiehi \cpu.ex.r_lr[0]$_DFFE_PP__1784  (.L_HI(net1784));
 sg13g2_tiehi \cpu.ex.r_lr[10]$_DFFE_PP__1785  (.L_HI(net1785));
 sg13g2_tiehi \cpu.ex.r_lr[11]$_DFFE_PP__1786  (.L_HI(net1786));
 sg13g2_tiehi \cpu.ex.r_lr[12]$_DFFE_PP__1787  (.L_HI(net1787));
 sg13g2_tiehi \cpu.ex.r_lr[13]$_DFFE_PP__1788  (.L_HI(net1788));
 sg13g2_tiehi \cpu.ex.r_lr[14]$_DFFE_PP__1789  (.L_HI(net1789));
 sg13g2_tiehi \cpu.ex.r_lr[1]$_DFFE_PP__1790  (.L_HI(net1790));
 sg13g2_tiehi \cpu.ex.r_lr[2]$_DFFE_PP__1791  (.L_HI(net1791));
 sg13g2_tiehi \cpu.ex.r_lr[3]$_DFFE_PP__1792  (.L_HI(net1792));
 sg13g2_tiehi \cpu.ex.r_lr[4]$_DFFE_PP__1793  (.L_HI(net1793));
 sg13g2_tiehi \cpu.ex.r_lr[5]$_DFFE_PP__1794  (.L_HI(net1794));
 sg13g2_tiehi \cpu.ex.r_lr[6]$_DFFE_PP__1795  (.L_HI(net1795));
 sg13g2_tiehi \cpu.ex.r_lr[7]$_DFFE_PP__1796  (.L_HI(net1796));
 sg13g2_tiehi \cpu.ex.r_lr[8]$_DFFE_PP__1797  (.L_HI(net1797));
 sg13g2_tiehi \cpu.ex.r_lr[9]$_DFFE_PP__1798  (.L_HI(net1798));
 sg13g2_tiehi \cpu.ex.r_mult[0]$_DFF_P__1799  (.L_HI(net1799));
 sg13g2_tiehi \cpu.ex.r_mult[10]$_DFF_P__1800  (.L_HI(net1800));
 sg13g2_tiehi \cpu.ex.r_mult[11]$_DFF_P__1801  (.L_HI(net1801));
 sg13g2_tiehi \cpu.ex.r_mult[12]$_DFF_P__1802  (.L_HI(net1802));
 sg13g2_tiehi \cpu.ex.r_mult[13]$_DFF_P__1803  (.L_HI(net1803));
 sg13g2_tiehi \cpu.ex.r_mult[14]$_DFF_P__1804  (.L_HI(net1804));
 sg13g2_tiehi \cpu.ex.r_mult[15]$_DFF_P__1805  (.L_HI(net1805));
 sg13g2_tiehi \cpu.ex.r_mult[16]$_DFFE_PP__1806  (.L_HI(net1806));
 sg13g2_tiehi \cpu.ex.r_mult[17]$_DFFE_PP__1807  (.L_HI(net1807));
 sg13g2_tiehi \cpu.ex.r_mult[18]$_DFFE_PP__1808  (.L_HI(net1808));
 sg13g2_tiehi \cpu.ex.r_mult[19]$_DFFE_PP__1809  (.L_HI(net1809));
 sg13g2_tiehi \cpu.ex.r_mult[1]$_DFF_P__1810  (.L_HI(net1810));
 sg13g2_tiehi \cpu.ex.r_mult[20]$_DFFE_PP__1811  (.L_HI(net1811));
 sg13g2_tiehi \cpu.ex.r_mult[21]$_DFFE_PP__1812  (.L_HI(net1812));
 sg13g2_tiehi \cpu.ex.r_mult[22]$_DFFE_PP__1813  (.L_HI(net1813));
 sg13g2_tiehi \cpu.ex.r_mult[23]$_DFFE_PP__1814  (.L_HI(net1814));
 sg13g2_tiehi \cpu.ex.r_mult[24]$_DFFE_PP__1815  (.L_HI(net1815));
 sg13g2_tiehi \cpu.ex.r_mult[25]$_DFFE_PP__1816  (.L_HI(net1816));
 sg13g2_tiehi \cpu.ex.r_mult[26]$_DFFE_PP__1817  (.L_HI(net1817));
 sg13g2_tiehi \cpu.ex.r_mult[27]$_DFFE_PP__1818  (.L_HI(net1818));
 sg13g2_tiehi \cpu.ex.r_mult[28]$_DFFE_PP__1819  (.L_HI(net1819));
 sg13g2_tiehi \cpu.ex.r_mult[29]$_DFFE_PP__1820  (.L_HI(net1820));
 sg13g2_tiehi \cpu.ex.r_mult[2]$_DFF_P__1821  (.L_HI(net1821));
 sg13g2_tiehi \cpu.ex.r_mult[30]$_DFFE_PP__1822  (.L_HI(net1822));
 sg13g2_tiehi \cpu.ex.r_mult[31]$_DFFE_PP__1823  (.L_HI(net1823));
 sg13g2_tiehi \cpu.ex.r_mult[3]$_DFF_P__1824  (.L_HI(net1824));
 sg13g2_tiehi \cpu.ex.r_mult[4]$_DFF_P__1825  (.L_HI(net1825));
 sg13g2_tiehi \cpu.ex.r_mult[5]$_DFF_P__1826  (.L_HI(net1826));
 sg13g2_tiehi \cpu.ex.r_mult[6]$_DFF_P__1827  (.L_HI(net1827));
 sg13g2_tiehi \cpu.ex.r_mult[7]$_DFF_P__1828  (.L_HI(net1828));
 sg13g2_tiehi \cpu.ex.r_mult[8]$_DFF_P__1829  (.L_HI(net1829));
 sg13g2_tiehi \cpu.ex.r_mult[9]$_DFF_P__1830  (.L_HI(net1830));
 sg13g2_tiehi \cpu.ex.r_mult_off[0]$_DFF_P__1831  (.L_HI(net1831));
 sg13g2_tiehi \cpu.ex.r_mult_off[1]$_DFF_P__1832  (.L_HI(net1832));
 sg13g2_tiehi \cpu.ex.r_mult_off[2]$_DFF_P__1833  (.L_HI(net1833));
 sg13g2_tiehi \cpu.ex.r_mult_off[3]$_DFF_P__1834  (.L_HI(net1834));
 sg13g2_tiehi \cpu.ex.r_mult_running$_DFF_P__1835  (.L_HI(net1835));
 sg13g2_tiehi \cpu.ex.r_pc[0]$_DFFE_PP__1836  (.L_HI(net1836));
 sg13g2_tiehi \cpu.ex.r_pc[10]$_DFFE_PP__1837  (.L_HI(net1837));
 sg13g2_tiehi \cpu.ex.r_pc[11]$_DFFE_PP__1838  (.L_HI(net1838));
 sg13g2_tiehi \cpu.ex.r_pc[12]$_DFFE_PP__1839  (.L_HI(net1839));
 sg13g2_tiehi \cpu.ex.r_pc[13]$_DFFE_PP__1840  (.L_HI(net1840));
 sg13g2_tiehi \cpu.ex.r_pc[14]$_DFFE_PP__1841  (.L_HI(net1841));
 sg13g2_tiehi \cpu.ex.r_pc[1]$_DFFE_PP__1842  (.L_HI(net1842));
 sg13g2_tiehi \cpu.ex.r_pc[2]$_DFFE_PP__1843  (.L_HI(net1843));
 sg13g2_tiehi \cpu.ex.r_pc[3]$_DFFE_PP__1844  (.L_HI(net1844));
 sg13g2_tiehi \cpu.ex.r_pc[4]$_DFFE_PP__1845  (.L_HI(net1845));
 sg13g2_tiehi \cpu.ex.r_pc[5]$_DFFE_PP__1846  (.L_HI(net1846));
 sg13g2_tiehi \cpu.ex.r_pc[6]$_DFFE_PP__1847  (.L_HI(net1847));
 sg13g2_tiehi \cpu.ex.r_pc[7]$_DFFE_PP__1848  (.L_HI(net1848));
 sg13g2_tiehi \cpu.ex.r_pc[8]$_DFFE_PP__1849  (.L_HI(net1849));
 sg13g2_tiehi \cpu.ex.r_pc[9]$_DFFE_PP__1850  (.L_HI(net1850));
 sg13g2_tiehi \cpu.ex.r_prev_ie$_SDFFE_PN0P__1851  (.L_HI(net1851));
 sg13g2_tiehi \cpu.ex.r_read_stall$_SDFFE_PN0P__1852  (.L_HI(net1852));
 sg13g2_tiehi \cpu.ex.r_set_cc$_DFFE_PP__1853  (.L_HI(net1853));
 sg13g2_tiehi \cpu.ex.r_sp[0]$_DFFE_PP__1854  (.L_HI(net1854));
 sg13g2_tiehi \cpu.ex.r_sp[10]$_DFFE_PP__1855  (.L_HI(net1855));
 sg13g2_tiehi \cpu.ex.r_sp[11]$_DFFE_PP__1856  (.L_HI(net1856));
 sg13g2_tiehi \cpu.ex.r_sp[12]$_DFFE_PP__1857  (.L_HI(net1857));
 sg13g2_tiehi \cpu.ex.r_sp[13]$_DFFE_PP__1858  (.L_HI(net1858));
 sg13g2_tiehi \cpu.ex.r_sp[14]$_DFFE_PP__1859  (.L_HI(net1859));
 sg13g2_tiehi \cpu.ex.r_sp[1]$_DFFE_PP__1860  (.L_HI(net1860));
 sg13g2_tiehi \cpu.ex.r_sp[2]$_DFFE_PP__1861  (.L_HI(net1861));
 sg13g2_tiehi \cpu.ex.r_sp[3]$_DFFE_PP__1862  (.L_HI(net1862));
 sg13g2_tiehi \cpu.ex.r_sp[4]$_DFFE_PP__1863  (.L_HI(net1863));
 sg13g2_tiehi \cpu.ex.r_sp[5]$_DFFE_PP__1864  (.L_HI(net1864));
 sg13g2_tiehi \cpu.ex.r_sp[6]$_DFFE_PP__1865  (.L_HI(net1865));
 sg13g2_tiehi \cpu.ex.r_sp[7]$_DFFE_PP__1866  (.L_HI(net1866));
 sg13g2_tiehi \cpu.ex.r_sp[8]$_DFFE_PP__1867  (.L_HI(net1867));
 sg13g2_tiehi \cpu.ex.r_sp[9]$_DFFE_PP__1868  (.L_HI(net1868));
 sg13g2_tiehi \cpu.ex.r_stmp[0]$_SDFFCE_PN0P__1869  (.L_HI(net1869));
 sg13g2_tiehi \cpu.ex.r_stmp[10]$_DFFE_PP__1870  (.L_HI(net1870));
 sg13g2_tiehi \cpu.ex.r_stmp[11]$_DFFE_PP__1871  (.L_HI(net1871));
 sg13g2_tiehi \cpu.ex.r_stmp[12]$_DFFE_PP__1872  (.L_HI(net1872));
 sg13g2_tiehi \cpu.ex.r_stmp[13]$_DFFE_PP__1873  (.L_HI(net1873));
 sg13g2_tiehi \cpu.ex.r_stmp[14]$_DFFE_PP__1874  (.L_HI(net1874));
 sg13g2_tiehi \cpu.ex.r_stmp[15]$_DFFE_PP__1875  (.L_HI(net1875));
 sg13g2_tiehi \cpu.ex.r_stmp[1]$_DFFE_PP__1876  (.L_HI(net1876));
 sg13g2_tiehi \cpu.ex.r_stmp[2]$_DFFE_PP__1877  (.L_HI(net1877));
 sg13g2_tiehi \cpu.ex.r_stmp[3]$_DFFE_PP__1878  (.L_HI(net1878));
 sg13g2_tiehi \cpu.ex.r_stmp[4]$_DFFE_PP__1879  (.L_HI(net1879));
 sg13g2_tiehi \cpu.ex.r_stmp[5]$_DFFE_PP__1880  (.L_HI(net1880));
 sg13g2_tiehi \cpu.ex.r_stmp[6]$_DFFE_PP__1881  (.L_HI(net1881));
 sg13g2_tiehi \cpu.ex.r_stmp[7]$_DFFE_PP__1882  (.L_HI(net1882));
 sg13g2_tiehi \cpu.ex.r_stmp[8]$_DFFE_PP__1883  (.L_HI(net1883));
 sg13g2_tiehi \cpu.ex.r_stmp[9]$_DFFE_PP__1884  (.L_HI(net1884));
 sg13g2_tiehi \cpu.ex.r_wb[0]$_DFFE_PP__1885  (.L_HI(net1885));
 sg13g2_tiehi \cpu.ex.r_wb[10]$_DFFE_PP__1886  (.L_HI(net1886));
 sg13g2_tiehi \cpu.ex.r_wb[11]$_DFFE_PP__1887  (.L_HI(net1887));
 sg13g2_tiehi \cpu.ex.r_wb[12]$_DFFE_PP__1888  (.L_HI(net1888));
 sg13g2_tiehi \cpu.ex.r_wb[13]$_DFFE_PP__1889  (.L_HI(net1889));
 sg13g2_tiehi \cpu.ex.r_wb[14]$_DFFE_PP__1890  (.L_HI(net1890));
 sg13g2_tiehi \cpu.ex.r_wb[15]$_DFFE_PP__1891  (.L_HI(net1891));
 sg13g2_tiehi \cpu.ex.r_wb[1]$_DFFE_PP__1892  (.L_HI(net1892));
 sg13g2_tiehi \cpu.ex.r_wb[2]$_DFFE_PP__1893  (.L_HI(net1893));
 sg13g2_tiehi \cpu.ex.r_wb[3]$_DFFE_PP__1894  (.L_HI(net1894));
 sg13g2_tiehi \cpu.ex.r_wb[4]$_DFFE_PP__1895  (.L_HI(net1895));
 sg13g2_tiehi \cpu.ex.r_wb[5]$_DFFE_PP__1896  (.L_HI(net1896));
 sg13g2_tiehi \cpu.ex.r_wb[6]$_DFFE_PP__1897  (.L_HI(net1897));
 sg13g2_tiehi \cpu.ex.r_wb[7]$_DFFE_PP__1898  (.L_HI(net1898));
 sg13g2_tiehi \cpu.ex.r_wb[8]$_DFFE_PP__1899  (.L_HI(net1899));
 sg13g2_tiehi \cpu.ex.r_wb[9]$_DFFE_PP__1900  (.L_HI(net1900));
 sg13g2_tiehi \cpu.ex.r_wb_addr[0]$_SDFFCE_PN0P__1901  (.L_HI(net1901));
 sg13g2_tiehi \cpu.ex.r_wb_addr[1]$_SDFFCE_PN0P__1902  (.L_HI(net1902));
 sg13g2_tiehi \cpu.ex.r_wb_addr[2]$_SDFFCE_PP0P__1903  (.L_HI(net1903));
 sg13g2_tiehi \cpu.ex.r_wb_addr[3]$_SDFFCE_PP0P__1904  (.L_HI(net1904));
 sg13g2_tiehi \cpu.ex.r_wb_swapsp$_DFFE_PP__1905  (.L_HI(net1905));
 sg13g2_tiehi \cpu.ex.r_wb_valid$_DFF_P__1906  (.L_HI(net1906));
 sg13g2_tiehi \cpu.ex.r_wdata[0]$_DFFE_PP__1907  (.L_HI(net1907));
 sg13g2_tiehi \cpu.ex.r_wdata[10]$_DFFE_PP__1908  (.L_HI(net1908));
 sg13g2_tiehi \cpu.ex.r_wdata[11]$_DFFE_PP__1909  (.L_HI(net1909));
 sg13g2_tiehi \cpu.ex.r_wdata[12]$_DFFE_PP__1910  (.L_HI(net1910));
 sg13g2_tiehi \cpu.ex.r_wdata[13]$_DFFE_PP__1911  (.L_HI(net1911));
 sg13g2_tiehi \cpu.ex.r_wdata[14]$_DFFE_PP__1912  (.L_HI(net1912));
 sg13g2_tiehi \cpu.ex.r_wdata[15]$_DFFE_PP__1913  (.L_HI(net1913));
 sg13g2_tiehi \cpu.ex.r_wdata[1]$_DFFE_PP__1914  (.L_HI(net1914));
 sg13g2_tiehi \cpu.ex.r_wdata[2]$_DFFE_PP__1915  (.L_HI(net1915));
 sg13g2_tiehi \cpu.ex.r_wdata[3]$_DFFE_PP__1916  (.L_HI(net1916));
 sg13g2_tiehi \cpu.ex.r_wdata[4]$_DFFE_PP__1917  (.L_HI(net1917));
 sg13g2_tiehi \cpu.ex.r_wdata[5]$_DFFE_PP__1918  (.L_HI(net1918));
 sg13g2_tiehi \cpu.ex.r_wdata[6]$_DFFE_PP__1919  (.L_HI(net1919));
 sg13g2_tiehi \cpu.ex.r_wdata[7]$_DFFE_PP__1920  (.L_HI(net1920));
 sg13g2_tiehi \cpu.ex.r_wdata[8]$_DFFE_PP__1921  (.L_HI(net1921));
 sg13g2_tiehi \cpu.ex.r_wdata[9]$_DFFE_PP__1922  (.L_HI(net1922));
 sg13g2_tiehi \cpu.ex.r_wmask[0]$_SDFFE_PP0P__1923  (.L_HI(net1923));
 sg13g2_tiehi \cpu.ex.r_wmask[1]$_SDFFE_PP0P__1924  (.L_HI(net1924));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[0]$_DFFE_PP__1925  (.L_HI(net1925));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[1]$_DFFE_PP__1926  (.L_HI(net1926));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[2]$_DFFE_PP__1927  (.L_HI(net1927));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[3]$_DFFE_PP__1928  (.L_HI(net1928));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_ins$_SDFFE_PN0P__1929  (.L_HI(net1929));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_sup$_SDFFE_PN0P__1930  (.L_HI(net1930));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_type$_SDFFE_PN0P__1931  (.L_HI(net1931));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[0]$_SDFFE_PN0P__1932  (.L_HI(net1932));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[10]$_SDFFE_PN0P__1933  (.L_HI(net1933));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[11]$_SDFFE_PN0P__1934  (.L_HI(net1934));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[12]$_SDFFE_PN0P__1935  (.L_HI(net1935));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[13]$_SDFFE_PN0P__1936  (.L_HI(net1936));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[14]$_SDFFE_PN0P__1937  (.L_HI(net1937));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[15]$_SDFFE_PN0P__1938  (.L_HI(net1938));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[16]$_SDFFE_PN0P__1939  (.L_HI(net1939));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[17]$_SDFFE_PN0P__1940  (.L_HI(net1940));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[18]$_SDFFE_PN0P__1941  (.L_HI(net1941));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[19]$_SDFFE_PN0P__1942  (.L_HI(net1942));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[1]$_SDFFE_PN0P__1943  (.L_HI(net1943));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[20]$_SDFFE_PN0P__1944  (.L_HI(net1944));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[21]$_SDFFE_PN0P__1945  (.L_HI(net1945));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[22]$_SDFFE_PN0P__1946  (.L_HI(net1946));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[23]$_SDFFE_PN0P__1947  (.L_HI(net1947));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[24]$_SDFFE_PN0P__1948  (.L_HI(net1948));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[25]$_SDFFE_PN0P__1949  (.L_HI(net1949));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[26]$_SDFFE_PN0P__1950  (.L_HI(net1950));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[27]$_SDFFE_PN0P__1951  (.L_HI(net1951));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[28]$_SDFFE_PN0P__1952  (.L_HI(net1952));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[29]$_SDFFE_PN0P__1953  (.L_HI(net1953));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[2]$_SDFFE_PN0P__1954  (.L_HI(net1954));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[30]$_SDFFE_PN0P__1955  (.L_HI(net1955));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[31]$_SDFFE_PN0P__1956  (.L_HI(net1956));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[3]$_SDFFE_PN0P__1957  (.L_HI(net1957));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[4]$_SDFFE_PN0P__1958  (.L_HI(net1958));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[5]$_SDFFE_PN0P__1959  (.L_HI(net1959));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[6]$_SDFFE_PN0P__1960  (.L_HI(net1960));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[7]$_SDFFE_PN0P__1961  (.L_HI(net1961));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[8]$_SDFFE_PN0P__1962  (.L_HI(net1962));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[9]$_SDFFE_PN0P__1963  (.L_HI(net1963));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[0]$_SDFFE_PN0P__1964  (.L_HI(net1964));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[10]$_SDFFE_PN0P__1965  (.L_HI(net1965));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[11]$_SDFFE_PN0P__1966  (.L_HI(net1966));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[12]$_SDFFE_PN0P__1967  (.L_HI(net1967));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[13]$_SDFFE_PN0P__1968  (.L_HI(net1968));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[14]$_SDFFE_PN0P__1969  (.L_HI(net1969));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[15]$_SDFFE_PN0P__1970  (.L_HI(net1970));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[16]$_SDFFE_PN0P__1971  (.L_HI(net1971));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[17]$_SDFFE_PN0P__1972  (.L_HI(net1972));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[18]$_SDFFE_PN0P__1973  (.L_HI(net1973));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[19]$_SDFFE_PN0P__1974  (.L_HI(net1974));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[1]$_SDFFE_PN0P__1975  (.L_HI(net1975));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[20]$_SDFFE_PN0P__1976  (.L_HI(net1976));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[21]$_SDFFE_PN0P__1977  (.L_HI(net1977));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[22]$_SDFFE_PN0P__1978  (.L_HI(net1978));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[23]$_SDFFE_PN0P__1979  (.L_HI(net1979));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[24]$_SDFFE_PN0P__1980  (.L_HI(net1980));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[25]$_SDFFE_PN0P__1981  (.L_HI(net1981));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[26]$_SDFFE_PN0P__1982  (.L_HI(net1982));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[27]$_SDFFE_PN0P__1983  (.L_HI(net1983));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[28]$_SDFFE_PN0P__1984  (.L_HI(net1984));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[29]$_SDFFE_PN0P__1985  (.L_HI(net1985));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[2]$_SDFFE_PN0P__1986  (.L_HI(net1986));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[30]$_SDFFE_PN0P__1987  (.L_HI(net1987));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[31]$_SDFFE_PN0P__1988  (.L_HI(net1988));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[3]$_SDFFE_PN0P__1989  (.L_HI(net1989));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[4]$_SDFFE_PN0P__1990  (.L_HI(net1990));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[5]$_SDFFE_PN0P__1991  (.L_HI(net1991));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[6]$_SDFFE_PN0P__1992  (.L_HI(net1992));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[7]$_SDFFE_PN0P__1993  (.L_HI(net1993));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[8]$_SDFFE_PN0P__1994  (.L_HI(net1994));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[9]$_SDFFE_PN0P__1995  (.L_HI(net1995));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][0]$_DFFE_PP__1996  (.L_HI(net1996));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][10]$_DFFE_PP__1997  (.L_HI(net1997));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][11]$_DFFE_PP__1998  (.L_HI(net1998));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][1]$_DFFE_PP__1999  (.L_HI(net1999));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][2]$_DFFE_PP__2000  (.L_HI(net2000));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][3]$_DFFE_PP__2001  (.L_HI(net2001));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][4]$_DFFE_PP__2002  (.L_HI(net2002));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][5]$_DFFE_PP__2003  (.L_HI(net2003));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][6]$_DFFE_PP__2004  (.L_HI(net2004));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][7]$_DFFE_PP__2005  (.L_HI(net2005));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][8]$_DFFE_PP__2006  (.L_HI(net2006));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][9]$_DFFE_PP__2007  (.L_HI(net2007));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][0]$_DFFE_PP__2008  (.L_HI(net2008));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][10]$_DFFE_PP__2009  (.L_HI(net2009));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][11]$_DFFE_PP__2010  (.L_HI(net2010));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][1]$_DFFE_PP__2011  (.L_HI(net2011));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][2]$_DFFE_PP__2012  (.L_HI(net2012));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][3]$_DFFE_PP__2013  (.L_HI(net2013));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][4]$_DFFE_PP__2014  (.L_HI(net2014));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][5]$_DFFE_PP__2015  (.L_HI(net2015));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][6]$_DFFE_PP__2016  (.L_HI(net2016));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][7]$_DFFE_PP__2017  (.L_HI(net2017));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][8]$_DFFE_PP__2018  (.L_HI(net2018));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][9]$_DFFE_PP__2019  (.L_HI(net2019));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][0]$_DFFE_PP__2020  (.L_HI(net2020));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][10]$_DFFE_PP__2021  (.L_HI(net2021));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][11]$_DFFE_PP__2022  (.L_HI(net2022));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][1]$_DFFE_PP__2023  (.L_HI(net2023));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][2]$_DFFE_PP__2024  (.L_HI(net2024));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][3]$_DFFE_PP__2025  (.L_HI(net2025));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][4]$_DFFE_PP__2026  (.L_HI(net2026));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][5]$_DFFE_PP__2027  (.L_HI(net2027));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][6]$_DFFE_PP__2028  (.L_HI(net2028));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][7]$_DFFE_PP__2029  (.L_HI(net2029));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][8]$_DFFE_PP__2030  (.L_HI(net2030));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][9]$_DFFE_PP__2031  (.L_HI(net2031));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][0]$_DFFE_PP__2032  (.L_HI(net2032));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][10]$_DFFE_PP__2033  (.L_HI(net2033));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][11]$_DFFE_PP__2034  (.L_HI(net2034));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][1]$_DFFE_PP__2035  (.L_HI(net2035));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][2]$_DFFE_PP__2036  (.L_HI(net2036));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][3]$_DFFE_PP__2037  (.L_HI(net2037));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][4]$_DFFE_PP__2038  (.L_HI(net2038));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][5]$_DFFE_PP__2039  (.L_HI(net2039));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][6]$_DFFE_PP__2040  (.L_HI(net2040));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][7]$_DFFE_PP__2041  (.L_HI(net2041));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][8]$_DFFE_PP__2042  (.L_HI(net2042));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][9]$_DFFE_PP__2043  (.L_HI(net2043));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][0]$_DFFE_PP__2044  (.L_HI(net2044));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][10]$_DFFE_PP__2045  (.L_HI(net2045));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][11]$_DFFE_PP__2046  (.L_HI(net2046));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][1]$_DFFE_PP__2047  (.L_HI(net2047));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][2]$_DFFE_PP__2048  (.L_HI(net2048));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][3]$_DFFE_PP__2049  (.L_HI(net2049));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][4]$_DFFE_PP__2050  (.L_HI(net2050));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][5]$_DFFE_PP__2051  (.L_HI(net2051));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][6]$_DFFE_PP__2052  (.L_HI(net2052));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][7]$_DFFE_PP__2053  (.L_HI(net2053));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][8]$_DFFE_PP__2054  (.L_HI(net2054));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][9]$_DFFE_PP__2055  (.L_HI(net2055));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][0]$_DFFE_PP__2056  (.L_HI(net2056));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][10]$_DFFE_PP__2057  (.L_HI(net2057));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][11]$_DFFE_PP__2058  (.L_HI(net2058));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][1]$_DFFE_PP__2059  (.L_HI(net2059));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][2]$_DFFE_PP__2060  (.L_HI(net2060));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][3]$_DFFE_PP__2061  (.L_HI(net2061));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][4]$_DFFE_PP__2062  (.L_HI(net2062));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][5]$_DFFE_PP__2063  (.L_HI(net2063));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][6]$_DFFE_PP__2064  (.L_HI(net2064));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][7]$_DFFE_PP__2065  (.L_HI(net2065));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][8]$_DFFE_PP__2066  (.L_HI(net2066));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][9]$_DFFE_PP__2067  (.L_HI(net2067));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][0]$_DFFE_PP__2068  (.L_HI(net2068));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][10]$_DFFE_PP__2069  (.L_HI(net2069));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][11]$_DFFE_PP__2070  (.L_HI(net2070));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][1]$_DFFE_PP__2071  (.L_HI(net2071));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][2]$_DFFE_PP__2072  (.L_HI(net2072));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][3]$_DFFE_PP__2073  (.L_HI(net2073));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][4]$_DFFE_PP__2074  (.L_HI(net2074));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][5]$_DFFE_PP__2075  (.L_HI(net2075));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][6]$_DFFE_PP__2076  (.L_HI(net2076));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][7]$_DFFE_PP__2077  (.L_HI(net2077));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][8]$_DFFE_PP__2078  (.L_HI(net2078));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][9]$_DFFE_PP__2079  (.L_HI(net2079));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][0]$_DFFE_PP__2080  (.L_HI(net2080));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][10]$_DFFE_PP__2081  (.L_HI(net2081));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][11]$_DFFE_PP__2082  (.L_HI(net2082));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][1]$_DFFE_PP__2083  (.L_HI(net2083));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][2]$_DFFE_PP__2084  (.L_HI(net2084));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][3]$_DFFE_PP__2085  (.L_HI(net2085));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][4]$_DFFE_PP__2086  (.L_HI(net2086));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][5]$_DFFE_PP__2087  (.L_HI(net2087));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][6]$_DFFE_PP__2088  (.L_HI(net2088));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][7]$_DFFE_PP__2089  (.L_HI(net2089));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][8]$_DFFE_PP__2090  (.L_HI(net2090));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][9]$_DFFE_PP__2091  (.L_HI(net2091));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][0]$_DFFE_PP__2092  (.L_HI(net2092));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][10]$_DFFE_PP__2093  (.L_HI(net2093));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][11]$_DFFE_PP__2094  (.L_HI(net2094));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][1]$_DFFE_PP__2095  (.L_HI(net2095));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][2]$_DFFE_PP__2096  (.L_HI(net2096));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][3]$_DFFE_PP__2097  (.L_HI(net2097));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][4]$_DFFE_PP__2098  (.L_HI(net2098));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][5]$_DFFE_PP__2099  (.L_HI(net2099));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][6]$_DFFE_PP__2100  (.L_HI(net2100));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][7]$_DFFE_PP__2101  (.L_HI(net2101));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][8]$_DFFE_PP__2102  (.L_HI(net2102));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][9]$_DFFE_PP__2103  (.L_HI(net2103));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][0]$_DFFE_PP__2104  (.L_HI(net2104));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][10]$_DFFE_PP__2105  (.L_HI(net2105));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][11]$_DFFE_PP__2106  (.L_HI(net2106));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][1]$_DFFE_PP__2107  (.L_HI(net2107));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][2]$_DFFE_PP__2108  (.L_HI(net2108));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][3]$_DFFE_PP__2109  (.L_HI(net2109));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][4]$_DFFE_PP__2110  (.L_HI(net2110));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][5]$_DFFE_PP__2111  (.L_HI(net2111));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][6]$_DFFE_PP__2112  (.L_HI(net2112));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][7]$_DFFE_PP__2113  (.L_HI(net2113));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][8]$_DFFE_PP__2114  (.L_HI(net2114));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][9]$_DFFE_PP__2115  (.L_HI(net2115));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][0]$_DFFE_PP__2116  (.L_HI(net2116));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][10]$_DFFE_PP__2117  (.L_HI(net2117));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][11]$_DFFE_PP__2118  (.L_HI(net2118));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][1]$_DFFE_PP__2119  (.L_HI(net2119));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][2]$_DFFE_PP__2120  (.L_HI(net2120));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][3]$_DFFE_PP__2121  (.L_HI(net2121));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][4]$_DFFE_PP__2122  (.L_HI(net2122));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][5]$_DFFE_PP__2123  (.L_HI(net2123));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][6]$_DFFE_PP__2124  (.L_HI(net2124));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][7]$_DFFE_PP__2125  (.L_HI(net2125));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][8]$_DFFE_PP__2126  (.L_HI(net2126));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][9]$_DFFE_PP__2127  (.L_HI(net2127));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][0]$_DFFE_PP__2128  (.L_HI(net2128));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][10]$_DFFE_PP__2129  (.L_HI(net2129));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][11]$_DFFE_PP__2130  (.L_HI(net2130));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][1]$_DFFE_PP__2131  (.L_HI(net2131));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][2]$_DFFE_PP__2132  (.L_HI(net2132));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][3]$_DFFE_PP__2133  (.L_HI(net2133));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][4]$_DFFE_PP__2134  (.L_HI(net2134));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][5]$_DFFE_PP__2135  (.L_HI(net2135));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][6]$_DFFE_PP__2136  (.L_HI(net2136));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][7]$_DFFE_PP__2137  (.L_HI(net2137));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][8]$_DFFE_PP__2138  (.L_HI(net2138));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][9]$_DFFE_PP__2139  (.L_HI(net2139));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][0]$_DFFE_PP__2140  (.L_HI(net2140));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][10]$_DFFE_PP__2141  (.L_HI(net2141));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][11]$_DFFE_PP__2142  (.L_HI(net2142));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][1]$_DFFE_PP__2143  (.L_HI(net2143));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][2]$_DFFE_PP__2144  (.L_HI(net2144));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][3]$_DFFE_PP__2145  (.L_HI(net2145));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][4]$_DFFE_PP__2146  (.L_HI(net2146));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][5]$_DFFE_PP__2147  (.L_HI(net2147));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][6]$_DFFE_PP__2148  (.L_HI(net2148));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][7]$_DFFE_PP__2149  (.L_HI(net2149));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][8]$_DFFE_PP__2150  (.L_HI(net2150));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][9]$_DFFE_PP__2151  (.L_HI(net2151));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][0]$_DFFE_PP__2152  (.L_HI(net2152));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][10]$_DFFE_PP__2153  (.L_HI(net2153));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][11]$_DFFE_PP__2154  (.L_HI(net2154));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][1]$_DFFE_PP__2155  (.L_HI(net2155));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][2]$_DFFE_PP__2156  (.L_HI(net2156));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][3]$_DFFE_PP__2157  (.L_HI(net2157));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][4]$_DFFE_PP__2158  (.L_HI(net2158));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][5]$_DFFE_PP__2159  (.L_HI(net2159));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][6]$_DFFE_PP__2160  (.L_HI(net2160));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][7]$_DFFE_PP__2161  (.L_HI(net2161));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][8]$_DFFE_PP__2162  (.L_HI(net2162));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][9]$_DFFE_PP__2163  (.L_HI(net2163));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][0]$_DFFE_PP__2164  (.L_HI(net2164));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][10]$_DFFE_PP__2165  (.L_HI(net2165));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][11]$_DFFE_PP__2166  (.L_HI(net2166));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][1]$_DFFE_PP__2167  (.L_HI(net2167));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][2]$_DFFE_PP__2168  (.L_HI(net2168));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][3]$_DFFE_PP__2169  (.L_HI(net2169));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][4]$_DFFE_PP__2170  (.L_HI(net2170));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][5]$_DFFE_PP__2171  (.L_HI(net2171));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][6]$_DFFE_PP__2172  (.L_HI(net2172));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][7]$_DFFE_PP__2173  (.L_HI(net2173));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][8]$_DFFE_PP__2174  (.L_HI(net2174));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][9]$_DFFE_PP__2175  (.L_HI(net2175));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][0]$_DFFE_PP__2176  (.L_HI(net2176));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][10]$_DFFE_PP__2177  (.L_HI(net2177));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][11]$_DFFE_PP__2178  (.L_HI(net2178));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][1]$_DFFE_PP__2179  (.L_HI(net2179));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][2]$_DFFE_PP__2180  (.L_HI(net2180));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][3]$_DFFE_PP__2181  (.L_HI(net2181));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][4]$_DFFE_PP__2182  (.L_HI(net2182));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][5]$_DFFE_PP__2183  (.L_HI(net2183));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][6]$_DFFE_PP__2184  (.L_HI(net2184));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][7]$_DFFE_PP__2185  (.L_HI(net2185));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][8]$_DFFE_PP__2186  (.L_HI(net2186));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][9]$_DFFE_PP__2187  (.L_HI(net2187));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][0]$_DFFE_PP__2188  (.L_HI(net2188));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][10]$_DFFE_PP__2189  (.L_HI(net2189));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][11]$_DFFE_PP__2190  (.L_HI(net2190));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][1]$_DFFE_PP__2191  (.L_HI(net2191));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][2]$_DFFE_PP__2192  (.L_HI(net2192));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][3]$_DFFE_PP__2193  (.L_HI(net2193));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][4]$_DFFE_PP__2194  (.L_HI(net2194));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][5]$_DFFE_PP__2195  (.L_HI(net2195));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][6]$_DFFE_PP__2196  (.L_HI(net2196));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][7]$_DFFE_PP__2197  (.L_HI(net2197));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][8]$_DFFE_PP__2198  (.L_HI(net2198));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][9]$_DFFE_PP__2199  (.L_HI(net2199));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][0]$_DFFE_PP__2200  (.L_HI(net2200));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][10]$_DFFE_PP__2201  (.L_HI(net2201));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][11]$_DFFE_PP__2202  (.L_HI(net2202));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][1]$_DFFE_PP__2203  (.L_HI(net2203));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][2]$_DFFE_PP__2204  (.L_HI(net2204));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][3]$_DFFE_PP__2205  (.L_HI(net2205));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][4]$_DFFE_PP__2206  (.L_HI(net2206));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][5]$_DFFE_PP__2207  (.L_HI(net2207));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][6]$_DFFE_PP__2208  (.L_HI(net2208));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][7]$_DFFE_PP__2209  (.L_HI(net2209));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][8]$_DFFE_PP__2210  (.L_HI(net2210));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][9]$_DFFE_PP__2211  (.L_HI(net2211));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][0]$_DFFE_PP__2212  (.L_HI(net2212));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][10]$_DFFE_PP__2213  (.L_HI(net2213));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][11]$_DFFE_PP__2214  (.L_HI(net2214));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][1]$_DFFE_PP__2215  (.L_HI(net2215));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][2]$_DFFE_PP__2216  (.L_HI(net2216));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][3]$_DFFE_PP__2217  (.L_HI(net2217));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][4]$_DFFE_PP__2218  (.L_HI(net2218));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][5]$_DFFE_PP__2219  (.L_HI(net2219));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][6]$_DFFE_PP__2220  (.L_HI(net2220));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][7]$_DFFE_PP__2221  (.L_HI(net2221));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][8]$_DFFE_PP__2222  (.L_HI(net2222));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][9]$_DFFE_PP__2223  (.L_HI(net2223));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][0]$_DFFE_PP__2224  (.L_HI(net2224));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][10]$_DFFE_PP__2225  (.L_HI(net2225));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][11]$_DFFE_PP__2226  (.L_HI(net2226));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][1]$_DFFE_PP__2227  (.L_HI(net2227));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][2]$_DFFE_PP__2228  (.L_HI(net2228));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][3]$_DFFE_PP__2229  (.L_HI(net2229));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][4]$_DFFE_PP__2230  (.L_HI(net2230));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][5]$_DFFE_PP__2231  (.L_HI(net2231));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][6]$_DFFE_PP__2232  (.L_HI(net2232));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][7]$_DFFE_PP__2233  (.L_HI(net2233));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][8]$_DFFE_PP__2234  (.L_HI(net2234));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][9]$_DFFE_PP__2235  (.L_HI(net2235));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][0]$_DFFE_PP__2236  (.L_HI(net2236));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][10]$_DFFE_PP__2237  (.L_HI(net2237));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][11]$_DFFE_PP__2238  (.L_HI(net2238));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][1]$_DFFE_PP__2239  (.L_HI(net2239));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][2]$_DFFE_PP__2240  (.L_HI(net2240));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][3]$_DFFE_PP__2241  (.L_HI(net2241));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][4]$_DFFE_PP__2242  (.L_HI(net2242));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][5]$_DFFE_PP__2243  (.L_HI(net2243));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][6]$_DFFE_PP__2244  (.L_HI(net2244));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][7]$_DFFE_PP__2245  (.L_HI(net2245));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][8]$_DFFE_PP__2246  (.L_HI(net2246));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][9]$_DFFE_PP__2247  (.L_HI(net2247));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][0]$_DFFE_PP__2248  (.L_HI(net2248));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][10]$_DFFE_PP__2249  (.L_HI(net2249));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][11]$_DFFE_PP__2250  (.L_HI(net2250));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][1]$_DFFE_PP__2251  (.L_HI(net2251));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][2]$_DFFE_PP__2252  (.L_HI(net2252));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][3]$_DFFE_PP__2253  (.L_HI(net2253));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][4]$_DFFE_PP__2254  (.L_HI(net2254));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][5]$_DFFE_PP__2255  (.L_HI(net2255));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][6]$_DFFE_PP__2256  (.L_HI(net2256));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][7]$_DFFE_PP__2257  (.L_HI(net2257));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][8]$_DFFE_PP__2258  (.L_HI(net2258));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][9]$_DFFE_PP__2259  (.L_HI(net2259));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][0]$_DFFE_PP__2260  (.L_HI(net2260));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][10]$_DFFE_PP__2261  (.L_HI(net2261));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][11]$_DFFE_PP__2262  (.L_HI(net2262));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][1]$_DFFE_PP__2263  (.L_HI(net2263));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][2]$_DFFE_PP__2264  (.L_HI(net2264));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][3]$_DFFE_PP__2265  (.L_HI(net2265));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][4]$_DFFE_PP__2266  (.L_HI(net2266));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][5]$_DFFE_PP__2267  (.L_HI(net2267));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][6]$_DFFE_PP__2268  (.L_HI(net2268));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][7]$_DFFE_PP__2269  (.L_HI(net2269));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][8]$_DFFE_PP__2270  (.L_HI(net2270));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][9]$_DFFE_PP__2271  (.L_HI(net2271));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][0]$_DFFE_PP__2272  (.L_HI(net2272));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][10]$_DFFE_PP__2273  (.L_HI(net2273));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][11]$_DFFE_PP__2274  (.L_HI(net2274));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][1]$_DFFE_PP__2275  (.L_HI(net2275));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][2]$_DFFE_PP__2276  (.L_HI(net2276));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][3]$_DFFE_PP__2277  (.L_HI(net2277));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][4]$_DFFE_PP__2278  (.L_HI(net2278));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][5]$_DFFE_PP__2279  (.L_HI(net2279));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][6]$_DFFE_PP__2280  (.L_HI(net2280));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][7]$_DFFE_PP__2281  (.L_HI(net2281));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][8]$_DFFE_PP__2282  (.L_HI(net2282));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][9]$_DFFE_PP__2283  (.L_HI(net2283));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][0]$_DFFE_PP__2284  (.L_HI(net2284));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][10]$_DFFE_PP__2285  (.L_HI(net2285));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][11]$_DFFE_PP__2286  (.L_HI(net2286));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][1]$_DFFE_PP__2287  (.L_HI(net2287));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][2]$_DFFE_PP__2288  (.L_HI(net2288));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][3]$_DFFE_PP__2289  (.L_HI(net2289));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][4]$_DFFE_PP__2290  (.L_HI(net2290));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][5]$_DFFE_PP__2291  (.L_HI(net2291));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][6]$_DFFE_PP__2292  (.L_HI(net2292));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][7]$_DFFE_PP__2293  (.L_HI(net2293));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][8]$_DFFE_PP__2294  (.L_HI(net2294));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][9]$_DFFE_PP__2295  (.L_HI(net2295));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][0]$_DFFE_PP__2296  (.L_HI(net2296));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][10]$_DFFE_PP__2297  (.L_HI(net2297));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][11]$_DFFE_PP__2298  (.L_HI(net2298));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][1]$_DFFE_PP__2299  (.L_HI(net2299));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][2]$_DFFE_PP__2300  (.L_HI(net2300));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][3]$_DFFE_PP__2301  (.L_HI(net2301));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][4]$_DFFE_PP__2302  (.L_HI(net2302));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][5]$_DFFE_PP__2303  (.L_HI(net2303));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][6]$_DFFE_PP__2304  (.L_HI(net2304));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][7]$_DFFE_PP__2305  (.L_HI(net2305));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][8]$_DFFE_PP__2306  (.L_HI(net2306));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][9]$_DFFE_PP__2307  (.L_HI(net2307));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][0]$_DFFE_PP__2308  (.L_HI(net2308));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][10]$_DFFE_PP__2309  (.L_HI(net2309));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][11]$_DFFE_PP__2310  (.L_HI(net2310));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][1]$_DFFE_PP__2311  (.L_HI(net2311));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][2]$_DFFE_PP__2312  (.L_HI(net2312));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][3]$_DFFE_PP__2313  (.L_HI(net2313));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][4]$_DFFE_PP__2314  (.L_HI(net2314));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][5]$_DFFE_PP__2315  (.L_HI(net2315));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][6]$_DFFE_PP__2316  (.L_HI(net2316));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][7]$_DFFE_PP__2317  (.L_HI(net2317));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][8]$_DFFE_PP__2318  (.L_HI(net2318));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][9]$_DFFE_PP__2319  (.L_HI(net2319));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][0]$_DFFE_PP__2320  (.L_HI(net2320));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][10]$_DFFE_PP__2321  (.L_HI(net2321));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][11]$_DFFE_PP__2322  (.L_HI(net2322));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][1]$_DFFE_PP__2323  (.L_HI(net2323));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][2]$_DFFE_PP__2324  (.L_HI(net2324));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][3]$_DFFE_PP__2325  (.L_HI(net2325));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][4]$_DFFE_PP__2326  (.L_HI(net2326));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][5]$_DFFE_PP__2327  (.L_HI(net2327));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][6]$_DFFE_PP__2328  (.L_HI(net2328));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][7]$_DFFE_PP__2329  (.L_HI(net2329));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][8]$_DFFE_PP__2330  (.L_HI(net2330));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][9]$_DFFE_PP__2331  (.L_HI(net2331));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][0]$_DFFE_PP__2332  (.L_HI(net2332));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][10]$_DFFE_PP__2333  (.L_HI(net2333));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][11]$_DFFE_PP__2334  (.L_HI(net2334));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][1]$_DFFE_PP__2335  (.L_HI(net2335));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][2]$_DFFE_PP__2336  (.L_HI(net2336));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][3]$_DFFE_PP__2337  (.L_HI(net2337));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][4]$_DFFE_PP__2338  (.L_HI(net2338));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][5]$_DFFE_PP__2339  (.L_HI(net2339));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][6]$_DFFE_PP__2340  (.L_HI(net2340));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][7]$_DFFE_PP__2341  (.L_HI(net2341));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][8]$_DFFE_PP__2342  (.L_HI(net2342));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][9]$_DFFE_PP__2343  (.L_HI(net2343));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][0]$_DFFE_PP__2344  (.L_HI(net2344));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][10]$_DFFE_PP__2345  (.L_HI(net2345));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][11]$_DFFE_PP__2346  (.L_HI(net2346));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][1]$_DFFE_PP__2347  (.L_HI(net2347));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][2]$_DFFE_PP__2348  (.L_HI(net2348));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][3]$_DFFE_PP__2349  (.L_HI(net2349));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][4]$_DFFE_PP__2350  (.L_HI(net2350));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][5]$_DFFE_PP__2351  (.L_HI(net2351));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][6]$_DFFE_PP__2352  (.L_HI(net2352));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][7]$_DFFE_PP__2353  (.L_HI(net2353));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][8]$_DFFE_PP__2354  (.L_HI(net2354));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][9]$_DFFE_PP__2355  (.L_HI(net2355));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][0]$_DFFE_PP__2356  (.L_HI(net2356));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][10]$_DFFE_PP__2357  (.L_HI(net2357));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][11]$_DFFE_PP__2358  (.L_HI(net2358));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][1]$_DFFE_PP__2359  (.L_HI(net2359));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][2]$_DFFE_PP__2360  (.L_HI(net2360));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][3]$_DFFE_PP__2361  (.L_HI(net2361));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][4]$_DFFE_PP__2362  (.L_HI(net2362));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][5]$_DFFE_PP__2363  (.L_HI(net2363));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][6]$_DFFE_PP__2364  (.L_HI(net2364));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][7]$_DFFE_PP__2365  (.L_HI(net2365));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][8]$_DFFE_PP__2366  (.L_HI(net2366));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][9]$_DFFE_PP__2367  (.L_HI(net2367));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][0]$_DFFE_PP__2368  (.L_HI(net2368));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][10]$_DFFE_PP__2369  (.L_HI(net2369));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][11]$_DFFE_PP__2370  (.L_HI(net2370));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][1]$_DFFE_PP__2371  (.L_HI(net2371));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][2]$_DFFE_PP__2372  (.L_HI(net2372));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][3]$_DFFE_PP__2373  (.L_HI(net2373));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][4]$_DFFE_PP__2374  (.L_HI(net2374));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][5]$_DFFE_PP__2375  (.L_HI(net2375));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][6]$_DFFE_PP__2376  (.L_HI(net2376));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][7]$_DFFE_PP__2377  (.L_HI(net2377));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][8]$_DFFE_PP__2378  (.L_HI(net2378));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][9]$_DFFE_PP__2379  (.L_HI(net2379));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][0]$_DFFE_PP__2380  (.L_HI(net2380));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][10]$_DFFE_PP__2381  (.L_HI(net2381));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][11]$_DFFE_PP__2382  (.L_HI(net2382));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][1]$_DFFE_PP__2383  (.L_HI(net2383));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][2]$_DFFE_PP__2384  (.L_HI(net2384));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][3]$_DFFE_PP__2385  (.L_HI(net2385));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][4]$_DFFE_PP__2386  (.L_HI(net2386));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][5]$_DFFE_PP__2387  (.L_HI(net2387));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][6]$_DFFE_PP__2388  (.L_HI(net2388));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][7]$_DFFE_PP__2389  (.L_HI(net2389));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][8]$_DFFE_PP__2390  (.L_HI(net2390));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][9]$_DFFE_PP__2391  (.L_HI(net2391));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][0]$_DFFE_PP__2392  (.L_HI(net2392));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][10]$_DFFE_PP__2393  (.L_HI(net2393));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][11]$_DFFE_PP__2394  (.L_HI(net2394));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][1]$_DFFE_PP__2395  (.L_HI(net2395));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][2]$_DFFE_PP__2396  (.L_HI(net2396));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][3]$_DFFE_PP__2397  (.L_HI(net2397));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][4]$_DFFE_PP__2398  (.L_HI(net2398));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][5]$_DFFE_PP__2399  (.L_HI(net2399));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][6]$_DFFE_PP__2400  (.L_HI(net2400));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][7]$_DFFE_PP__2401  (.L_HI(net2401));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][8]$_DFFE_PP__2402  (.L_HI(net2402));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][9]$_DFFE_PP__2403  (.L_HI(net2403));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][0]$_DFFE_PP__2404  (.L_HI(net2404));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][10]$_DFFE_PP__2405  (.L_HI(net2405));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][11]$_DFFE_PP__2406  (.L_HI(net2406));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][1]$_DFFE_PP__2407  (.L_HI(net2407));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][2]$_DFFE_PP__2408  (.L_HI(net2408));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][3]$_DFFE_PP__2409  (.L_HI(net2409));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][4]$_DFFE_PP__2410  (.L_HI(net2410));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][5]$_DFFE_PP__2411  (.L_HI(net2411));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][6]$_DFFE_PP__2412  (.L_HI(net2412));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][7]$_DFFE_PP__2413  (.L_HI(net2413));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][8]$_DFFE_PP__2414  (.L_HI(net2414));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][9]$_DFFE_PP__2415  (.L_HI(net2415));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][0]$_DFFE_PP__2416  (.L_HI(net2416));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][10]$_DFFE_PP__2417  (.L_HI(net2417));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][11]$_DFFE_PP__2418  (.L_HI(net2418));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][1]$_DFFE_PP__2419  (.L_HI(net2419));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][2]$_DFFE_PP__2420  (.L_HI(net2420));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][3]$_DFFE_PP__2421  (.L_HI(net2421));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][4]$_DFFE_PP__2422  (.L_HI(net2422));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][5]$_DFFE_PP__2423  (.L_HI(net2423));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][6]$_DFFE_PP__2424  (.L_HI(net2424));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][7]$_DFFE_PP__2425  (.L_HI(net2425));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][8]$_DFFE_PP__2426  (.L_HI(net2426));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][9]$_DFFE_PP__2427  (.L_HI(net2427));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][0]$_DFFE_PP__2428  (.L_HI(net2428));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][10]$_DFFE_PP__2429  (.L_HI(net2429));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][11]$_DFFE_PP__2430  (.L_HI(net2430));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][1]$_DFFE_PP__2431  (.L_HI(net2431));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][2]$_DFFE_PP__2432  (.L_HI(net2432));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][3]$_DFFE_PP__2433  (.L_HI(net2433));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][4]$_DFFE_PP__2434  (.L_HI(net2434));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][5]$_DFFE_PP__2435  (.L_HI(net2435));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][6]$_DFFE_PP__2436  (.L_HI(net2436));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][7]$_DFFE_PP__2437  (.L_HI(net2437));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][8]$_DFFE_PP__2438  (.L_HI(net2438));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][9]$_DFFE_PP__2439  (.L_HI(net2439));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][0]$_DFFE_PP__2440  (.L_HI(net2440));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][10]$_DFFE_PP__2441  (.L_HI(net2441));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][11]$_DFFE_PP__2442  (.L_HI(net2442));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][1]$_DFFE_PP__2443  (.L_HI(net2443));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][2]$_DFFE_PP__2444  (.L_HI(net2444));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][3]$_DFFE_PP__2445  (.L_HI(net2445));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][4]$_DFFE_PP__2446  (.L_HI(net2446));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][5]$_DFFE_PP__2447  (.L_HI(net2447));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][6]$_DFFE_PP__2448  (.L_HI(net2448));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][7]$_DFFE_PP__2449  (.L_HI(net2449));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][8]$_DFFE_PP__2450  (.L_HI(net2450));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][9]$_DFFE_PP__2451  (.L_HI(net2451));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][0]$_DFFE_PP__2452  (.L_HI(net2452));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][10]$_DFFE_PP__2453  (.L_HI(net2453));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][11]$_DFFE_PP__2454  (.L_HI(net2454));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][1]$_DFFE_PP__2455  (.L_HI(net2455));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][2]$_DFFE_PP__2456  (.L_HI(net2456));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][3]$_DFFE_PP__2457  (.L_HI(net2457));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][4]$_DFFE_PP__2458  (.L_HI(net2458));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][5]$_DFFE_PP__2459  (.L_HI(net2459));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][6]$_DFFE_PP__2460  (.L_HI(net2460));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][7]$_DFFE_PP__2461  (.L_HI(net2461));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][8]$_DFFE_PP__2462  (.L_HI(net2462));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][9]$_DFFE_PP__2463  (.L_HI(net2463));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][0]$_DFFE_PP__2464  (.L_HI(net2464));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][10]$_DFFE_PP__2465  (.L_HI(net2465));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][11]$_DFFE_PP__2466  (.L_HI(net2466));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][1]$_DFFE_PP__2467  (.L_HI(net2467));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][2]$_DFFE_PP__2468  (.L_HI(net2468));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][3]$_DFFE_PP__2469  (.L_HI(net2469));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][4]$_DFFE_PP__2470  (.L_HI(net2470));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][5]$_DFFE_PP__2471  (.L_HI(net2471));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][6]$_DFFE_PP__2472  (.L_HI(net2472));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][7]$_DFFE_PP__2473  (.L_HI(net2473));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][8]$_DFFE_PP__2474  (.L_HI(net2474));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][9]$_DFFE_PP__2475  (.L_HI(net2475));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][0]$_DFFE_PP__2476  (.L_HI(net2476));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][10]$_DFFE_PP__2477  (.L_HI(net2477));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][11]$_DFFE_PP__2478  (.L_HI(net2478));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][1]$_DFFE_PP__2479  (.L_HI(net2479));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][2]$_DFFE_PP__2480  (.L_HI(net2480));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][3]$_DFFE_PP__2481  (.L_HI(net2481));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][4]$_DFFE_PP__2482  (.L_HI(net2482));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][5]$_DFFE_PP__2483  (.L_HI(net2483));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][6]$_DFFE_PP__2484  (.L_HI(net2484));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][7]$_DFFE_PP__2485  (.L_HI(net2485));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][8]$_DFFE_PP__2486  (.L_HI(net2486));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][9]$_DFFE_PP__2487  (.L_HI(net2487));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][0]$_DFFE_PP__2488  (.L_HI(net2488));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][10]$_DFFE_PP__2489  (.L_HI(net2489));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][11]$_DFFE_PP__2490  (.L_HI(net2490));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][1]$_DFFE_PP__2491  (.L_HI(net2491));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][2]$_DFFE_PP__2492  (.L_HI(net2492));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][3]$_DFFE_PP__2493  (.L_HI(net2493));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][4]$_DFFE_PP__2494  (.L_HI(net2494));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][5]$_DFFE_PP__2495  (.L_HI(net2495));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][6]$_DFFE_PP__2496  (.L_HI(net2496));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][7]$_DFFE_PP__2497  (.L_HI(net2497));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][8]$_DFFE_PP__2498  (.L_HI(net2498));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][9]$_DFFE_PP__2499  (.L_HI(net2499));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][0]$_DFFE_PP__2500  (.L_HI(net2500));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][10]$_DFFE_PP__2501  (.L_HI(net2501));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][11]$_DFFE_PP__2502  (.L_HI(net2502));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][1]$_DFFE_PP__2503  (.L_HI(net2503));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][2]$_DFFE_PP__2504  (.L_HI(net2504));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][3]$_DFFE_PP__2505  (.L_HI(net2505));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][4]$_DFFE_PP__2506  (.L_HI(net2506));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][5]$_DFFE_PP__2507  (.L_HI(net2507));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][6]$_DFFE_PP__2508  (.L_HI(net2508));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][7]$_DFFE_PP__2509  (.L_HI(net2509));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][8]$_DFFE_PP__2510  (.L_HI(net2510));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][9]$_DFFE_PP__2511  (.L_HI(net2511));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][0]$_DFFE_PP__2512  (.L_HI(net2512));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][10]$_DFFE_PP__2513  (.L_HI(net2513));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][11]$_DFFE_PP__2514  (.L_HI(net2514));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][1]$_DFFE_PP__2515  (.L_HI(net2515));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][2]$_DFFE_PP__2516  (.L_HI(net2516));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][3]$_DFFE_PP__2517  (.L_HI(net2517));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][4]$_DFFE_PP__2518  (.L_HI(net2518));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][5]$_DFFE_PP__2519  (.L_HI(net2519));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][6]$_DFFE_PP__2520  (.L_HI(net2520));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][7]$_DFFE_PP__2521  (.L_HI(net2521));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][8]$_DFFE_PP__2522  (.L_HI(net2522));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][9]$_DFFE_PP__2523  (.L_HI(net2523));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][0]$_DFFE_PP__2524  (.L_HI(net2524));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][10]$_DFFE_PP__2525  (.L_HI(net2525));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][11]$_DFFE_PP__2526  (.L_HI(net2526));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][1]$_DFFE_PP__2527  (.L_HI(net2527));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][2]$_DFFE_PP__2528  (.L_HI(net2528));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][3]$_DFFE_PP__2529  (.L_HI(net2529));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][4]$_DFFE_PP__2530  (.L_HI(net2530));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][5]$_DFFE_PP__2531  (.L_HI(net2531));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][6]$_DFFE_PP__2532  (.L_HI(net2532));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][7]$_DFFE_PP__2533  (.L_HI(net2533));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][8]$_DFFE_PP__2534  (.L_HI(net2534));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][9]$_DFFE_PP__2535  (.L_HI(net2535));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][0]$_DFFE_PP__2536  (.L_HI(net2536));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][10]$_DFFE_PP__2537  (.L_HI(net2537));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][11]$_DFFE_PP__2538  (.L_HI(net2538));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][1]$_DFFE_PP__2539  (.L_HI(net2539));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][2]$_DFFE_PP__2540  (.L_HI(net2540));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][3]$_DFFE_PP__2541  (.L_HI(net2541));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][4]$_DFFE_PP__2542  (.L_HI(net2542));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][5]$_DFFE_PP__2543  (.L_HI(net2543));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][6]$_DFFE_PP__2544  (.L_HI(net2544));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][7]$_DFFE_PP__2545  (.L_HI(net2545));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][8]$_DFFE_PP__2546  (.L_HI(net2546));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][9]$_DFFE_PP__2547  (.L_HI(net2547));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][0]$_DFFE_PP__2548  (.L_HI(net2548));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][10]$_DFFE_PP__2549  (.L_HI(net2549));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][11]$_DFFE_PP__2550  (.L_HI(net2550));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][1]$_DFFE_PP__2551  (.L_HI(net2551));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][2]$_DFFE_PP__2552  (.L_HI(net2552));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][3]$_DFFE_PP__2553  (.L_HI(net2553));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][4]$_DFFE_PP__2554  (.L_HI(net2554));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][5]$_DFFE_PP__2555  (.L_HI(net2555));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][6]$_DFFE_PP__2556  (.L_HI(net2556));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][7]$_DFFE_PP__2557  (.L_HI(net2557));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][8]$_DFFE_PP__2558  (.L_HI(net2558));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][9]$_DFFE_PP__2559  (.L_HI(net2559));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][0]$_DFFE_PP__2560  (.L_HI(net2560));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][10]$_DFFE_PP__2561  (.L_HI(net2561));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][11]$_DFFE_PP__2562  (.L_HI(net2562));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][1]$_DFFE_PP__2563  (.L_HI(net2563));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][2]$_DFFE_PP__2564  (.L_HI(net2564));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][3]$_DFFE_PP__2565  (.L_HI(net2565));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][4]$_DFFE_PP__2566  (.L_HI(net2566));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][5]$_DFFE_PP__2567  (.L_HI(net2567));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][6]$_DFFE_PP__2568  (.L_HI(net2568));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][7]$_DFFE_PP__2569  (.L_HI(net2569));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][8]$_DFFE_PP__2570  (.L_HI(net2570));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][9]$_DFFE_PP__2571  (.L_HI(net2571));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][0]$_DFFE_PP__2572  (.L_HI(net2572));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][10]$_DFFE_PP__2573  (.L_HI(net2573));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][11]$_DFFE_PP__2574  (.L_HI(net2574));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][1]$_DFFE_PP__2575  (.L_HI(net2575));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][2]$_DFFE_PP__2576  (.L_HI(net2576));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][3]$_DFFE_PP__2577  (.L_HI(net2577));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][4]$_DFFE_PP__2578  (.L_HI(net2578));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][5]$_DFFE_PP__2579  (.L_HI(net2579));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][6]$_DFFE_PP__2580  (.L_HI(net2580));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][7]$_DFFE_PP__2581  (.L_HI(net2581));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][8]$_DFFE_PP__2582  (.L_HI(net2582));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][9]$_DFFE_PP__2583  (.L_HI(net2583));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][0]$_DFFE_PP__2584  (.L_HI(net2584));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][10]$_DFFE_PP__2585  (.L_HI(net2585));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][11]$_DFFE_PP__2586  (.L_HI(net2586));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][1]$_DFFE_PP__2587  (.L_HI(net2587));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][2]$_DFFE_PP__2588  (.L_HI(net2588));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][3]$_DFFE_PP__2589  (.L_HI(net2589));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][4]$_DFFE_PP__2590  (.L_HI(net2590));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][5]$_DFFE_PP__2591  (.L_HI(net2591));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][6]$_DFFE_PP__2592  (.L_HI(net2592));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][7]$_DFFE_PP__2593  (.L_HI(net2593));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][8]$_DFFE_PP__2594  (.L_HI(net2594));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][9]$_DFFE_PP__2595  (.L_HI(net2595));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][0]$_DFFE_PP__2596  (.L_HI(net2596));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][10]$_DFFE_PP__2597  (.L_HI(net2597));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][11]$_DFFE_PP__2598  (.L_HI(net2598));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][1]$_DFFE_PP__2599  (.L_HI(net2599));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][2]$_DFFE_PP__2600  (.L_HI(net2600));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][3]$_DFFE_PP__2601  (.L_HI(net2601));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][4]$_DFFE_PP__2602  (.L_HI(net2602));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][5]$_DFFE_PP__2603  (.L_HI(net2603));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][6]$_DFFE_PP__2604  (.L_HI(net2604));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][7]$_DFFE_PP__2605  (.L_HI(net2605));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][8]$_DFFE_PP__2606  (.L_HI(net2606));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][9]$_DFFE_PP__2607  (.L_HI(net2607));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][0]$_DFFE_PP__2608  (.L_HI(net2608));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][10]$_DFFE_PP__2609  (.L_HI(net2609));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][11]$_DFFE_PP__2610  (.L_HI(net2610));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][1]$_DFFE_PP__2611  (.L_HI(net2611));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][2]$_DFFE_PP__2612  (.L_HI(net2612));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][3]$_DFFE_PP__2613  (.L_HI(net2613));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][4]$_DFFE_PP__2614  (.L_HI(net2614));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][5]$_DFFE_PP__2615  (.L_HI(net2615));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][6]$_DFFE_PP__2616  (.L_HI(net2616));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][7]$_DFFE_PP__2617  (.L_HI(net2617));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][8]$_DFFE_PP__2618  (.L_HI(net2618));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][9]$_DFFE_PP__2619  (.L_HI(net2619));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][0]$_DFFE_PP__2620  (.L_HI(net2620));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][10]$_DFFE_PP__2621  (.L_HI(net2621));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][11]$_DFFE_PP__2622  (.L_HI(net2622));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][1]$_DFFE_PP__2623  (.L_HI(net2623));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][2]$_DFFE_PP__2624  (.L_HI(net2624));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][3]$_DFFE_PP__2625  (.L_HI(net2625));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][4]$_DFFE_PP__2626  (.L_HI(net2626));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][5]$_DFFE_PP__2627  (.L_HI(net2627));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][6]$_DFFE_PP__2628  (.L_HI(net2628));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][7]$_DFFE_PP__2629  (.L_HI(net2629));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][8]$_DFFE_PP__2630  (.L_HI(net2630));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][9]$_DFFE_PP__2631  (.L_HI(net2631));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][0]$_DFFE_PP__2632  (.L_HI(net2632));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][10]$_DFFE_PP__2633  (.L_HI(net2633));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][11]$_DFFE_PP__2634  (.L_HI(net2634));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][1]$_DFFE_PP__2635  (.L_HI(net2635));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][2]$_DFFE_PP__2636  (.L_HI(net2636));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][3]$_DFFE_PP__2637  (.L_HI(net2637));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][4]$_DFFE_PP__2638  (.L_HI(net2638));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][5]$_DFFE_PP__2639  (.L_HI(net2639));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][6]$_DFFE_PP__2640  (.L_HI(net2640));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][7]$_DFFE_PP__2641  (.L_HI(net2641));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][8]$_DFFE_PP__2642  (.L_HI(net2642));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][9]$_DFFE_PP__2643  (.L_HI(net2643));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][0]$_DFFE_PP__2644  (.L_HI(net2644));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][10]$_DFFE_PP__2645  (.L_HI(net2645));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][11]$_DFFE_PP__2646  (.L_HI(net2646));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][1]$_DFFE_PP__2647  (.L_HI(net2647));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][2]$_DFFE_PP__2648  (.L_HI(net2648));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][3]$_DFFE_PP__2649  (.L_HI(net2649));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][4]$_DFFE_PP__2650  (.L_HI(net2650));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][5]$_DFFE_PP__2651  (.L_HI(net2651));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][6]$_DFFE_PP__2652  (.L_HI(net2652));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][7]$_DFFE_PP__2653  (.L_HI(net2653));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][8]$_DFFE_PP__2654  (.L_HI(net2654));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][9]$_DFFE_PP__2655  (.L_HI(net2655));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][0]$_DFFE_PP__2656  (.L_HI(net2656));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][10]$_DFFE_PP__2657  (.L_HI(net2657));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][11]$_DFFE_PP__2658  (.L_HI(net2658));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][1]$_DFFE_PP__2659  (.L_HI(net2659));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][2]$_DFFE_PP__2660  (.L_HI(net2660));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][3]$_DFFE_PP__2661  (.L_HI(net2661));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][4]$_DFFE_PP__2662  (.L_HI(net2662));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][5]$_DFFE_PP__2663  (.L_HI(net2663));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][6]$_DFFE_PP__2664  (.L_HI(net2664));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][7]$_DFFE_PP__2665  (.L_HI(net2665));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][8]$_DFFE_PP__2666  (.L_HI(net2666));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][9]$_DFFE_PP__2667  (.L_HI(net2667));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][0]$_DFFE_PP__2668  (.L_HI(net2668));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][10]$_DFFE_PP__2669  (.L_HI(net2669));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][11]$_DFFE_PP__2670  (.L_HI(net2670));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][1]$_DFFE_PP__2671  (.L_HI(net2671));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][2]$_DFFE_PP__2672  (.L_HI(net2672));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][3]$_DFFE_PP__2673  (.L_HI(net2673));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][4]$_DFFE_PP__2674  (.L_HI(net2674));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][5]$_DFFE_PP__2675  (.L_HI(net2675));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][6]$_DFFE_PP__2676  (.L_HI(net2676));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][7]$_DFFE_PP__2677  (.L_HI(net2677));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][8]$_DFFE_PP__2678  (.L_HI(net2678));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][9]$_DFFE_PP__2679  (.L_HI(net2679));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][0]$_DFFE_PP__2680  (.L_HI(net2680));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][10]$_DFFE_PP__2681  (.L_HI(net2681));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][11]$_DFFE_PP__2682  (.L_HI(net2682));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][1]$_DFFE_PP__2683  (.L_HI(net2683));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][2]$_DFFE_PP__2684  (.L_HI(net2684));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][3]$_DFFE_PP__2685  (.L_HI(net2685));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][4]$_DFFE_PP__2686  (.L_HI(net2686));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][5]$_DFFE_PP__2687  (.L_HI(net2687));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][6]$_DFFE_PP__2688  (.L_HI(net2688));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][7]$_DFFE_PP__2689  (.L_HI(net2689));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][8]$_DFFE_PP__2690  (.L_HI(net2690));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][9]$_DFFE_PP__2691  (.L_HI(net2691));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][0]$_DFFE_PP__2692  (.L_HI(net2692));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][10]$_DFFE_PP__2693  (.L_HI(net2693));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][11]$_DFFE_PP__2694  (.L_HI(net2694));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][1]$_DFFE_PP__2695  (.L_HI(net2695));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][2]$_DFFE_PP__2696  (.L_HI(net2696));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][3]$_DFFE_PP__2697  (.L_HI(net2697));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][4]$_DFFE_PP__2698  (.L_HI(net2698));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][5]$_DFFE_PP__2699  (.L_HI(net2699));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][6]$_DFFE_PP__2700  (.L_HI(net2700));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][7]$_DFFE_PP__2701  (.L_HI(net2701));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][8]$_DFFE_PP__2702  (.L_HI(net2702));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][9]$_DFFE_PP__2703  (.L_HI(net2703));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][0]$_DFFE_PP__2704  (.L_HI(net2704));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][10]$_DFFE_PP__2705  (.L_HI(net2705));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][11]$_DFFE_PP__2706  (.L_HI(net2706));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][1]$_DFFE_PP__2707  (.L_HI(net2707));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][2]$_DFFE_PP__2708  (.L_HI(net2708));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][3]$_DFFE_PP__2709  (.L_HI(net2709));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][4]$_DFFE_PP__2710  (.L_HI(net2710));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][5]$_DFFE_PP__2711  (.L_HI(net2711));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][6]$_DFFE_PP__2712  (.L_HI(net2712));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][7]$_DFFE_PP__2713  (.L_HI(net2713));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][8]$_DFFE_PP__2714  (.L_HI(net2714));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][9]$_DFFE_PP__2715  (.L_HI(net2715));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][0]$_DFFE_PP__2716  (.L_HI(net2716));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][10]$_DFFE_PP__2717  (.L_HI(net2717));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][11]$_DFFE_PP__2718  (.L_HI(net2718));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][1]$_DFFE_PP__2719  (.L_HI(net2719));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][2]$_DFFE_PP__2720  (.L_HI(net2720));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][3]$_DFFE_PP__2721  (.L_HI(net2721));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][4]$_DFFE_PP__2722  (.L_HI(net2722));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][5]$_DFFE_PP__2723  (.L_HI(net2723));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][6]$_DFFE_PP__2724  (.L_HI(net2724));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][7]$_DFFE_PP__2725  (.L_HI(net2725));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][8]$_DFFE_PP__2726  (.L_HI(net2726));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][9]$_DFFE_PP__2727  (.L_HI(net2727));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][0]$_DFFE_PP__2728  (.L_HI(net2728));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][10]$_DFFE_PP__2729  (.L_HI(net2729));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][11]$_DFFE_PP__2730  (.L_HI(net2730));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][1]$_DFFE_PP__2731  (.L_HI(net2731));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][2]$_DFFE_PP__2732  (.L_HI(net2732));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][3]$_DFFE_PP__2733  (.L_HI(net2733));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][4]$_DFFE_PP__2734  (.L_HI(net2734));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][5]$_DFFE_PP__2735  (.L_HI(net2735));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][6]$_DFFE_PP__2736  (.L_HI(net2736));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][7]$_DFFE_PP__2737  (.L_HI(net2737));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][8]$_DFFE_PP__2738  (.L_HI(net2738));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][9]$_DFFE_PP__2739  (.L_HI(net2739));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][0]$_DFFE_PP__2740  (.L_HI(net2740));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][10]$_DFFE_PP__2741  (.L_HI(net2741));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][11]$_DFFE_PP__2742  (.L_HI(net2742));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][1]$_DFFE_PP__2743  (.L_HI(net2743));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][2]$_DFFE_PP__2744  (.L_HI(net2744));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][3]$_DFFE_PP__2745  (.L_HI(net2745));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][4]$_DFFE_PP__2746  (.L_HI(net2746));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][5]$_DFFE_PP__2747  (.L_HI(net2747));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][6]$_DFFE_PP__2748  (.L_HI(net2748));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][7]$_DFFE_PP__2749  (.L_HI(net2749));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][8]$_DFFE_PP__2750  (.L_HI(net2750));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][9]$_DFFE_PP__2751  (.L_HI(net2751));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][0]$_DFFE_PP__2752  (.L_HI(net2752));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][10]$_DFFE_PP__2753  (.L_HI(net2753));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][11]$_DFFE_PP__2754  (.L_HI(net2754));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][1]$_DFFE_PP__2755  (.L_HI(net2755));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][2]$_DFFE_PP__2756  (.L_HI(net2756));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][3]$_DFFE_PP__2757  (.L_HI(net2757));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][4]$_DFFE_PP__2758  (.L_HI(net2758));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][5]$_DFFE_PP__2759  (.L_HI(net2759));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][6]$_DFFE_PP__2760  (.L_HI(net2760));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][7]$_DFFE_PP__2761  (.L_HI(net2761));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][8]$_DFFE_PP__2762  (.L_HI(net2762));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][9]$_DFFE_PP__2763  (.L_HI(net2763));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[0]$_DFFE_PP__2764  (.L_HI(net2764));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[10]$_DFFE_PP__2765  (.L_HI(net2765));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[11]$_DFFE_PP__2766  (.L_HI(net2766));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[12]$_DFFE_PP__2767  (.L_HI(net2767));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[13]$_DFFE_PP__2768  (.L_HI(net2768));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[14]$_DFFE_PP__2769  (.L_HI(net2769));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[15]$_DFFE_PP__2770  (.L_HI(net2770));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[16]$_DFFE_PP__2771  (.L_HI(net2771));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[17]$_DFFE_PP__2772  (.L_HI(net2772));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[18]$_DFFE_PP__2773  (.L_HI(net2773));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[19]$_DFFE_PP__2774  (.L_HI(net2774));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[1]$_DFFE_PP__2775  (.L_HI(net2775));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[20]$_DFFE_PP__2776  (.L_HI(net2776));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[21]$_DFFE_PP__2777  (.L_HI(net2777));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[22]$_DFFE_PP__2778  (.L_HI(net2778));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[23]$_DFFE_PP__2779  (.L_HI(net2779));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[24]$_DFFE_PP__2780  (.L_HI(net2780));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[25]$_DFFE_PP__2781  (.L_HI(net2781));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[26]$_DFFE_PP__2782  (.L_HI(net2782));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[27]$_DFFE_PP__2783  (.L_HI(net2783));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[28]$_DFFE_PP__2784  (.L_HI(net2784));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[29]$_DFFE_PP__2785  (.L_HI(net2785));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[2]$_DFFE_PP__2786  (.L_HI(net2786));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[30]$_DFFE_PP__2787  (.L_HI(net2787));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[31]$_DFFE_PP__2788  (.L_HI(net2788));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[3]$_DFFE_PP__2789  (.L_HI(net2789));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[4]$_DFFE_PP__2790  (.L_HI(net2790));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[5]$_DFFE_PP__2791  (.L_HI(net2791));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[6]$_DFFE_PP__2792  (.L_HI(net2792));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[7]$_DFFE_PP__2793  (.L_HI(net2793));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[8]$_DFFE_PP__2794  (.L_HI(net2794));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[9]$_DFFE_PP__2795  (.L_HI(net2795));
 sg13g2_tiehi \cpu.gpio.r_enable_in[0]$_SDFFE_PN0P__2796  (.L_HI(net2796));
 sg13g2_tiehi \cpu.gpio.r_enable_in[1]$_SDFFE_PN0P__2797  (.L_HI(net2797));
 sg13g2_tiehi \cpu.gpio.r_enable_in[2]$_SDFFE_PN0P__2798  (.L_HI(net2798));
 sg13g2_tiehi \cpu.gpio.r_enable_in[3]$_SDFFE_PN0P__2799  (.L_HI(net2799));
 sg13g2_tiehi \cpu.gpio.r_enable_in[4]$_SDFFE_PN0P__2800  (.L_HI(net2800));
 sg13g2_tiehi \cpu.gpio.r_enable_in[5]$_SDFFE_PN0P__2801  (.L_HI(net2801));
 sg13g2_tiehi \cpu.gpio.r_enable_in[6]$_SDFFE_PN0P__2802  (.L_HI(net2802));
 sg13g2_tiehi \cpu.gpio.r_enable_in[7]$_SDFFE_PN0P__2803  (.L_HI(net2803));
 sg13g2_tiehi \cpu.gpio.r_enable_io[0]$_SDFFE_PN0P__2804  (.L_HI(net2804));
 sg13g2_tiehi \cpu.gpio.r_enable_io[1]$_SDFFE_PN0P__2805  (.L_HI(net2805));
 sg13g2_tiehi \cpu.gpio.r_enable_io[2]$_SDFFE_PN0P__2806  (.L_HI(net2806));
 sg13g2_tiehi \cpu.gpio.r_enable_io[3]$_SDFFE_PN0P__2807  (.L_HI(net2807));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[0]$_SDFFE_PN0P__2808  (.L_HI(net2808));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[1]$_SDFFE_PN0P__2809  (.L_HI(net2809));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[2]$_SDFFE_PN0P__2810  (.L_HI(net2810));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[3]$_SDFFE_PN0P__2811  (.L_HI(net2811));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[0]$_DFFE_PP__2812  (.L_HI(net2812));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[1]$_DFFE_PP__2813  (.L_HI(net2813));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[2]$_DFFE_PP__2814  (.L_HI(net2814));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[3]$_DFFE_PP__2815  (.L_HI(net2815));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[0]$_DFFE_PP__2816  (.L_HI(net2816));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[1]$_DFFE_PP__2817  (.L_HI(net2817));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[2]$_DFFE_PP__2818  (.L_HI(net2818));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[3]$_DFFE_PP__2819  (.L_HI(net2819));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[4]$_DFFE_PP__2820  (.L_HI(net2820));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][0]$_DFFE_PP__2821  (.L_HI(net2821));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][1]$_DFFE_PP__2822  (.L_HI(net2822));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][2]$_DFFE_PP__2823  (.L_HI(net2823));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][3]$_DFFE_PP__2824  (.L_HI(net2824));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][0]$_DFFE_PP__2825  (.L_HI(net2825));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][1]$_DFFE_PP__2826  (.L_HI(net2826));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][2]$_DFFE_PP__2827  (.L_HI(net2827));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][3]$_DFFE_PP__2828  (.L_HI(net2828));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][0]$_DFFE_PP__2829  (.L_HI(net2829));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][1]$_DFFE_PP__2830  (.L_HI(net2830));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][2]$_DFFE_PP__2831  (.L_HI(net2831));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][3]$_DFFE_PP__2832  (.L_HI(net2832));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][0]$_DFFE_PP__2833  (.L_HI(net2833));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][1]$_DFFE_PP__2834  (.L_HI(net2834));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][2]$_DFFE_PP__2835  (.L_HI(net2835));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][3]$_DFFE_PP__2836  (.L_HI(net2836));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][0]$_DFFE_PP__2837  (.L_HI(net2837));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][1]$_DFFE_PP__2838  (.L_HI(net2838));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][2]$_DFFE_PP__2839  (.L_HI(net2839));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][3]$_DFFE_PP__2840  (.L_HI(net2840));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][0]$_DFFE_PP__2841  (.L_HI(net2841));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][1]$_DFFE_PP__2842  (.L_HI(net2842));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][2]$_DFFE_PP__2843  (.L_HI(net2843));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][3]$_DFFE_PP__2844  (.L_HI(net2844));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][0]$_DFFE_PP__2845  (.L_HI(net2845));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][1]$_DFFE_PP__2846  (.L_HI(net2846));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][2]$_DFFE_PP__2847  (.L_HI(net2847));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][3]$_DFFE_PP__2848  (.L_HI(net2848));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][0]$_DFFE_PP__2849  (.L_HI(net2849));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][1]$_DFFE_PP__2850  (.L_HI(net2850));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][2]$_DFFE_PP__2851  (.L_HI(net2851));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][3]$_DFFE_PP__2852  (.L_HI(net2852));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][0]$_DFFE_PP__2853  (.L_HI(net2853));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][1]$_DFFE_PP__2854  (.L_HI(net2854));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][2]$_DFFE_PP__2855  (.L_HI(net2855));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][3]$_DFFE_PP__2856  (.L_HI(net2856));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][0]$_SDFFE_PN1P__2857  (.L_HI(net2857));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][1]$_SDFFE_PN0P__2858  (.L_HI(net2858));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][2]$_SDFFE_PN0P__2859  (.L_HI(net2859));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][3]$_SDFFE_PN0P__2860  (.L_HI(net2860));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][0]$_DFFE_PP__2861  (.L_HI(net2861));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][1]$_DFFE_PP__2862  (.L_HI(net2862));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][2]$_DFFE_PP__2863  (.L_HI(net2863));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][3]$_DFFE_PP__2864  (.L_HI(net2864));
 sg13g2_tiehi \cpu.gpio.r_uart_rx_src[0]$_SDFFE_PN0P__2865  (.L_HI(net2865));
 sg13g2_tiehi \cpu.gpio.r_uart_rx_src[1]$_SDFFE_PN0P__2866  (.L_HI(net2866));
 sg13g2_tiehi \cpu.gpio.r_uart_rx_src[2]$_SDFFE_PN0P__2867  (.L_HI(net2867));
 sg13g2_tiehi \cpu.icache.r_data[0][0]$_DFFE_PP__2868  (.L_HI(net2868));
 sg13g2_tiehi \cpu.icache.r_data[0][10]$_DFFE_PP__2869  (.L_HI(net2869));
 sg13g2_tiehi \cpu.icache.r_data[0][11]$_DFFE_PP__2870  (.L_HI(net2870));
 sg13g2_tiehi \cpu.icache.r_data[0][12]$_DFFE_PP__2871  (.L_HI(net2871));
 sg13g2_tiehi \cpu.icache.r_data[0][13]$_DFFE_PP__2872  (.L_HI(net2872));
 sg13g2_tiehi \cpu.icache.r_data[0][14]$_DFFE_PP__2873  (.L_HI(net2873));
 sg13g2_tiehi \cpu.icache.r_data[0][15]$_DFFE_PP__2874  (.L_HI(net2874));
 sg13g2_tiehi \cpu.icache.r_data[0][16]$_DFFE_PP__2875  (.L_HI(net2875));
 sg13g2_tiehi \cpu.icache.r_data[0][17]$_DFFE_PP__2876  (.L_HI(net2876));
 sg13g2_tiehi \cpu.icache.r_data[0][18]$_DFFE_PP__2877  (.L_HI(net2877));
 sg13g2_tiehi \cpu.icache.r_data[0][19]$_DFFE_PP__2878  (.L_HI(net2878));
 sg13g2_tiehi \cpu.icache.r_data[0][1]$_DFFE_PP__2879  (.L_HI(net2879));
 sg13g2_tiehi \cpu.icache.r_data[0][20]$_DFFE_PP__2880  (.L_HI(net2880));
 sg13g2_tiehi \cpu.icache.r_data[0][21]$_DFFE_PP__2881  (.L_HI(net2881));
 sg13g2_tiehi \cpu.icache.r_data[0][22]$_DFFE_PP__2882  (.L_HI(net2882));
 sg13g2_tiehi \cpu.icache.r_data[0][23]$_DFFE_PP__2883  (.L_HI(net2883));
 sg13g2_tiehi \cpu.icache.r_data[0][24]$_DFFE_PP__2884  (.L_HI(net2884));
 sg13g2_tiehi \cpu.icache.r_data[0][25]$_DFFE_PP__2885  (.L_HI(net2885));
 sg13g2_tiehi \cpu.icache.r_data[0][26]$_DFFE_PP__2886  (.L_HI(net2886));
 sg13g2_tiehi \cpu.icache.r_data[0][27]$_DFFE_PP__2887  (.L_HI(net2887));
 sg13g2_tiehi \cpu.icache.r_data[0][28]$_DFFE_PP__2888  (.L_HI(net2888));
 sg13g2_tiehi \cpu.icache.r_data[0][29]$_DFFE_PP__2889  (.L_HI(net2889));
 sg13g2_tiehi \cpu.icache.r_data[0][2]$_DFFE_PP__2890  (.L_HI(net2890));
 sg13g2_tiehi \cpu.icache.r_data[0][30]$_DFFE_PP__2891  (.L_HI(net2891));
 sg13g2_tiehi \cpu.icache.r_data[0][31]$_DFFE_PP__2892  (.L_HI(net2892));
 sg13g2_tiehi \cpu.icache.r_data[0][3]$_DFFE_PP__2893  (.L_HI(net2893));
 sg13g2_tiehi \cpu.icache.r_data[0][4]$_DFFE_PP__2894  (.L_HI(net2894));
 sg13g2_tiehi \cpu.icache.r_data[0][5]$_DFFE_PP__2895  (.L_HI(net2895));
 sg13g2_tiehi \cpu.icache.r_data[0][6]$_DFFE_PP__2896  (.L_HI(net2896));
 sg13g2_tiehi \cpu.icache.r_data[0][7]$_DFFE_PP__2897  (.L_HI(net2897));
 sg13g2_tiehi \cpu.icache.r_data[0][8]$_DFFE_PP__2898  (.L_HI(net2898));
 sg13g2_tiehi \cpu.icache.r_data[0][9]$_DFFE_PP__2899  (.L_HI(net2899));
 sg13g2_tiehi \cpu.icache.r_data[1][0]$_DFFE_PP__2900  (.L_HI(net2900));
 sg13g2_tiehi \cpu.icache.r_data[1][10]$_DFFE_PP__2901  (.L_HI(net2901));
 sg13g2_tiehi \cpu.icache.r_data[1][11]$_DFFE_PP__2902  (.L_HI(net2902));
 sg13g2_tiehi \cpu.icache.r_data[1][12]$_DFFE_PP__2903  (.L_HI(net2903));
 sg13g2_tiehi \cpu.icache.r_data[1][13]$_DFFE_PP__2904  (.L_HI(net2904));
 sg13g2_tiehi \cpu.icache.r_data[1][14]$_DFFE_PP__2905  (.L_HI(net2905));
 sg13g2_tiehi \cpu.icache.r_data[1][15]$_DFFE_PP__2906  (.L_HI(net2906));
 sg13g2_tiehi \cpu.icache.r_data[1][16]$_DFFE_PP__2907  (.L_HI(net2907));
 sg13g2_tiehi \cpu.icache.r_data[1][17]$_DFFE_PP__2908  (.L_HI(net2908));
 sg13g2_tiehi \cpu.icache.r_data[1][18]$_DFFE_PP__2909  (.L_HI(net2909));
 sg13g2_tiehi \cpu.icache.r_data[1][19]$_DFFE_PP__2910  (.L_HI(net2910));
 sg13g2_tiehi \cpu.icache.r_data[1][1]$_DFFE_PP__2911  (.L_HI(net2911));
 sg13g2_tiehi \cpu.icache.r_data[1][20]$_DFFE_PP__2912  (.L_HI(net2912));
 sg13g2_tiehi \cpu.icache.r_data[1][21]$_DFFE_PP__2913  (.L_HI(net2913));
 sg13g2_tiehi \cpu.icache.r_data[1][22]$_DFFE_PP__2914  (.L_HI(net2914));
 sg13g2_tiehi \cpu.icache.r_data[1][23]$_DFFE_PP__2915  (.L_HI(net2915));
 sg13g2_tiehi \cpu.icache.r_data[1][24]$_DFFE_PP__2916  (.L_HI(net2916));
 sg13g2_tiehi \cpu.icache.r_data[1][25]$_DFFE_PP__2917  (.L_HI(net2917));
 sg13g2_tiehi \cpu.icache.r_data[1][26]$_DFFE_PP__2918  (.L_HI(net2918));
 sg13g2_tiehi \cpu.icache.r_data[1][27]$_DFFE_PP__2919  (.L_HI(net2919));
 sg13g2_tiehi \cpu.icache.r_data[1][28]$_DFFE_PP__2920  (.L_HI(net2920));
 sg13g2_tiehi \cpu.icache.r_data[1][29]$_DFFE_PP__2921  (.L_HI(net2921));
 sg13g2_tiehi \cpu.icache.r_data[1][2]$_DFFE_PP__2922  (.L_HI(net2922));
 sg13g2_tiehi \cpu.icache.r_data[1][30]$_DFFE_PP__2923  (.L_HI(net2923));
 sg13g2_tiehi \cpu.icache.r_data[1][31]$_DFFE_PP__2924  (.L_HI(net2924));
 sg13g2_tiehi \cpu.icache.r_data[1][3]$_DFFE_PP__2925  (.L_HI(net2925));
 sg13g2_tiehi \cpu.icache.r_data[1][4]$_DFFE_PP__2926  (.L_HI(net2926));
 sg13g2_tiehi \cpu.icache.r_data[1][5]$_DFFE_PP__2927  (.L_HI(net2927));
 sg13g2_tiehi \cpu.icache.r_data[1][6]$_DFFE_PP__2928  (.L_HI(net2928));
 sg13g2_tiehi \cpu.icache.r_data[1][7]$_DFFE_PP__2929  (.L_HI(net2929));
 sg13g2_tiehi \cpu.icache.r_data[1][8]$_DFFE_PP__2930  (.L_HI(net2930));
 sg13g2_tiehi \cpu.icache.r_data[1][9]$_DFFE_PP__2931  (.L_HI(net2931));
 sg13g2_tiehi \cpu.icache.r_data[2][0]$_DFFE_PP__2932  (.L_HI(net2932));
 sg13g2_tiehi \cpu.icache.r_data[2][10]$_DFFE_PP__2933  (.L_HI(net2933));
 sg13g2_tiehi \cpu.icache.r_data[2][11]$_DFFE_PP__2934  (.L_HI(net2934));
 sg13g2_tiehi \cpu.icache.r_data[2][12]$_DFFE_PP__2935  (.L_HI(net2935));
 sg13g2_tiehi \cpu.icache.r_data[2][13]$_DFFE_PP__2936  (.L_HI(net2936));
 sg13g2_tiehi \cpu.icache.r_data[2][14]$_DFFE_PP__2937  (.L_HI(net2937));
 sg13g2_tiehi \cpu.icache.r_data[2][15]$_DFFE_PP__2938  (.L_HI(net2938));
 sg13g2_tiehi \cpu.icache.r_data[2][16]$_DFFE_PP__2939  (.L_HI(net2939));
 sg13g2_tiehi \cpu.icache.r_data[2][17]$_DFFE_PP__2940  (.L_HI(net2940));
 sg13g2_tiehi \cpu.icache.r_data[2][18]$_DFFE_PP__2941  (.L_HI(net2941));
 sg13g2_tiehi \cpu.icache.r_data[2][19]$_DFFE_PP__2942  (.L_HI(net2942));
 sg13g2_tiehi \cpu.icache.r_data[2][1]$_DFFE_PP__2943  (.L_HI(net2943));
 sg13g2_tiehi \cpu.icache.r_data[2][20]$_DFFE_PP__2944  (.L_HI(net2944));
 sg13g2_tiehi \cpu.icache.r_data[2][21]$_DFFE_PP__2945  (.L_HI(net2945));
 sg13g2_tiehi \cpu.icache.r_data[2][22]$_DFFE_PP__2946  (.L_HI(net2946));
 sg13g2_tiehi \cpu.icache.r_data[2][23]$_DFFE_PP__2947  (.L_HI(net2947));
 sg13g2_tiehi \cpu.icache.r_data[2][24]$_DFFE_PP__2948  (.L_HI(net2948));
 sg13g2_tiehi \cpu.icache.r_data[2][25]$_DFFE_PP__2949  (.L_HI(net2949));
 sg13g2_tiehi \cpu.icache.r_data[2][26]$_DFFE_PP__2950  (.L_HI(net2950));
 sg13g2_tiehi \cpu.icache.r_data[2][27]$_DFFE_PP__2951  (.L_HI(net2951));
 sg13g2_tiehi \cpu.icache.r_data[2][28]$_DFFE_PP__2952  (.L_HI(net2952));
 sg13g2_tiehi \cpu.icache.r_data[2][29]$_DFFE_PP__2953  (.L_HI(net2953));
 sg13g2_tiehi \cpu.icache.r_data[2][2]$_DFFE_PP__2954  (.L_HI(net2954));
 sg13g2_tiehi \cpu.icache.r_data[2][30]$_DFFE_PP__2955  (.L_HI(net2955));
 sg13g2_tiehi \cpu.icache.r_data[2][31]$_DFFE_PP__2956  (.L_HI(net2956));
 sg13g2_tiehi \cpu.icache.r_data[2][3]$_DFFE_PP__2957  (.L_HI(net2957));
 sg13g2_tiehi \cpu.icache.r_data[2][4]$_DFFE_PP__2958  (.L_HI(net2958));
 sg13g2_tiehi \cpu.icache.r_data[2][5]$_DFFE_PP__2959  (.L_HI(net2959));
 sg13g2_tiehi \cpu.icache.r_data[2][6]$_DFFE_PP__2960  (.L_HI(net2960));
 sg13g2_tiehi \cpu.icache.r_data[2][7]$_DFFE_PP__2961  (.L_HI(net2961));
 sg13g2_tiehi \cpu.icache.r_data[2][8]$_DFFE_PP__2962  (.L_HI(net2962));
 sg13g2_tiehi \cpu.icache.r_data[2][9]$_DFFE_PP__2963  (.L_HI(net2963));
 sg13g2_tiehi \cpu.icache.r_data[3][0]$_DFFE_PP__2964  (.L_HI(net2964));
 sg13g2_tiehi \cpu.icache.r_data[3][10]$_DFFE_PP__2965  (.L_HI(net2965));
 sg13g2_tiehi \cpu.icache.r_data[3][11]$_DFFE_PP__2966  (.L_HI(net2966));
 sg13g2_tiehi \cpu.icache.r_data[3][12]$_DFFE_PP__2967  (.L_HI(net2967));
 sg13g2_tiehi \cpu.icache.r_data[3][13]$_DFFE_PP__2968  (.L_HI(net2968));
 sg13g2_tiehi \cpu.icache.r_data[3][14]$_DFFE_PP__2969  (.L_HI(net2969));
 sg13g2_tiehi \cpu.icache.r_data[3][15]$_DFFE_PP__2970  (.L_HI(net2970));
 sg13g2_tiehi \cpu.icache.r_data[3][16]$_DFFE_PP__2971  (.L_HI(net2971));
 sg13g2_tiehi \cpu.icache.r_data[3][17]$_DFFE_PP__2972  (.L_HI(net2972));
 sg13g2_tiehi \cpu.icache.r_data[3][18]$_DFFE_PP__2973  (.L_HI(net2973));
 sg13g2_tiehi \cpu.icache.r_data[3][19]$_DFFE_PP__2974  (.L_HI(net2974));
 sg13g2_tiehi \cpu.icache.r_data[3][1]$_DFFE_PP__2975  (.L_HI(net2975));
 sg13g2_tiehi \cpu.icache.r_data[3][20]$_DFFE_PP__2976  (.L_HI(net2976));
 sg13g2_tiehi \cpu.icache.r_data[3][21]$_DFFE_PP__2977  (.L_HI(net2977));
 sg13g2_tiehi \cpu.icache.r_data[3][22]$_DFFE_PP__2978  (.L_HI(net2978));
 sg13g2_tiehi \cpu.icache.r_data[3][23]$_DFFE_PP__2979  (.L_HI(net2979));
 sg13g2_tiehi \cpu.icache.r_data[3][24]$_DFFE_PP__2980  (.L_HI(net2980));
 sg13g2_tiehi \cpu.icache.r_data[3][25]$_DFFE_PP__2981  (.L_HI(net2981));
 sg13g2_tiehi \cpu.icache.r_data[3][26]$_DFFE_PP__2982  (.L_HI(net2982));
 sg13g2_tiehi \cpu.icache.r_data[3][27]$_DFFE_PP__2983  (.L_HI(net2983));
 sg13g2_tiehi \cpu.icache.r_data[3][28]$_DFFE_PP__2984  (.L_HI(net2984));
 sg13g2_tiehi \cpu.icache.r_data[3][29]$_DFFE_PP__2985  (.L_HI(net2985));
 sg13g2_tiehi \cpu.icache.r_data[3][2]$_DFFE_PP__2986  (.L_HI(net2986));
 sg13g2_tiehi \cpu.icache.r_data[3][30]$_DFFE_PP__2987  (.L_HI(net2987));
 sg13g2_tiehi \cpu.icache.r_data[3][31]$_DFFE_PP__2988  (.L_HI(net2988));
 sg13g2_tiehi \cpu.icache.r_data[3][3]$_DFFE_PP__2989  (.L_HI(net2989));
 sg13g2_tiehi \cpu.icache.r_data[3][4]$_DFFE_PP__2990  (.L_HI(net2990));
 sg13g2_tiehi \cpu.icache.r_data[3][5]$_DFFE_PP__2991  (.L_HI(net2991));
 sg13g2_tiehi \cpu.icache.r_data[3][6]$_DFFE_PP__2992  (.L_HI(net2992));
 sg13g2_tiehi \cpu.icache.r_data[3][7]$_DFFE_PP__2993  (.L_HI(net2993));
 sg13g2_tiehi \cpu.icache.r_data[3][8]$_DFFE_PP__2994  (.L_HI(net2994));
 sg13g2_tiehi \cpu.icache.r_data[3][9]$_DFFE_PP__2995  (.L_HI(net2995));
 sg13g2_tiehi \cpu.icache.r_data[4][0]$_DFFE_PP__2996  (.L_HI(net2996));
 sg13g2_tiehi \cpu.icache.r_data[4][10]$_DFFE_PP__2997  (.L_HI(net2997));
 sg13g2_tiehi \cpu.icache.r_data[4][11]$_DFFE_PP__2998  (.L_HI(net2998));
 sg13g2_tiehi \cpu.icache.r_data[4][12]$_DFFE_PP__2999  (.L_HI(net2999));
 sg13g2_tiehi \cpu.icache.r_data[4][13]$_DFFE_PP__3000  (.L_HI(net3000));
 sg13g2_tiehi \cpu.icache.r_data[4][14]$_DFFE_PP__3001  (.L_HI(net3001));
 sg13g2_tiehi \cpu.icache.r_data[4][15]$_DFFE_PP__3002  (.L_HI(net3002));
 sg13g2_tiehi \cpu.icache.r_data[4][16]$_DFFE_PP__3003  (.L_HI(net3003));
 sg13g2_tiehi \cpu.icache.r_data[4][17]$_DFFE_PP__3004  (.L_HI(net3004));
 sg13g2_tiehi \cpu.icache.r_data[4][18]$_DFFE_PP__3005  (.L_HI(net3005));
 sg13g2_tiehi \cpu.icache.r_data[4][19]$_DFFE_PP__3006  (.L_HI(net3006));
 sg13g2_tiehi \cpu.icache.r_data[4][1]$_DFFE_PP__3007  (.L_HI(net3007));
 sg13g2_tiehi \cpu.icache.r_data[4][20]$_DFFE_PP__3008  (.L_HI(net3008));
 sg13g2_tiehi \cpu.icache.r_data[4][21]$_DFFE_PP__3009  (.L_HI(net3009));
 sg13g2_tiehi \cpu.icache.r_data[4][22]$_DFFE_PP__3010  (.L_HI(net3010));
 sg13g2_tiehi \cpu.icache.r_data[4][23]$_DFFE_PP__3011  (.L_HI(net3011));
 sg13g2_tiehi \cpu.icache.r_data[4][24]$_DFFE_PP__3012  (.L_HI(net3012));
 sg13g2_tiehi \cpu.icache.r_data[4][25]$_DFFE_PP__3013  (.L_HI(net3013));
 sg13g2_tiehi \cpu.icache.r_data[4][26]$_DFFE_PP__3014  (.L_HI(net3014));
 sg13g2_tiehi \cpu.icache.r_data[4][27]$_DFFE_PP__3015  (.L_HI(net3015));
 sg13g2_tiehi \cpu.icache.r_data[4][28]$_DFFE_PP__3016  (.L_HI(net3016));
 sg13g2_tiehi \cpu.icache.r_data[4][29]$_DFFE_PP__3017  (.L_HI(net3017));
 sg13g2_tiehi \cpu.icache.r_data[4][2]$_DFFE_PP__3018  (.L_HI(net3018));
 sg13g2_tiehi \cpu.icache.r_data[4][30]$_DFFE_PP__3019  (.L_HI(net3019));
 sg13g2_tiehi \cpu.icache.r_data[4][31]$_DFFE_PP__3020  (.L_HI(net3020));
 sg13g2_tiehi \cpu.icache.r_data[4][3]$_DFFE_PP__3021  (.L_HI(net3021));
 sg13g2_tiehi \cpu.icache.r_data[4][4]$_DFFE_PP__3022  (.L_HI(net3022));
 sg13g2_tiehi \cpu.icache.r_data[4][5]$_DFFE_PP__3023  (.L_HI(net3023));
 sg13g2_tiehi \cpu.icache.r_data[4][6]$_DFFE_PP__3024  (.L_HI(net3024));
 sg13g2_tiehi \cpu.icache.r_data[4][7]$_DFFE_PP__3025  (.L_HI(net3025));
 sg13g2_tiehi \cpu.icache.r_data[4][8]$_DFFE_PP__3026  (.L_HI(net3026));
 sg13g2_tiehi \cpu.icache.r_data[4][9]$_DFFE_PP__3027  (.L_HI(net3027));
 sg13g2_tiehi \cpu.icache.r_data[5][0]$_DFFE_PP__3028  (.L_HI(net3028));
 sg13g2_tiehi \cpu.icache.r_data[5][10]$_DFFE_PP__3029  (.L_HI(net3029));
 sg13g2_tiehi \cpu.icache.r_data[5][11]$_DFFE_PP__3030  (.L_HI(net3030));
 sg13g2_tiehi \cpu.icache.r_data[5][12]$_DFFE_PP__3031  (.L_HI(net3031));
 sg13g2_tiehi \cpu.icache.r_data[5][13]$_DFFE_PP__3032  (.L_HI(net3032));
 sg13g2_tiehi \cpu.icache.r_data[5][14]$_DFFE_PP__3033  (.L_HI(net3033));
 sg13g2_tiehi \cpu.icache.r_data[5][15]$_DFFE_PP__3034  (.L_HI(net3034));
 sg13g2_tiehi \cpu.icache.r_data[5][16]$_DFFE_PP__3035  (.L_HI(net3035));
 sg13g2_tiehi \cpu.icache.r_data[5][17]$_DFFE_PP__3036  (.L_HI(net3036));
 sg13g2_tiehi \cpu.icache.r_data[5][18]$_DFFE_PP__3037  (.L_HI(net3037));
 sg13g2_tiehi \cpu.icache.r_data[5][19]$_DFFE_PP__3038  (.L_HI(net3038));
 sg13g2_tiehi \cpu.icache.r_data[5][1]$_DFFE_PP__3039  (.L_HI(net3039));
 sg13g2_tiehi \cpu.icache.r_data[5][20]$_DFFE_PP__3040  (.L_HI(net3040));
 sg13g2_tiehi \cpu.icache.r_data[5][21]$_DFFE_PP__3041  (.L_HI(net3041));
 sg13g2_tiehi \cpu.icache.r_data[5][22]$_DFFE_PP__3042  (.L_HI(net3042));
 sg13g2_tiehi \cpu.icache.r_data[5][23]$_DFFE_PP__3043  (.L_HI(net3043));
 sg13g2_tiehi \cpu.icache.r_data[5][24]$_DFFE_PP__3044  (.L_HI(net3044));
 sg13g2_tiehi \cpu.icache.r_data[5][25]$_DFFE_PP__3045  (.L_HI(net3045));
 sg13g2_tiehi \cpu.icache.r_data[5][26]$_DFFE_PP__3046  (.L_HI(net3046));
 sg13g2_tiehi \cpu.icache.r_data[5][27]$_DFFE_PP__3047  (.L_HI(net3047));
 sg13g2_tiehi \cpu.icache.r_data[5][28]$_DFFE_PP__3048  (.L_HI(net3048));
 sg13g2_tiehi \cpu.icache.r_data[5][29]$_DFFE_PP__3049  (.L_HI(net3049));
 sg13g2_tiehi \cpu.icache.r_data[5][2]$_DFFE_PP__3050  (.L_HI(net3050));
 sg13g2_tiehi \cpu.icache.r_data[5][30]$_DFFE_PP__3051  (.L_HI(net3051));
 sg13g2_tiehi \cpu.icache.r_data[5][31]$_DFFE_PP__3052  (.L_HI(net3052));
 sg13g2_tiehi \cpu.icache.r_data[5][3]$_DFFE_PP__3053  (.L_HI(net3053));
 sg13g2_tiehi \cpu.icache.r_data[5][4]$_DFFE_PP__3054  (.L_HI(net3054));
 sg13g2_tiehi \cpu.icache.r_data[5][5]$_DFFE_PP__3055  (.L_HI(net3055));
 sg13g2_tiehi \cpu.icache.r_data[5][6]$_DFFE_PP__3056  (.L_HI(net3056));
 sg13g2_tiehi \cpu.icache.r_data[5][7]$_DFFE_PP__3057  (.L_HI(net3057));
 sg13g2_tiehi \cpu.icache.r_data[5][8]$_DFFE_PP__3058  (.L_HI(net3058));
 sg13g2_tiehi \cpu.icache.r_data[5][9]$_DFFE_PP__3059  (.L_HI(net3059));
 sg13g2_tiehi \cpu.icache.r_data[6][0]$_DFFE_PP__3060  (.L_HI(net3060));
 sg13g2_tiehi \cpu.icache.r_data[6][10]$_DFFE_PP__3061  (.L_HI(net3061));
 sg13g2_tiehi \cpu.icache.r_data[6][11]$_DFFE_PP__3062  (.L_HI(net3062));
 sg13g2_tiehi \cpu.icache.r_data[6][12]$_DFFE_PP__3063  (.L_HI(net3063));
 sg13g2_tiehi \cpu.icache.r_data[6][13]$_DFFE_PP__3064  (.L_HI(net3064));
 sg13g2_tiehi \cpu.icache.r_data[6][14]$_DFFE_PP__3065  (.L_HI(net3065));
 sg13g2_tiehi \cpu.icache.r_data[6][15]$_DFFE_PP__3066  (.L_HI(net3066));
 sg13g2_tiehi \cpu.icache.r_data[6][16]$_DFFE_PP__3067  (.L_HI(net3067));
 sg13g2_tiehi \cpu.icache.r_data[6][17]$_DFFE_PP__3068  (.L_HI(net3068));
 sg13g2_tiehi \cpu.icache.r_data[6][18]$_DFFE_PP__3069  (.L_HI(net3069));
 sg13g2_tiehi \cpu.icache.r_data[6][19]$_DFFE_PP__3070  (.L_HI(net3070));
 sg13g2_tiehi \cpu.icache.r_data[6][1]$_DFFE_PP__3071  (.L_HI(net3071));
 sg13g2_tiehi \cpu.icache.r_data[6][20]$_DFFE_PP__3072  (.L_HI(net3072));
 sg13g2_tiehi \cpu.icache.r_data[6][21]$_DFFE_PP__3073  (.L_HI(net3073));
 sg13g2_tiehi \cpu.icache.r_data[6][22]$_DFFE_PP__3074  (.L_HI(net3074));
 sg13g2_tiehi \cpu.icache.r_data[6][23]$_DFFE_PP__3075  (.L_HI(net3075));
 sg13g2_tiehi \cpu.icache.r_data[6][24]$_DFFE_PP__3076  (.L_HI(net3076));
 sg13g2_tiehi \cpu.icache.r_data[6][25]$_DFFE_PP__3077  (.L_HI(net3077));
 sg13g2_tiehi \cpu.icache.r_data[6][26]$_DFFE_PP__3078  (.L_HI(net3078));
 sg13g2_tiehi \cpu.icache.r_data[6][27]$_DFFE_PP__3079  (.L_HI(net3079));
 sg13g2_tiehi \cpu.icache.r_data[6][28]$_DFFE_PP__3080  (.L_HI(net3080));
 sg13g2_tiehi \cpu.icache.r_data[6][29]$_DFFE_PP__3081  (.L_HI(net3081));
 sg13g2_tiehi \cpu.icache.r_data[6][2]$_DFFE_PP__3082  (.L_HI(net3082));
 sg13g2_tiehi \cpu.icache.r_data[6][30]$_DFFE_PP__3083  (.L_HI(net3083));
 sg13g2_tiehi \cpu.icache.r_data[6][31]$_DFFE_PP__3084  (.L_HI(net3084));
 sg13g2_tiehi \cpu.icache.r_data[6][3]$_DFFE_PP__3085  (.L_HI(net3085));
 sg13g2_tiehi \cpu.icache.r_data[6][4]$_DFFE_PP__3086  (.L_HI(net3086));
 sg13g2_tiehi \cpu.icache.r_data[6][5]$_DFFE_PP__3087  (.L_HI(net3087));
 sg13g2_tiehi \cpu.icache.r_data[6][6]$_DFFE_PP__3088  (.L_HI(net3088));
 sg13g2_tiehi \cpu.icache.r_data[6][7]$_DFFE_PP__3089  (.L_HI(net3089));
 sg13g2_tiehi \cpu.icache.r_data[6][8]$_DFFE_PP__3090  (.L_HI(net3090));
 sg13g2_tiehi \cpu.icache.r_data[6][9]$_DFFE_PP__3091  (.L_HI(net3091));
 sg13g2_tiehi \cpu.icache.r_data[7][0]$_DFFE_PP__3092  (.L_HI(net3092));
 sg13g2_tiehi \cpu.icache.r_data[7][10]$_DFFE_PP__3093  (.L_HI(net3093));
 sg13g2_tiehi \cpu.icache.r_data[7][11]$_DFFE_PP__3094  (.L_HI(net3094));
 sg13g2_tiehi \cpu.icache.r_data[7][12]$_DFFE_PP__3095  (.L_HI(net3095));
 sg13g2_tiehi \cpu.icache.r_data[7][13]$_DFFE_PP__3096  (.L_HI(net3096));
 sg13g2_tiehi \cpu.icache.r_data[7][14]$_DFFE_PP__3097  (.L_HI(net3097));
 sg13g2_tiehi \cpu.icache.r_data[7][15]$_DFFE_PP__3098  (.L_HI(net3098));
 sg13g2_tiehi \cpu.icache.r_data[7][16]$_DFFE_PP__3099  (.L_HI(net3099));
 sg13g2_tiehi \cpu.icache.r_data[7][17]$_DFFE_PP__3100  (.L_HI(net3100));
 sg13g2_tiehi \cpu.icache.r_data[7][18]$_DFFE_PP__3101  (.L_HI(net3101));
 sg13g2_tiehi \cpu.icache.r_data[7][19]$_DFFE_PP__3102  (.L_HI(net3102));
 sg13g2_tiehi \cpu.icache.r_data[7][1]$_DFFE_PP__3103  (.L_HI(net3103));
 sg13g2_tiehi \cpu.icache.r_data[7][20]$_DFFE_PP__3104  (.L_HI(net3104));
 sg13g2_tiehi \cpu.icache.r_data[7][21]$_DFFE_PP__3105  (.L_HI(net3105));
 sg13g2_tiehi \cpu.icache.r_data[7][22]$_DFFE_PP__3106  (.L_HI(net3106));
 sg13g2_tiehi \cpu.icache.r_data[7][23]$_DFFE_PP__3107  (.L_HI(net3107));
 sg13g2_tiehi \cpu.icache.r_data[7][24]$_DFFE_PP__3108  (.L_HI(net3108));
 sg13g2_tiehi \cpu.icache.r_data[7][25]$_DFFE_PP__3109  (.L_HI(net3109));
 sg13g2_tiehi \cpu.icache.r_data[7][26]$_DFFE_PP__3110  (.L_HI(net3110));
 sg13g2_tiehi \cpu.icache.r_data[7][27]$_DFFE_PP__3111  (.L_HI(net3111));
 sg13g2_tiehi \cpu.icache.r_data[7][28]$_DFFE_PP__3112  (.L_HI(net3112));
 sg13g2_tiehi \cpu.icache.r_data[7][29]$_DFFE_PP__3113  (.L_HI(net3113));
 sg13g2_tiehi \cpu.icache.r_data[7][2]$_DFFE_PP__3114  (.L_HI(net3114));
 sg13g2_tiehi \cpu.icache.r_data[7][30]$_DFFE_PP__3115  (.L_HI(net3115));
 sg13g2_tiehi \cpu.icache.r_data[7][31]$_DFFE_PP__3116  (.L_HI(net3116));
 sg13g2_tiehi \cpu.icache.r_data[7][3]$_DFFE_PP__3117  (.L_HI(net3117));
 sg13g2_tiehi \cpu.icache.r_data[7][4]$_DFFE_PP__3118  (.L_HI(net3118));
 sg13g2_tiehi \cpu.icache.r_data[7][5]$_DFFE_PP__3119  (.L_HI(net3119));
 sg13g2_tiehi \cpu.icache.r_data[7][6]$_DFFE_PP__3120  (.L_HI(net3120));
 sg13g2_tiehi \cpu.icache.r_data[7][7]$_DFFE_PP__3121  (.L_HI(net3121));
 sg13g2_tiehi \cpu.icache.r_data[7][8]$_DFFE_PP__3122  (.L_HI(net3122));
 sg13g2_tiehi \cpu.icache.r_data[7][9]$_DFFE_PP__3123  (.L_HI(net3123));
 sg13g2_tiehi \cpu.icache.r_offset[0]$_SDFF_PN0__3124  (.L_HI(net3124));
 sg13g2_tiehi \cpu.icache.r_offset[1]$_SDFF_PN0__3125  (.L_HI(net3125));
 sg13g2_tiehi \cpu.icache.r_offset[2]$_SDFF_PN0__3126  (.L_HI(net3126));
 sg13g2_tiehi \cpu.icache.r_tag[0][0]$_DFFE_PP__3127  (.L_HI(net3127));
 sg13g2_tiehi \cpu.icache.r_tag[0][10]$_DFFE_PP__3128  (.L_HI(net3128));
 sg13g2_tiehi \cpu.icache.r_tag[0][11]$_DFFE_PP__3129  (.L_HI(net3129));
 sg13g2_tiehi \cpu.icache.r_tag[0][12]$_DFFE_PP__3130  (.L_HI(net3130));
 sg13g2_tiehi \cpu.icache.r_tag[0][13]$_DFFE_PP__3131  (.L_HI(net3131));
 sg13g2_tiehi \cpu.icache.r_tag[0][14]$_DFFE_PP__3132  (.L_HI(net3132));
 sg13g2_tiehi \cpu.icache.r_tag[0][15]$_DFFE_PP__3133  (.L_HI(net3133));
 sg13g2_tiehi \cpu.icache.r_tag[0][16]$_DFFE_PP__3134  (.L_HI(net3134));
 sg13g2_tiehi \cpu.icache.r_tag[0][17]$_DFFE_PP__3135  (.L_HI(net3135));
 sg13g2_tiehi \cpu.icache.r_tag[0][18]$_DFFE_PP__3136  (.L_HI(net3136));
 sg13g2_tiehi \cpu.icache.r_tag[0][1]$_DFFE_PP__3137  (.L_HI(net3137));
 sg13g2_tiehi \cpu.icache.r_tag[0][2]$_DFFE_PP__3138  (.L_HI(net3138));
 sg13g2_tiehi \cpu.icache.r_tag[0][3]$_DFFE_PP__3139  (.L_HI(net3139));
 sg13g2_tiehi \cpu.icache.r_tag[0][4]$_DFFE_PP__3140  (.L_HI(net3140));
 sg13g2_tiehi \cpu.icache.r_tag[0][5]$_DFFE_PP__3141  (.L_HI(net3141));
 sg13g2_tiehi \cpu.icache.r_tag[0][6]$_DFFE_PP__3142  (.L_HI(net3142));
 sg13g2_tiehi \cpu.icache.r_tag[0][7]$_DFFE_PP__3143  (.L_HI(net3143));
 sg13g2_tiehi \cpu.icache.r_tag[0][8]$_DFFE_PP__3144  (.L_HI(net3144));
 sg13g2_tiehi \cpu.icache.r_tag[0][9]$_DFFE_PP__3145  (.L_HI(net3145));
 sg13g2_tiehi \cpu.icache.r_tag[1][0]$_DFFE_PP__3146  (.L_HI(net3146));
 sg13g2_tiehi \cpu.icache.r_tag[1][10]$_DFFE_PP__3147  (.L_HI(net3147));
 sg13g2_tiehi \cpu.icache.r_tag[1][11]$_DFFE_PP__3148  (.L_HI(net3148));
 sg13g2_tiehi \cpu.icache.r_tag[1][12]$_DFFE_PP__3149  (.L_HI(net3149));
 sg13g2_tiehi \cpu.icache.r_tag[1][13]$_DFFE_PP__3150  (.L_HI(net3150));
 sg13g2_tiehi \cpu.icache.r_tag[1][14]$_DFFE_PP__3151  (.L_HI(net3151));
 sg13g2_tiehi \cpu.icache.r_tag[1][15]$_DFFE_PP__3152  (.L_HI(net3152));
 sg13g2_tiehi \cpu.icache.r_tag[1][16]$_DFFE_PP__3153  (.L_HI(net3153));
 sg13g2_tiehi \cpu.icache.r_tag[1][17]$_DFFE_PP__3154  (.L_HI(net3154));
 sg13g2_tiehi \cpu.icache.r_tag[1][18]$_DFFE_PP__3155  (.L_HI(net3155));
 sg13g2_tiehi \cpu.icache.r_tag[1][1]$_DFFE_PP__3156  (.L_HI(net3156));
 sg13g2_tiehi \cpu.icache.r_tag[1][2]$_DFFE_PP__3157  (.L_HI(net3157));
 sg13g2_tiehi \cpu.icache.r_tag[1][3]$_DFFE_PP__3158  (.L_HI(net3158));
 sg13g2_tiehi \cpu.icache.r_tag[1][4]$_DFFE_PP__3159  (.L_HI(net3159));
 sg13g2_tiehi \cpu.icache.r_tag[1][5]$_DFFE_PP__3160  (.L_HI(net3160));
 sg13g2_tiehi \cpu.icache.r_tag[1][6]$_DFFE_PP__3161  (.L_HI(net3161));
 sg13g2_tiehi \cpu.icache.r_tag[1][7]$_DFFE_PP__3162  (.L_HI(net3162));
 sg13g2_tiehi \cpu.icache.r_tag[1][8]$_DFFE_PP__3163  (.L_HI(net3163));
 sg13g2_tiehi \cpu.icache.r_tag[1][9]$_DFFE_PP__3164  (.L_HI(net3164));
 sg13g2_tiehi \cpu.icache.r_tag[2][0]$_DFFE_PP__3165  (.L_HI(net3165));
 sg13g2_tiehi \cpu.icache.r_tag[2][10]$_DFFE_PP__3166  (.L_HI(net3166));
 sg13g2_tiehi \cpu.icache.r_tag[2][11]$_DFFE_PP__3167  (.L_HI(net3167));
 sg13g2_tiehi \cpu.icache.r_tag[2][12]$_DFFE_PP__3168  (.L_HI(net3168));
 sg13g2_tiehi \cpu.icache.r_tag[2][13]$_DFFE_PP__3169  (.L_HI(net3169));
 sg13g2_tiehi \cpu.icache.r_tag[2][14]$_DFFE_PP__3170  (.L_HI(net3170));
 sg13g2_tiehi \cpu.icache.r_tag[2][15]$_DFFE_PP__3171  (.L_HI(net3171));
 sg13g2_tiehi \cpu.icache.r_tag[2][16]$_DFFE_PP__3172  (.L_HI(net3172));
 sg13g2_tiehi \cpu.icache.r_tag[2][17]$_DFFE_PP__3173  (.L_HI(net3173));
 sg13g2_tiehi \cpu.icache.r_tag[2][18]$_DFFE_PP__3174  (.L_HI(net3174));
 sg13g2_tiehi \cpu.icache.r_tag[2][1]$_DFFE_PP__3175  (.L_HI(net3175));
 sg13g2_tiehi \cpu.icache.r_tag[2][2]$_DFFE_PP__3176  (.L_HI(net3176));
 sg13g2_tiehi \cpu.icache.r_tag[2][3]$_DFFE_PP__3177  (.L_HI(net3177));
 sg13g2_tiehi \cpu.icache.r_tag[2][4]$_DFFE_PP__3178  (.L_HI(net3178));
 sg13g2_tiehi \cpu.icache.r_tag[2][5]$_DFFE_PP__3179  (.L_HI(net3179));
 sg13g2_tiehi \cpu.icache.r_tag[2][6]$_DFFE_PP__3180  (.L_HI(net3180));
 sg13g2_tiehi \cpu.icache.r_tag[2][7]$_DFFE_PP__3181  (.L_HI(net3181));
 sg13g2_tiehi \cpu.icache.r_tag[2][8]$_DFFE_PP__3182  (.L_HI(net3182));
 sg13g2_tiehi \cpu.icache.r_tag[2][9]$_DFFE_PP__3183  (.L_HI(net3183));
 sg13g2_tiehi \cpu.icache.r_tag[3][0]$_DFFE_PP__3184  (.L_HI(net3184));
 sg13g2_tiehi \cpu.icache.r_tag[3][10]$_DFFE_PP__3185  (.L_HI(net3185));
 sg13g2_tiehi \cpu.icache.r_tag[3][11]$_DFFE_PP__3186  (.L_HI(net3186));
 sg13g2_tiehi \cpu.icache.r_tag[3][12]$_DFFE_PP__3187  (.L_HI(net3187));
 sg13g2_tiehi \cpu.icache.r_tag[3][13]$_DFFE_PP__3188  (.L_HI(net3188));
 sg13g2_tiehi \cpu.icache.r_tag[3][14]$_DFFE_PP__3189  (.L_HI(net3189));
 sg13g2_tiehi \cpu.icache.r_tag[3][15]$_DFFE_PP__3190  (.L_HI(net3190));
 sg13g2_tiehi \cpu.icache.r_tag[3][16]$_DFFE_PP__3191  (.L_HI(net3191));
 sg13g2_tiehi \cpu.icache.r_tag[3][17]$_DFFE_PP__3192  (.L_HI(net3192));
 sg13g2_tiehi \cpu.icache.r_tag[3][18]$_DFFE_PP__3193  (.L_HI(net3193));
 sg13g2_tiehi \cpu.icache.r_tag[3][1]$_DFFE_PP__3194  (.L_HI(net3194));
 sg13g2_tiehi \cpu.icache.r_tag[3][2]$_DFFE_PP__3195  (.L_HI(net3195));
 sg13g2_tiehi \cpu.icache.r_tag[3][3]$_DFFE_PP__3196  (.L_HI(net3196));
 sg13g2_tiehi \cpu.icache.r_tag[3][4]$_DFFE_PP__3197  (.L_HI(net3197));
 sg13g2_tiehi \cpu.icache.r_tag[3][5]$_DFFE_PP__3198  (.L_HI(net3198));
 sg13g2_tiehi \cpu.icache.r_tag[3][6]$_DFFE_PP__3199  (.L_HI(net3199));
 sg13g2_tiehi \cpu.icache.r_tag[3][7]$_DFFE_PP__3200  (.L_HI(net3200));
 sg13g2_tiehi \cpu.icache.r_tag[3][8]$_DFFE_PP__3201  (.L_HI(net3201));
 sg13g2_tiehi \cpu.icache.r_tag[3][9]$_DFFE_PP__3202  (.L_HI(net3202));
 sg13g2_tiehi \cpu.icache.r_tag[4][0]$_DFFE_PP__3203  (.L_HI(net3203));
 sg13g2_tiehi \cpu.icache.r_tag[4][10]$_DFFE_PP__3204  (.L_HI(net3204));
 sg13g2_tiehi \cpu.icache.r_tag[4][11]$_DFFE_PP__3205  (.L_HI(net3205));
 sg13g2_tiehi \cpu.icache.r_tag[4][12]$_DFFE_PP__3206  (.L_HI(net3206));
 sg13g2_tiehi \cpu.icache.r_tag[4][13]$_DFFE_PP__3207  (.L_HI(net3207));
 sg13g2_tiehi \cpu.icache.r_tag[4][14]$_DFFE_PP__3208  (.L_HI(net3208));
 sg13g2_tiehi \cpu.icache.r_tag[4][15]$_DFFE_PP__3209  (.L_HI(net3209));
 sg13g2_tiehi \cpu.icache.r_tag[4][16]$_DFFE_PP__3210  (.L_HI(net3210));
 sg13g2_tiehi \cpu.icache.r_tag[4][17]$_DFFE_PP__3211  (.L_HI(net3211));
 sg13g2_tiehi \cpu.icache.r_tag[4][18]$_DFFE_PP__3212  (.L_HI(net3212));
 sg13g2_tiehi \cpu.icache.r_tag[4][1]$_DFFE_PP__3213  (.L_HI(net3213));
 sg13g2_tiehi \cpu.icache.r_tag[4][2]$_DFFE_PP__3214  (.L_HI(net3214));
 sg13g2_tiehi \cpu.icache.r_tag[4][3]$_DFFE_PP__3215  (.L_HI(net3215));
 sg13g2_tiehi \cpu.icache.r_tag[4][4]$_DFFE_PP__3216  (.L_HI(net3216));
 sg13g2_tiehi \cpu.icache.r_tag[4][5]$_DFFE_PP__3217  (.L_HI(net3217));
 sg13g2_tiehi \cpu.icache.r_tag[4][6]$_DFFE_PP__3218  (.L_HI(net3218));
 sg13g2_tiehi \cpu.icache.r_tag[4][7]$_DFFE_PP__3219  (.L_HI(net3219));
 sg13g2_tiehi \cpu.icache.r_tag[4][8]$_DFFE_PP__3220  (.L_HI(net3220));
 sg13g2_tiehi \cpu.icache.r_tag[4][9]$_DFFE_PP__3221  (.L_HI(net3221));
 sg13g2_tiehi \cpu.icache.r_tag[5][0]$_DFFE_PP__3222  (.L_HI(net3222));
 sg13g2_tiehi \cpu.icache.r_tag[5][10]$_DFFE_PP__3223  (.L_HI(net3223));
 sg13g2_tiehi \cpu.icache.r_tag[5][11]$_DFFE_PP__3224  (.L_HI(net3224));
 sg13g2_tiehi \cpu.icache.r_tag[5][12]$_DFFE_PP__3225  (.L_HI(net3225));
 sg13g2_tiehi \cpu.icache.r_tag[5][13]$_DFFE_PP__3226  (.L_HI(net3226));
 sg13g2_tiehi \cpu.icache.r_tag[5][14]$_DFFE_PP__3227  (.L_HI(net3227));
 sg13g2_tiehi \cpu.icache.r_tag[5][15]$_DFFE_PP__3228  (.L_HI(net3228));
 sg13g2_tiehi \cpu.icache.r_tag[5][16]$_DFFE_PP__3229  (.L_HI(net3229));
 sg13g2_tiehi \cpu.icache.r_tag[5][17]$_DFFE_PP__3230  (.L_HI(net3230));
 sg13g2_tiehi \cpu.icache.r_tag[5][18]$_DFFE_PP__3231  (.L_HI(net3231));
 sg13g2_tiehi \cpu.icache.r_tag[5][1]$_DFFE_PP__3232  (.L_HI(net3232));
 sg13g2_tiehi \cpu.icache.r_tag[5][2]$_DFFE_PP__3233  (.L_HI(net3233));
 sg13g2_tiehi \cpu.icache.r_tag[5][3]$_DFFE_PP__3234  (.L_HI(net3234));
 sg13g2_tiehi \cpu.icache.r_tag[5][4]$_DFFE_PP__3235  (.L_HI(net3235));
 sg13g2_tiehi \cpu.icache.r_tag[5][5]$_DFFE_PP__3236  (.L_HI(net3236));
 sg13g2_tiehi \cpu.icache.r_tag[5][6]$_DFFE_PP__3237  (.L_HI(net3237));
 sg13g2_tiehi \cpu.icache.r_tag[5][7]$_DFFE_PP__3238  (.L_HI(net3238));
 sg13g2_tiehi \cpu.icache.r_tag[5][8]$_DFFE_PP__3239  (.L_HI(net3239));
 sg13g2_tiehi \cpu.icache.r_tag[5][9]$_DFFE_PP__3240  (.L_HI(net3240));
 sg13g2_tiehi \cpu.icache.r_tag[6][0]$_DFFE_PP__3241  (.L_HI(net3241));
 sg13g2_tiehi \cpu.icache.r_tag[6][10]$_DFFE_PP__3242  (.L_HI(net3242));
 sg13g2_tiehi \cpu.icache.r_tag[6][11]$_DFFE_PP__3243  (.L_HI(net3243));
 sg13g2_tiehi \cpu.icache.r_tag[6][12]$_DFFE_PP__3244  (.L_HI(net3244));
 sg13g2_tiehi \cpu.icache.r_tag[6][13]$_DFFE_PP__3245  (.L_HI(net3245));
 sg13g2_tiehi \cpu.icache.r_tag[6][14]$_DFFE_PP__3246  (.L_HI(net3246));
 sg13g2_tiehi \cpu.icache.r_tag[6][15]$_DFFE_PP__3247  (.L_HI(net3247));
 sg13g2_tiehi \cpu.icache.r_tag[6][16]$_DFFE_PP__3248  (.L_HI(net3248));
 sg13g2_tiehi \cpu.icache.r_tag[6][17]$_DFFE_PP__3249  (.L_HI(net3249));
 sg13g2_tiehi \cpu.icache.r_tag[6][18]$_DFFE_PP__3250  (.L_HI(net3250));
 sg13g2_tiehi \cpu.icache.r_tag[6][1]$_DFFE_PP__3251  (.L_HI(net3251));
 sg13g2_tiehi \cpu.icache.r_tag[6][2]$_DFFE_PP__3252  (.L_HI(net3252));
 sg13g2_tiehi \cpu.icache.r_tag[6][3]$_DFFE_PP__3253  (.L_HI(net3253));
 sg13g2_tiehi \cpu.icache.r_tag[6][4]$_DFFE_PP__3254  (.L_HI(net3254));
 sg13g2_tiehi \cpu.icache.r_tag[6][5]$_DFFE_PP__3255  (.L_HI(net3255));
 sg13g2_tiehi \cpu.icache.r_tag[6][6]$_DFFE_PP__3256  (.L_HI(net3256));
 sg13g2_tiehi \cpu.icache.r_tag[6][7]$_DFFE_PP__3257  (.L_HI(net3257));
 sg13g2_tiehi \cpu.icache.r_tag[6][8]$_DFFE_PP__3258  (.L_HI(net3258));
 sg13g2_tiehi \cpu.icache.r_tag[6][9]$_DFFE_PP__3259  (.L_HI(net3259));
 sg13g2_tiehi \cpu.icache.r_tag[7][0]$_DFFE_PP__3260  (.L_HI(net3260));
 sg13g2_tiehi \cpu.icache.r_tag[7][10]$_DFFE_PP__3261  (.L_HI(net3261));
 sg13g2_tiehi \cpu.icache.r_tag[7][11]$_DFFE_PP__3262  (.L_HI(net3262));
 sg13g2_tiehi \cpu.icache.r_tag[7][12]$_DFFE_PP__3263  (.L_HI(net3263));
 sg13g2_tiehi \cpu.icache.r_tag[7][13]$_DFFE_PP__3264  (.L_HI(net3264));
 sg13g2_tiehi \cpu.icache.r_tag[7][14]$_DFFE_PP__3265  (.L_HI(net3265));
 sg13g2_tiehi \cpu.icache.r_tag[7][15]$_DFFE_PP__3266  (.L_HI(net3266));
 sg13g2_tiehi \cpu.icache.r_tag[7][16]$_DFFE_PP__3267  (.L_HI(net3267));
 sg13g2_tiehi \cpu.icache.r_tag[7][17]$_DFFE_PP__3268  (.L_HI(net3268));
 sg13g2_tiehi \cpu.icache.r_tag[7][18]$_DFFE_PP__3269  (.L_HI(net3269));
 sg13g2_tiehi \cpu.icache.r_tag[7][1]$_DFFE_PP__3270  (.L_HI(net3270));
 sg13g2_tiehi \cpu.icache.r_tag[7][2]$_DFFE_PP__3271  (.L_HI(net3271));
 sg13g2_tiehi \cpu.icache.r_tag[7][3]$_DFFE_PP__3272  (.L_HI(net3272));
 sg13g2_tiehi \cpu.icache.r_tag[7][4]$_DFFE_PP__3273  (.L_HI(net3273));
 sg13g2_tiehi \cpu.icache.r_tag[7][5]$_DFFE_PP__3274  (.L_HI(net3274));
 sg13g2_tiehi \cpu.icache.r_tag[7][6]$_DFFE_PP__3275  (.L_HI(net3275));
 sg13g2_tiehi \cpu.icache.r_tag[7][7]$_DFFE_PP__3276  (.L_HI(net3276));
 sg13g2_tiehi \cpu.icache.r_tag[7][8]$_DFFE_PP__3277  (.L_HI(net3277));
 sg13g2_tiehi \cpu.icache.r_tag[7][9]$_DFFE_PP__3278  (.L_HI(net3278));
 sg13g2_tiehi \cpu.icache.r_valid[0]$_SDFFE_PP0P__3279  (.L_HI(net3279));
 sg13g2_tiehi \cpu.icache.r_valid[1]$_SDFFE_PP0P__3280  (.L_HI(net3280));
 sg13g2_tiehi \cpu.icache.r_valid[2]$_SDFFE_PP0P__3281  (.L_HI(net3281));
 sg13g2_tiehi \cpu.icache.r_valid[3]$_SDFFE_PP0P__3282  (.L_HI(net3282));
 sg13g2_tiehi \cpu.icache.r_valid[4]$_SDFFE_PP0P__3283  (.L_HI(net3283));
 sg13g2_tiehi \cpu.icache.r_valid[5]$_SDFFE_PP0P__3284  (.L_HI(net3284));
 sg13g2_tiehi \cpu.icache.r_valid[6]$_SDFFE_PP0P__3285  (.L_HI(net3285));
 sg13g2_tiehi \cpu.icache.r_valid[7]$_SDFFE_PP0P__3286  (.L_HI(net3286));
 sg13g2_tiehi \cpu.intr.r_clock$_SDFFE_PN0P__3287  (.L_HI(net3287));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[0]$_DFFE_PP__3288  (.L_HI(net3288));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[10]$_DFFE_PP__3289  (.L_HI(net3289));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[11]$_DFFE_PP__3290  (.L_HI(net3290));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[12]$_DFFE_PP__3291  (.L_HI(net3291));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[13]$_DFFE_PP__3292  (.L_HI(net3292));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[14]$_DFFE_PP__3293  (.L_HI(net3293));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[15]$_DFFE_PP__3294  (.L_HI(net3294));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[16]$_DFFE_PP__3295  (.L_HI(net3295));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[17]$_DFFE_PP__3296  (.L_HI(net3296));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[18]$_DFFE_PP__3297  (.L_HI(net3297));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[19]$_DFFE_PP__3298  (.L_HI(net3298));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[1]$_DFFE_PP__3299  (.L_HI(net3299));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[20]$_DFFE_PP__3300  (.L_HI(net3300));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[21]$_DFFE_PP__3301  (.L_HI(net3301));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[22]$_DFFE_PP__3302  (.L_HI(net3302));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[23]$_DFFE_PP__3303  (.L_HI(net3303));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[24]$_DFFE_PP__3304  (.L_HI(net3304));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[25]$_DFFE_PP__3305  (.L_HI(net3305));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[26]$_DFFE_PP__3306  (.L_HI(net3306));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[27]$_DFFE_PP__3307  (.L_HI(net3307));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[28]$_DFFE_PP__3308  (.L_HI(net3308));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[29]$_DFFE_PP__3309  (.L_HI(net3309));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[2]$_DFFE_PP__3310  (.L_HI(net3310));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[30]$_DFFE_PP__3311  (.L_HI(net3311));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[31]$_DFFE_PP__3312  (.L_HI(net3312));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[3]$_DFFE_PP__3313  (.L_HI(net3313));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[4]$_DFFE_PP__3314  (.L_HI(net3314));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[5]$_DFFE_PP__3315  (.L_HI(net3315));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[6]$_DFFE_PP__3316  (.L_HI(net3316));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[7]$_DFFE_PP__3317  (.L_HI(net3317));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[8]$_DFFE_PP__3318  (.L_HI(net3318));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[9]$_DFFE_PP__3319  (.L_HI(net3319));
 sg13g2_tiehi \cpu.intr.r_clock_count[0]$_DFF_P__3320  (.L_HI(net3320));
 sg13g2_tiehi \cpu.intr.r_clock_count[10]$_DFF_P__3321  (.L_HI(net3321));
 sg13g2_tiehi \cpu.intr.r_clock_count[11]$_DFF_P__3322  (.L_HI(net3322));
 sg13g2_tiehi \cpu.intr.r_clock_count[12]$_DFF_P__3323  (.L_HI(net3323));
 sg13g2_tiehi \cpu.intr.r_clock_count[13]$_DFF_P__3324  (.L_HI(net3324));
 sg13g2_tiehi \cpu.intr.r_clock_count[14]$_DFF_P__3325  (.L_HI(net3325));
 sg13g2_tiehi \cpu.intr.r_clock_count[15]$_DFF_P__3326  (.L_HI(net3326));
 sg13g2_tiehi \cpu.intr.r_clock_count[16]$_DFFE_PN__3327  (.L_HI(net3327));
 sg13g2_tiehi \cpu.intr.r_clock_count[17]$_DFFE_PN__3328  (.L_HI(net3328));
 sg13g2_tiehi \cpu.intr.r_clock_count[18]$_DFFE_PN__3329  (.L_HI(net3329));
 sg13g2_tiehi \cpu.intr.r_clock_count[19]$_DFFE_PN__3330  (.L_HI(net3330));
 sg13g2_tiehi \cpu.intr.r_clock_count[1]$_DFF_P__3331  (.L_HI(net3331));
 sg13g2_tiehi \cpu.intr.r_clock_count[20]$_DFFE_PN__3332  (.L_HI(net3332));
 sg13g2_tiehi \cpu.intr.r_clock_count[21]$_DFFE_PN__3333  (.L_HI(net3333));
 sg13g2_tiehi \cpu.intr.r_clock_count[22]$_DFFE_PN__3334  (.L_HI(net3334));
 sg13g2_tiehi \cpu.intr.r_clock_count[23]$_DFFE_PN__3335  (.L_HI(net3335));
 sg13g2_tiehi \cpu.intr.r_clock_count[24]$_DFFE_PN__3336  (.L_HI(net3336));
 sg13g2_tiehi \cpu.intr.r_clock_count[25]$_DFFE_PN__3337  (.L_HI(net3337));
 sg13g2_tiehi \cpu.intr.r_clock_count[26]$_DFFE_PN__3338  (.L_HI(net3338));
 sg13g2_tiehi \cpu.intr.r_clock_count[27]$_DFFE_PN__3339  (.L_HI(net3339));
 sg13g2_tiehi \cpu.intr.r_clock_count[28]$_DFFE_PN__3340  (.L_HI(net3340));
 sg13g2_tiehi \cpu.intr.r_clock_count[29]$_DFFE_PN__3341  (.L_HI(net3341));
 sg13g2_tiehi \cpu.intr.r_clock_count[2]$_DFF_P__3342  (.L_HI(net3342));
 sg13g2_tiehi \cpu.intr.r_clock_count[30]$_DFFE_PN__3343  (.L_HI(net3343));
 sg13g2_tiehi \cpu.intr.r_clock_count[31]$_DFFE_PN__3344  (.L_HI(net3344));
 sg13g2_tiehi \cpu.intr.r_clock_count[3]$_DFF_P__3345  (.L_HI(net3345));
 sg13g2_tiehi \cpu.intr.r_clock_count[4]$_DFF_P__3346  (.L_HI(net3346));
 sg13g2_tiehi \cpu.intr.r_clock_count[5]$_DFF_P__3347  (.L_HI(net3347));
 sg13g2_tiehi \cpu.intr.r_clock_count[6]$_DFF_P__3348  (.L_HI(net3348));
 sg13g2_tiehi \cpu.intr.r_clock_count[7]$_DFF_P__3349  (.L_HI(net3349));
 sg13g2_tiehi \cpu.intr.r_clock_count[8]$_DFF_P__3350  (.L_HI(net3350));
 sg13g2_tiehi \cpu.intr.r_clock_count[9]$_DFF_P__3351  (.L_HI(net3351));
 sg13g2_tiehi \cpu.intr.r_enable[0]$_SDFFE_PN0P__3352  (.L_HI(net3352));
 sg13g2_tiehi \cpu.intr.r_enable[1]$_SDFFE_PN0P__3353  (.L_HI(net3353));
 sg13g2_tiehi \cpu.intr.r_enable[2]$_SDFFE_PN0P__3354  (.L_HI(net3354));
 sg13g2_tiehi \cpu.intr.r_enable[3]$_SDFFE_PN0P__3355  (.L_HI(net3355));
 sg13g2_tiehi \cpu.intr.r_enable[4]$_SDFFE_PN0P__3356  (.L_HI(net3356));
 sg13g2_tiehi \cpu.intr.r_enable[5]$_SDFFE_PN0P__3357  (.L_HI(net3357));
 sg13g2_tiehi \cpu.intr.r_timer$_SDFFE_PN0P__3358  (.L_HI(net3358));
 sg13g2_tiehi \cpu.intr.r_timer_count[0]$_DFF_P__3359  (.L_HI(net3359));
 sg13g2_tiehi \cpu.intr.r_timer_count[10]$_DFF_P__3360  (.L_HI(net3360));
 sg13g2_tiehi \cpu.intr.r_timer_count[11]$_DFF_P__3361  (.L_HI(net3361));
 sg13g2_tiehi \cpu.intr.r_timer_count[12]$_DFF_P__3362  (.L_HI(net3362));
 sg13g2_tiehi \cpu.intr.r_timer_count[13]$_DFF_P__3363  (.L_HI(net3363));
 sg13g2_tiehi \cpu.intr.r_timer_count[14]$_DFF_P__3364  (.L_HI(net3364));
 sg13g2_tiehi \cpu.intr.r_timer_count[15]$_DFF_P__3365  (.L_HI(net3365));
 sg13g2_tiehi \cpu.intr.r_timer_count[16]$_DFF_P__3366  (.L_HI(net3366));
 sg13g2_tiehi \cpu.intr.r_timer_count[17]$_DFF_P__3367  (.L_HI(net3367));
 sg13g2_tiehi \cpu.intr.r_timer_count[18]$_DFF_P__3368  (.L_HI(net3368));
 sg13g2_tiehi \cpu.intr.r_timer_count[19]$_DFF_P__3369  (.L_HI(net3369));
 sg13g2_tiehi \cpu.intr.r_timer_count[1]$_DFF_P__3370  (.L_HI(net3370));
 sg13g2_tiehi \cpu.intr.r_timer_count[20]$_DFF_P__3371  (.L_HI(net3371));
 sg13g2_tiehi \cpu.intr.r_timer_count[21]$_DFF_P__3372  (.L_HI(net3372));
 sg13g2_tiehi \cpu.intr.r_timer_count[22]$_DFF_P__3373  (.L_HI(net3373));
 sg13g2_tiehi \cpu.intr.r_timer_count[23]$_DFF_P__3374  (.L_HI(net3374));
 sg13g2_tiehi \cpu.intr.r_timer_count[2]$_DFF_P__3375  (.L_HI(net3375));
 sg13g2_tiehi \cpu.intr.r_timer_count[3]$_DFF_P__3376  (.L_HI(net3376));
 sg13g2_tiehi \cpu.intr.r_timer_count[4]$_DFF_P__3377  (.L_HI(net3377));
 sg13g2_tiehi \cpu.intr.r_timer_count[5]$_DFF_P__3378  (.L_HI(net3378));
 sg13g2_tiehi \cpu.intr.r_timer_count[6]$_DFF_P__3379  (.L_HI(net3379));
 sg13g2_tiehi \cpu.intr.r_timer_count[7]$_DFF_P__3380  (.L_HI(net3380));
 sg13g2_tiehi \cpu.intr.r_timer_count[8]$_DFF_P__3381  (.L_HI(net3381));
 sg13g2_tiehi \cpu.intr.r_timer_count[9]$_DFF_P__3382  (.L_HI(net3382));
 sg13g2_tiehi \cpu.intr.r_timer_reload[0]$_DFFE_PP__3383  (.L_HI(net3383));
 sg13g2_tiehi \cpu.intr.r_timer_reload[10]$_DFFE_PP__3384  (.L_HI(net3384));
 sg13g2_tiehi \cpu.intr.r_timer_reload[11]$_DFFE_PP__3385  (.L_HI(net3385));
 sg13g2_tiehi \cpu.intr.r_timer_reload[12]$_DFFE_PP__3386  (.L_HI(net3386));
 sg13g2_tiehi \cpu.intr.r_timer_reload[13]$_DFFE_PP__3387  (.L_HI(net3387));
 sg13g2_tiehi \cpu.intr.r_timer_reload[14]$_DFFE_PP__3388  (.L_HI(net3388));
 sg13g2_tiehi \cpu.intr.r_timer_reload[15]$_DFFE_PP__3389  (.L_HI(net3389));
 sg13g2_tiehi \cpu.intr.r_timer_reload[16]$_DFFE_PP__3390  (.L_HI(net3390));
 sg13g2_tiehi \cpu.intr.r_timer_reload[17]$_DFFE_PP__3391  (.L_HI(net3391));
 sg13g2_tiehi \cpu.intr.r_timer_reload[18]$_DFFE_PP__3392  (.L_HI(net3392));
 sg13g2_tiehi \cpu.intr.r_timer_reload[19]$_DFFE_PP__3393  (.L_HI(net3393));
 sg13g2_tiehi \cpu.intr.r_timer_reload[1]$_DFFE_PP__3394  (.L_HI(net3394));
 sg13g2_tiehi \cpu.intr.r_timer_reload[20]$_DFFE_PP__3395  (.L_HI(net3395));
 sg13g2_tiehi \cpu.intr.r_timer_reload[21]$_DFFE_PP__3396  (.L_HI(net3396));
 sg13g2_tiehi \cpu.intr.r_timer_reload[22]$_DFFE_PP__3397  (.L_HI(net3397));
 sg13g2_tiehi \cpu.intr.r_timer_reload[23]$_DFFE_PP__3398  (.L_HI(net3398));
 sg13g2_tiehi \cpu.intr.r_timer_reload[2]$_DFFE_PP__3399  (.L_HI(net3399));
 sg13g2_tiehi \cpu.intr.r_timer_reload[3]$_DFFE_PP__3400  (.L_HI(net3400));
 sg13g2_tiehi \cpu.intr.r_timer_reload[4]$_DFFE_PP__3401  (.L_HI(net3401));
 sg13g2_tiehi \cpu.intr.r_timer_reload[5]$_DFFE_PP__3402  (.L_HI(net3402));
 sg13g2_tiehi \cpu.intr.r_timer_reload[6]$_DFFE_PP__3403  (.L_HI(net3403));
 sg13g2_tiehi \cpu.intr.r_timer_reload[7]$_DFFE_PP__3404  (.L_HI(net3404));
 sg13g2_tiehi \cpu.intr.r_timer_reload[8]$_DFFE_PP__3405  (.L_HI(net3405));
 sg13g2_tiehi \cpu.intr.r_timer_reload[9]$_DFFE_PP__3406  (.L_HI(net3406));
 sg13g2_tiehi \cpu.qspi.r_count[0]$_DFFE_PP__3407  (.L_HI(net3407));
 sg13g2_tiehi \cpu.qspi.r_count[1]$_DFFE_PP__3408  (.L_HI(net3408));
 sg13g2_tiehi \cpu.qspi.r_count[2]$_DFFE_PP__3409  (.L_HI(net3409));
 sg13g2_tiehi \cpu.qspi.r_count[3]$_DFFE_PP__3410  (.L_HI(net3410));
 sg13g2_tiehi \cpu.qspi.r_count[4]$_DFFE_PP__3411  (.L_HI(net3411));
 sg13g2_tiehi \cpu.qspi.r_cs[0]$_SDFFE_PN1P__3412  (.L_HI(net3412));
 sg13g2_tiehi \cpu.qspi.r_cs[1]$_SDFFE_PN1P__3413  (.L_HI(net3413));
 sg13g2_tiehi \cpu.qspi.r_cs[2]$_SDFFE_PN1P__3414  (.L_HI(net3414));
 sg13g2_tiehi \cpu.qspi.r_ind$_SDFFE_PN0N__3415  (.L_HI(net3415));
 sg13g2_tiehi \cpu.qspi.r_mask[0]$_SDFFE_PN0P__3416  (.L_HI(net3416));
 sg13g2_tiehi \cpu.qspi.r_mask[1]$_SDFFE_PN1P__3417  (.L_HI(net3417));
 sg13g2_tiehi \cpu.qspi.r_mask[2]$_SDFFE_PN0P__3418  (.L_HI(net3418));
 sg13g2_tiehi \cpu.qspi.r_quad[0]$_SDFFE_PN1P__3419  (.L_HI(net3419));
 sg13g2_tiehi \cpu.qspi.r_quad[1]$_SDFFE_PN0P__3420  (.L_HI(net3420));
 sg13g2_tiehi \cpu.qspi.r_quad[2]$_SDFFE_PN1P__3421  (.L_HI(net3421));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][0]$_SDFFCE_PN0P__3422  (.L_HI(net3422));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][1]$_SDFFCE_PN0P__3423  (.L_HI(net3423));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][2]$_SDFFCE_PN1P__3424  (.L_HI(net3424));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][3]$_SDFFCE_PN0P__3425  (.L_HI(net3425));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][0]$_SDFFCE_PN0P__3426  (.L_HI(net3426));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][1]$_SDFFCE_PN0P__3427  (.L_HI(net3427));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][2]$_SDFFCE_PN1P__3428  (.L_HI(net3428));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][3]$_SDFFCE_PN0P__3429  (.L_HI(net3429));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][0]$_SDFFCE_PN0P__3430  (.L_HI(net3430));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][1]$_SDFFCE_PN0P__3431  (.L_HI(net3431));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][2]$_SDFFCE_PN1P__3432  (.L_HI(net3432));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][3]$_SDFFCE_PN0P__3433  (.L_HI(net3433));
 sg13g2_tiehi \cpu.qspi.r_rom_mode[0]$_SDFFE_PN1P__3434  (.L_HI(net3434));
 sg13g2_tiehi \cpu.qspi.r_rom_mode[1]$_SDFFE_PN1P__3435  (.L_HI(net3435));
 sg13g2_tiehi \cpu.qspi.r_rstrobe_d$_DFF_P__3436  (.L_HI(net3436));
 sg13g2_tiehi \cpu.qspi.r_state[0]$_DFF_P__3437  (.L_HI(net3437));
 sg13g2_tiehi \cpu.qspi.r_state[10]$_DFF_P__3438  (.L_HI(net3438));
 sg13g2_tiehi \cpu.qspi.r_state[11]$_DFF_P__3439  (.L_HI(net3439));
 sg13g2_tiehi \cpu.qspi.r_state[12]$_DFF_P__3440  (.L_HI(net3440));
 sg13g2_tiehi \cpu.qspi.r_state[13]$_DFF_P__3441  (.L_HI(net3441));
 sg13g2_tiehi \cpu.qspi.r_state[14]$_DFF_P__3442  (.L_HI(net3442));
 sg13g2_tiehi \cpu.qspi.r_state[15]$_DFF_P__3443  (.L_HI(net3443));
 sg13g2_tiehi \cpu.qspi.r_state[16]$_DFF_P__3444  (.L_HI(net3444));
 sg13g2_tiehi \cpu.qspi.r_state[17]$_DFF_P__3445  (.L_HI(net3445));
 sg13g2_tiehi \cpu.qspi.r_state[1]$_DFF_P__3446  (.L_HI(net3446));
 sg13g2_tiehi \cpu.qspi.r_state[2]$_DFF_P__3447  (.L_HI(net3447));
 sg13g2_tiehi \cpu.qspi.r_state[3]$_DFF_P__3448  (.L_HI(net3448));
 sg13g2_tiehi \cpu.qspi.r_state[4]$_DFF_P__3449  (.L_HI(net3449));
 sg13g2_tiehi \cpu.qspi.r_state[5]$_DFF_P__3450  (.L_HI(net3450));
 sg13g2_tiehi \cpu.qspi.r_state[6]$_DFF_P__3451  (.L_HI(net3451));
 sg13g2_tiehi \cpu.qspi.r_state[7]$_DFF_P__3452  (.L_HI(net3452));
 sg13g2_tiehi \cpu.qspi.r_state[8]$_DFF_P__3453  (.L_HI(net3453));
 sg13g2_tiehi \cpu.qspi.r_state[9]$_DFF_P__3454  (.L_HI(net3454));
 sg13g2_tiehi \cpu.qspi.r_uio_oe[0]$_SDFFE_PN0P__3455  (.L_HI(net3455));
 sg13g2_tiehi \cpu.qspi.r_uio_oe[1]$_SDFFE_PN0P__3456  (.L_HI(net3456));
 sg13g2_tiehi \cpu.qspi.r_uio_out[0]$_DFFE_PP__3457  (.L_HI(net3457));
 sg13g2_tiehi \cpu.qspi.r_uio_out[1]$_DFFE_PP__3458  (.L_HI(net3458));
 sg13g2_tiehi \cpu.qspi.r_uio_out[2]$_DFFE_PP__3459  (.L_HI(net3459));
 sg13g2_tiehi \cpu.qspi.r_uio_out[3]$_DFFE_PP__3460  (.L_HI(net3460));
 sg13g2_tiehi \cpu.qspi.r_wstrobe_d$_DFF_P__3461  (.L_HI(net3461));
 sg13g2_tiehi \cpu.qspi.r_wstrobe_i$_DFF_P__3462  (.L_HI(net3462));
 sg13g2_tiehi \cpu.r_clk_invert$_DFFE_PN__3463  (.L_HI(net3463));
 sg13g2_tiehi \cpu.spi.r_bits[0]$_SDFFE_PN1P__3464  (.L_HI(net3464));
 sg13g2_tiehi \cpu.spi.r_bits[1]$_SDFFE_PN1P__3465  (.L_HI(net3465));
 sg13g2_tiehi \cpu.spi.r_bits[2]$_SDFFE_PN1P__3466  (.L_HI(net3466));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][0]$_SDFFE_PN0P__3467  (.L_HI(net3467));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][1]$_SDFFE_PN0P__3468  (.L_HI(net3468));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][2]$_SDFFE_PN0P__3469  (.L_HI(net3469));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][3]$_SDFFE_PN0P__3470  (.L_HI(net3470));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][4]$_SDFFE_PN0P__3471  (.L_HI(net3471));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][5]$_SDFFE_PN0P__3472  (.L_HI(net3472));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][6]$_SDFFE_PN0P__3473  (.L_HI(net3473));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][7]$_SDFFE_PN0P__3474  (.L_HI(net3474));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][0]$_SDFFE_PN0P__3475  (.L_HI(net3475));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][1]$_SDFFE_PN0P__3476  (.L_HI(net3476));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][2]$_SDFFE_PN0P__3477  (.L_HI(net3477));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][3]$_SDFFE_PN0P__3478  (.L_HI(net3478));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][4]$_SDFFE_PN0P__3479  (.L_HI(net3479));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][5]$_SDFFE_PN0P__3480  (.L_HI(net3480));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][6]$_SDFFE_PN0P__3481  (.L_HI(net3481));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][7]$_SDFFE_PN0P__3482  (.L_HI(net3482));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][0]$_SDFFE_PN0P__3483  (.L_HI(net3483));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][1]$_SDFFE_PN0P__3484  (.L_HI(net3484));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][2]$_SDFFE_PN0P__3485  (.L_HI(net3485));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][3]$_SDFFE_PN0P__3486  (.L_HI(net3486));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][4]$_SDFFE_PN0P__3487  (.L_HI(net3487));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][5]$_SDFFE_PN0P__3488  (.L_HI(net3488));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][6]$_SDFFE_PN0P__3489  (.L_HI(net3489));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][7]$_SDFFE_PN0P__3490  (.L_HI(net3490));
 sg13g2_tiehi \cpu.spi.r_count[0]$_SDFFE_PN0P__3491  (.L_HI(net3491));
 sg13g2_tiehi \cpu.spi.r_count[1]$_SDFFE_PN0P__3492  (.L_HI(net3492));
 sg13g2_tiehi \cpu.spi.r_count[2]$_SDFFE_PN0P__3493  (.L_HI(net3493));
 sg13g2_tiehi \cpu.spi.r_count[3]$_SDFFE_PN0P__3494  (.L_HI(net3494));
 sg13g2_tiehi \cpu.spi.r_count[4]$_SDFFE_PN0P__3495  (.L_HI(net3495));
 sg13g2_tiehi \cpu.spi.r_count[5]$_SDFFE_PN0P__3496  (.L_HI(net3496));
 sg13g2_tiehi \cpu.spi.r_count[6]$_SDFFE_PN0P__3497  (.L_HI(net3497));
 sg13g2_tiehi \cpu.spi.r_count[7]$_SDFFE_PN0P__3498  (.L_HI(net3498));
 sg13g2_tiehi \cpu.spi.r_cs[0]$_SDFFE_PN1P__3499  (.L_HI(net3499));
 sg13g2_tiehi \cpu.spi.r_cs[1]$_SDFFE_PN1P__3500  (.L_HI(net3500));
 sg13g2_tiehi \cpu.spi.r_cs[2]$_SDFFE_PN1P__3501  (.L_HI(net3501));
 sg13g2_tiehi \cpu.spi.r_in[0]$_DFFE_PP__3502  (.L_HI(net3502));
 sg13g2_tiehi \cpu.spi.r_in[1]$_DFFE_PP__3503  (.L_HI(net3503));
 sg13g2_tiehi \cpu.spi.r_in[2]$_DFFE_PP__3504  (.L_HI(net3504));
 sg13g2_tiehi \cpu.spi.r_in[3]$_DFFE_PP__3505  (.L_HI(net3505));
 sg13g2_tiehi \cpu.spi.r_in[4]$_DFFE_PP__3506  (.L_HI(net3506));
 sg13g2_tiehi \cpu.spi.r_in[5]$_DFFE_PP__3507  (.L_HI(net3507));
 sg13g2_tiehi \cpu.spi.r_in[6]$_DFFE_PP__3508  (.L_HI(net3508));
 sg13g2_tiehi \cpu.spi.r_in[7]$_DFFE_PP__3509  (.L_HI(net3509));
 sg13g2_tiehi \cpu.spi.r_interrupt$_SDFFE_PN0P__3510  (.L_HI(net3510));
 sg13g2_tiehi \cpu.spi.r_mode[0][0]$_SDFFE_PN0P__3511  (.L_HI(net3511));
 sg13g2_tiehi \cpu.spi.r_mode[0][1]$_SDFFE_PN0P__3512  (.L_HI(net3512));
 sg13g2_tiehi \cpu.spi.r_mode[1][0]$_SDFFE_PN0P__3513  (.L_HI(net3513));
 sg13g2_tiehi \cpu.spi.r_mode[1][1]$_SDFFE_PN0P__3514  (.L_HI(net3514));
 sg13g2_tiehi \cpu.spi.r_mode[2][0]$_SDFFE_PN0P__3515  (.L_HI(net3515));
 sg13g2_tiehi \cpu.spi.r_mode[2][1]$_SDFFE_PN0P__3516  (.L_HI(net3516));
 sg13g2_tiehi \cpu.spi.r_out[0]$_DFFE_PP__3517  (.L_HI(net3517));
 sg13g2_tiehi \cpu.spi.r_out[1]$_DFFE_PP__3518  (.L_HI(net3518));
 sg13g2_tiehi \cpu.spi.r_out[2]$_DFFE_PP__3519  (.L_HI(net3519));
 sg13g2_tiehi \cpu.spi.r_out[3]$_DFFE_PP__3520  (.L_HI(net3520));
 sg13g2_tiehi \cpu.spi.r_out[4]$_DFFE_PP__3521  (.L_HI(net3521));
 sg13g2_tiehi \cpu.spi.r_out[5]$_DFFE_PP__3522  (.L_HI(net3522));
 sg13g2_tiehi \cpu.spi.r_out[6]$_DFFE_PP__3523  (.L_HI(net3523));
 sg13g2_tiehi \cpu.spi.r_out[7]$_DFFE_PP__3524  (.L_HI(net3524));
 sg13g2_tiehi \cpu.spi.r_ready$_SDFFE_PN1P__3525  (.L_HI(net3525));
 sg13g2_tiehi \cpu.spi.r_searching$_SDFFE_PN0P__3526  (.L_HI(net3526));
 sg13g2_tiehi \cpu.spi.r_sel[0]$_DFFE_PP__3527  (.L_HI(net3527));
 sg13g2_tiehi \cpu.spi.r_sel[1]$_DFFE_PP__3528  (.L_HI(net3528));
 sg13g2_tiehi \cpu.spi.r_src[0]$_SDFFE_PN0P__3529  (.L_HI(net3529));
 sg13g2_tiehi \cpu.spi.r_src[1]$_SDFFE_PN0P__3530  (.L_HI(net3530));
 sg13g2_tiehi \cpu.spi.r_src[2]$_SDFFE_PN0P__3531  (.L_HI(net3531));
 sg13g2_tiehi \cpu.spi.r_state[0]$_DFF_P__3532  (.L_HI(net3532));
 sg13g2_tiehi \cpu.spi.r_state[1]$_DFF_P__3533  (.L_HI(net3533));
 sg13g2_tiehi \cpu.spi.r_state[2]$_DFF_P__3534  (.L_HI(net3534));
 sg13g2_tiehi \cpu.spi.r_state[3]$_DFF_P__3535  (.L_HI(net3535));
 sg13g2_tiehi \cpu.spi.r_state[4]$_DFF_P__3536  (.L_HI(net3536));
 sg13g2_tiehi \cpu.spi.r_state[5]$_DFF_P__3537  (.L_HI(net3537));
 sg13g2_tiehi \cpu.spi.r_state[6]$_DFF_P__3538  (.L_HI(net3538));
 sg13g2_tiehi \cpu.spi.r_timeout[0]$_DFFE_PP__3539  (.L_HI(net3539));
 sg13g2_tiehi \cpu.spi.r_timeout[1]$_DFFE_PP__3540  (.L_HI(net3540));
 sg13g2_tiehi \cpu.spi.r_timeout[2]$_DFFE_PP__3541  (.L_HI(net3541));
 sg13g2_tiehi \cpu.spi.r_timeout[3]$_DFFE_PP__3542  (.L_HI(net3542));
 sg13g2_tiehi \cpu.spi.r_timeout[4]$_DFFE_PP__3543  (.L_HI(net3543));
 sg13g2_tiehi \cpu.spi.r_timeout[5]$_DFFE_PP__3544  (.L_HI(net3544));
 sg13g2_tiehi \cpu.spi.r_timeout[6]$_DFFE_PP__3545  (.L_HI(net3545));
 sg13g2_tiehi \cpu.spi.r_timeout[7]$_DFFE_PP__3546  (.L_HI(net3546));
 sg13g2_tiehi \cpu.spi.r_timeout_count[0]$_DFFE_PP__3547  (.L_HI(net3547));
 sg13g2_tiehi \cpu.spi.r_timeout_count[1]$_DFFE_PP__3548  (.L_HI(net3548));
 sg13g2_tiehi \cpu.spi.r_timeout_count[2]$_DFFE_PP__3549  (.L_HI(net3549));
 sg13g2_tiehi \cpu.spi.r_timeout_count[3]$_DFFE_PP__3550  (.L_HI(net3550));
 sg13g2_tiehi \cpu.spi.r_timeout_count[4]$_DFFE_PP__3551  (.L_HI(net3551));
 sg13g2_tiehi \cpu.spi.r_timeout_count[5]$_DFFE_PP__3552  (.L_HI(net3552));
 sg13g2_tiehi \cpu.spi.r_timeout_count[6]$_DFFE_PP__3553  (.L_HI(net3553));
 sg13g2_tiehi \cpu.spi.r_timeout_count[7]$_DFFE_PP__3554  (.L_HI(net3554));
 sg13g2_tiehi \cpu.uart.r_div[0]$_DFF_P__3555  (.L_HI(net3555));
 sg13g2_tiehi \cpu.uart.r_div[10]$_DFF_P__3556  (.L_HI(net3556));
 sg13g2_tiehi \cpu.uart.r_div[11]$_DFF_P__3557  (.L_HI(net3557));
 sg13g2_tiehi \cpu.uart.r_div[1]$_DFF_P__3558  (.L_HI(net3558));
 sg13g2_tiehi \cpu.uart.r_div[2]$_DFF_P__3559  (.L_HI(net3559));
 sg13g2_tiehi \cpu.uart.r_div[3]$_DFF_P__3560  (.L_HI(net3560));
 sg13g2_tiehi \cpu.uart.r_div[4]$_DFF_P__3561  (.L_HI(net3561));
 sg13g2_tiehi \cpu.uart.r_div[5]$_DFF_P__3562  (.L_HI(net3562));
 sg13g2_tiehi \cpu.uart.r_div[6]$_DFF_P__3563  (.L_HI(net3563));
 sg13g2_tiehi \cpu.uart.r_div[7]$_DFF_P__3564  (.L_HI(net3564));
 sg13g2_tiehi \cpu.uart.r_div[8]$_DFF_P__3565  (.L_HI(net3565));
 sg13g2_tiehi \cpu.uart.r_div[9]$_DFF_P__3566  (.L_HI(net3566));
 sg13g2_tiehi \cpu.uart.r_div_value[0]$_SDFFE_PN1P__3567  (.L_HI(net3567));
 sg13g2_tiehi \cpu.uart.r_div_value[10]$_SDFFE_PN0P__3568  (.L_HI(net3568));
 sg13g2_tiehi \cpu.uart.r_div_value[11]$_SDFFE_PN0P__3569  (.L_HI(net3569));
 sg13g2_tiehi \cpu.uart.r_div_value[1]$_SDFFE_PN0P__3570  (.L_HI(net3570));
 sg13g2_tiehi \cpu.uart.r_div_value[2]$_SDFFE_PN0P__3571  (.L_HI(net3571));
 sg13g2_tiehi \cpu.uart.r_div_value[3]$_SDFFE_PN0P__3572  (.L_HI(net3572));
 sg13g2_tiehi \cpu.uart.r_div_value[4]$_SDFFE_PN0P__3573  (.L_HI(net3573));
 sg13g2_tiehi \cpu.uart.r_div_value[5]$_SDFFE_PN0P__3574  (.L_HI(net3574));
 sg13g2_tiehi \cpu.uart.r_div_value[6]$_SDFFE_PN0P__3575  (.L_HI(net3575));
 sg13g2_tiehi \cpu.uart.r_div_value[7]$_SDFFE_PN0P__3576  (.L_HI(net3576));
 sg13g2_tiehi \cpu.uart.r_div_value[8]$_SDFFE_PN0P__3577  (.L_HI(net3577));
 sg13g2_tiehi \cpu.uart.r_div_value[9]$_SDFFE_PN0P__3578  (.L_HI(net3578));
 sg13g2_tiehi \cpu.uart.r_ib[0]$_DFFE_PP__3579  (.L_HI(net3579));
 sg13g2_tiehi \cpu.uart.r_ib[1]$_DFFE_PP__3580  (.L_HI(net3580));
 sg13g2_tiehi \cpu.uart.r_ib[2]$_DFFE_PP__3581  (.L_HI(net3581));
 sg13g2_tiehi \cpu.uart.r_ib[3]$_DFFE_PP__3582  (.L_HI(net3582));
 sg13g2_tiehi \cpu.uart.r_ib[4]$_DFFE_PP__3583  (.L_HI(net3583));
 sg13g2_tiehi \cpu.uart.r_ib[5]$_DFFE_PP__3584  (.L_HI(net3584));
 sg13g2_tiehi \cpu.uart.r_ib[6]$_DFFE_PP__3585  (.L_HI(net3585));
 sg13g2_tiehi \cpu.uart.r_in[0]$_DFFE_PP__3586  (.L_HI(net3586));
 sg13g2_tiehi \cpu.uart.r_in[1]$_DFFE_PP__3587  (.L_HI(net3587));
 sg13g2_tiehi \cpu.uart.r_in[2]$_DFFE_PP__3588  (.L_HI(net3588));
 sg13g2_tiehi \cpu.uart.r_in[3]$_DFFE_PP__3589  (.L_HI(net3589));
 sg13g2_tiehi \cpu.uart.r_in[4]$_DFFE_PP__3590  (.L_HI(net3590));
 sg13g2_tiehi \cpu.uart.r_in[5]$_DFFE_PP__3591  (.L_HI(net3591));
 sg13g2_tiehi \cpu.uart.r_in[6]$_DFFE_PP__3592  (.L_HI(net3592));
 sg13g2_tiehi \cpu.uart.r_in[7]$_DFFE_PP__3593  (.L_HI(net3593));
 sg13g2_tiehi \cpu.uart.r_out[0]$_DFFE_PP__3594  (.L_HI(net3594));
 sg13g2_tiehi \cpu.uart.r_out[1]$_DFFE_PP__3595  (.L_HI(net3595));
 sg13g2_tiehi \cpu.uart.r_out[2]$_DFFE_PP__3596  (.L_HI(net3596));
 sg13g2_tiehi \cpu.uart.r_out[3]$_DFFE_PP__3597  (.L_HI(net3597));
 sg13g2_tiehi \cpu.uart.r_out[4]$_DFFE_PP__3598  (.L_HI(net3598));
 sg13g2_tiehi \cpu.uart.r_out[5]$_DFFE_PP__3599  (.L_HI(net3599));
 sg13g2_tiehi \cpu.uart.r_out[6]$_DFFE_PP__3600  (.L_HI(net3600));
 sg13g2_tiehi \cpu.uart.r_out[7]$_DFFE_PP__3601  (.L_HI(net3601));
 sg13g2_tiehi \cpu.uart.r_r$_DFF_P__3602  (.L_HI(net3602));
 sg13g2_tiehi \cpu.uart.r_r_int$_SDFFE_PN0P__3603  (.L_HI(net3603));
 sg13g2_tiehi \cpu.uart.r_r_invert$_SDFFE_PN0P__3604  (.L_HI(net3604));
 sg13g2_tiehi \cpu.uart.r_rcnt[0]$_DFFE_PP__3605  (.L_HI(net3605));
 sg13g2_tiehi \cpu.uart.r_rcnt[1]$_DFFE_PP__3606  (.L_HI(net3606));
 sg13g2_tiehi \cpu.uart.r_rstate[0]$_SDFFE_PN0P__3607  (.L_HI(net3607));
 sg13g2_tiehi \cpu.uart.r_rstate[1]$_SDFFE_PN0P__3608  (.L_HI(net3608));
 sg13g2_tiehi \cpu.uart.r_rstate[2]$_SDFFE_PN0P__3609  (.L_HI(net3609));
 sg13g2_tiehi \cpu.uart.r_rstate[3]$_SDFFE_PN0P__3610  (.L_HI(net3610));
 sg13g2_tiehi \cpu.uart.r_x$_DFFE_PP__3611  (.L_HI(net3611));
 sg13g2_tiehi \cpu.uart.r_x_int$_SDFFE_PN0P__3612  (.L_HI(net3612));
 sg13g2_tiehi \cpu.uart.r_x_invert$_SDFFE_PN0P__3613  (.L_HI(net3613));
 sg13g2_tiehi \cpu.uart.r_xcnt[0]$_DFFE_PP__3614  (.L_HI(net3614));
 sg13g2_tiehi \cpu.uart.r_xcnt[1]$_DFFE_PP__3615  (.L_HI(net3615));
 sg13g2_tiehi \cpu.uart.r_xstate[0]$_SDFFE_PN0P__3616  (.L_HI(net3616));
 sg13g2_tiehi \cpu.uart.r_xstate[1]$_SDFFE_PN0P__3617  (.L_HI(net3617));
 sg13g2_tiehi \cpu.uart.r_xstate[2]$_SDFFE_PN0P__3618  (.L_HI(net3618));
 sg13g2_tiehi \cpu.uart.r_xstate[3]$_SDFFE_PN0P__3619  (.L_HI(net3619));
 sg13g2_tiehi \r_reset$_DFF_P__3620  (.L_HI(net3620));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_8 clkbuf_leaf_78_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_8 clkbuf_leaf_79_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_8 clkbuf_leaf_80_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_8 clkbuf_leaf_81_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_8 clkbuf_leaf_82_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_8 clkbuf_leaf_83_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_8 clkbuf_leaf_84_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_8 clkbuf_leaf_85_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_8 clkbuf_leaf_86_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_8 clkbuf_leaf_87_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_8 clkbuf_leaf_88_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_8 clkbuf_leaf_89_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_8 clkbuf_leaf_90_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_8 clkbuf_leaf_91_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_8 clkbuf_leaf_92_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_8 clkbuf_leaf_93_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_8 clkbuf_leaf_94_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_8 clkbuf_leaf_95_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_8 clkbuf_leaf_96_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_8 clkbuf_leaf_97_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_8 clkbuf_leaf_98_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_8 clkbuf_leaf_99_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_8 clkbuf_leaf_100_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_8 clkbuf_leaf_101_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_8 clkbuf_leaf_102_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_8 clkbuf_leaf_103_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_8 clkbuf_leaf_104_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_8 clkbuf_leaf_105_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_8 clkbuf_leaf_106_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_8 clkbuf_leaf_107_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_8 clkbuf_leaf_108_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_8 clkbuf_leaf_109_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_8 clkbuf_leaf_110_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_8 clkbuf_leaf_111_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_8 clkbuf_leaf_112_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_8 clkbuf_leaf_113_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_8 clkbuf_leaf_114_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_8 clkbuf_leaf_115_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_8 clkbuf_leaf_116_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_8 clkbuf_leaf_117_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_8 clkbuf_leaf_118_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_8 clkbuf_leaf_119_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_8 clkbuf_leaf_120_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_8 clkbuf_leaf_121_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_8 clkbuf_leaf_122_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_8 clkbuf_leaf_123_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_8 clkbuf_leaf_124_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_8 clkbuf_leaf_125_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_8 clkbuf_leaf_126_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_8 clkbuf_leaf_127_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_8 clkbuf_leaf_128_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_8 clkbuf_leaf_129_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_8 clkbuf_leaf_130_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_8 clkbuf_leaf_131_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_8 clkbuf_leaf_132_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_8 clkbuf_leaf_133_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_8 clkbuf_leaf_134_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_8 clkbuf_leaf_135_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_8 clkbuf_leaf_136_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_8 clkbuf_leaf_137_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_8 clkbuf_leaf_138_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_8 clkbuf_leaf_139_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_8 clkbuf_leaf_140_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_8 clkbuf_leaf_141_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_8 clkbuf_leaf_142_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_8 clkbuf_leaf_143_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_8 clkbuf_leaf_144_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_144_clk));
 sg13g2_buf_8 clkbuf_leaf_145_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_8 clkbuf_leaf_146_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_146_clk));
 sg13g2_buf_8 clkbuf_leaf_147_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_147_clk));
 sg13g2_buf_8 clkbuf_leaf_148_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_148_clk));
 sg13g2_buf_8 clkbuf_leaf_149_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_149_clk));
 sg13g2_buf_8 clkbuf_leaf_150_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_150_clk));
 sg13g2_buf_8 clkbuf_leaf_151_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_151_clk));
 sg13g2_buf_8 clkbuf_leaf_152_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_152_clk));
 sg13g2_buf_8 clkbuf_leaf_153_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_153_clk));
 sg13g2_buf_8 clkbuf_leaf_154_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_154_clk));
 sg13g2_buf_8 clkbuf_leaf_155_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_155_clk));
 sg13g2_buf_8 clkbuf_leaf_156_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_156_clk));
 sg13g2_buf_8 clkbuf_leaf_157_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_157_clk));
 sg13g2_buf_8 clkbuf_leaf_158_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_158_clk));
 sg13g2_buf_8 clkbuf_leaf_159_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_159_clk));
 sg13g2_buf_8 clkbuf_leaf_160_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_160_clk));
 sg13g2_buf_8 clkbuf_leaf_161_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_161_clk));
 sg13g2_buf_8 clkbuf_leaf_162_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_162_clk));
 sg13g2_buf_8 clkbuf_leaf_163_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_163_clk));
 sg13g2_buf_8 clkbuf_leaf_164_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_164_clk));
 sg13g2_buf_8 clkbuf_leaf_165_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_165_clk));
 sg13g2_buf_8 clkbuf_leaf_166_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_166_clk));
 sg13g2_buf_8 clkbuf_leaf_167_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_167_clk));
 sg13g2_buf_8 clkbuf_leaf_168_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_168_clk));
 sg13g2_buf_8 clkbuf_leaf_169_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_169_clk));
 sg13g2_buf_8 clkbuf_leaf_170_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_170_clk));
 sg13g2_buf_8 clkbuf_leaf_171_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_171_clk));
 sg13g2_buf_8 clkbuf_leaf_172_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_172_clk));
 sg13g2_buf_8 clkbuf_leaf_173_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_173_clk));
 sg13g2_buf_8 clkbuf_leaf_174_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_174_clk));
 sg13g2_buf_8 clkbuf_leaf_175_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_175_clk));
 sg13g2_buf_8 clkbuf_leaf_176_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_176_clk));
 sg13g2_buf_8 clkbuf_leaf_177_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_177_clk));
 sg13g2_buf_8 clkbuf_leaf_178_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_178_clk));
 sg13g2_buf_8 clkbuf_leaf_179_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_179_clk));
 sg13g2_buf_8 clkbuf_leaf_180_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_180_clk));
 sg13g2_buf_8 clkbuf_leaf_181_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_181_clk));
 sg13g2_buf_8 clkbuf_leaf_182_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_182_clk));
 sg13g2_buf_8 clkbuf_leaf_183_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_183_clk));
 sg13g2_buf_8 clkbuf_leaf_184_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_184_clk));
 sg13g2_buf_8 clkbuf_leaf_185_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_185_clk));
 sg13g2_buf_8 clkbuf_leaf_186_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_186_clk));
 sg13g2_buf_8 clkbuf_leaf_187_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_187_clk));
 sg13g2_buf_8 clkbuf_leaf_188_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_188_clk));
 sg13g2_buf_8 clkbuf_leaf_189_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_189_clk));
 sg13g2_buf_8 clkbuf_leaf_190_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_190_clk));
 sg13g2_buf_8 clkbuf_leaf_191_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_191_clk));
 sg13g2_buf_8 clkbuf_leaf_192_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_192_clk));
 sg13g2_buf_8 clkbuf_leaf_193_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_193_clk));
 sg13g2_buf_8 clkbuf_leaf_194_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_194_clk));
 sg13g2_buf_8 clkbuf_leaf_195_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_195_clk));
 sg13g2_buf_8 clkbuf_leaf_196_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_196_clk));
 sg13g2_buf_8 clkbuf_leaf_197_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_197_clk));
 sg13g2_buf_8 clkbuf_leaf_198_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_198_clk));
 sg13g2_buf_8 clkbuf_leaf_199_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_199_clk));
 sg13g2_buf_8 clkbuf_leaf_200_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_200_clk));
 sg13g2_buf_8 clkbuf_leaf_201_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_201_clk));
 sg13g2_buf_8 clkbuf_leaf_202_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_202_clk));
 sg13g2_buf_8 clkbuf_leaf_203_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_203_clk));
 sg13g2_buf_8 clkbuf_leaf_204_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_204_clk));
 sg13g2_buf_8 clkbuf_leaf_205_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_205_clk));
 sg13g2_buf_8 clkbuf_leaf_206_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_206_clk));
 sg13g2_buf_8 clkbuf_leaf_207_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_207_clk));
 sg13g2_buf_8 clkbuf_leaf_208_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_208_clk));
 sg13g2_buf_8 clkbuf_leaf_209_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_209_clk));
 sg13g2_buf_8 clkbuf_leaf_210_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_210_clk));
 sg13g2_buf_8 clkbuf_leaf_211_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_211_clk));
 sg13g2_buf_8 clkbuf_leaf_212_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_212_clk));
 sg13g2_buf_8 clkbuf_leaf_213_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_213_clk));
 sg13g2_buf_8 clkbuf_leaf_214_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_214_clk));
 sg13g2_buf_8 clkbuf_leaf_215_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_215_clk));
 sg13g2_buf_8 clkbuf_leaf_216_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_216_clk));
 sg13g2_buf_8 clkbuf_leaf_217_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_217_clk));
 sg13g2_buf_8 clkbuf_leaf_218_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_218_clk));
 sg13g2_buf_8 clkbuf_leaf_219_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_219_clk));
 sg13g2_buf_8 clkbuf_leaf_220_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_220_clk));
 sg13g2_buf_8 clkbuf_leaf_221_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_221_clk));
 sg13g2_buf_8 clkbuf_leaf_222_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_222_clk));
 sg13g2_buf_8 clkbuf_leaf_223_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_223_clk));
 sg13g2_buf_8 clkbuf_leaf_224_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_224_clk));
 sg13g2_buf_8 clkbuf_leaf_225_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_225_clk));
 sg13g2_buf_8 clkbuf_leaf_226_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_226_clk));
 sg13g2_buf_8 clkbuf_leaf_227_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_227_clk));
 sg13g2_buf_8 clkbuf_leaf_228_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_228_clk));
 sg13g2_buf_8 clkbuf_leaf_229_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_229_clk));
 sg13g2_buf_8 clkbuf_leaf_230_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_230_clk));
 sg13g2_buf_8 clkbuf_leaf_231_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_231_clk));
 sg13g2_buf_8 clkbuf_leaf_232_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_232_clk));
 sg13g2_buf_8 clkbuf_leaf_233_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_233_clk));
 sg13g2_buf_8 clkbuf_leaf_234_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_234_clk));
 sg13g2_buf_8 clkbuf_leaf_235_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_235_clk));
 sg13g2_buf_8 clkbuf_leaf_236_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_236_clk));
 sg13g2_buf_8 clkbuf_leaf_237_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_237_clk));
 sg13g2_buf_8 clkbuf_leaf_238_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_238_clk));
 sg13g2_buf_8 clkbuf_leaf_239_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_239_clk));
 sg13g2_buf_8 clkbuf_leaf_240_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_240_clk));
 sg13g2_buf_8 clkbuf_leaf_241_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_241_clk));
 sg13g2_buf_8 clkbuf_leaf_242_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_242_clk));
 sg13g2_buf_8 clkbuf_leaf_243_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_243_clk));
 sg13g2_buf_8 clkbuf_leaf_244_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_244_clk));
 sg13g2_buf_8 clkbuf_leaf_245_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_245_clk));
 sg13g2_buf_8 clkbuf_leaf_246_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_246_clk));
 sg13g2_buf_8 clkbuf_leaf_247_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_247_clk));
 sg13g2_buf_8 clkbuf_leaf_248_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_248_clk));
 sg13g2_buf_8 clkbuf_leaf_249_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_249_clk));
 sg13g2_buf_8 clkbuf_leaf_250_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_250_clk));
 sg13g2_buf_8 clkbuf_leaf_251_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_251_clk));
 sg13g2_buf_8 clkbuf_leaf_252_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_252_clk));
 sg13g2_buf_8 clkbuf_leaf_253_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_253_clk));
 sg13g2_buf_8 clkbuf_leaf_254_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_254_clk));
 sg13g2_buf_8 clkbuf_leaf_255_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_255_clk));
 sg13g2_buf_8 clkbuf_leaf_256_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_256_clk));
 sg13g2_buf_8 clkbuf_leaf_257_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_257_clk));
 sg13g2_buf_8 clkbuf_leaf_258_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_258_clk));
 sg13g2_buf_8 clkbuf_leaf_259_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_259_clk));
 sg13g2_buf_8 clkbuf_leaf_260_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_260_clk));
 sg13g2_buf_8 clkbuf_leaf_261_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_261_clk));
 sg13g2_buf_8 clkbuf_leaf_262_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_262_clk));
 sg13g2_buf_8 clkbuf_leaf_263_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_263_clk));
 sg13g2_buf_8 clkbuf_leaf_264_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_264_clk));
 sg13g2_buf_8 clkbuf_leaf_265_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_265_clk));
 sg13g2_buf_8 clkbuf_leaf_266_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_266_clk));
 sg13g2_buf_8 clkbuf_leaf_267_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_267_clk));
 sg13g2_buf_8 clkbuf_leaf_268_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_268_clk));
 sg13g2_buf_8 clkbuf_leaf_269_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_269_clk));
 sg13g2_buf_8 clkbuf_leaf_270_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_270_clk));
 sg13g2_buf_8 clkbuf_leaf_271_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_271_clk));
 sg13g2_buf_8 clkbuf_leaf_272_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_272_clk));
 sg13g2_buf_8 clkbuf_leaf_273_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_273_clk));
 sg13g2_buf_8 clkbuf_leaf_274_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_274_clk));
 sg13g2_buf_8 clkbuf_leaf_275_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_275_clk));
 sg13g2_buf_8 clkbuf_leaf_276_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_276_clk));
 sg13g2_buf_8 clkbuf_leaf_277_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_277_clk));
 sg13g2_buf_8 clkbuf_leaf_278_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_278_clk));
 sg13g2_buf_8 clkbuf_leaf_279_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_279_clk));
 sg13g2_buf_8 clkbuf_leaf_280_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_280_clk));
 sg13g2_buf_8 clkbuf_leaf_281_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_281_clk));
 sg13g2_buf_8 clkbuf_leaf_282_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_282_clk));
 sg13g2_buf_8 clkbuf_leaf_283_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_283_clk));
 sg13g2_buf_8 clkbuf_leaf_284_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_284_clk));
 sg13g2_buf_8 clkbuf_leaf_285_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_285_clk));
 sg13g2_buf_8 clkbuf_leaf_286_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_286_clk));
 sg13g2_buf_8 clkbuf_leaf_287_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_287_clk));
 sg13g2_buf_8 clkbuf_leaf_288_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_288_clk));
 sg13g2_buf_8 clkbuf_leaf_289_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_289_clk));
 sg13g2_buf_8 clkbuf_leaf_290_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_290_clk));
 sg13g2_buf_8 clkbuf_leaf_291_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_291_clk));
 sg13g2_buf_8 clkbuf_leaf_292_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_292_clk));
 sg13g2_buf_8 clkbuf_leaf_293_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_293_clk));
 sg13g2_buf_8 clkbuf_leaf_294_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_294_clk));
 sg13g2_buf_8 clkbuf_leaf_295_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_295_clk));
 sg13g2_buf_8 clkbuf_leaf_296_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_296_clk));
 sg13g2_buf_8 clkbuf_leaf_297_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_297_clk));
 sg13g2_buf_8 clkbuf_leaf_298_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_298_clk));
 sg13g2_buf_8 clkbuf_leaf_299_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_299_clk));
 sg13g2_buf_8 clkbuf_leaf_300_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_300_clk));
 sg13g2_buf_8 clkbuf_leaf_301_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_301_clk));
 sg13g2_buf_8 clkbuf_leaf_302_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_302_clk));
 sg13g2_buf_8 clkbuf_leaf_303_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_303_clk));
 sg13g2_buf_8 clkbuf_leaf_304_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_304_clk));
 sg13g2_buf_8 clkbuf_leaf_305_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_305_clk));
 sg13g2_buf_8 clkbuf_leaf_306_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_306_clk));
 sg13g2_buf_8 clkbuf_leaf_307_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_307_clk));
 sg13g2_buf_8 clkbuf_leaf_308_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_308_clk));
 sg13g2_buf_8 clkbuf_leaf_309_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_309_clk));
 sg13g2_buf_8 clkbuf_leaf_310_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_310_clk));
 sg13g2_buf_4 clkbuf_0_clk (.X(clknet_0_clk),
    .A(clk));
 sg13g2_buf_8 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sg13g2_buf_8 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sg13g2_buf_8 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sg13g2_buf_8 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sg13g2_buf_8 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sg13g2_buf_8 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sg13g2_buf_8 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sg13g2_buf_8 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_0__f_clk (.X(clknet_6_0__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_1__f_clk (.X(clknet_6_1__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_2__f_clk (.X(clknet_6_2__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_3__f_clk (.X(clknet_6_3__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_4__f_clk (.X(clknet_6_4__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_5__f_clk (.X(clknet_6_5__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_6__f_clk (.X(clknet_6_6__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_7__f_clk (.X(clknet_6_7__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_8__f_clk (.X(clknet_6_8__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_9__f_clk (.X(clknet_6_9__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_10__f_clk (.X(clknet_6_10__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_11__f_clk (.X(clknet_6_11__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_12__f_clk (.X(clknet_6_12__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_13__f_clk (.X(clknet_6_13__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_14__f_clk (.X(clknet_6_14__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_15__f_clk (.X(clknet_6_15__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_16__f_clk (.X(clknet_6_16__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_17__f_clk (.X(clknet_6_17__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_18__f_clk (.X(clknet_6_18__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_19__f_clk (.X(clknet_6_19__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_20__f_clk (.X(clknet_6_20__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_21__f_clk (.X(clknet_6_21__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_22__f_clk (.X(clknet_6_22__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_23__f_clk (.X(clknet_6_23__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_24__f_clk (.X(clknet_6_24__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_25__f_clk (.X(clknet_6_25__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_26__f_clk (.X(clknet_6_26__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_27__f_clk (.X(clknet_6_27__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_28__f_clk (.X(clknet_6_28__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_29__f_clk (.X(clknet_6_29__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_30__f_clk (.X(clknet_6_30__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_31__f_clk (.X(clknet_6_31__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_32__f_clk (.X(clknet_6_32__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_33__f_clk (.X(clknet_6_33__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_34__f_clk (.X(clknet_6_34__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_35__f_clk (.X(clknet_6_35__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_36__f_clk (.X(clknet_6_36__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_37__f_clk (.X(clknet_6_37__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_38__f_clk (.X(clknet_6_38__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_39__f_clk (.X(clknet_6_39__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_40__f_clk (.X(clknet_6_40__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_41__f_clk (.X(clknet_6_41__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_42__f_clk (.X(clknet_6_42__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_43__f_clk (.X(clknet_6_43__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_44__f_clk (.X(clknet_6_44__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_45__f_clk (.X(clknet_6_45__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_46__f_clk (.X(clknet_6_46__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_47__f_clk (.X(clknet_6_47__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_48__f_clk (.X(clknet_6_48__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_49__f_clk (.X(clknet_6_49__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_50__f_clk (.X(clknet_6_50__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_51__f_clk (.X(clknet_6_51__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_52__f_clk (.X(clknet_6_52__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_53__f_clk (.X(clknet_6_53__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_54__f_clk (.X(clknet_6_54__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_55__f_clk (.X(clknet_6_55__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_56__f_clk (.X(clknet_6_56__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_57__f_clk (.X(clknet_6_57__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_58__f_clk (.X(clknet_6_58__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_59__f_clk (.X(clknet_6_59__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_60__f_clk (.X(clknet_6_60__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_61__f_clk (.X(clknet_6_61__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_62__f_clk (.X(clknet_6_62__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_63__f_clk (.X(clknet_6_63__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_6_7__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_6_15__leaf_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_6_23__leaf_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_6_31__leaf_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_6_39__leaf_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_6_47__leaf_clk));
 sg13g2_buf_8 clkload6 (.A(clknet_6_55__leaf_clk));
 sg13g2_buf_8 clkload7 (.A(clknet_6_59__leaf_clk));
 sg13g2_buf_8 clkload8 (.A(clknet_6_63__leaf_clk));
 sg13g2_inv_2 clkload9 (.A(clknet_leaf_310_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_00190_));
 sg13g2_antennanp ANTENNA_2 (.A(_00197_));
 sg13g2_antennanp ANTENNA_3 (.A(_00197_));
 sg13g2_antennanp ANTENNA_4 (.A(_00197_));
 sg13g2_antennanp ANTENNA_5 (.A(_00197_));
 sg13g2_antennanp ANTENNA_6 (.A(_00228_));
 sg13g2_antennanp ANTENNA_7 (.A(_00228_));
 sg13g2_antennanp ANTENNA_8 (.A(_00235_));
 sg13g2_antennanp ANTENNA_9 (.A(_00930_));
 sg13g2_antennanp ANTENNA_10 (.A(_01052_));
 sg13g2_antennanp ANTENNA_11 (.A(_01052_));
 sg13g2_antennanp ANTENNA_12 (.A(_02943_));
 sg13g2_antennanp ANTENNA_13 (.A(_02943_));
 sg13g2_antennanp ANTENNA_14 (.A(_02943_));
 sg13g2_antennanp ANTENNA_15 (.A(_02943_));
 sg13g2_antennanp ANTENNA_16 (.A(_02950_));
 sg13g2_antennanp ANTENNA_17 (.A(_02950_));
 sg13g2_antennanp ANTENNA_18 (.A(_02950_));
 sg13g2_antennanp ANTENNA_19 (.A(_02950_));
 sg13g2_antennanp ANTENNA_20 (.A(_02950_));
 sg13g2_antennanp ANTENNA_21 (.A(_02950_));
 sg13g2_antennanp ANTENNA_22 (.A(_02953_));
 sg13g2_antennanp ANTENNA_23 (.A(_02953_));
 sg13g2_antennanp ANTENNA_24 (.A(_02953_));
 sg13g2_antennanp ANTENNA_25 (.A(_02953_));
 sg13g2_antennanp ANTENNA_26 (.A(_02960_));
 sg13g2_antennanp ANTENNA_27 (.A(_02960_));
 sg13g2_antennanp ANTENNA_28 (.A(_02960_));
 sg13g2_antennanp ANTENNA_29 (.A(_02965_));
 sg13g2_antennanp ANTENNA_30 (.A(_02965_));
 sg13g2_antennanp ANTENNA_31 (.A(_02965_));
 sg13g2_antennanp ANTENNA_32 (.A(_02965_));
 sg13g2_antennanp ANTENNA_33 (.A(_02965_));
 sg13g2_antennanp ANTENNA_34 (.A(_02965_));
 sg13g2_antennanp ANTENNA_35 (.A(_02965_));
 sg13g2_antennanp ANTENNA_36 (.A(_02973_));
 sg13g2_antennanp ANTENNA_37 (.A(_02973_));
 sg13g2_antennanp ANTENNA_38 (.A(_02973_));
 sg13g2_antennanp ANTENNA_39 (.A(_02973_));
 sg13g2_antennanp ANTENNA_40 (.A(_02973_));
 sg13g2_antennanp ANTENNA_41 (.A(_02973_));
 sg13g2_antennanp ANTENNA_42 (.A(_02973_));
 sg13g2_antennanp ANTENNA_43 (.A(_02973_));
 sg13g2_antennanp ANTENNA_44 (.A(_02973_));
 sg13g2_antennanp ANTENNA_45 (.A(_02973_));
 sg13g2_antennanp ANTENNA_46 (.A(_02973_));
 sg13g2_antennanp ANTENNA_47 (.A(_02973_));
 sg13g2_antennanp ANTENNA_48 (.A(_02973_));
 sg13g2_antennanp ANTENNA_49 (.A(_02973_));
 sg13g2_antennanp ANTENNA_50 (.A(_03429_));
 sg13g2_antennanp ANTENNA_51 (.A(_03429_));
 sg13g2_antennanp ANTENNA_52 (.A(_03429_));
 sg13g2_antennanp ANTENNA_53 (.A(_03429_));
 sg13g2_antennanp ANTENNA_54 (.A(_03429_));
 sg13g2_antennanp ANTENNA_55 (.A(_03435_));
 sg13g2_antennanp ANTENNA_56 (.A(_03435_));
 sg13g2_antennanp ANTENNA_57 (.A(_03435_));
 sg13g2_antennanp ANTENNA_58 (.A(_03435_));
 sg13g2_antennanp ANTENNA_59 (.A(_03435_));
 sg13g2_antennanp ANTENNA_60 (.A(_03435_));
 sg13g2_antennanp ANTENNA_61 (.A(_03435_));
 sg13g2_antennanp ANTENNA_62 (.A(_03435_));
 sg13g2_antennanp ANTENNA_63 (.A(_03435_));
 sg13g2_antennanp ANTENNA_64 (.A(_04212_));
 sg13g2_antennanp ANTENNA_65 (.A(_04212_));
 sg13g2_antennanp ANTENNA_66 (.A(_04212_));
 sg13g2_antennanp ANTENNA_67 (.A(_04212_));
 sg13g2_antennanp ANTENNA_68 (.A(_04212_));
 sg13g2_antennanp ANTENNA_69 (.A(_04212_));
 sg13g2_antennanp ANTENNA_70 (.A(_04212_));
 sg13g2_antennanp ANTENNA_71 (.A(_04742_));
 sg13g2_antennanp ANTENNA_72 (.A(_04742_));
 sg13g2_antennanp ANTENNA_73 (.A(_04742_));
 sg13g2_antennanp ANTENNA_74 (.A(_04742_));
 sg13g2_antennanp ANTENNA_75 (.A(_04887_));
 sg13g2_antennanp ANTENNA_76 (.A(_04887_));
 sg13g2_antennanp ANTENNA_77 (.A(_04887_));
 sg13g2_antennanp ANTENNA_78 (.A(_04887_));
 sg13g2_antennanp ANTENNA_79 (.A(_04894_));
 sg13g2_antennanp ANTENNA_80 (.A(_05013_));
 sg13g2_antennanp ANTENNA_81 (.A(_05015_));
 sg13g2_antennanp ANTENNA_82 (.A(_05169_));
 sg13g2_antennanp ANTENNA_83 (.A(_05280_));
 sg13g2_antennanp ANTENNA_84 (.A(_05311_));
 sg13g2_antennanp ANTENNA_85 (.A(_05311_));
 sg13g2_antennanp ANTENNA_86 (.A(_05311_));
 sg13g2_antennanp ANTENNA_87 (.A(_05311_));
 sg13g2_antennanp ANTENNA_88 (.A(_05372_));
 sg13g2_antennanp ANTENNA_89 (.A(_05432_));
 sg13g2_antennanp ANTENNA_90 (.A(_05442_));
 sg13g2_antennanp ANTENNA_91 (.A(_05442_));
 sg13g2_antennanp ANTENNA_92 (.A(_05508_));
 sg13g2_antennanp ANTENNA_93 (.A(_05646_));
 sg13g2_antennanp ANTENNA_94 (.A(_05650_));
 sg13g2_antennanp ANTENNA_95 (.A(_05654_));
 sg13g2_antennanp ANTENNA_96 (.A(_05654_));
 sg13g2_antennanp ANTENNA_97 (.A(_05763_));
 sg13g2_antennanp ANTENNA_98 (.A(_05763_));
 sg13g2_antennanp ANTENNA_99 (.A(_05763_));
 sg13g2_antennanp ANTENNA_100 (.A(_05763_));
 sg13g2_antennanp ANTENNA_101 (.A(_05763_));
 sg13g2_antennanp ANTENNA_102 (.A(_05766_));
 sg13g2_antennanp ANTENNA_103 (.A(_05766_));
 sg13g2_antennanp ANTENNA_104 (.A(_05766_));
 sg13g2_antennanp ANTENNA_105 (.A(_05770_));
 sg13g2_antennanp ANTENNA_106 (.A(_05770_));
 sg13g2_antennanp ANTENNA_107 (.A(_05770_));
 sg13g2_antennanp ANTENNA_108 (.A(_05770_));
 sg13g2_antennanp ANTENNA_109 (.A(_05770_));
 sg13g2_antennanp ANTENNA_110 (.A(_05775_));
 sg13g2_antennanp ANTENNA_111 (.A(_05775_));
 sg13g2_antennanp ANTENNA_112 (.A(_05775_));
 sg13g2_antennanp ANTENNA_113 (.A(_05785_));
 sg13g2_antennanp ANTENNA_114 (.A(_05785_));
 sg13g2_antennanp ANTENNA_115 (.A(_05785_));
 sg13g2_antennanp ANTENNA_116 (.A(_05785_));
 sg13g2_antennanp ANTENNA_117 (.A(_05785_));
 sg13g2_antennanp ANTENNA_118 (.A(_05835_));
 sg13g2_antennanp ANTENNA_119 (.A(_05835_));
 sg13g2_antennanp ANTENNA_120 (.A(_05835_));
 sg13g2_antennanp ANTENNA_121 (.A(_05835_));
 sg13g2_antennanp ANTENNA_122 (.A(_05835_));
 sg13g2_antennanp ANTENNA_123 (.A(_05835_));
 sg13g2_antennanp ANTENNA_124 (.A(_06843_));
 sg13g2_antennanp ANTENNA_125 (.A(_06843_));
 sg13g2_antennanp ANTENNA_126 (.A(_06843_));
 sg13g2_antennanp ANTENNA_127 (.A(_07398_));
 sg13g2_antennanp ANTENNA_128 (.A(_07433_));
 sg13g2_antennanp ANTENNA_129 (.A(_07434_));
 sg13g2_antennanp ANTENNA_130 (.A(_08297_));
 sg13g2_antennanp ANTENNA_131 (.A(_08297_));
 sg13g2_antennanp ANTENNA_132 (.A(_08502_));
 sg13g2_antennanp ANTENNA_133 (.A(_08502_));
 sg13g2_antennanp ANTENNA_134 (.A(_08502_));
 sg13g2_antennanp ANTENNA_135 (.A(_08502_));
 sg13g2_antennanp ANTENNA_136 (.A(_08502_));
 sg13g2_antennanp ANTENNA_137 (.A(_08502_));
 sg13g2_antennanp ANTENNA_138 (.A(_08502_));
 sg13g2_antennanp ANTENNA_139 (.A(_08502_));
 sg13g2_antennanp ANTENNA_140 (.A(_08502_));
 sg13g2_antennanp ANTENNA_141 (.A(_08502_));
 sg13g2_antennanp ANTENNA_142 (.A(_08502_));
 sg13g2_antennanp ANTENNA_143 (.A(_08502_));
 sg13g2_antennanp ANTENNA_144 (.A(_08533_));
 sg13g2_antennanp ANTENNA_145 (.A(_08533_));
 sg13g2_antennanp ANTENNA_146 (.A(_08533_));
 sg13g2_antennanp ANTENNA_147 (.A(_08533_));
 sg13g2_antennanp ANTENNA_148 (.A(_08533_));
 sg13g2_antennanp ANTENNA_149 (.A(_08533_));
 sg13g2_antennanp ANTENNA_150 (.A(_08558_));
 sg13g2_antennanp ANTENNA_151 (.A(_08558_));
 sg13g2_antennanp ANTENNA_152 (.A(_08558_));
 sg13g2_antennanp ANTENNA_153 (.A(_08558_));
 sg13g2_antennanp ANTENNA_154 (.A(_08558_));
 sg13g2_antennanp ANTENNA_155 (.A(_08558_));
 sg13g2_antennanp ANTENNA_156 (.A(_08558_));
 sg13g2_antennanp ANTENNA_157 (.A(_08558_));
 sg13g2_antennanp ANTENNA_158 (.A(_08558_));
 sg13g2_antennanp ANTENNA_159 (.A(_08558_));
 sg13g2_antennanp ANTENNA_160 (.A(_08558_));
 sg13g2_antennanp ANTENNA_161 (.A(_08558_));
 sg13g2_antennanp ANTENNA_162 (.A(_08634_));
 sg13g2_antennanp ANTENNA_163 (.A(_08634_));
 sg13g2_antennanp ANTENNA_164 (.A(_08634_));
 sg13g2_antennanp ANTENNA_165 (.A(_08634_));
 sg13g2_antennanp ANTENNA_166 (.A(_08634_));
 sg13g2_antennanp ANTENNA_167 (.A(_08634_));
 sg13g2_antennanp ANTENNA_168 (.A(_08634_));
 sg13g2_antennanp ANTENNA_169 (.A(_08634_));
 sg13g2_antennanp ANTENNA_170 (.A(_08634_));
 sg13g2_antennanp ANTENNA_171 (.A(_08679_));
 sg13g2_antennanp ANTENNA_172 (.A(_08679_));
 sg13g2_antennanp ANTENNA_173 (.A(_08679_));
 sg13g2_antennanp ANTENNA_174 (.A(_08679_));
 sg13g2_antennanp ANTENNA_175 (.A(_08679_));
 sg13g2_antennanp ANTENNA_176 (.A(_08689_));
 sg13g2_antennanp ANTENNA_177 (.A(_08689_));
 sg13g2_antennanp ANTENNA_178 (.A(_08689_));
 sg13g2_antennanp ANTENNA_179 (.A(_08689_));
 sg13g2_antennanp ANTENNA_180 (.A(_08698_));
 sg13g2_antennanp ANTENNA_181 (.A(_08698_));
 sg13g2_antennanp ANTENNA_182 (.A(_08698_));
 sg13g2_antennanp ANTENNA_183 (.A(_08728_));
 sg13g2_antennanp ANTENNA_184 (.A(_08728_));
 sg13g2_antennanp ANTENNA_185 (.A(_08728_));
 sg13g2_antennanp ANTENNA_186 (.A(_08728_));
 sg13g2_antennanp ANTENNA_187 (.A(_08759_));
 sg13g2_antennanp ANTENNA_188 (.A(_08759_));
 sg13g2_antennanp ANTENNA_189 (.A(_08759_));
 sg13g2_antennanp ANTENNA_190 (.A(_08759_));
 sg13g2_antennanp ANTENNA_191 (.A(_08779_));
 sg13g2_antennanp ANTENNA_192 (.A(_08779_));
 sg13g2_antennanp ANTENNA_193 (.A(_08779_));
 sg13g2_antennanp ANTENNA_194 (.A(_08853_));
 sg13g2_antennanp ANTENNA_195 (.A(_08918_));
 sg13g2_antennanp ANTENNA_196 (.A(_08918_));
 sg13g2_antennanp ANTENNA_197 (.A(_08918_));
 sg13g2_antennanp ANTENNA_198 (.A(_08938_));
 sg13g2_antennanp ANTENNA_199 (.A(_08959_));
 sg13g2_antennanp ANTENNA_200 (.A(_08970_));
 sg13g2_antennanp ANTENNA_201 (.A(_08970_));
 sg13g2_antennanp ANTENNA_202 (.A(_08970_));
 sg13g2_antennanp ANTENNA_203 (.A(_09158_));
 sg13g2_antennanp ANTENNA_204 (.A(_09158_));
 sg13g2_antennanp ANTENNA_205 (.A(_09158_));
 sg13g2_antennanp ANTENNA_206 (.A(_09167_));
 sg13g2_antennanp ANTENNA_207 (.A(_09277_));
 sg13g2_antennanp ANTENNA_208 (.A(_09277_));
 sg13g2_antennanp ANTENNA_209 (.A(_09277_));
 sg13g2_antennanp ANTENNA_210 (.A(_09277_));
 sg13g2_antennanp ANTENNA_211 (.A(_09277_));
 sg13g2_antennanp ANTENNA_212 (.A(_09277_));
 sg13g2_antennanp ANTENNA_213 (.A(_09277_));
 sg13g2_antennanp ANTENNA_214 (.A(_09277_));
 sg13g2_antennanp ANTENNA_215 (.A(_09277_));
 sg13g2_antennanp ANTENNA_216 (.A(_09277_));
 sg13g2_antennanp ANTENNA_217 (.A(_09320_));
 sg13g2_antennanp ANTENNA_218 (.A(_09320_));
 sg13g2_antennanp ANTENNA_219 (.A(_09320_));
 sg13g2_antennanp ANTENNA_220 (.A(_09320_));
 sg13g2_antennanp ANTENNA_221 (.A(_09320_));
 sg13g2_antennanp ANTENNA_222 (.A(_09320_));
 sg13g2_antennanp ANTENNA_223 (.A(_09320_));
 sg13g2_antennanp ANTENNA_224 (.A(_09320_));
 sg13g2_antennanp ANTENNA_225 (.A(_09336_));
 sg13g2_antennanp ANTENNA_226 (.A(_09336_));
 sg13g2_antennanp ANTENNA_227 (.A(_09349_));
 sg13g2_antennanp ANTENNA_228 (.A(_09349_));
 sg13g2_antennanp ANTENNA_229 (.A(_09349_));
 sg13g2_antennanp ANTENNA_230 (.A(_09349_));
 sg13g2_antennanp ANTENNA_231 (.A(_09349_));
 sg13g2_antennanp ANTENNA_232 (.A(_09349_));
 sg13g2_antennanp ANTENNA_233 (.A(_09349_));
 sg13g2_antennanp ANTENNA_234 (.A(_09349_));
 sg13g2_antennanp ANTENNA_235 (.A(_09351_));
 sg13g2_antennanp ANTENNA_236 (.A(_09351_));
 sg13g2_antennanp ANTENNA_237 (.A(_09351_));
 sg13g2_antennanp ANTENNA_238 (.A(_09351_));
 sg13g2_antennanp ANTENNA_239 (.A(_09351_));
 sg13g2_antennanp ANTENNA_240 (.A(_09351_));
 sg13g2_antennanp ANTENNA_241 (.A(_09351_));
 sg13g2_antennanp ANTENNA_242 (.A(_09351_));
 sg13g2_antennanp ANTENNA_243 (.A(_09351_));
 sg13g2_antennanp ANTENNA_244 (.A(_09351_));
 sg13g2_antennanp ANTENNA_245 (.A(_09351_));
 sg13g2_antennanp ANTENNA_246 (.A(_09351_));
 sg13g2_antennanp ANTENNA_247 (.A(_09380_));
 sg13g2_antennanp ANTENNA_248 (.A(_09380_));
 sg13g2_antennanp ANTENNA_249 (.A(_09380_));
 sg13g2_antennanp ANTENNA_250 (.A(_09380_));
 sg13g2_antennanp ANTENNA_251 (.A(_09385_));
 sg13g2_antennanp ANTENNA_252 (.A(_09385_));
 sg13g2_antennanp ANTENNA_253 (.A(_09385_));
 sg13g2_antennanp ANTENNA_254 (.A(_09385_));
 sg13g2_antennanp ANTENNA_255 (.A(_09385_));
 sg13g2_antennanp ANTENNA_256 (.A(_09385_));
 sg13g2_antennanp ANTENNA_257 (.A(_09385_));
 sg13g2_antennanp ANTENNA_258 (.A(_09385_));
 sg13g2_antennanp ANTENNA_259 (.A(_09385_));
 sg13g2_antennanp ANTENNA_260 (.A(_09386_));
 sg13g2_antennanp ANTENNA_261 (.A(_09386_));
 sg13g2_antennanp ANTENNA_262 (.A(_09386_));
 sg13g2_antennanp ANTENNA_263 (.A(_09386_));
 sg13g2_antennanp ANTENNA_264 (.A(_09386_));
 sg13g2_antennanp ANTENNA_265 (.A(_09386_));
 sg13g2_antennanp ANTENNA_266 (.A(_09386_));
 sg13g2_antennanp ANTENNA_267 (.A(_09386_));
 sg13g2_antennanp ANTENNA_268 (.A(_09386_));
 sg13g2_antennanp ANTENNA_269 (.A(_09386_));
 sg13g2_antennanp ANTENNA_270 (.A(_09388_));
 sg13g2_antennanp ANTENNA_271 (.A(_09388_));
 sg13g2_antennanp ANTENNA_272 (.A(_09388_));
 sg13g2_antennanp ANTENNA_273 (.A(_09389_));
 sg13g2_antennanp ANTENNA_274 (.A(_09389_));
 sg13g2_antennanp ANTENNA_275 (.A(_09389_));
 sg13g2_antennanp ANTENNA_276 (.A(_09389_));
 sg13g2_antennanp ANTENNA_277 (.A(_09389_));
 sg13g2_antennanp ANTENNA_278 (.A(_09389_));
 sg13g2_antennanp ANTENNA_279 (.A(_09390_));
 sg13g2_antennanp ANTENNA_280 (.A(_09390_));
 sg13g2_antennanp ANTENNA_281 (.A(_09390_));
 sg13g2_antennanp ANTENNA_282 (.A(_09390_));
 sg13g2_antennanp ANTENNA_283 (.A(_09444_));
 sg13g2_antennanp ANTENNA_284 (.A(_09444_));
 sg13g2_antennanp ANTENNA_285 (.A(_09444_));
 sg13g2_antennanp ANTENNA_286 (.A(_09444_));
 sg13g2_antennanp ANTENNA_287 (.A(_09444_));
 sg13g2_antennanp ANTENNA_288 (.A(_09444_));
 sg13g2_antennanp ANTENNA_289 (.A(_09444_));
 sg13g2_antennanp ANTENNA_290 (.A(_09444_));
 sg13g2_antennanp ANTENNA_291 (.A(_09444_));
 sg13g2_antennanp ANTENNA_292 (.A(_09444_));
 sg13g2_antennanp ANTENNA_293 (.A(_09445_));
 sg13g2_antennanp ANTENNA_294 (.A(_09445_));
 sg13g2_antennanp ANTENNA_295 (.A(_09445_));
 sg13g2_antennanp ANTENNA_296 (.A(_09445_));
 sg13g2_antennanp ANTENNA_297 (.A(_09445_));
 sg13g2_antennanp ANTENNA_298 (.A(_09445_));
 sg13g2_antennanp ANTENNA_299 (.A(_09445_));
 sg13g2_antennanp ANTENNA_300 (.A(_09445_));
 sg13g2_antennanp ANTENNA_301 (.A(_09445_));
 sg13g2_antennanp ANTENNA_302 (.A(_09554_));
 sg13g2_antennanp ANTENNA_303 (.A(_09554_));
 sg13g2_antennanp ANTENNA_304 (.A(_09562_));
 sg13g2_antennanp ANTENNA_305 (.A(_09562_));
 sg13g2_antennanp ANTENNA_306 (.A(_09587_));
 sg13g2_antennanp ANTENNA_307 (.A(_09608_));
 sg13g2_antennanp ANTENNA_308 (.A(_09665_));
 sg13g2_antennanp ANTENNA_309 (.A(_09695_));
 sg13g2_antennanp ANTENNA_310 (.A(_09721_));
 sg13g2_antennanp ANTENNA_311 (.A(_09742_));
 sg13g2_antennanp ANTENNA_312 (.A(_09765_));
 sg13g2_antennanp ANTENNA_313 (.A(_09794_));
 sg13g2_antennanp ANTENNA_314 (.A(_09796_));
 sg13g2_antennanp ANTENNA_315 (.A(_09836_));
 sg13g2_antennanp ANTENNA_316 (.A(_09836_));
 sg13g2_antennanp ANTENNA_317 (.A(_09836_));
 sg13g2_antennanp ANTENNA_318 (.A(_09836_));
 sg13g2_antennanp ANTENNA_319 (.A(_09836_));
 sg13g2_antennanp ANTENNA_320 (.A(_09836_));
 sg13g2_antennanp ANTENNA_321 (.A(_09836_));
 sg13g2_antennanp ANTENNA_322 (.A(_09836_));
 sg13g2_antennanp ANTENNA_323 (.A(_09836_));
 sg13g2_antennanp ANTENNA_324 (.A(_09912_));
 sg13g2_antennanp ANTENNA_325 (.A(_09990_));
 sg13g2_antennanp ANTENNA_326 (.A(_09990_));
 sg13g2_antennanp ANTENNA_327 (.A(_09990_));
 sg13g2_antennanp ANTENNA_328 (.A(_09990_));
 sg13g2_antennanp ANTENNA_329 (.A(_09990_));
 sg13g2_antennanp ANTENNA_330 (.A(_09990_));
 sg13g2_antennanp ANTENNA_331 (.A(_09990_));
 sg13g2_antennanp ANTENNA_332 (.A(_09990_));
 sg13g2_antennanp ANTENNA_333 (.A(_10172_));
 sg13g2_antennanp ANTENNA_334 (.A(_10172_));
 sg13g2_antennanp ANTENNA_335 (.A(_10172_));
 sg13g2_antennanp ANTENNA_336 (.A(_10172_));
 sg13g2_antennanp ANTENNA_337 (.A(_10240_));
 sg13g2_antennanp ANTENNA_338 (.A(_10240_));
 sg13g2_antennanp ANTENNA_339 (.A(_10240_));
 sg13g2_antennanp ANTENNA_340 (.A(_10240_));
 sg13g2_antennanp ANTENNA_341 (.A(_10246_));
 sg13g2_antennanp ANTENNA_342 (.A(_10246_));
 sg13g2_antennanp ANTENNA_343 (.A(_10246_));
 sg13g2_antennanp ANTENNA_344 (.A(_10246_));
 sg13g2_antennanp ANTENNA_345 (.A(_10246_));
 sg13g2_antennanp ANTENNA_346 (.A(_10246_));
 sg13g2_antennanp ANTENNA_347 (.A(_10246_));
 sg13g2_antennanp ANTENNA_348 (.A(_10307_));
 sg13g2_antennanp ANTENNA_349 (.A(_10307_));
 sg13g2_antennanp ANTENNA_350 (.A(_10307_));
 sg13g2_antennanp ANTENNA_351 (.A(_10307_));
 sg13g2_antennanp ANTENNA_352 (.A(_10307_));
 sg13g2_antennanp ANTENNA_353 (.A(_10307_));
 sg13g2_antennanp ANTENNA_354 (.A(_10307_));
 sg13g2_antennanp ANTENNA_355 (.A(_10307_));
 sg13g2_antennanp ANTENNA_356 (.A(_10312_));
 sg13g2_antennanp ANTENNA_357 (.A(_10312_));
 sg13g2_antennanp ANTENNA_358 (.A(_10312_));
 sg13g2_antennanp ANTENNA_359 (.A(_10312_));
 sg13g2_antennanp ANTENNA_360 (.A(_10312_));
 sg13g2_antennanp ANTENNA_361 (.A(_10312_));
 sg13g2_antennanp ANTENNA_362 (.A(_10312_));
 sg13g2_antennanp ANTENNA_363 (.A(_10312_));
 sg13g2_antennanp ANTENNA_364 (.A(_10319_));
 sg13g2_antennanp ANTENNA_365 (.A(_10319_));
 sg13g2_antennanp ANTENNA_366 (.A(_10319_));
 sg13g2_antennanp ANTENNA_367 (.A(_10319_));
 sg13g2_antennanp ANTENNA_368 (.A(_10319_));
 sg13g2_antennanp ANTENNA_369 (.A(_10319_));
 sg13g2_antennanp ANTENNA_370 (.A(_10319_));
 sg13g2_antennanp ANTENNA_371 (.A(_10319_));
 sg13g2_antennanp ANTENNA_372 (.A(_10326_));
 sg13g2_antennanp ANTENNA_373 (.A(_10326_));
 sg13g2_antennanp ANTENNA_374 (.A(_10326_));
 sg13g2_antennanp ANTENNA_375 (.A(_10326_));
 sg13g2_antennanp ANTENNA_376 (.A(_10326_));
 sg13g2_antennanp ANTENNA_377 (.A(_10326_));
 sg13g2_antennanp ANTENNA_378 (.A(_10326_));
 sg13g2_antennanp ANTENNA_379 (.A(_10326_));
 sg13g2_antennanp ANTENNA_380 (.A(_10339_));
 sg13g2_antennanp ANTENNA_381 (.A(_10339_));
 sg13g2_antennanp ANTENNA_382 (.A(_10339_));
 sg13g2_antennanp ANTENNA_383 (.A(_10339_));
 sg13g2_antennanp ANTENNA_384 (.A(_10339_));
 sg13g2_antennanp ANTENNA_385 (.A(_10339_));
 sg13g2_antennanp ANTENNA_386 (.A(_10339_));
 sg13g2_antennanp ANTENNA_387 (.A(_10344_));
 sg13g2_antennanp ANTENNA_388 (.A(_10344_));
 sg13g2_antennanp ANTENNA_389 (.A(_10344_));
 sg13g2_antennanp ANTENNA_390 (.A(_10344_));
 sg13g2_antennanp ANTENNA_391 (.A(_10344_));
 sg13g2_antennanp ANTENNA_392 (.A(_10344_));
 sg13g2_antennanp ANTENNA_393 (.A(_10344_));
 sg13g2_antennanp ANTENNA_394 (.A(_10344_));
 sg13g2_antennanp ANTENNA_395 (.A(_10562_));
 sg13g2_antennanp ANTENNA_396 (.A(_10562_));
 sg13g2_antennanp ANTENNA_397 (.A(_10612_));
 sg13g2_antennanp ANTENNA_398 (.A(_10612_));
 sg13g2_antennanp ANTENNA_399 (.A(_10645_));
 sg13g2_antennanp ANTENNA_400 (.A(_10645_));
 sg13g2_antennanp ANTENNA_401 (.A(_11129_));
 sg13g2_antennanp ANTENNA_402 (.A(_11383_));
 sg13g2_antennanp ANTENNA_403 (.A(_11383_));
 sg13g2_antennanp ANTENNA_404 (.A(_11383_));
 sg13g2_antennanp ANTENNA_405 (.A(_11383_));
 sg13g2_antennanp ANTENNA_406 (.A(_11383_));
 sg13g2_antennanp ANTENNA_407 (.A(_11383_));
 sg13g2_antennanp ANTENNA_408 (.A(_11383_));
 sg13g2_antennanp ANTENNA_409 (.A(_11383_));
 sg13g2_antennanp ANTENNA_410 (.A(_11383_));
 sg13g2_antennanp ANTENNA_411 (.A(_11383_));
 sg13g2_antennanp ANTENNA_412 (.A(_11383_));
 sg13g2_antennanp ANTENNA_413 (.A(_11383_));
 sg13g2_antennanp ANTENNA_414 (.A(_11383_));
 sg13g2_antennanp ANTENNA_415 (.A(_11383_));
 sg13g2_antennanp ANTENNA_416 (.A(_11383_));
 sg13g2_antennanp ANTENNA_417 (.A(_11383_));
 sg13g2_antennanp ANTENNA_418 (.A(_11383_));
 sg13g2_antennanp ANTENNA_419 (.A(_11383_));
 sg13g2_antennanp ANTENNA_420 (.A(_11383_));
 sg13g2_antennanp ANTENNA_421 (.A(_11383_));
 sg13g2_antennanp ANTENNA_422 (.A(_11407_));
 sg13g2_antennanp ANTENNA_423 (.A(_11407_));
 sg13g2_antennanp ANTENNA_424 (.A(_11407_));
 sg13g2_antennanp ANTENNA_425 (.A(_11407_));
 sg13g2_antennanp ANTENNA_426 (.A(_12004_));
 sg13g2_antennanp ANTENNA_427 (.A(_12004_));
 sg13g2_antennanp ANTENNA_428 (.A(_12004_));
 sg13g2_antennanp ANTENNA_429 (.A(_12004_));
 sg13g2_antennanp ANTENNA_430 (.A(_12058_));
 sg13g2_antennanp ANTENNA_431 (.A(_12058_));
 sg13g2_antennanp ANTENNA_432 (.A(_12058_));
 sg13g2_antennanp ANTENNA_433 (.A(_12058_));
 sg13g2_antennanp ANTENNA_434 (.A(_12058_));
 sg13g2_antennanp ANTENNA_435 (.A(_12058_));
 sg13g2_antennanp ANTENNA_436 (.A(_12058_));
 sg13g2_antennanp ANTENNA_437 (.A(_12058_));
 sg13g2_antennanp ANTENNA_438 (.A(_12058_));
 sg13g2_antennanp ANTENNA_439 (.A(_12127_));
 sg13g2_antennanp ANTENNA_440 (.A(_12127_));
 sg13g2_antennanp ANTENNA_441 (.A(_12127_));
 sg13g2_antennanp ANTENNA_442 (.A(_12127_));
 sg13g2_antennanp ANTENNA_443 (.A(_12127_));
 sg13g2_antennanp ANTENNA_444 (.A(_12127_));
 sg13g2_antennanp ANTENNA_445 (.A(_12127_));
 sg13g2_antennanp ANTENNA_446 (.A(_12127_));
 sg13g2_antennanp ANTENNA_447 (.A(_12127_));
 sg13g2_antennanp ANTENNA_448 (.A(_12152_));
 sg13g2_antennanp ANTENNA_449 (.A(_12152_));
 sg13g2_antennanp ANTENNA_450 (.A(_12152_));
 sg13g2_antennanp ANTENNA_451 (.A(_12152_));
 sg13g2_antennanp ANTENNA_452 (.A(_12152_));
 sg13g2_antennanp ANTENNA_453 (.A(_12152_));
 sg13g2_antennanp ANTENNA_454 (.A(_12152_));
 sg13g2_antennanp ANTENNA_455 (.A(_12152_));
 sg13g2_antennanp ANTENNA_456 (.A(_12218_));
 sg13g2_antennanp ANTENNA_457 (.A(_12218_));
 sg13g2_antennanp ANTENNA_458 (.A(_12218_));
 sg13g2_antennanp ANTENNA_459 (.A(_12218_));
 sg13g2_antennanp ANTENNA_460 (.A(_12218_));
 sg13g2_antennanp ANTENNA_461 (.A(_12218_));
 sg13g2_antennanp ANTENNA_462 (.A(_12218_));
 sg13g2_antennanp ANTENNA_463 (.A(_12218_));
 sg13g2_antennanp ANTENNA_464 (.A(_12218_));
 sg13g2_antennanp ANTENNA_465 (.A(_12223_));
 sg13g2_antennanp ANTENNA_466 (.A(_12223_));
 sg13g2_antennanp ANTENNA_467 (.A(_12223_));
 sg13g2_antennanp ANTENNA_468 (.A(_12223_));
 sg13g2_antennanp ANTENNA_469 (.A(_12223_));
 sg13g2_antennanp ANTENNA_470 (.A(_12223_));
 sg13g2_antennanp ANTENNA_471 (.A(_12223_));
 sg13g2_antennanp ANTENNA_472 (.A(_12223_));
 sg13g2_antennanp ANTENNA_473 (.A(_12223_));
 sg13g2_antennanp ANTENNA_474 (.A(_12229_));
 sg13g2_antennanp ANTENNA_475 (.A(_12229_));
 sg13g2_antennanp ANTENNA_476 (.A(_12229_));
 sg13g2_antennanp ANTENNA_477 (.A(_12229_));
 sg13g2_antennanp ANTENNA_478 (.A(_12229_));
 sg13g2_antennanp ANTENNA_479 (.A(_12229_));
 sg13g2_antennanp ANTENNA_480 (.A(_12229_));
 sg13g2_antennanp ANTENNA_481 (.A(_12229_));
 sg13g2_antennanp ANTENNA_482 (.A(_12229_));
 sg13g2_antennanp ANTENNA_483 (.A(_12558_));
 sg13g2_antennanp ANTENNA_484 (.A(_12558_));
 sg13g2_antennanp ANTENNA_485 (.A(_12558_));
 sg13g2_antennanp ANTENNA_486 (.A(_12558_));
 sg13g2_antennanp ANTENNA_487 (.A(_12558_));
 sg13g2_antennanp ANTENNA_488 (.A(_12726_));
 sg13g2_antennanp ANTENNA_489 (.A(_12726_));
 sg13g2_antennanp ANTENNA_490 (.A(_12726_));
 sg13g2_antennanp ANTENNA_491 (.A(clk));
 sg13g2_antennanp ANTENNA_492 (.A(clk));
 sg13g2_antennanp ANTENNA_493 (.A(\cpu.ex.pc[3] ));
 sg13g2_antennanp ANTENNA_494 (.A(\cpu.gpio.uart_rx ));
 sg13g2_antennanp ANTENNA_495 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_496 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_497 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_498 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_499 (.A(net3));
 sg13g2_antennanp ANTENNA_500 (.A(net3));
 sg13g2_antennanp ANTENNA_501 (.A(net3));
 sg13g2_antennanp ANTENNA_502 (.A(net12));
 sg13g2_antennanp ANTENNA_503 (.A(net12));
 sg13g2_antennanp ANTENNA_504 (.A(net12));
 sg13g2_antennanp ANTENNA_505 (.A(net13));
 sg13g2_antennanp ANTENNA_506 (.A(net13));
 sg13g2_antennanp ANTENNA_507 (.A(net13));
 sg13g2_antennanp ANTENNA_508 (.A(net14));
 sg13g2_antennanp ANTENNA_509 (.A(net14));
 sg13g2_antennanp ANTENNA_510 (.A(net14));
 sg13g2_antennanp ANTENNA_511 (.A(net437));
 sg13g2_antennanp ANTENNA_512 (.A(net437));
 sg13g2_antennanp ANTENNA_513 (.A(net437));
 sg13g2_antennanp ANTENNA_514 (.A(net437));
 sg13g2_antennanp ANTENNA_515 (.A(net437));
 sg13g2_antennanp ANTENNA_516 (.A(net437));
 sg13g2_antennanp ANTENNA_517 (.A(net437));
 sg13g2_antennanp ANTENNA_518 (.A(net437));
 sg13g2_antennanp ANTENNA_519 (.A(net437));
 sg13g2_antennanp ANTENNA_520 (.A(net437));
 sg13g2_antennanp ANTENNA_521 (.A(net437));
 sg13g2_antennanp ANTENNA_522 (.A(net437));
 sg13g2_antennanp ANTENNA_523 (.A(net437));
 sg13g2_antennanp ANTENNA_524 (.A(net437));
 sg13g2_antennanp ANTENNA_525 (.A(net437));
 sg13g2_antennanp ANTENNA_526 (.A(net524));
 sg13g2_antennanp ANTENNA_527 (.A(net524));
 sg13g2_antennanp ANTENNA_528 (.A(net524));
 sg13g2_antennanp ANTENNA_529 (.A(net524));
 sg13g2_antennanp ANTENNA_530 (.A(net524));
 sg13g2_antennanp ANTENNA_531 (.A(net524));
 sg13g2_antennanp ANTENNA_532 (.A(net524));
 sg13g2_antennanp ANTENNA_533 (.A(net524));
 sg13g2_antennanp ANTENNA_534 (.A(net524));
 sg13g2_antennanp ANTENNA_535 (.A(net524));
 sg13g2_antennanp ANTENNA_536 (.A(net524));
 sg13g2_antennanp ANTENNA_537 (.A(net524));
 sg13g2_antennanp ANTENNA_538 (.A(net524));
 sg13g2_antennanp ANTENNA_539 (.A(net542));
 sg13g2_antennanp ANTENNA_540 (.A(net542));
 sg13g2_antennanp ANTENNA_541 (.A(net542));
 sg13g2_antennanp ANTENNA_542 (.A(net542));
 sg13g2_antennanp ANTENNA_543 (.A(net542));
 sg13g2_antennanp ANTENNA_544 (.A(net542));
 sg13g2_antennanp ANTENNA_545 (.A(net542));
 sg13g2_antennanp ANTENNA_546 (.A(net542));
 sg13g2_antennanp ANTENNA_547 (.A(net656));
 sg13g2_antennanp ANTENNA_548 (.A(net656));
 sg13g2_antennanp ANTENNA_549 (.A(net656));
 sg13g2_antennanp ANTENNA_550 (.A(net656));
 sg13g2_antennanp ANTENNA_551 (.A(net656));
 sg13g2_antennanp ANTENNA_552 (.A(net656));
 sg13g2_antennanp ANTENNA_553 (.A(net656));
 sg13g2_antennanp ANTENNA_554 (.A(net656));
 sg13g2_antennanp ANTENNA_555 (.A(net656));
 sg13g2_antennanp ANTENNA_556 (.A(net656));
 sg13g2_antennanp ANTENNA_557 (.A(net656));
 sg13g2_antennanp ANTENNA_558 (.A(net656));
 sg13g2_antennanp ANTENNA_559 (.A(net656));
 sg13g2_antennanp ANTENNA_560 (.A(net656));
 sg13g2_antennanp ANTENNA_561 (.A(net656));
 sg13g2_antennanp ANTENNA_562 (.A(net656));
 sg13g2_antennanp ANTENNA_563 (.A(net656));
 sg13g2_antennanp ANTENNA_564 (.A(net656));
 sg13g2_antennanp ANTENNA_565 (.A(net656));
 sg13g2_antennanp ANTENNA_566 (.A(net656));
 sg13g2_antennanp ANTENNA_567 (.A(net656));
 sg13g2_antennanp ANTENNA_568 (.A(net656));
 sg13g2_antennanp ANTENNA_569 (.A(net685));
 sg13g2_antennanp ANTENNA_570 (.A(net685));
 sg13g2_antennanp ANTENNA_571 (.A(net685));
 sg13g2_antennanp ANTENNA_572 (.A(net685));
 sg13g2_antennanp ANTENNA_573 (.A(net685));
 sg13g2_antennanp ANTENNA_574 (.A(net685));
 sg13g2_antennanp ANTENNA_575 (.A(net685));
 sg13g2_antennanp ANTENNA_576 (.A(net685));
 sg13g2_antennanp ANTENNA_577 (.A(net685));
 sg13g2_antennanp ANTENNA_578 (.A(net707));
 sg13g2_antennanp ANTENNA_579 (.A(net707));
 sg13g2_antennanp ANTENNA_580 (.A(net707));
 sg13g2_antennanp ANTENNA_581 (.A(net707));
 sg13g2_antennanp ANTENNA_582 (.A(net707));
 sg13g2_antennanp ANTENNA_583 (.A(net707));
 sg13g2_antennanp ANTENNA_584 (.A(net707));
 sg13g2_antennanp ANTENNA_585 (.A(net707));
 sg13g2_antennanp ANTENNA_586 (.A(net707));
 sg13g2_antennanp ANTENNA_587 (.A(net707));
 sg13g2_antennanp ANTENNA_588 (.A(net707));
 sg13g2_antennanp ANTENNA_589 (.A(net707));
 sg13g2_antennanp ANTENNA_590 (.A(net707));
 sg13g2_antennanp ANTENNA_591 (.A(net707));
 sg13g2_antennanp ANTENNA_592 (.A(net707));
 sg13g2_antennanp ANTENNA_593 (.A(net707));
 sg13g2_antennanp ANTENNA_594 (.A(net707));
 sg13g2_antennanp ANTENNA_595 (.A(net707));
 sg13g2_antennanp ANTENNA_596 (.A(net707));
 sg13g2_antennanp ANTENNA_597 (.A(net707));
 sg13g2_antennanp ANTENNA_598 (.A(net707));
 sg13g2_antennanp ANTENNA_599 (.A(net707));
 sg13g2_antennanp ANTENNA_600 (.A(net707));
 sg13g2_antennanp ANTENNA_601 (.A(net707));
 sg13g2_antennanp ANTENNA_602 (.A(net803));
 sg13g2_antennanp ANTENNA_603 (.A(net803));
 sg13g2_antennanp ANTENNA_604 (.A(net803));
 sg13g2_antennanp ANTENNA_605 (.A(net803));
 sg13g2_antennanp ANTENNA_606 (.A(net803));
 sg13g2_antennanp ANTENNA_607 (.A(net803));
 sg13g2_antennanp ANTENNA_608 (.A(net803));
 sg13g2_antennanp ANTENNA_609 (.A(net803));
 sg13g2_antennanp ANTENNA_610 (.A(net803));
 sg13g2_antennanp ANTENNA_611 (.A(net803));
 sg13g2_antennanp ANTENNA_612 (.A(net803));
 sg13g2_antennanp ANTENNA_613 (.A(net803));
 sg13g2_antennanp ANTENNA_614 (.A(net803));
 sg13g2_antennanp ANTENNA_615 (.A(net803));
 sg13g2_antennanp ANTENNA_616 (.A(net803));
 sg13g2_antennanp ANTENNA_617 (.A(net803));
 sg13g2_antennanp ANTENNA_618 (.A(net887));
 sg13g2_antennanp ANTENNA_619 (.A(net887));
 sg13g2_antennanp ANTENNA_620 (.A(net887));
 sg13g2_antennanp ANTENNA_621 (.A(net887));
 sg13g2_antennanp ANTENNA_622 (.A(net887));
 sg13g2_antennanp ANTENNA_623 (.A(net887));
 sg13g2_antennanp ANTENNA_624 (.A(net887));
 sg13g2_antennanp ANTENNA_625 (.A(net887));
 sg13g2_antennanp ANTENNA_626 (.A(net887));
 sg13g2_antennanp ANTENNA_627 (.A(net889));
 sg13g2_antennanp ANTENNA_628 (.A(net889));
 sg13g2_antennanp ANTENNA_629 (.A(net889));
 sg13g2_antennanp ANTENNA_630 (.A(net889));
 sg13g2_antennanp ANTENNA_631 (.A(net889));
 sg13g2_antennanp ANTENNA_632 (.A(net889));
 sg13g2_antennanp ANTENNA_633 (.A(net889));
 sg13g2_antennanp ANTENNA_634 (.A(net889));
 sg13g2_antennanp ANTENNA_635 (.A(net928));
 sg13g2_antennanp ANTENNA_636 (.A(net928));
 sg13g2_antennanp ANTENNA_637 (.A(net928));
 sg13g2_antennanp ANTENNA_638 (.A(net928));
 sg13g2_antennanp ANTENNA_639 (.A(net928));
 sg13g2_antennanp ANTENNA_640 (.A(net928));
 sg13g2_antennanp ANTENNA_641 (.A(net928));
 sg13g2_antennanp ANTENNA_642 (.A(net928));
 sg13g2_antennanp ANTENNA_643 (.A(net928));
 sg13g2_antennanp ANTENNA_644 (.A(net941));
 sg13g2_antennanp ANTENNA_645 (.A(net941));
 sg13g2_antennanp ANTENNA_646 (.A(net941));
 sg13g2_antennanp ANTENNA_647 (.A(net941));
 sg13g2_antennanp ANTENNA_648 (.A(net941));
 sg13g2_antennanp ANTENNA_649 (.A(net941));
 sg13g2_antennanp ANTENNA_650 (.A(net941));
 sg13g2_antennanp ANTENNA_651 (.A(net941));
 sg13g2_antennanp ANTENNA_652 (.A(net941));
 sg13g2_antennanp ANTENNA_653 (.A(net980));
 sg13g2_antennanp ANTENNA_654 (.A(net980));
 sg13g2_antennanp ANTENNA_655 (.A(net980));
 sg13g2_antennanp ANTENNA_656 (.A(net980));
 sg13g2_antennanp ANTENNA_657 (.A(net980));
 sg13g2_antennanp ANTENNA_658 (.A(net980));
 sg13g2_antennanp ANTENNA_659 (.A(net980));
 sg13g2_antennanp ANTENNA_660 (.A(net980));
 sg13g2_antennanp ANTENNA_661 (.A(net980));
 sg13g2_antennanp ANTENNA_662 (.A(net983));
 sg13g2_antennanp ANTENNA_663 (.A(net983));
 sg13g2_antennanp ANTENNA_664 (.A(net983));
 sg13g2_antennanp ANTENNA_665 (.A(net983));
 sg13g2_antennanp ANTENNA_666 (.A(net983));
 sg13g2_antennanp ANTENNA_667 (.A(net983));
 sg13g2_antennanp ANTENNA_668 (.A(net983));
 sg13g2_antennanp ANTENNA_669 (.A(net983));
 sg13g2_antennanp ANTENNA_670 (.A(net983));
 sg13g2_antennanp ANTENNA_671 (.A(net983));
 sg13g2_antennanp ANTENNA_672 (.A(net983));
 sg13g2_antennanp ANTENNA_673 (.A(net983));
 sg13g2_antennanp ANTENNA_674 (.A(net983));
 sg13g2_antennanp ANTENNA_675 (.A(net983));
 sg13g2_antennanp ANTENNA_676 (.A(net983));
 sg13g2_antennanp ANTENNA_677 (.A(net983));
 sg13g2_antennanp ANTENNA_678 (.A(net983));
 sg13g2_antennanp ANTENNA_679 (.A(net983));
 sg13g2_antennanp ANTENNA_680 (.A(net983));
 sg13g2_antennanp ANTENNA_681 (.A(net984));
 sg13g2_antennanp ANTENNA_682 (.A(net984));
 sg13g2_antennanp ANTENNA_683 (.A(net984));
 sg13g2_antennanp ANTENNA_684 (.A(net984));
 sg13g2_antennanp ANTENNA_685 (.A(net984));
 sg13g2_antennanp ANTENNA_686 (.A(net984));
 sg13g2_antennanp ANTENNA_687 (.A(net984));
 sg13g2_antennanp ANTENNA_688 (.A(net984));
 sg13g2_antennanp ANTENNA_689 (.A(net984));
 sg13g2_antennanp ANTENNA_690 (.A(net984));
 sg13g2_antennanp ANTENNA_691 (.A(net984));
 sg13g2_antennanp ANTENNA_692 (.A(net984));
 sg13g2_antennanp ANTENNA_693 (.A(net984));
 sg13g2_antennanp ANTENNA_694 (.A(net984));
 sg13g2_antennanp ANTENNA_695 (.A(net984));
 sg13g2_antennanp ANTENNA_696 (.A(net984));
 sg13g2_antennanp ANTENNA_697 (.A(net984));
 sg13g2_antennanp ANTENNA_698 (.A(net984));
 sg13g2_antennanp ANTENNA_699 (.A(net984));
 sg13g2_antennanp ANTENNA_700 (.A(net984));
 sg13g2_antennanp ANTENNA_701 (.A(net984));
 sg13g2_antennanp ANTENNA_702 (.A(net984));
 sg13g2_antennanp ANTENNA_703 (.A(net984));
 sg13g2_antennanp ANTENNA_704 (.A(net984));
 sg13g2_antennanp ANTENNA_705 (.A(net984));
 sg13g2_antennanp ANTENNA_706 (.A(net984));
 sg13g2_antennanp ANTENNA_707 (.A(net984));
 sg13g2_antennanp ANTENNA_708 (.A(net984));
 sg13g2_antennanp ANTENNA_709 (.A(net984));
 sg13g2_antennanp ANTENNA_710 (.A(net984));
 sg13g2_antennanp ANTENNA_711 (.A(net984));
 sg13g2_antennanp ANTENNA_712 (.A(net1006));
 sg13g2_antennanp ANTENNA_713 (.A(net1006));
 sg13g2_antennanp ANTENNA_714 (.A(net1006));
 sg13g2_antennanp ANTENNA_715 (.A(net1006));
 sg13g2_antennanp ANTENNA_716 (.A(net1006));
 sg13g2_antennanp ANTENNA_717 (.A(net1006));
 sg13g2_antennanp ANTENNA_718 (.A(net1006));
 sg13g2_antennanp ANTENNA_719 (.A(net1006));
 sg13g2_antennanp ANTENNA_720 (.A(net1006));
 sg13g2_antennanp ANTENNA_721 (.A(net1006));
 sg13g2_antennanp ANTENNA_722 (.A(net1006));
 sg13g2_antennanp ANTENNA_723 (.A(net1006));
 sg13g2_antennanp ANTENNA_724 (.A(net1006));
 sg13g2_antennanp ANTENNA_725 (.A(net1006));
 sg13g2_antennanp ANTENNA_726 (.A(net1006));
 sg13g2_antennanp ANTENNA_727 (.A(net1006));
 sg13g2_antennanp ANTENNA_728 (.A(net1006));
 sg13g2_antennanp ANTENNA_729 (.A(net1006));
 sg13g2_antennanp ANTENNA_730 (.A(net1006));
 sg13g2_antennanp ANTENNA_731 (.A(net1006));
 sg13g2_antennanp ANTENNA_732 (.A(net1006));
 sg13g2_antennanp ANTENNA_733 (.A(net1006));
 sg13g2_antennanp ANTENNA_734 (.A(net1006));
 sg13g2_antennanp ANTENNA_735 (.A(net1006));
 sg13g2_antennanp ANTENNA_736 (.A(net1006));
 sg13g2_antennanp ANTENNA_737 (.A(net1006));
 sg13g2_antennanp ANTENNA_738 (.A(net1075));
 sg13g2_antennanp ANTENNA_739 (.A(net1075));
 sg13g2_antennanp ANTENNA_740 (.A(net1075));
 sg13g2_antennanp ANTENNA_741 (.A(net1075));
 sg13g2_antennanp ANTENNA_742 (.A(net1075));
 sg13g2_antennanp ANTENNA_743 (.A(net1075));
 sg13g2_antennanp ANTENNA_744 (.A(net1075));
 sg13g2_antennanp ANTENNA_745 (.A(net1075));
 sg13g2_antennanp ANTENNA_746 (.A(net1075));
 sg13g2_antennanp ANTENNA_747 (.A(_00190_));
 sg13g2_antennanp ANTENNA_748 (.A(_00197_));
 sg13g2_antennanp ANTENNA_749 (.A(_00197_));
 sg13g2_antennanp ANTENNA_750 (.A(_00197_));
 sg13g2_antennanp ANTENNA_751 (.A(_00197_));
 sg13g2_antennanp ANTENNA_752 (.A(_00228_));
 sg13g2_antennanp ANTENNA_753 (.A(_00235_));
 sg13g2_antennanp ANTENNA_754 (.A(_00930_));
 sg13g2_antennanp ANTENNA_755 (.A(_01052_));
 sg13g2_antennanp ANTENNA_756 (.A(_01052_));
 sg13g2_antennanp ANTENNA_757 (.A(_02950_));
 sg13g2_antennanp ANTENNA_758 (.A(_02950_));
 sg13g2_antennanp ANTENNA_759 (.A(_02950_));
 sg13g2_antennanp ANTENNA_760 (.A(_02950_));
 sg13g2_antennanp ANTENNA_761 (.A(_02950_));
 sg13g2_antennanp ANTENNA_762 (.A(_02950_));
 sg13g2_antennanp ANTENNA_763 (.A(_02953_));
 sg13g2_antennanp ANTENNA_764 (.A(_02953_));
 sg13g2_antennanp ANTENNA_765 (.A(_02953_));
 sg13g2_antennanp ANTENNA_766 (.A(_02953_));
 sg13g2_antennanp ANTENNA_767 (.A(_02965_));
 sg13g2_antennanp ANTENNA_768 (.A(_02965_));
 sg13g2_antennanp ANTENNA_769 (.A(_02965_));
 sg13g2_antennanp ANTENNA_770 (.A(_02965_));
 sg13g2_antennanp ANTENNA_771 (.A(_02965_));
 sg13g2_antennanp ANTENNA_772 (.A(_02965_));
 sg13g2_antennanp ANTENNA_773 (.A(_02965_));
 sg13g2_antennanp ANTENNA_774 (.A(_02965_));
 sg13g2_antennanp ANTENNA_775 (.A(_02965_));
 sg13g2_antennanp ANTENNA_776 (.A(_03429_));
 sg13g2_antennanp ANTENNA_777 (.A(_03429_));
 sg13g2_antennanp ANTENNA_778 (.A(_03429_));
 sg13g2_antennanp ANTENNA_779 (.A(_03429_));
 sg13g2_antennanp ANTENNA_780 (.A(_03435_));
 sg13g2_antennanp ANTENNA_781 (.A(_03435_));
 sg13g2_antennanp ANTENNA_782 (.A(_03435_));
 sg13g2_antennanp ANTENNA_783 (.A(_03435_));
 sg13g2_antennanp ANTENNA_784 (.A(_03435_));
 sg13g2_antennanp ANTENNA_785 (.A(_03435_));
 sg13g2_antennanp ANTENNA_786 (.A(_03435_));
 sg13g2_antennanp ANTENNA_787 (.A(_03435_));
 sg13g2_antennanp ANTENNA_788 (.A(_03435_));
 sg13g2_antennanp ANTENNA_789 (.A(_04212_));
 sg13g2_antennanp ANTENNA_790 (.A(_04212_));
 sg13g2_antennanp ANTENNA_791 (.A(_04212_));
 sg13g2_antennanp ANTENNA_792 (.A(_04212_));
 sg13g2_antennanp ANTENNA_793 (.A(_04212_));
 sg13g2_antennanp ANTENNA_794 (.A(_04742_));
 sg13g2_antennanp ANTENNA_795 (.A(_04742_));
 sg13g2_antennanp ANTENNA_796 (.A(_04742_));
 sg13g2_antennanp ANTENNA_797 (.A(_04742_));
 sg13g2_antennanp ANTENNA_798 (.A(_04887_));
 sg13g2_antennanp ANTENNA_799 (.A(_04887_));
 sg13g2_antennanp ANTENNA_800 (.A(_04887_));
 sg13g2_antennanp ANTENNA_801 (.A(_04887_));
 sg13g2_antennanp ANTENNA_802 (.A(_04894_));
 sg13g2_antennanp ANTENNA_803 (.A(_05013_));
 sg13g2_antennanp ANTENNA_804 (.A(_05013_));
 sg13g2_antennanp ANTENNA_805 (.A(_05015_));
 sg13g2_antennanp ANTENNA_806 (.A(_05169_));
 sg13g2_antennanp ANTENNA_807 (.A(_05280_));
 sg13g2_antennanp ANTENNA_808 (.A(_05372_));
 sg13g2_antennanp ANTENNA_809 (.A(_05432_));
 sg13g2_antennanp ANTENNA_810 (.A(_05442_));
 sg13g2_antennanp ANTENNA_811 (.A(_05442_));
 sg13g2_antennanp ANTENNA_812 (.A(_05508_));
 sg13g2_antennanp ANTENNA_813 (.A(_05646_));
 sg13g2_antennanp ANTENNA_814 (.A(_05650_));
 sg13g2_antennanp ANTENNA_815 (.A(_05654_));
 sg13g2_antennanp ANTENNA_816 (.A(_05654_));
 sg13g2_antennanp ANTENNA_817 (.A(_05742_));
 sg13g2_antennanp ANTENNA_818 (.A(_05760_));
 sg13g2_antennanp ANTENNA_819 (.A(_05760_));
 sg13g2_antennanp ANTENNA_820 (.A(_05763_));
 sg13g2_antennanp ANTENNA_821 (.A(_05763_));
 sg13g2_antennanp ANTENNA_822 (.A(_05763_));
 sg13g2_antennanp ANTENNA_823 (.A(_05763_));
 sg13g2_antennanp ANTENNA_824 (.A(_05763_));
 sg13g2_antennanp ANTENNA_825 (.A(_05763_));
 sg13g2_antennanp ANTENNA_826 (.A(_05763_));
 sg13g2_antennanp ANTENNA_827 (.A(_05766_));
 sg13g2_antennanp ANTENNA_828 (.A(_05766_));
 sg13g2_antennanp ANTENNA_829 (.A(_05766_));
 sg13g2_antennanp ANTENNA_830 (.A(_05766_));
 sg13g2_antennanp ANTENNA_831 (.A(_05775_));
 sg13g2_antennanp ANTENNA_832 (.A(_05775_));
 sg13g2_antennanp ANTENNA_833 (.A(_05775_));
 sg13g2_antennanp ANTENNA_834 (.A(_05785_));
 sg13g2_antennanp ANTENNA_835 (.A(_05785_));
 sg13g2_antennanp ANTENNA_836 (.A(_05785_));
 sg13g2_antennanp ANTENNA_837 (.A(_05835_));
 sg13g2_antennanp ANTENNA_838 (.A(_05835_));
 sg13g2_antennanp ANTENNA_839 (.A(_05835_));
 sg13g2_antennanp ANTENNA_840 (.A(_05835_));
 sg13g2_antennanp ANTENNA_841 (.A(_06843_));
 sg13g2_antennanp ANTENNA_842 (.A(_06843_));
 sg13g2_antennanp ANTENNA_843 (.A(_06843_));
 sg13g2_antennanp ANTENNA_844 (.A(_07398_));
 sg13g2_antennanp ANTENNA_845 (.A(_07433_));
 sg13g2_antennanp ANTENNA_846 (.A(_07434_));
 sg13g2_antennanp ANTENNA_847 (.A(_08297_));
 sg13g2_antennanp ANTENNA_848 (.A(_08297_));
 sg13g2_antennanp ANTENNA_849 (.A(_08502_));
 sg13g2_antennanp ANTENNA_850 (.A(_08502_));
 sg13g2_antennanp ANTENNA_851 (.A(_08502_));
 sg13g2_antennanp ANTENNA_852 (.A(_08502_));
 sg13g2_antennanp ANTENNA_853 (.A(_08502_));
 sg13g2_antennanp ANTENNA_854 (.A(_08502_));
 sg13g2_antennanp ANTENNA_855 (.A(_08502_));
 sg13g2_antennanp ANTENNA_856 (.A(_08502_));
 sg13g2_antennanp ANTENNA_857 (.A(_08502_));
 sg13g2_antennanp ANTENNA_858 (.A(_08502_));
 sg13g2_antennanp ANTENNA_859 (.A(_08502_));
 sg13g2_antennanp ANTENNA_860 (.A(_08502_));
 sg13g2_antennanp ANTENNA_861 (.A(_08533_));
 sg13g2_antennanp ANTENNA_862 (.A(_08533_));
 sg13g2_antennanp ANTENNA_863 (.A(_08533_));
 sg13g2_antennanp ANTENNA_864 (.A(_08533_));
 sg13g2_antennanp ANTENNA_865 (.A(_08533_));
 sg13g2_antennanp ANTENNA_866 (.A(_08533_));
 sg13g2_antennanp ANTENNA_867 (.A(_08558_));
 sg13g2_antennanp ANTENNA_868 (.A(_08558_));
 sg13g2_antennanp ANTENNA_869 (.A(_08558_));
 sg13g2_antennanp ANTENNA_870 (.A(_08634_));
 sg13g2_antennanp ANTENNA_871 (.A(_08634_));
 sg13g2_antennanp ANTENNA_872 (.A(_08634_));
 sg13g2_antennanp ANTENNA_873 (.A(_08634_));
 sg13g2_antennanp ANTENNA_874 (.A(_08634_));
 sg13g2_antennanp ANTENNA_875 (.A(_08634_));
 sg13g2_antennanp ANTENNA_876 (.A(_08634_));
 sg13g2_antennanp ANTENNA_877 (.A(_08634_));
 sg13g2_antennanp ANTENNA_878 (.A(_08634_));
 sg13g2_antennanp ANTENNA_879 (.A(_08679_));
 sg13g2_antennanp ANTENNA_880 (.A(_08679_));
 sg13g2_antennanp ANTENNA_881 (.A(_08679_));
 sg13g2_antennanp ANTENNA_882 (.A(_08679_));
 sg13g2_antennanp ANTENNA_883 (.A(_08679_));
 sg13g2_antennanp ANTENNA_884 (.A(_08689_));
 sg13g2_antennanp ANTENNA_885 (.A(_08689_));
 sg13g2_antennanp ANTENNA_886 (.A(_08689_));
 sg13g2_antennanp ANTENNA_887 (.A(_08689_));
 sg13g2_antennanp ANTENNA_888 (.A(_08689_));
 sg13g2_antennanp ANTENNA_889 (.A(_08698_));
 sg13g2_antennanp ANTENNA_890 (.A(_08698_));
 sg13g2_antennanp ANTENNA_891 (.A(_08698_));
 sg13g2_antennanp ANTENNA_892 (.A(_08728_));
 sg13g2_antennanp ANTENNA_893 (.A(_08728_));
 sg13g2_antennanp ANTENNA_894 (.A(_08728_));
 sg13g2_antennanp ANTENNA_895 (.A(_08728_));
 sg13g2_antennanp ANTENNA_896 (.A(_08759_));
 sg13g2_antennanp ANTENNA_897 (.A(_08759_));
 sg13g2_antennanp ANTENNA_898 (.A(_08759_));
 sg13g2_antennanp ANTENNA_899 (.A(_08759_));
 sg13g2_antennanp ANTENNA_900 (.A(_08853_));
 sg13g2_antennanp ANTENNA_901 (.A(_08938_));
 sg13g2_antennanp ANTENNA_902 (.A(_08959_));
 sg13g2_antennanp ANTENNA_903 (.A(_08970_));
 sg13g2_antennanp ANTENNA_904 (.A(_08970_));
 sg13g2_antennanp ANTENNA_905 (.A(_08970_));
 sg13g2_antennanp ANTENNA_906 (.A(_08970_));
 sg13g2_antennanp ANTENNA_907 (.A(_09167_));
 sg13g2_antennanp ANTENNA_908 (.A(_09277_));
 sg13g2_antennanp ANTENNA_909 (.A(_09277_));
 sg13g2_antennanp ANTENNA_910 (.A(_09277_));
 sg13g2_antennanp ANTENNA_911 (.A(_09277_));
 sg13g2_antennanp ANTENNA_912 (.A(_09277_));
 sg13g2_antennanp ANTENNA_913 (.A(_09277_));
 sg13g2_antennanp ANTENNA_914 (.A(_09320_));
 sg13g2_antennanp ANTENNA_915 (.A(_09320_));
 sg13g2_antennanp ANTENNA_916 (.A(_09320_));
 sg13g2_antennanp ANTENNA_917 (.A(_09320_));
 sg13g2_antennanp ANTENNA_918 (.A(_09320_));
 sg13g2_antennanp ANTENNA_919 (.A(_09320_));
 sg13g2_antennanp ANTENNA_920 (.A(_09320_));
 sg13g2_antennanp ANTENNA_921 (.A(_09320_));
 sg13g2_antennanp ANTENNA_922 (.A(_09336_));
 sg13g2_antennanp ANTENNA_923 (.A(_09336_));
 sg13g2_antennanp ANTENNA_924 (.A(_09349_));
 sg13g2_antennanp ANTENNA_925 (.A(_09349_));
 sg13g2_antennanp ANTENNA_926 (.A(_09349_));
 sg13g2_antennanp ANTENNA_927 (.A(_09349_));
 sg13g2_antennanp ANTENNA_928 (.A(_09349_));
 sg13g2_antennanp ANTENNA_929 (.A(_09349_));
 sg13g2_antennanp ANTENNA_930 (.A(_09349_));
 sg13g2_antennanp ANTENNA_931 (.A(_09349_));
 sg13g2_antennanp ANTENNA_932 (.A(_09349_));
 sg13g2_antennanp ANTENNA_933 (.A(_09349_));
 sg13g2_antennanp ANTENNA_934 (.A(_09351_));
 sg13g2_antennanp ANTENNA_935 (.A(_09351_));
 sg13g2_antennanp ANTENNA_936 (.A(_09351_));
 sg13g2_antennanp ANTENNA_937 (.A(_09351_));
 sg13g2_antennanp ANTENNA_938 (.A(_09351_));
 sg13g2_antennanp ANTENNA_939 (.A(_09351_));
 sg13g2_antennanp ANTENNA_940 (.A(_09351_));
 sg13g2_antennanp ANTENNA_941 (.A(_09351_));
 sg13g2_antennanp ANTENNA_942 (.A(_09351_));
 sg13g2_antennanp ANTENNA_943 (.A(_09351_));
 sg13g2_antennanp ANTENNA_944 (.A(_09351_));
 sg13g2_antennanp ANTENNA_945 (.A(_09351_));
 sg13g2_antennanp ANTENNA_946 (.A(_09380_));
 sg13g2_antennanp ANTENNA_947 (.A(_09380_));
 sg13g2_antennanp ANTENNA_948 (.A(_09380_));
 sg13g2_antennanp ANTENNA_949 (.A(_09380_));
 sg13g2_antennanp ANTENNA_950 (.A(_09386_));
 sg13g2_antennanp ANTENNA_951 (.A(_09386_));
 sg13g2_antennanp ANTENNA_952 (.A(_09386_));
 sg13g2_antennanp ANTENNA_953 (.A(_09386_));
 sg13g2_antennanp ANTENNA_954 (.A(_09386_));
 sg13g2_antennanp ANTENNA_955 (.A(_09386_));
 sg13g2_antennanp ANTENNA_956 (.A(_09386_));
 sg13g2_antennanp ANTENNA_957 (.A(_09386_));
 sg13g2_antennanp ANTENNA_958 (.A(_09388_));
 sg13g2_antennanp ANTENNA_959 (.A(_09388_));
 sg13g2_antennanp ANTENNA_960 (.A(_09388_));
 sg13g2_antennanp ANTENNA_961 (.A(_09388_));
 sg13g2_antennanp ANTENNA_962 (.A(_09388_));
 sg13g2_antennanp ANTENNA_963 (.A(_09388_));
 sg13g2_antennanp ANTENNA_964 (.A(_09389_));
 sg13g2_antennanp ANTENNA_965 (.A(_09389_));
 sg13g2_antennanp ANTENNA_966 (.A(_09389_));
 sg13g2_antennanp ANTENNA_967 (.A(_09389_));
 sg13g2_antennanp ANTENNA_968 (.A(_09389_));
 sg13g2_antennanp ANTENNA_969 (.A(_09389_));
 sg13g2_antennanp ANTENNA_970 (.A(_09389_));
 sg13g2_antennanp ANTENNA_971 (.A(_09389_));
 sg13g2_antennanp ANTENNA_972 (.A(_09389_));
 sg13g2_antennanp ANTENNA_973 (.A(_09390_));
 sg13g2_antennanp ANTENNA_974 (.A(_09390_));
 sg13g2_antennanp ANTENNA_975 (.A(_09390_));
 sg13g2_antennanp ANTENNA_976 (.A(_09444_));
 sg13g2_antennanp ANTENNA_977 (.A(_09444_));
 sg13g2_antennanp ANTENNA_978 (.A(_09444_));
 sg13g2_antennanp ANTENNA_979 (.A(_09444_));
 sg13g2_antennanp ANTENNA_980 (.A(_09444_));
 sg13g2_antennanp ANTENNA_981 (.A(_09444_));
 sg13g2_antennanp ANTENNA_982 (.A(_09444_));
 sg13g2_antennanp ANTENNA_983 (.A(_09444_));
 sg13g2_antennanp ANTENNA_984 (.A(_09444_));
 sg13g2_antennanp ANTENNA_985 (.A(_09444_));
 sg13g2_antennanp ANTENNA_986 (.A(_09444_));
 sg13g2_antennanp ANTENNA_987 (.A(_09444_));
 sg13g2_antennanp ANTENNA_988 (.A(_09445_));
 sg13g2_antennanp ANTENNA_989 (.A(_09445_));
 sg13g2_antennanp ANTENNA_990 (.A(_09445_));
 sg13g2_antennanp ANTENNA_991 (.A(_09445_));
 sg13g2_antennanp ANTENNA_992 (.A(_09445_));
 sg13g2_antennanp ANTENNA_993 (.A(_09445_));
 sg13g2_antennanp ANTENNA_994 (.A(_09554_));
 sg13g2_antennanp ANTENNA_995 (.A(_09562_));
 sg13g2_antennanp ANTENNA_996 (.A(_09587_));
 sg13g2_antennanp ANTENNA_997 (.A(_09608_));
 sg13g2_antennanp ANTENNA_998 (.A(_09665_));
 sg13g2_antennanp ANTENNA_999 (.A(_09695_));
 sg13g2_antennanp ANTENNA_1000 (.A(_09721_));
 sg13g2_antennanp ANTENNA_1001 (.A(_09742_));
 sg13g2_antennanp ANTENNA_1002 (.A(_09765_));
 sg13g2_antennanp ANTENNA_1003 (.A(_09794_));
 sg13g2_antennanp ANTENNA_1004 (.A(_09796_));
 sg13g2_antennanp ANTENNA_1005 (.A(_09836_));
 sg13g2_antennanp ANTENNA_1006 (.A(_09836_));
 sg13g2_antennanp ANTENNA_1007 (.A(_09836_));
 sg13g2_antennanp ANTENNA_1008 (.A(_09836_));
 sg13g2_antennanp ANTENNA_1009 (.A(_09836_));
 sg13g2_antennanp ANTENNA_1010 (.A(_09836_));
 sg13g2_antennanp ANTENNA_1011 (.A(_09836_));
 sg13g2_antennanp ANTENNA_1012 (.A(_09836_));
 sg13g2_antennanp ANTENNA_1013 (.A(_09836_));
 sg13g2_antennanp ANTENNA_1014 (.A(_09912_));
 sg13g2_antennanp ANTENNA_1015 (.A(_09990_));
 sg13g2_antennanp ANTENNA_1016 (.A(_09990_));
 sg13g2_antennanp ANTENNA_1017 (.A(_09990_));
 sg13g2_antennanp ANTENNA_1018 (.A(_09990_));
 sg13g2_antennanp ANTENNA_1019 (.A(_09990_));
 sg13g2_antennanp ANTENNA_1020 (.A(_09990_));
 sg13g2_antennanp ANTENNA_1021 (.A(_09990_));
 sg13g2_antennanp ANTENNA_1022 (.A(_09990_));
 sg13g2_antennanp ANTENNA_1023 (.A(_09990_));
 sg13g2_antennanp ANTENNA_1024 (.A(_09990_));
 sg13g2_antennanp ANTENNA_1025 (.A(_10172_));
 sg13g2_antennanp ANTENNA_1026 (.A(_10172_));
 sg13g2_antennanp ANTENNA_1027 (.A(_10172_));
 sg13g2_antennanp ANTENNA_1028 (.A(_10172_));
 sg13g2_antennanp ANTENNA_1029 (.A(_10172_));
 sg13g2_antennanp ANTENNA_1030 (.A(_10172_));
 sg13g2_antennanp ANTENNA_1031 (.A(_10172_));
 sg13g2_antennanp ANTENNA_1032 (.A(_10172_));
 sg13g2_antennanp ANTENNA_1033 (.A(_10240_));
 sg13g2_antennanp ANTENNA_1034 (.A(_10240_));
 sg13g2_antennanp ANTENNA_1035 (.A(_10240_));
 sg13g2_antennanp ANTENNA_1036 (.A(_10240_));
 sg13g2_antennanp ANTENNA_1037 (.A(_10246_));
 sg13g2_antennanp ANTENNA_1038 (.A(_10246_));
 sg13g2_antennanp ANTENNA_1039 (.A(_10246_));
 sg13g2_antennanp ANTENNA_1040 (.A(_10246_));
 sg13g2_antennanp ANTENNA_1041 (.A(_10246_));
 sg13g2_antennanp ANTENNA_1042 (.A(_10302_));
 sg13g2_antennanp ANTENNA_1043 (.A(_10302_));
 sg13g2_antennanp ANTENNA_1044 (.A(_10302_));
 sg13g2_antennanp ANTENNA_1045 (.A(_10302_));
 sg13g2_antennanp ANTENNA_1046 (.A(_10302_));
 sg13g2_antennanp ANTENNA_1047 (.A(_10302_));
 sg13g2_antennanp ANTENNA_1048 (.A(_10302_));
 sg13g2_antennanp ANTENNA_1049 (.A(_10302_));
 sg13g2_antennanp ANTENNA_1050 (.A(_10302_));
 sg13g2_antennanp ANTENNA_1051 (.A(_10302_));
 sg13g2_antennanp ANTENNA_1052 (.A(_10302_));
 sg13g2_antennanp ANTENNA_1053 (.A(_10302_));
 sg13g2_antennanp ANTENNA_1054 (.A(_10302_));
 sg13g2_antennanp ANTENNA_1055 (.A(_10302_));
 sg13g2_antennanp ANTENNA_1056 (.A(_10302_));
 sg13g2_antennanp ANTENNA_1057 (.A(_10302_));
 sg13g2_antennanp ANTENNA_1058 (.A(_10302_));
 sg13g2_antennanp ANTENNA_1059 (.A(_10302_));
 sg13g2_antennanp ANTENNA_1060 (.A(_10302_));
 sg13g2_antennanp ANTENNA_1061 (.A(_10302_));
 sg13g2_antennanp ANTENNA_1062 (.A(_10307_));
 sg13g2_antennanp ANTENNA_1063 (.A(_10307_));
 sg13g2_antennanp ANTENNA_1064 (.A(_10307_));
 sg13g2_antennanp ANTENNA_1065 (.A(_10307_));
 sg13g2_antennanp ANTENNA_1066 (.A(_10307_));
 sg13g2_antennanp ANTENNA_1067 (.A(_10307_));
 sg13g2_antennanp ANTENNA_1068 (.A(_10307_));
 sg13g2_antennanp ANTENNA_1069 (.A(_10307_));
 sg13g2_antennanp ANTENNA_1070 (.A(_10312_));
 sg13g2_antennanp ANTENNA_1071 (.A(_10312_));
 sg13g2_antennanp ANTENNA_1072 (.A(_10312_));
 sg13g2_antennanp ANTENNA_1073 (.A(_10312_));
 sg13g2_antennanp ANTENNA_1074 (.A(_10312_));
 sg13g2_antennanp ANTENNA_1075 (.A(_10312_));
 sg13g2_antennanp ANTENNA_1076 (.A(_10312_));
 sg13g2_antennanp ANTENNA_1077 (.A(_10312_));
 sg13g2_antennanp ANTENNA_1078 (.A(_10326_));
 sg13g2_antennanp ANTENNA_1079 (.A(_10326_));
 sg13g2_antennanp ANTENNA_1080 (.A(_10326_));
 sg13g2_antennanp ANTENNA_1081 (.A(_10326_));
 sg13g2_antennanp ANTENNA_1082 (.A(_10326_));
 sg13g2_antennanp ANTENNA_1083 (.A(_10326_));
 sg13g2_antennanp ANTENNA_1084 (.A(_10326_));
 sg13g2_antennanp ANTENNA_1085 (.A(_10326_));
 sg13g2_antennanp ANTENNA_1086 (.A(_10339_));
 sg13g2_antennanp ANTENNA_1087 (.A(_10339_));
 sg13g2_antennanp ANTENNA_1088 (.A(_10339_));
 sg13g2_antennanp ANTENNA_1089 (.A(_10339_));
 sg13g2_antennanp ANTENNA_1090 (.A(_10339_));
 sg13g2_antennanp ANTENNA_1091 (.A(_10339_));
 sg13g2_antennanp ANTENNA_1092 (.A(_10339_));
 sg13g2_antennanp ANTENNA_1093 (.A(_10339_));
 sg13g2_antennanp ANTENNA_1094 (.A(_10344_));
 sg13g2_antennanp ANTENNA_1095 (.A(_10344_));
 sg13g2_antennanp ANTENNA_1096 (.A(_10344_));
 sg13g2_antennanp ANTENNA_1097 (.A(_10344_));
 sg13g2_antennanp ANTENNA_1098 (.A(_10344_));
 sg13g2_antennanp ANTENNA_1099 (.A(_10344_));
 sg13g2_antennanp ANTENNA_1100 (.A(_10344_));
 sg13g2_antennanp ANTENNA_1101 (.A(_10344_));
 sg13g2_antennanp ANTENNA_1102 (.A(_10562_));
 sg13g2_antennanp ANTENNA_1103 (.A(_10562_));
 sg13g2_antennanp ANTENNA_1104 (.A(_10645_));
 sg13g2_antennanp ANTENNA_1105 (.A(_10645_));
 sg13g2_antennanp ANTENNA_1106 (.A(_11129_));
 sg13g2_antennanp ANTENNA_1107 (.A(_11129_));
 sg13g2_antennanp ANTENNA_1108 (.A(_12058_));
 sg13g2_antennanp ANTENNA_1109 (.A(_12058_));
 sg13g2_antennanp ANTENNA_1110 (.A(_12058_));
 sg13g2_antennanp ANTENNA_1111 (.A(_12058_));
 sg13g2_antennanp ANTENNA_1112 (.A(_12058_));
 sg13g2_antennanp ANTENNA_1113 (.A(_12058_));
 sg13g2_antennanp ANTENNA_1114 (.A(_12058_));
 sg13g2_antennanp ANTENNA_1115 (.A(_12058_));
 sg13g2_antennanp ANTENNA_1116 (.A(_12058_));
 sg13g2_antennanp ANTENNA_1117 (.A(_12127_));
 sg13g2_antennanp ANTENNA_1118 (.A(_12127_));
 sg13g2_antennanp ANTENNA_1119 (.A(_12127_));
 sg13g2_antennanp ANTENNA_1120 (.A(_12127_));
 sg13g2_antennanp ANTENNA_1121 (.A(_12127_));
 sg13g2_antennanp ANTENNA_1122 (.A(_12127_));
 sg13g2_antennanp ANTENNA_1123 (.A(_12127_));
 sg13g2_antennanp ANTENNA_1124 (.A(_12127_));
 sg13g2_antennanp ANTENNA_1125 (.A(_12127_));
 sg13g2_antennanp ANTENNA_1126 (.A(_12152_));
 sg13g2_antennanp ANTENNA_1127 (.A(_12152_));
 sg13g2_antennanp ANTENNA_1128 (.A(_12152_));
 sg13g2_antennanp ANTENNA_1129 (.A(_12152_));
 sg13g2_antennanp ANTENNA_1130 (.A(_12152_));
 sg13g2_antennanp ANTENNA_1131 (.A(_12152_));
 sg13g2_antennanp ANTENNA_1132 (.A(_12152_));
 sg13g2_antennanp ANTENNA_1133 (.A(_12152_));
 sg13g2_antennanp ANTENNA_1134 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1135 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1136 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1137 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1138 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1139 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1140 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1141 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1142 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1143 (.A(_12223_));
 sg13g2_antennanp ANTENNA_1144 (.A(_12223_));
 sg13g2_antennanp ANTENNA_1145 (.A(_12223_));
 sg13g2_antennanp ANTENNA_1146 (.A(_12223_));
 sg13g2_antennanp ANTENNA_1147 (.A(_12223_));
 sg13g2_antennanp ANTENNA_1148 (.A(_12223_));
 sg13g2_antennanp ANTENNA_1149 (.A(_12223_));
 sg13g2_antennanp ANTENNA_1150 (.A(_12223_));
 sg13g2_antennanp ANTENNA_1151 (.A(_12223_));
 sg13g2_antennanp ANTENNA_1152 (.A(_12229_));
 sg13g2_antennanp ANTENNA_1153 (.A(_12229_));
 sg13g2_antennanp ANTENNA_1154 (.A(_12229_));
 sg13g2_antennanp ANTENNA_1155 (.A(_12229_));
 sg13g2_antennanp ANTENNA_1156 (.A(_12229_));
 sg13g2_antennanp ANTENNA_1157 (.A(_12229_));
 sg13g2_antennanp ANTENNA_1158 (.A(_12229_));
 sg13g2_antennanp ANTENNA_1159 (.A(_12229_));
 sg13g2_antennanp ANTENNA_1160 (.A(_12229_));
 sg13g2_antennanp ANTENNA_1161 (.A(_12558_));
 sg13g2_antennanp ANTENNA_1162 (.A(_12558_));
 sg13g2_antennanp ANTENNA_1163 (.A(_12558_));
 sg13g2_antennanp ANTENNA_1164 (.A(_12558_));
 sg13g2_antennanp ANTENNA_1165 (.A(_12558_));
 sg13g2_antennanp ANTENNA_1166 (.A(_12726_));
 sg13g2_antennanp ANTENNA_1167 (.A(_12726_));
 sg13g2_antennanp ANTENNA_1168 (.A(_12726_));
 sg13g2_antennanp ANTENNA_1169 (.A(clk));
 sg13g2_antennanp ANTENNA_1170 (.A(clk));
 sg13g2_antennanp ANTENNA_1171 (.A(\cpu.ex.pc[3] ));
 sg13g2_antennanp ANTENNA_1172 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_1173 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_1174 (.A(net3));
 sg13g2_antennanp ANTENNA_1175 (.A(net3));
 sg13g2_antennanp ANTENNA_1176 (.A(net3));
 sg13g2_antennanp ANTENNA_1177 (.A(net12));
 sg13g2_antennanp ANTENNA_1178 (.A(net12));
 sg13g2_antennanp ANTENNA_1179 (.A(net12));
 sg13g2_antennanp ANTENNA_1180 (.A(net13));
 sg13g2_antennanp ANTENNA_1181 (.A(net13));
 sg13g2_antennanp ANTENNA_1182 (.A(net13));
 sg13g2_antennanp ANTENNA_1183 (.A(net14));
 sg13g2_antennanp ANTENNA_1184 (.A(net14));
 sg13g2_antennanp ANTENNA_1185 (.A(net14));
 sg13g2_antennanp ANTENNA_1186 (.A(net524));
 sg13g2_antennanp ANTENNA_1187 (.A(net524));
 sg13g2_antennanp ANTENNA_1188 (.A(net524));
 sg13g2_antennanp ANTENNA_1189 (.A(net524));
 sg13g2_antennanp ANTENNA_1190 (.A(net524));
 sg13g2_antennanp ANTENNA_1191 (.A(net524));
 sg13g2_antennanp ANTENNA_1192 (.A(net524));
 sg13g2_antennanp ANTENNA_1193 (.A(net524));
 sg13g2_antennanp ANTENNA_1194 (.A(net524));
 sg13g2_antennanp ANTENNA_1195 (.A(net524));
 sg13g2_antennanp ANTENNA_1196 (.A(net524));
 sg13g2_antennanp ANTENNA_1197 (.A(net524));
 sg13g2_antennanp ANTENNA_1198 (.A(net524));
 sg13g2_antennanp ANTENNA_1199 (.A(net542));
 sg13g2_antennanp ANTENNA_1200 (.A(net542));
 sg13g2_antennanp ANTENNA_1201 (.A(net542));
 sg13g2_antennanp ANTENNA_1202 (.A(net542));
 sg13g2_antennanp ANTENNA_1203 (.A(net542));
 sg13g2_antennanp ANTENNA_1204 (.A(net542));
 sg13g2_antennanp ANTENNA_1205 (.A(net542));
 sg13g2_antennanp ANTENNA_1206 (.A(net542));
 sg13g2_antennanp ANTENNA_1207 (.A(net542));
 sg13g2_antennanp ANTENNA_1208 (.A(net542));
 sg13g2_antennanp ANTENNA_1209 (.A(net542));
 sg13g2_antennanp ANTENNA_1210 (.A(net542));
 sg13g2_antennanp ANTENNA_1211 (.A(net542));
 sg13g2_antennanp ANTENNA_1212 (.A(net656));
 sg13g2_antennanp ANTENNA_1213 (.A(net656));
 sg13g2_antennanp ANTENNA_1214 (.A(net656));
 sg13g2_antennanp ANTENNA_1215 (.A(net656));
 sg13g2_antennanp ANTENNA_1216 (.A(net656));
 sg13g2_antennanp ANTENNA_1217 (.A(net656));
 sg13g2_antennanp ANTENNA_1218 (.A(net656));
 sg13g2_antennanp ANTENNA_1219 (.A(net656));
 sg13g2_antennanp ANTENNA_1220 (.A(net656));
 sg13g2_antennanp ANTENNA_1221 (.A(net656));
 sg13g2_antennanp ANTENNA_1222 (.A(net656));
 sg13g2_antennanp ANTENNA_1223 (.A(net656));
 sg13g2_antennanp ANTENNA_1224 (.A(net656));
 sg13g2_antennanp ANTENNA_1225 (.A(net656));
 sg13g2_antennanp ANTENNA_1226 (.A(net656));
 sg13g2_antennanp ANTENNA_1227 (.A(net656));
 sg13g2_antennanp ANTENNA_1228 (.A(net656));
 sg13g2_antennanp ANTENNA_1229 (.A(net656));
 sg13g2_antennanp ANTENNA_1230 (.A(net656));
 sg13g2_antennanp ANTENNA_1231 (.A(net707));
 sg13g2_antennanp ANTENNA_1232 (.A(net707));
 sg13g2_antennanp ANTENNA_1233 (.A(net707));
 sg13g2_antennanp ANTENNA_1234 (.A(net707));
 sg13g2_antennanp ANTENNA_1235 (.A(net707));
 sg13g2_antennanp ANTENNA_1236 (.A(net707));
 sg13g2_antennanp ANTENNA_1237 (.A(net707));
 sg13g2_antennanp ANTENNA_1238 (.A(net707));
 sg13g2_antennanp ANTENNA_1239 (.A(net707));
 sg13g2_antennanp ANTENNA_1240 (.A(net707));
 sg13g2_antennanp ANTENNA_1241 (.A(net707));
 sg13g2_antennanp ANTENNA_1242 (.A(net707));
 sg13g2_antennanp ANTENNA_1243 (.A(net707));
 sg13g2_antennanp ANTENNA_1244 (.A(net707));
 sg13g2_antennanp ANTENNA_1245 (.A(net707));
 sg13g2_antennanp ANTENNA_1246 (.A(net707));
 sg13g2_antennanp ANTENNA_1247 (.A(net707));
 sg13g2_antennanp ANTENNA_1248 (.A(net707));
 sg13g2_antennanp ANTENNA_1249 (.A(net707));
 sg13g2_antennanp ANTENNA_1250 (.A(net707));
 sg13g2_antennanp ANTENNA_1251 (.A(net707));
 sg13g2_antennanp ANTENNA_1252 (.A(net707));
 sg13g2_antennanp ANTENNA_1253 (.A(net707));
 sg13g2_antennanp ANTENNA_1254 (.A(net803));
 sg13g2_antennanp ANTENNA_1255 (.A(net803));
 sg13g2_antennanp ANTENNA_1256 (.A(net803));
 sg13g2_antennanp ANTENNA_1257 (.A(net803));
 sg13g2_antennanp ANTENNA_1258 (.A(net803));
 sg13g2_antennanp ANTENNA_1259 (.A(net803));
 sg13g2_antennanp ANTENNA_1260 (.A(net803));
 sg13g2_antennanp ANTENNA_1261 (.A(net803));
 sg13g2_antennanp ANTENNA_1262 (.A(net803));
 sg13g2_antennanp ANTENNA_1263 (.A(net803));
 sg13g2_antennanp ANTENNA_1264 (.A(net803));
 sg13g2_antennanp ANTENNA_1265 (.A(net803));
 sg13g2_antennanp ANTENNA_1266 (.A(net803));
 sg13g2_antennanp ANTENNA_1267 (.A(net803));
 sg13g2_antennanp ANTENNA_1268 (.A(net803));
 sg13g2_antennanp ANTENNA_1269 (.A(net803));
 sg13g2_antennanp ANTENNA_1270 (.A(net887));
 sg13g2_antennanp ANTENNA_1271 (.A(net887));
 sg13g2_antennanp ANTENNA_1272 (.A(net887));
 sg13g2_antennanp ANTENNA_1273 (.A(net887));
 sg13g2_antennanp ANTENNA_1274 (.A(net887));
 sg13g2_antennanp ANTENNA_1275 (.A(net887));
 sg13g2_antennanp ANTENNA_1276 (.A(net887));
 sg13g2_antennanp ANTENNA_1277 (.A(net887));
 sg13g2_antennanp ANTENNA_1278 (.A(net887));
 sg13g2_antennanp ANTENNA_1279 (.A(net928));
 sg13g2_antennanp ANTENNA_1280 (.A(net928));
 sg13g2_antennanp ANTENNA_1281 (.A(net928));
 sg13g2_antennanp ANTENNA_1282 (.A(net928));
 sg13g2_antennanp ANTENNA_1283 (.A(net928));
 sg13g2_antennanp ANTENNA_1284 (.A(net928));
 sg13g2_antennanp ANTENNA_1285 (.A(net928));
 sg13g2_antennanp ANTENNA_1286 (.A(net928));
 sg13g2_antennanp ANTENNA_1287 (.A(net928));
 sg13g2_antennanp ANTENNA_1288 (.A(net941));
 sg13g2_antennanp ANTENNA_1289 (.A(net941));
 sg13g2_antennanp ANTENNA_1290 (.A(net941));
 sg13g2_antennanp ANTENNA_1291 (.A(net941));
 sg13g2_antennanp ANTENNA_1292 (.A(net941));
 sg13g2_antennanp ANTENNA_1293 (.A(net941));
 sg13g2_antennanp ANTENNA_1294 (.A(net941));
 sg13g2_antennanp ANTENNA_1295 (.A(net941));
 sg13g2_antennanp ANTENNA_1296 (.A(net941));
 sg13g2_antennanp ANTENNA_1297 (.A(net982));
 sg13g2_antennanp ANTENNA_1298 (.A(net982));
 sg13g2_antennanp ANTENNA_1299 (.A(net982));
 sg13g2_antennanp ANTENNA_1300 (.A(net982));
 sg13g2_antennanp ANTENNA_1301 (.A(net982));
 sg13g2_antennanp ANTENNA_1302 (.A(net982));
 sg13g2_antennanp ANTENNA_1303 (.A(net982));
 sg13g2_antennanp ANTENNA_1304 (.A(net982));
 sg13g2_antennanp ANTENNA_1305 (.A(net982));
 sg13g2_antennanp ANTENNA_1306 (.A(net984));
 sg13g2_antennanp ANTENNA_1307 (.A(net984));
 sg13g2_antennanp ANTENNA_1308 (.A(net984));
 sg13g2_antennanp ANTENNA_1309 (.A(net984));
 sg13g2_antennanp ANTENNA_1310 (.A(net984));
 sg13g2_antennanp ANTENNA_1311 (.A(net984));
 sg13g2_antennanp ANTENNA_1312 (.A(net984));
 sg13g2_antennanp ANTENNA_1313 (.A(net984));
 sg13g2_antennanp ANTENNA_1314 (.A(net984));
 sg13g2_antennanp ANTENNA_1315 (.A(net984));
 sg13g2_antennanp ANTENNA_1316 (.A(net984));
 sg13g2_antennanp ANTENNA_1317 (.A(net984));
 sg13g2_antennanp ANTENNA_1318 (.A(net984));
 sg13g2_antennanp ANTENNA_1319 (.A(net984));
 sg13g2_antennanp ANTENNA_1320 (.A(net984));
 sg13g2_antennanp ANTENNA_1321 (.A(net984));
 sg13g2_antennanp ANTENNA_1322 (.A(net984));
 sg13g2_antennanp ANTENNA_1323 (.A(net984));
 sg13g2_antennanp ANTENNA_1324 (.A(net984));
 sg13g2_antennanp ANTENNA_1325 (.A(net984));
 sg13g2_antennanp ANTENNA_1326 (.A(net984));
 sg13g2_antennanp ANTENNA_1327 (.A(net984));
 sg13g2_antennanp ANTENNA_1328 (.A(net984));
 sg13g2_antennanp ANTENNA_1329 (.A(net984));
 sg13g2_antennanp ANTENNA_1330 (.A(net984));
 sg13g2_antennanp ANTENNA_1331 (.A(net984));
 sg13g2_antennanp ANTENNA_1332 (.A(net984));
 sg13g2_antennanp ANTENNA_1333 (.A(net984));
 sg13g2_antennanp ANTENNA_1334 (.A(net984));
 sg13g2_antennanp ANTENNA_1335 (.A(net984));
 sg13g2_antennanp ANTENNA_1336 (.A(net984));
 sg13g2_antennanp ANTENNA_1337 (.A(net984));
 sg13g2_antennanp ANTENNA_1338 (.A(net984));
 sg13g2_antennanp ANTENNA_1339 (.A(net984));
 sg13g2_antennanp ANTENNA_1340 (.A(net1004));
 sg13g2_antennanp ANTENNA_1341 (.A(net1004));
 sg13g2_antennanp ANTENNA_1342 (.A(net1004));
 sg13g2_antennanp ANTENNA_1343 (.A(net1004));
 sg13g2_antennanp ANTENNA_1344 (.A(net1004));
 sg13g2_antennanp ANTENNA_1345 (.A(net1004));
 sg13g2_antennanp ANTENNA_1346 (.A(net1004));
 sg13g2_antennanp ANTENNA_1347 (.A(net1004));
 sg13g2_antennanp ANTENNA_1348 (.A(net1004));
 sg13g2_antennanp ANTENNA_1349 (.A(net1004));
 sg13g2_antennanp ANTENNA_1350 (.A(net1004));
 sg13g2_antennanp ANTENNA_1351 (.A(net1004));
 sg13g2_antennanp ANTENNA_1352 (.A(net1004));
 sg13g2_antennanp ANTENNA_1353 (.A(net1004));
 sg13g2_antennanp ANTENNA_1354 (.A(net1004));
 sg13g2_antennanp ANTENNA_1355 (.A(net1004));
 sg13g2_antennanp ANTENNA_1356 (.A(net1004));
 sg13g2_antennanp ANTENNA_1357 (.A(net1004));
 sg13g2_antennanp ANTENNA_1358 (.A(net1004));
 sg13g2_antennanp ANTENNA_1359 (.A(net1004));
 sg13g2_antennanp ANTENNA_1360 (.A(net1004));
 sg13g2_antennanp ANTENNA_1361 (.A(net1004));
 sg13g2_antennanp ANTENNA_1362 (.A(net1004));
 sg13g2_antennanp ANTENNA_1363 (.A(net1004));
 sg13g2_antennanp ANTENNA_1364 (.A(net1004));
 sg13g2_antennanp ANTENNA_1365 (.A(net1004));
 sg13g2_antennanp ANTENNA_1366 (.A(net1004));
 sg13g2_antennanp ANTENNA_1367 (.A(net1004));
 sg13g2_antennanp ANTENNA_1368 (.A(net1004));
 sg13g2_antennanp ANTENNA_1369 (.A(net1004));
 sg13g2_antennanp ANTENNA_1370 (.A(net1004));
 sg13g2_antennanp ANTENNA_1371 (.A(net1004));
 sg13g2_antennanp ANTENNA_1372 (.A(net1004));
 sg13g2_antennanp ANTENNA_1373 (.A(net1075));
 sg13g2_antennanp ANTENNA_1374 (.A(net1075));
 sg13g2_antennanp ANTENNA_1375 (.A(net1075));
 sg13g2_antennanp ANTENNA_1376 (.A(net1075));
 sg13g2_antennanp ANTENNA_1377 (.A(net1075));
 sg13g2_antennanp ANTENNA_1378 (.A(net1075));
 sg13g2_antennanp ANTENNA_1379 (.A(net1075));
 sg13g2_antennanp ANTENNA_1380 (.A(net1075));
 sg13g2_antennanp ANTENNA_1381 (.A(net1075));
 sg13g2_antennanp ANTENNA_1382 (.A(_00190_));
 sg13g2_antennanp ANTENNA_1383 (.A(_00197_));
 sg13g2_antennanp ANTENNA_1384 (.A(_00197_));
 sg13g2_antennanp ANTENNA_1385 (.A(_00197_));
 sg13g2_antennanp ANTENNA_1386 (.A(_00197_));
 sg13g2_antennanp ANTENNA_1387 (.A(_00228_));
 sg13g2_antennanp ANTENNA_1388 (.A(_00228_));
 sg13g2_antennanp ANTENNA_1389 (.A(_00235_));
 sg13g2_antennanp ANTENNA_1390 (.A(_00235_));
 sg13g2_antennanp ANTENNA_1391 (.A(_00930_));
 sg13g2_antennanp ANTENNA_1392 (.A(_01052_));
 sg13g2_antennanp ANTENNA_1393 (.A(_01052_));
 sg13g2_antennanp ANTENNA_1394 (.A(_02950_));
 sg13g2_antennanp ANTENNA_1395 (.A(_02950_));
 sg13g2_antennanp ANTENNA_1396 (.A(_02950_));
 sg13g2_antennanp ANTENNA_1397 (.A(_02950_));
 sg13g2_antennanp ANTENNA_1398 (.A(_02950_));
 sg13g2_antennanp ANTENNA_1399 (.A(_02950_));
 sg13g2_antennanp ANTENNA_1400 (.A(_02950_));
 sg13g2_antennanp ANTENNA_1401 (.A(_02950_));
 sg13g2_antennanp ANTENNA_1402 (.A(_02950_));
 sg13g2_antennanp ANTENNA_1403 (.A(_02950_));
 sg13g2_antennanp ANTENNA_1404 (.A(_02953_));
 sg13g2_antennanp ANTENNA_1405 (.A(_02953_));
 sg13g2_antennanp ANTENNA_1406 (.A(_02953_));
 sg13g2_antennanp ANTENNA_1407 (.A(_02953_));
 sg13g2_antennanp ANTENNA_1408 (.A(_02965_));
 sg13g2_antennanp ANTENNA_1409 (.A(_02965_));
 sg13g2_antennanp ANTENNA_1410 (.A(_02965_));
 sg13g2_antennanp ANTENNA_1411 (.A(_02965_));
 sg13g2_antennanp ANTENNA_1412 (.A(_02965_));
 sg13g2_antennanp ANTENNA_1413 (.A(_02965_));
 sg13g2_antennanp ANTENNA_1414 (.A(_02965_));
 sg13g2_antennanp ANTENNA_1415 (.A(_02965_));
 sg13g2_antennanp ANTENNA_1416 (.A(_02965_));
 sg13g2_antennanp ANTENNA_1417 (.A(_03429_));
 sg13g2_antennanp ANTENNA_1418 (.A(_03429_));
 sg13g2_antennanp ANTENNA_1419 (.A(_03429_));
 sg13g2_antennanp ANTENNA_1420 (.A(_03429_));
 sg13g2_antennanp ANTENNA_1421 (.A(_03435_));
 sg13g2_antennanp ANTENNA_1422 (.A(_03435_));
 sg13g2_antennanp ANTENNA_1423 (.A(_03435_));
 sg13g2_antennanp ANTENNA_1424 (.A(_03435_));
 sg13g2_antennanp ANTENNA_1425 (.A(_03435_));
 sg13g2_antennanp ANTENNA_1426 (.A(_03435_));
 sg13g2_antennanp ANTENNA_1427 (.A(_03435_));
 sg13g2_antennanp ANTENNA_1428 (.A(_03435_));
 sg13g2_antennanp ANTENNA_1429 (.A(_03435_));
 sg13g2_antennanp ANTENNA_1430 (.A(_04212_));
 sg13g2_antennanp ANTENNA_1431 (.A(_04212_));
 sg13g2_antennanp ANTENNA_1432 (.A(_04212_));
 sg13g2_antennanp ANTENNA_1433 (.A(_04212_));
 sg13g2_antennanp ANTENNA_1434 (.A(_04212_));
 sg13g2_antennanp ANTENNA_1435 (.A(_04742_));
 sg13g2_antennanp ANTENNA_1436 (.A(_04742_));
 sg13g2_antennanp ANTENNA_1437 (.A(_04742_));
 sg13g2_antennanp ANTENNA_1438 (.A(_04742_));
 sg13g2_antennanp ANTENNA_1439 (.A(_04887_));
 sg13g2_antennanp ANTENNA_1440 (.A(_04887_));
 sg13g2_antennanp ANTENNA_1441 (.A(_04887_));
 sg13g2_antennanp ANTENNA_1442 (.A(_04887_));
 sg13g2_antennanp ANTENNA_1443 (.A(_04894_));
 sg13g2_antennanp ANTENNA_1444 (.A(_05013_));
 sg13g2_antennanp ANTENNA_1445 (.A(_05013_));
 sg13g2_antennanp ANTENNA_1446 (.A(_05015_));
 sg13g2_antennanp ANTENNA_1447 (.A(_05169_));
 sg13g2_antennanp ANTENNA_1448 (.A(_05278_));
 sg13g2_antennanp ANTENNA_1449 (.A(_05280_));
 sg13g2_antennanp ANTENNA_1450 (.A(_05372_));
 sg13g2_antennanp ANTENNA_1451 (.A(_05432_));
 sg13g2_antennanp ANTENNA_1452 (.A(_05442_));
 sg13g2_antennanp ANTENNA_1453 (.A(_05508_));
 sg13g2_antennanp ANTENNA_1454 (.A(_05646_));
 sg13g2_antennanp ANTENNA_1455 (.A(_05650_));
 sg13g2_antennanp ANTENNA_1456 (.A(_05654_));
 sg13g2_antennanp ANTENNA_1457 (.A(_05654_));
 sg13g2_antennanp ANTENNA_1458 (.A(_05742_));
 sg13g2_antennanp ANTENNA_1459 (.A(_05760_));
 sg13g2_antennanp ANTENNA_1460 (.A(_05760_));
 sg13g2_antennanp ANTENNA_1461 (.A(_05763_));
 sg13g2_antennanp ANTENNA_1462 (.A(_05763_));
 sg13g2_antennanp ANTENNA_1463 (.A(_05763_));
 sg13g2_antennanp ANTENNA_1464 (.A(_05763_));
 sg13g2_antennanp ANTENNA_1465 (.A(_05763_));
 sg13g2_antennanp ANTENNA_1466 (.A(_05763_));
 sg13g2_antennanp ANTENNA_1467 (.A(_05763_));
 sg13g2_antennanp ANTENNA_1468 (.A(_05766_));
 sg13g2_antennanp ANTENNA_1469 (.A(_05766_));
 sg13g2_antennanp ANTENNA_1470 (.A(_05766_));
 sg13g2_antennanp ANTENNA_1471 (.A(_05766_));
 sg13g2_antennanp ANTENNA_1472 (.A(_05770_));
 sg13g2_antennanp ANTENNA_1473 (.A(_05770_));
 sg13g2_antennanp ANTENNA_1474 (.A(_05770_));
 sg13g2_antennanp ANTENNA_1475 (.A(_05775_));
 sg13g2_antennanp ANTENNA_1476 (.A(_05775_));
 sg13g2_antennanp ANTENNA_1477 (.A(_05775_));
 sg13g2_antennanp ANTENNA_1478 (.A(_05785_));
 sg13g2_antennanp ANTENNA_1479 (.A(_05785_));
 sg13g2_antennanp ANTENNA_1480 (.A(_05785_));
 sg13g2_antennanp ANTENNA_1481 (.A(_05835_));
 sg13g2_antennanp ANTENNA_1482 (.A(_05835_));
 sg13g2_antennanp ANTENNA_1483 (.A(_05835_));
 sg13g2_antennanp ANTENNA_1484 (.A(_05835_));
 sg13g2_antennanp ANTENNA_1485 (.A(_06843_));
 sg13g2_antennanp ANTENNA_1486 (.A(_06843_));
 sg13g2_antennanp ANTENNA_1487 (.A(_06843_));
 sg13g2_antennanp ANTENNA_1488 (.A(_07398_));
 sg13g2_antennanp ANTENNA_1489 (.A(_07433_));
 sg13g2_antennanp ANTENNA_1490 (.A(_07434_));
 sg13g2_antennanp ANTENNA_1491 (.A(_08297_));
 sg13g2_antennanp ANTENNA_1492 (.A(_08297_));
 sg13g2_antennanp ANTENNA_1493 (.A(_08502_));
 sg13g2_antennanp ANTENNA_1494 (.A(_08502_));
 sg13g2_antennanp ANTENNA_1495 (.A(_08502_));
 sg13g2_antennanp ANTENNA_1496 (.A(_08502_));
 sg13g2_antennanp ANTENNA_1497 (.A(_08502_));
 sg13g2_antennanp ANTENNA_1498 (.A(_08502_));
 sg13g2_antennanp ANTENNA_1499 (.A(_08502_));
 sg13g2_antennanp ANTENNA_1500 (.A(_08533_));
 sg13g2_antennanp ANTENNA_1501 (.A(_08533_));
 sg13g2_antennanp ANTENNA_1502 (.A(_08533_));
 sg13g2_antennanp ANTENNA_1503 (.A(_08533_));
 sg13g2_antennanp ANTENNA_1504 (.A(_08533_));
 sg13g2_antennanp ANTENNA_1505 (.A(_08533_));
 sg13g2_antennanp ANTENNA_1506 (.A(_08558_));
 sg13g2_antennanp ANTENNA_1507 (.A(_08558_));
 sg13g2_antennanp ANTENNA_1508 (.A(_08558_));
 sg13g2_antennanp ANTENNA_1509 (.A(_08558_));
 sg13g2_antennanp ANTENNA_1510 (.A(_08558_));
 sg13g2_antennanp ANTENNA_1511 (.A(_08558_));
 sg13g2_antennanp ANTENNA_1512 (.A(_08558_));
 sg13g2_antennanp ANTENNA_1513 (.A(_08558_));
 sg13g2_antennanp ANTENNA_1514 (.A(_08558_));
 sg13g2_antennanp ANTENNA_1515 (.A(_08634_));
 sg13g2_antennanp ANTENNA_1516 (.A(_08634_));
 sg13g2_antennanp ANTENNA_1517 (.A(_08634_));
 sg13g2_antennanp ANTENNA_1518 (.A(_08634_));
 sg13g2_antennanp ANTENNA_1519 (.A(_08634_));
 sg13g2_antennanp ANTENNA_1520 (.A(_08634_));
 sg13g2_antennanp ANTENNA_1521 (.A(_08634_));
 sg13g2_antennanp ANTENNA_1522 (.A(_08634_));
 sg13g2_antennanp ANTENNA_1523 (.A(_08634_));
 sg13g2_antennanp ANTENNA_1524 (.A(_08679_));
 sg13g2_antennanp ANTENNA_1525 (.A(_08679_));
 sg13g2_antennanp ANTENNA_1526 (.A(_08679_));
 sg13g2_antennanp ANTENNA_1527 (.A(_08689_));
 sg13g2_antennanp ANTENNA_1528 (.A(_08689_));
 sg13g2_antennanp ANTENNA_1529 (.A(_08689_));
 sg13g2_antennanp ANTENNA_1530 (.A(_08689_));
 sg13g2_antennanp ANTENNA_1531 (.A(_08689_));
 sg13g2_antennanp ANTENNA_1532 (.A(_08698_));
 sg13g2_antennanp ANTENNA_1533 (.A(_08698_));
 sg13g2_antennanp ANTENNA_1534 (.A(_08698_));
 sg13g2_antennanp ANTENNA_1535 (.A(_08728_));
 sg13g2_antennanp ANTENNA_1536 (.A(_08728_));
 sg13g2_antennanp ANTENNA_1537 (.A(_08728_));
 sg13g2_antennanp ANTENNA_1538 (.A(_08728_));
 sg13g2_antennanp ANTENNA_1539 (.A(_08759_));
 sg13g2_antennanp ANTENNA_1540 (.A(_08759_));
 sg13g2_antennanp ANTENNA_1541 (.A(_08759_));
 sg13g2_antennanp ANTENNA_1542 (.A(_08759_));
 sg13g2_antennanp ANTENNA_1543 (.A(_08853_));
 sg13g2_antennanp ANTENNA_1544 (.A(_08938_));
 sg13g2_antennanp ANTENNA_1545 (.A(_08959_));
 sg13g2_antennanp ANTENNA_1546 (.A(_08970_));
 sg13g2_antennanp ANTENNA_1547 (.A(_08970_));
 sg13g2_antennanp ANTENNA_1548 (.A(_08970_));
 sg13g2_antennanp ANTENNA_1549 (.A(_08970_));
 sg13g2_antennanp ANTENNA_1550 (.A(_09167_));
 sg13g2_antennanp ANTENNA_1551 (.A(_09336_));
 sg13g2_antennanp ANTENNA_1552 (.A(_09336_));
 sg13g2_antennanp ANTENNA_1553 (.A(_09349_));
 sg13g2_antennanp ANTENNA_1554 (.A(_09349_));
 sg13g2_antennanp ANTENNA_1555 (.A(_09349_));
 sg13g2_antennanp ANTENNA_1556 (.A(_09349_));
 sg13g2_antennanp ANTENNA_1557 (.A(_09349_));
 sg13g2_antennanp ANTENNA_1558 (.A(_09349_));
 sg13g2_antennanp ANTENNA_1559 (.A(_09349_));
 sg13g2_antennanp ANTENNA_1560 (.A(_09349_));
 sg13g2_antennanp ANTENNA_1561 (.A(_09349_));
 sg13g2_antennanp ANTENNA_1562 (.A(_09349_));
 sg13g2_antennanp ANTENNA_1563 (.A(_09380_));
 sg13g2_antennanp ANTENNA_1564 (.A(_09380_));
 sg13g2_antennanp ANTENNA_1565 (.A(_09380_));
 sg13g2_antennanp ANTENNA_1566 (.A(_09380_));
 sg13g2_antennanp ANTENNA_1567 (.A(_09386_));
 sg13g2_antennanp ANTENNA_1568 (.A(_09386_));
 sg13g2_antennanp ANTENNA_1569 (.A(_09386_));
 sg13g2_antennanp ANTENNA_1570 (.A(_09386_));
 sg13g2_antennanp ANTENNA_1571 (.A(_09386_));
 sg13g2_antennanp ANTENNA_1572 (.A(_09386_));
 sg13g2_antennanp ANTENNA_1573 (.A(_09386_));
 sg13g2_antennanp ANTENNA_1574 (.A(_09386_));
 sg13g2_antennanp ANTENNA_1575 (.A(_09388_));
 sg13g2_antennanp ANTENNA_1576 (.A(_09388_));
 sg13g2_antennanp ANTENNA_1577 (.A(_09388_));
 sg13g2_antennanp ANTENNA_1578 (.A(_09388_));
 sg13g2_antennanp ANTENNA_1579 (.A(_09388_));
 sg13g2_antennanp ANTENNA_1580 (.A(_09388_));
 sg13g2_antennanp ANTENNA_1581 (.A(_09389_));
 sg13g2_antennanp ANTENNA_1582 (.A(_09389_));
 sg13g2_antennanp ANTENNA_1583 (.A(_09389_));
 sg13g2_antennanp ANTENNA_1584 (.A(_09389_));
 sg13g2_antennanp ANTENNA_1585 (.A(_09390_));
 sg13g2_antennanp ANTENNA_1586 (.A(_09390_));
 sg13g2_antennanp ANTENNA_1587 (.A(_09390_));
 sg13g2_antennanp ANTENNA_1588 (.A(_09444_));
 sg13g2_antennanp ANTENNA_1589 (.A(_09444_));
 sg13g2_antennanp ANTENNA_1590 (.A(_09444_));
 sg13g2_antennanp ANTENNA_1591 (.A(_09444_));
 sg13g2_antennanp ANTENNA_1592 (.A(_09444_));
 sg13g2_antennanp ANTENNA_1593 (.A(_09444_));
 sg13g2_antennanp ANTENNA_1594 (.A(_09445_));
 sg13g2_antennanp ANTENNA_1595 (.A(_09445_));
 sg13g2_antennanp ANTENNA_1596 (.A(_09445_));
 sg13g2_antennanp ANTENNA_1597 (.A(_09445_));
 sg13g2_antennanp ANTENNA_1598 (.A(_09554_));
 sg13g2_antennanp ANTENNA_1599 (.A(_09554_));
 sg13g2_antennanp ANTENNA_1600 (.A(_09562_));
 sg13g2_antennanp ANTENNA_1601 (.A(_09587_));
 sg13g2_antennanp ANTENNA_1602 (.A(_09608_));
 sg13g2_antennanp ANTENNA_1603 (.A(_09665_));
 sg13g2_antennanp ANTENNA_1604 (.A(_09695_));
 sg13g2_antennanp ANTENNA_1605 (.A(_09721_));
 sg13g2_antennanp ANTENNA_1606 (.A(_09742_));
 sg13g2_antennanp ANTENNA_1607 (.A(_09765_));
 sg13g2_antennanp ANTENNA_1608 (.A(_09765_));
 sg13g2_antennanp ANTENNA_1609 (.A(_09794_));
 sg13g2_antennanp ANTENNA_1610 (.A(_09796_));
 sg13g2_antennanp ANTENNA_1611 (.A(_09912_));
 sg13g2_antennanp ANTENNA_1612 (.A(_10246_));
 sg13g2_antennanp ANTENNA_1613 (.A(_10246_));
 sg13g2_antennanp ANTENNA_1614 (.A(_10246_));
 sg13g2_antennanp ANTENNA_1615 (.A(_10302_));
 sg13g2_antennanp ANTENNA_1616 (.A(_10302_));
 sg13g2_antennanp ANTENNA_1617 (.A(_10302_));
 sg13g2_antennanp ANTENNA_1618 (.A(_10302_));
 sg13g2_antennanp ANTENNA_1619 (.A(_10302_));
 sg13g2_antennanp ANTENNA_1620 (.A(_10302_));
 sg13g2_antennanp ANTENNA_1621 (.A(_10302_));
 sg13g2_antennanp ANTENNA_1622 (.A(_10302_));
 sg13g2_antennanp ANTENNA_1623 (.A(_10307_));
 sg13g2_antennanp ANTENNA_1624 (.A(_10307_));
 sg13g2_antennanp ANTENNA_1625 (.A(_10307_));
 sg13g2_antennanp ANTENNA_1626 (.A(_10307_));
 sg13g2_antennanp ANTENNA_1627 (.A(_10307_));
 sg13g2_antennanp ANTENNA_1628 (.A(_10307_));
 sg13g2_antennanp ANTENNA_1629 (.A(_10307_));
 sg13g2_antennanp ANTENNA_1630 (.A(_10307_));
 sg13g2_antennanp ANTENNA_1631 (.A(_10312_));
 sg13g2_antennanp ANTENNA_1632 (.A(_10312_));
 sg13g2_antennanp ANTENNA_1633 (.A(_10312_));
 sg13g2_antennanp ANTENNA_1634 (.A(_10312_));
 sg13g2_antennanp ANTENNA_1635 (.A(_10312_));
 sg13g2_antennanp ANTENNA_1636 (.A(_10312_));
 sg13g2_antennanp ANTENNA_1637 (.A(_10312_));
 sg13g2_antennanp ANTENNA_1638 (.A(_10312_));
 sg13g2_antennanp ANTENNA_1639 (.A(_10326_));
 sg13g2_antennanp ANTENNA_1640 (.A(_10326_));
 sg13g2_antennanp ANTENNA_1641 (.A(_10326_));
 sg13g2_antennanp ANTENNA_1642 (.A(_10326_));
 sg13g2_antennanp ANTENNA_1643 (.A(_10326_));
 sg13g2_antennanp ANTENNA_1644 (.A(_10326_));
 sg13g2_antennanp ANTENNA_1645 (.A(_10326_));
 sg13g2_antennanp ANTENNA_1646 (.A(_10326_));
 sg13g2_antennanp ANTENNA_1647 (.A(_10339_));
 sg13g2_antennanp ANTENNA_1648 (.A(_10339_));
 sg13g2_antennanp ANTENNA_1649 (.A(_10339_));
 sg13g2_antennanp ANTENNA_1650 (.A(_10339_));
 sg13g2_antennanp ANTENNA_1651 (.A(_10339_));
 sg13g2_antennanp ANTENNA_1652 (.A(_10339_));
 sg13g2_antennanp ANTENNA_1653 (.A(_10339_));
 sg13g2_antennanp ANTENNA_1654 (.A(_10344_));
 sg13g2_antennanp ANTENNA_1655 (.A(_10344_));
 sg13g2_antennanp ANTENNA_1656 (.A(_10344_));
 sg13g2_antennanp ANTENNA_1657 (.A(_10344_));
 sg13g2_antennanp ANTENNA_1658 (.A(_10344_));
 sg13g2_antennanp ANTENNA_1659 (.A(_10344_));
 sg13g2_antennanp ANTENNA_1660 (.A(_10344_));
 sg13g2_antennanp ANTENNA_1661 (.A(_10344_));
 sg13g2_antennanp ANTENNA_1662 (.A(_10645_));
 sg13g2_antennanp ANTENNA_1663 (.A(_10645_));
 sg13g2_antennanp ANTENNA_1664 (.A(_11129_));
 sg13g2_antennanp ANTENNA_1665 (.A(_12058_));
 sg13g2_antennanp ANTENNA_1666 (.A(_12058_));
 sg13g2_antennanp ANTENNA_1667 (.A(_12058_));
 sg13g2_antennanp ANTENNA_1668 (.A(_12058_));
 sg13g2_antennanp ANTENNA_1669 (.A(_12058_));
 sg13g2_antennanp ANTENNA_1670 (.A(_12058_));
 sg13g2_antennanp ANTENNA_1671 (.A(_12058_));
 sg13g2_antennanp ANTENNA_1672 (.A(_12058_));
 sg13g2_antennanp ANTENNA_1673 (.A(_12058_));
 sg13g2_antennanp ANTENNA_1674 (.A(_12127_));
 sg13g2_antennanp ANTENNA_1675 (.A(_12127_));
 sg13g2_antennanp ANTENNA_1676 (.A(_12127_));
 sg13g2_antennanp ANTENNA_1677 (.A(_12127_));
 sg13g2_antennanp ANTENNA_1678 (.A(_12127_));
 sg13g2_antennanp ANTENNA_1679 (.A(_12127_));
 sg13g2_antennanp ANTENNA_1680 (.A(_12127_));
 sg13g2_antennanp ANTENNA_1681 (.A(_12127_));
 sg13g2_antennanp ANTENNA_1682 (.A(_12127_));
 sg13g2_antennanp ANTENNA_1683 (.A(_12152_));
 sg13g2_antennanp ANTENNA_1684 (.A(_12152_));
 sg13g2_antennanp ANTENNA_1685 (.A(_12152_));
 sg13g2_antennanp ANTENNA_1686 (.A(_12152_));
 sg13g2_antennanp ANTENNA_1687 (.A(_12152_));
 sg13g2_antennanp ANTENNA_1688 (.A(_12152_));
 sg13g2_antennanp ANTENNA_1689 (.A(_12152_));
 sg13g2_antennanp ANTENNA_1690 (.A(_12152_));
 sg13g2_antennanp ANTENNA_1691 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1692 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1693 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1694 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1695 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1696 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1697 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1698 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1699 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1700 (.A(_12223_));
 sg13g2_antennanp ANTENNA_1701 (.A(_12223_));
 sg13g2_antennanp ANTENNA_1702 (.A(_12223_));
 sg13g2_antennanp ANTENNA_1703 (.A(_12223_));
 sg13g2_antennanp ANTENNA_1704 (.A(_12223_));
 sg13g2_antennanp ANTENNA_1705 (.A(_12223_));
 sg13g2_antennanp ANTENNA_1706 (.A(_12223_));
 sg13g2_antennanp ANTENNA_1707 (.A(_12223_));
 sg13g2_antennanp ANTENNA_1708 (.A(_12223_));
 sg13g2_antennanp ANTENNA_1709 (.A(_12223_));
 sg13g2_antennanp ANTENNA_1710 (.A(_12223_));
 sg13g2_antennanp ANTENNA_1711 (.A(_12223_));
 sg13g2_antennanp ANTENNA_1712 (.A(_12223_));
 sg13g2_antennanp ANTENNA_1713 (.A(_12223_));
 sg13g2_antennanp ANTENNA_1714 (.A(_12223_));
 sg13g2_antennanp ANTENNA_1715 (.A(_12223_));
 sg13g2_antennanp ANTENNA_1716 (.A(_12223_));
 sg13g2_antennanp ANTENNA_1717 (.A(_12223_));
 sg13g2_antennanp ANTENNA_1718 (.A(_12229_));
 sg13g2_antennanp ANTENNA_1719 (.A(_12229_));
 sg13g2_antennanp ANTENNA_1720 (.A(_12229_));
 sg13g2_antennanp ANTENNA_1721 (.A(_12229_));
 sg13g2_antennanp ANTENNA_1722 (.A(_12229_));
 sg13g2_antennanp ANTENNA_1723 (.A(_12229_));
 sg13g2_antennanp ANTENNA_1724 (.A(_12229_));
 sg13g2_antennanp ANTENNA_1725 (.A(_12229_));
 sg13g2_antennanp ANTENNA_1726 (.A(_12229_));
 sg13g2_antennanp ANTENNA_1727 (.A(_12558_));
 sg13g2_antennanp ANTENNA_1728 (.A(_12558_));
 sg13g2_antennanp ANTENNA_1729 (.A(_12558_));
 sg13g2_antennanp ANTENNA_1730 (.A(_12558_));
 sg13g2_antennanp ANTENNA_1731 (.A(_12558_));
 sg13g2_antennanp ANTENNA_1732 (.A(_12726_));
 sg13g2_antennanp ANTENNA_1733 (.A(_12726_));
 sg13g2_antennanp ANTENNA_1734 (.A(_12726_));
 sg13g2_antennanp ANTENNA_1735 (.A(_12726_));
 sg13g2_antennanp ANTENNA_1736 (.A(clk));
 sg13g2_antennanp ANTENNA_1737 (.A(clk));
 sg13g2_antennanp ANTENNA_1738 (.A(\cpu.ex.pc[3] ));
 sg13g2_antennanp ANTENNA_1739 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_1740 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_1741 (.A(net12));
 sg13g2_antennanp ANTENNA_1742 (.A(net12));
 sg13g2_antennanp ANTENNA_1743 (.A(net12));
 sg13g2_antennanp ANTENNA_1744 (.A(net13));
 sg13g2_antennanp ANTENNA_1745 (.A(net13));
 sg13g2_antennanp ANTENNA_1746 (.A(net13));
 sg13g2_antennanp ANTENNA_1747 (.A(net437));
 sg13g2_antennanp ANTENNA_1748 (.A(net437));
 sg13g2_antennanp ANTENNA_1749 (.A(net437));
 sg13g2_antennanp ANTENNA_1750 (.A(net437));
 sg13g2_antennanp ANTENNA_1751 (.A(net437));
 sg13g2_antennanp ANTENNA_1752 (.A(net437));
 sg13g2_antennanp ANTENNA_1753 (.A(net437));
 sg13g2_antennanp ANTENNA_1754 (.A(net437));
 sg13g2_antennanp ANTENNA_1755 (.A(net437));
 sg13g2_antennanp ANTENNA_1756 (.A(net524));
 sg13g2_antennanp ANTENNA_1757 (.A(net524));
 sg13g2_antennanp ANTENNA_1758 (.A(net524));
 sg13g2_antennanp ANTENNA_1759 (.A(net524));
 sg13g2_antennanp ANTENNA_1760 (.A(net524));
 sg13g2_antennanp ANTENNA_1761 (.A(net524));
 sg13g2_antennanp ANTENNA_1762 (.A(net524));
 sg13g2_antennanp ANTENNA_1763 (.A(net524));
 sg13g2_antennanp ANTENNA_1764 (.A(net524));
 sg13g2_antennanp ANTENNA_1765 (.A(net524));
 sg13g2_antennanp ANTENNA_1766 (.A(net524));
 sg13g2_antennanp ANTENNA_1767 (.A(net524));
 sg13g2_antennanp ANTENNA_1768 (.A(net524));
 sg13g2_antennanp ANTENNA_1769 (.A(net542));
 sg13g2_antennanp ANTENNA_1770 (.A(net542));
 sg13g2_antennanp ANTENNA_1771 (.A(net542));
 sg13g2_antennanp ANTENNA_1772 (.A(net542));
 sg13g2_antennanp ANTENNA_1773 (.A(net542));
 sg13g2_antennanp ANTENNA_1774 (.A(net542));
 sg13g2_antennanp ANTENNA_1775 (.A(net542));
 sg13g2_antennanp ANTENNA_1776 (.A(net542));
 sg13g2_antennanp ANTENNA_1777 (.A(net542));
 sg13g2_antennanp ANTENNA_1778 (.A(net542));
 sg13g2_antennanp ANTENNA_1779 (.A(net542));
 sg13g2_antennanp ANTENNA_1780 (.A(net542));
 sg13g2_antennanp ANTENNA_1781 (.A(net542));
 sg13g2_antennanp ANTENNA_1782 (.A(net542));
 sg13g2_antennanp ANTENNA_1783 (.A(net542));
 sg13g2_antennanp ANTENNA_1784 (.A(net542));
 sg13g2_antennanp ANTENNA_1785 (.A(net542));
 sg13g2_antennanp ANTENNA_1786 (.A(net542));
 sg13g2_antennanp ANTENNA_1787 (.A(net656));
 sg13g2_antennanp ANTENNA_1788 (.A(net656));
 sg13g2_antennanp ANTENNA_1789 (.A(net656));
 sg13g2_antennanp ANTENNA_1790 (.A(net656));
 sg13g2_antennanp ANTENNA_1791 (.A(net656));
 sg13g2_antennanp ANTENNA_1792 (.A(net656));
 sg13g2_antennanp ANTENNA_1793 (.A(net656));
 sg13g2_antennanp ANTENNA_1794 (.A(net656));
 sg13g2_antennanp ANTENNA_1795 (.A(net656));
 sg13g2_antennanp ANTENNA_1796 (.A(net685));
 sg13g2_antennanp ANTENNA_1797 (.A(net685));
 sg13g2_antennanp ANTENNA_1798 (.A(net685));
 sg13g2_antennanp ANTENNA_1799 (.A(net685));
 sg13g2_antennanp ANTENNA_1800 (.A(net685));
 sg13g2_antennanp ANTENNA_1801 (.A(net685));
 sg13g2_antennanp ANTENNA_1802 (.A(net685));
 sg13g2_antennanp ANTENNA_1803 (.A(net685));
 sg13g2_antennanp ANTENNA_1804 (.A(net685));
 sg13g2_antennanp ANTENNA_1805 (.A(net707));
 sg13g2_antennanp ANTENNA_1806 (.A(net707));
 sg13g2_antennanp ANTENNA_1807 (.A(net707));
 sg13g2_antennanp ANTENNA_1808 (.A(net707));
 sg13g2_antennanp ANTENNA_1809 (.A(net707));
 sg13g2_antennanp ANTENNA_1810 (.A(net707));
 sg13g2_antennanp ANTENNA_1811 (.A(net707));
 sg13g2_antennanp ANTENNA_1812 (.A(net707));
 sg13g2_antennanp ANTENNA_1813 (.A(net707));
 sg13g2_antennanp ANTENNA_1814 (.A(net803));
 sg13g2_antennanp ANTENNA_1815 (.A(net803));
 sg13g2_antennanp ANTENNA_1816 (.A(net803));
 sg13g2_antennanp ANTENNA_1817 (.A(net803));
 sg13g2_antennanp ANTENNA_1818 (.A(net803));
 sg13g2_antennanp ANTENNA_1819 (.A(net803));
 sg13g2_antennanp ANTENNA_1820 (.A(net803));
 sg13g2_antennanp ANTENNA_1821 (.A(net803));
 sg13g2_antennanp ANTENNA_1822 (.A(net888));
 sg13g2_antennanp ANTENNA_1823 (.A(net888));
 sg13g2_antennanp ANTENNA_1824 (.A(net888));
 sg13g2_antennanp ANTENNA_1825 (.A(net888));
 sg13g2_antennanp ANTENNA_1826 (.A(net888));
 sg13g2_antennanp ANTENNA_1827 (.A(net888));
 sg13g2_antennanp ANTENNA_1828 (.A(net888));
 sg13g2_antennanp ANTENNA_1829 (.A(net888));
 sg13g2_antennanp ANTENNA_1830 (.A(net888));
 sg13g2_antennanp ANTENNA_1831 (.A(net928));
 sg13g2_antennanp ANTENNA_1832 (.A(net928));
 sg13g2_antennanp ANTENNA_1833 (.A(net928));
 sg13g2_antennanp ANTENNA_1834 (.A(net928));
 sg13g2_antennanp ANTENNA_1835 (.A(net928));
 sg13g2_antennanp ANTENNA_1836 (.A(net928));
 sg13g2_antennanp ANTENNA_1837 (.A(net928));
 sg13g2_antennanp ANTENNA_1838 (.A(net928));
 sg13g2_antennanp ANTENNA_1839 (.A(net928));
 sg13g2_antennanp ANTENNA_1840 (.A(net984));
 sg13g2_antennanp ANTENNA_1841 (.A(net984));
 sg13g2_antennanp ANTENNA_1842 (.A(net984));
 sg13g2_antennanp ANTENNA_1843 (.A(net984));
 sg13g2_antennanp ANTENNA_1844 (.A(net984));
 sg13g2_antennanp ANTENNA_1845 (.A(net984));
 sg13g2_antennanp ANTENNA_1846 (.A(net984));
 sg13g2_antennanp ANTENNA_1847 (.A(net984));
 sg13g2_antennanp ANTENNA_1848 (.A(net984));
 sg13g2_antennanp ANTENNA_1849 (.A(net984));
 sg13g2_antennanp ANTENNA_1850 (.A(net984));
 sg13g2_antennanp ANTENNA_1851 (.A(net984));
 sg13g2_antennanp ANTENNA_1852 (.A(net984));
 sg13g2_antennanp ANTENNA_1853 (.A(net984));
 sg13g2_antennanp ANTENNA_1854 (.A(net984));
 sg13g2_antennanp ANTENNA_1855 (.A(net984));
 sg13g2_antennanp ANTENNA_1856 (.A(net984));
 sg13g2_antennanp ANTENNA_1857 (.A(net984));
 sg13g2_antennanp ANTENNA_1858 (.A(net984));
 sg13g2_antennanp ANTENNA_1859 (.A(net984));
 sg13g2_antennanp ANTENNA_1860 (.A(net984));
 sg13g2_antennanp ANTENNA_1861 (.A(net984));
 sg13g2_antennanp ANTENNA_1862 (.A(net984));
 sg13g2_antennanp ANTENNA_1863 (.A(net984));
 sg13g2_antennanp ANTENNA_1864 (.A(net984));
 sg13g2_antennanp ANTENNA_1865 (.A(net984));
 sg13g2_antennanp ANTENNA_1866 (.A(net984));
 sg13g2_antennanp ANTENNA_1867 (.A(net984));
 sg13g2_antennanp ANTENNA_1868 (.A(net984));
 sg13g2_antennanp ANTENNA_1869 (.A(net984));
 sg13g2_antennanp ANTENNA_1870 (.A(net984));
 sg13g2_antennanp ANTENNA_1871 (.A(net984));
 sg13g2_antennanp ANTENNA_1872 (.A(net984));
 sg13g2_antennanp ANTENNA_1873 (.A(net984));
 sg13g2_antennanp ANTENNA_1874 (.A(net1004));
 sg13g2_antennanp ANTENNA_1875 (.A(net1004));
 sg13g2_antennanp ANTENNA_1876 (.A(net1004));
 sg13g2_antennanp ANTENNA_1877 (.A(net1004));
 sg13g2_antennanp ANTENNA_1878 (.A(net1004));
 sg13g2_antennanp ANTENNA_1879 (.A(net1004));
 sg13g2_antennanp ANTENNA_1880 (.A(net1004));
 sg13g2_antennanp ANTENNA_1881 (.A(net1004));
 sg13g2_antennanp ANTENNA_1882 (.A(net1004));
 sg13g2_antennanp ANTENNA_1883 (.A(net1004));
 sg13g2_antennanp ANTENNA_1884 (.A(net1004));
 sg13g2_antennanp ANTENNA_1885 (.A(net1004));
 sg13g2_antennanp ANTENNA_1886 (.A(net1004));
 sg13g2_antennanp ANTENNA_1887 (.A(net1004));
 sg13g2_antennanp ANTENNA_1888 (.A(net1004));
 sg13g2_antennanp ANTENNA_1889 (.A(net1004));
 sg13g2_antennanp ANTENNA_1890 (.A(net1004));
 sg13g2_antennanp ANTENNA_1891 (.A(net1004));
 sg13g2_antennanp ANTENNA_1892 (.A(net1004));
 sg13g2_antennanp ANTENNA_1893 (.A(net1004));
 sg13g2_antennanp ANTENNA_1894 (.A(net1004));
 sg13g2_antennanp ANTENNA_1895 (.A(net1004));
 sg13g2_antennanp ANTENNA_1896 (.A(net1004));
 sg13g2_antennanp ANTENNA_1897 (.A(net1004));
 sg13g2_antennanp ANTENNA_1898 (.A(net1004));
 sg13g2_antennanp ANTENNA_1899 (.A(net1004));
 sg13g2_antennanp ANTENNA_1900 (.A(net1004));
 sg13g2_antennanp ANTENNA_1901 (.A(net1004));
 sg13g2_antennanp ANTENNA_1902 (.A(net1004));
 sg13g2_antennanp ANTENNA_1903 (.A(net1004));
 sg13g2_antennanp ANTENNA_1904 (.A(net1004));
 sg13g2_antennanp ANTENNA_1905 (.A(net1004));
 sg13g2_antennanp ANTENNA_1906 (.A(net1004));
 sg13g2_antennanp ANTENNA_1907 (.A(net1075));
 sg13g2_antennanp ANTENNA_1908 (.A(net1075));
 sg13g2_antennanp ANTENNA_1909 (.A(net1075));
 sg13g2_antennanp ANTENNA_1910 (.A(net1075));
 sg13g2_antennanp ANTENNA_1911 (.A(net1075));
 sg13g2_antennanp ANTENNA_1912 (.A(net1075));
 sg13g2_antennanp ANTENNA_1913 (.A(net1075));
 sg13g2_antennanp ANTENNA_1914 (.A(net1075));
 sg13g2_antennanp ANTENNA_1915 (.A(net1075));
 sg13g2_antennanp ANTENNA_1916 (.A(_00190_));
 sg13g2_antennanp ANTENNA_1917 (.A(_00197_));
 sg13g2_antennanp ANTENNA_1918 (.A(_00197_));
 sg13g2_antennanp ANTENNA_1919 (.A(_00197_));
 sg13g2_antennanp ANTENNA_1920 (.A(_00197_));
 sg13g2_antennanp ANTENNA_1921 (.A(_00228_));
 sg13g2_antennanp ANTENNA_1922 (.A(_00228_));
 sg13g2_antennanp ANTENNA_1923 (.A(_00235_));
 sg13g2_antennanp ANTENNA_1924 (.A(_00235_));
 sg13g2_antennanp ANTENNA_1925 (.A(_00930_));
 sg13g2_antennanp ANTENNA_1926 (.A(_01052_));
 sg13g2_antennanp ANTENNA_1927 (.A(_01052_));
 sg13g2_antennanp ANTENNA_1928 (.A(_02950_));
 sg13g2_antennanp ANTENNA_1929 (.A(_02950_));
 sg13g2_antennanp ANTENNA_1930 (.A(_02950_));
 sg13g2_antennanp ANTENNA_1931 (.A(_02950_));
 sg13g2_antennanp ANTENNA_1932 (.A(_02950_));
 sg13g2_antennanp ANTENNA_1933 (.A(_02950_));
 sg13g2_antennanp ANTENNA_1934 (.A(_02950_));
 sg13g2_antennanp ANTENNA_1935 (.A(_02950_));
 sg13g2_antennanp ANTENNA_1936 (.A(_02950_));
 sg13g2_antennanp ANTENNA_1937 (.A(_02950_));
 sg13g2_antennanp ANTENNA_1938 (.A(_02965_));
 sg13g2_antennanp ANTENNA_1939 (.A(_02965_));
 sg13g2_antennanp ANTENNA_1940 (.A(_02965_));
 sg13g2_antennanp ANTENNA_1941 (.A(_02965_));
 sg13g2_antennanp ANTENNA_1942 (.A(_02965_));
 sg13g2_antennanp ANTENNA_1943 (.A(_02965_));
 sg13g2_antennanp ANTENNA_1944 (.A(_02965_));
 sg13g2_antennanp ANTENNA_1945 (.A(_02965_));
 sg13g2_antennanp ANTENNA_1946 (.A(_02965_));
 sg13g2_antennanp ANTENNA_1947 (.A(_02965_));
 sg13g2_antennanp ANTENNA_1948 (.A(_03429_));
 sg13g2_antennanp ANTENNA_1949 (.A(_03429_));
 sg13g2_antennanp ANTENNA_1950 (.A(_03429_));
 sg13g2_antennanp ANTENNA_1951 (.A(_03429_));
 sg13g2_antennanp ANTENNA_1952 (.A(_03435_));
 sg13g2_antennanp ANTENNA_1953 (.A(_03435_));
 sg13g2_antennanp ANTENNA_1954 (.A(_03435_));
 sg13g2_antennanp ANTENNA_1955 (.A(_03435_));
 sg13g2_antennanp ANTENNA_1956 (.A(_03435_));
 sg13g2_antennanp ANTENNA_1957 (.A(_03435_));
 sg13g2_antennanp ANTENNA_1958 (.A(_03435_));
 sg13g2_antennanp ANTENNA_1959 (.A(_03435_));
 sg13g2_antennanp ANTENNA_1960 (.A(_03435_));
 sg13g2_antennanp ANTENNA_1961 (.A(_04742_));
 sg13g2_antennanp ANTENNA_1962 (.A(_04742_));
 sg13g2_antennanp ANTENNA_1963 (.A(_04742_));
 sg13g2_antennanp ANTENNA_1964 (.A(_04742_));
 sg13g2_antennanp ANTENNA_1965 (.A(_04887_));
 sg13g2_antennanp ANTENNA_1966 (.A(_04887_));
 sg13g2_antennanp ANTENNA_1967 (.A(_04887_));
 sg13g2_antennanp ANTENNA_1968 (.A(_04887_));
 sg13g2_antennanp ANTENNA_1969 (.A(_04894_));
 sg13g2_antennanp ANTENNA_1970 (.A(_05013_));
 sg13g2_antennanp ANTENNA_1971 (.A(_05015_));
 sg13g2_antennanp ANTENNA_1972 (.A(_05168_));
 sg13g2_antennanp ANTENNA_1973 (.A(_05169_));
 sg13g2_antennanp ANTENNA_1974 (.A(_05245_));
 sg13g2_antennanp ANTENNA_1975 (.A(_05278_));
 sg13g2_antennanp ANTENNA_1976 (.A(_05280_));
 sg13g2_antennanp ANTENNA_1977 (.A(_05372_));
 sg13g2_antennanp ANTENNA_1978 (.A(_05432_));
 sg13g2_antennanp ANTENNA_1979 (.A(_05508_));
 sg13g2_antennanp ANTENNA_1980 (.A(_05646_));
 sg13g2_antennanp ANTENNA_1981 (.A(_05650_));
 sg13g2_antennanp ANTENNA_1982 (.A(_05654_));
 sg13g2_antennanp ANTENNA_1983 (.A(_05763_));
 sg13g2_antennanp ANTENNA_1984 (.A(_05763_));
 sg13g2_antennanp ANTENNA_1985 (.A(_05763_));
 sg13g2_antennanp ANTENNA_1986 (.A(_05763_));
 sg13g2_antennanp ANTENNA_1987 (.A(_05763_));
 sg13g2_antennanp ANTENNA_1988 (.A(_05763_));
 sg13g2_antennanp ANTENNA_1989 (.A(_05763_));
 sg13g2_antennanp ANTENNA_1990 (.A(_05766_));
 sg13g2_antennanp ANTENNA_1991 (.A(_05766_));
 sg13g2_antennanp ANTENNA_1992 (.A(_05766_));
 sg13g2_antennanp ANTENNA_1993 (.A(_05766_));
 sg13g2_antennanp ANTENNA_1994 (.A(_05770_));
 sg13g2_antennanp ANTENNA_1995 (.A(_05770_));
 sg13g2_antennanp ANTENNA_1996 (.A(_05770_));
 sg13g2_antennanp ANTENNA_1997 (.A(_05770_));
 sg13g2_antennanp ANTENNA_1998 (.A(_05770_));
 sg13g2_antennanp ANTENNA_1999 (.A(_05770_));
 sg13g2_antennanp ANTENNA_2000 (.A(_05770_));
 sg13g2_antennanp ANTENNA_2001 (.A(_05770_));
 sg13g2_antennanp ANTENNA_2002 (.A(_05775_));
 sg13g2_antennanp ANTENNA_2003 (.A(_05775_));
 sg13g2_antennanp ANTENNA_2004 (.A(_05775_));
 sg13g2_antennanp ANTENNA_2005 (.A(_05785_));
 sg13g2_antennanp ANTENNA_2006 (.A(_05785_));
 sg13g2_antennanp ANTENNA_2007 (.A(_05785_));
 sg13g2_antennanp ANTENNA_2008 (.A(_05785_));
 sg13g2_antennanp ANTENNA_2009 (.A(_05835_));
 sg13g2_antennanp ANTENNA_2010 (.A(_05835_));
 sg13g2_antennanp ANTENNA_2011 (.A(_05835_));
 sg13g2_antennanp ANTENNA_2012 (.A(_05835_));
 sg13g2_antennanp ANTENNA_2013 (.A(_06843_));
 sg13g2_antennanp ANTENNA_2014 (.A(_06843_));
 sg13g2_antennanp ANTENNA_2015 (.A(_06843_));
 sg13g2_antennanp ANTENNA_2016 (.A(_07398_));
 sg13g2_antennanp ANTENNA_2017 (.A(_07434_));
 sg13g2_antennanp ANTENNA_2018 (.A(_08297_));
 sg13g2_antennanp ANTENNA_2019 (.A(_08297_));
 sg13g2_antennanp ANTENNA_2020 (.A(_08502_));
 sg13g2_antennanp ANTENNA_2021 (.A(_08502_));
 sg13g2_antennanp ANTENNA_2022 (.A(_08502_));
 sg13g2_antennanp ANTENNA_2023 (.A(_08502_));
 sg13g2_antennanp ANTENNA_2024 (.A(_08502_));
 sg13g2_antennanp ANTENNA_2025 (.A(_08502_));
 sg13g2_antennanp ANTENNA_2026 (.A(_08502_));
 sg13g2_antennanp ANTENNA_2027 (.A(_08533_));
 sg13g2_antennanp ANTENNA_2028 (.A(_08533_));
 sg13g2_antennanp ANTENNA_2029 (.A(_08533_));
 sg13g2_antennanp ANTENNA_2030 (.A(_08533_));
 sg13g2_antennanp ANTENNA_2031 (.A(_08533_));
 sg13g2_antennanp ANTENNA_2032 (.A(_08533_));
 sg13g2_antennanp ANTENNA_2033 (.A(_08558_));
 sg13g2_antennanp ANTENNA_2034 (.A(_08558_));
 sg13g2_antennanp ANTENNA_2035 (.A(_08558_));
 sg13g2_antennanp ANTENNA_2036 (.A(_08558_));
 sg13g2_antennanp ANTENNA_2037 (.A(_08634_));
 sg13g2_antennanp ANTENNA_2038 (.A(_08634_));
 sg13g2_antennanp ANTENNA_2039 (.A(_08634_));
 sg13g2_antennanp ANTENNA_2040 (.A(_08634_));
 sg13g2_antennanp ANTENNA_2041 (.A(_08634_));
 sg13g2_antennanp ANTENNA_2042 (.A(_08634_));
 sg13g2_antennanp ANTENNA_2043 (.A(_08634_));
 sg13g2_antennanp ANTENNA_2044 (.A(_08634_));
 sg13g2_antennanp ANTENNA_2045 (.A(_08634_));
 sg13g2_antennanp ANTENNA_2046 (.A(_08679_));
 sg13g2_antennanp ANTENNA_2047 (.A(_08679_));
 sg13g2_antennanp ANTENNA_2048 (.A(_08679_));
 sg13g2_antennanp ANTENNA_2049 (.A(_08728_));
 sg13g2_antennanp ANTENNA_2050 (.A(_08728_));
 sg13g2_antennanp ANTENNA_2051 (.A(_08728_));
 sg13g2_antennanp ANTENNA_2052 (.A(_08853_));
 sg13g2_antennanp ANTENNA_2053 (.A(_08918_));
 sg13g2_antennanp ANTENNA_2054 (.A(_08918_));
 sg13g2_antennanp ANTENNA_2055 (.A(_08918_));
 sg13g2_antennanp ANTENNA_2056 (.A(_08918_));
 sg13g2_antennanp ANTENNA_2057 (.A(_08918_));
 sg13g2_antennanp ANTENNA_2058 (.A(_08918_));
 sg13g2_antennanp ANTENNA_2059 (.A(_08918_));
 sg13g2_antennanp ANTENNA_2060 (.A(_08918_));
 sg13g2_antennanp ANTENNA_2061 (.A(_08918_));
 sg13g2_antennanp ANTENNA_2062 (.A(_08918_));
 sg13g2_antennanp ANTENNA_2063 (.A(_08938_));
 sg13g2_antennanp ANTENNA_2064 (.A(_08959_));
 sg13g2_antennanp ANTENNA_2065 (.A(_08970_));
 sg13g2_antennanp ANTENNA_2066 (.A(_08970_));
 sg13g2_antennanp ANTENNA_2067 (.A(_08970_));
 sg13g2_antennanp ANTENNA_2068 (.A(_08970_));
 sg13g2_antennanp ANTENNA_2069 (.A(_09167_));
 sg13g2_antennanp ANTENNA_2070 (.A(_09336_));
 sg13g2_antennanp ANTENNA_2071 (.A(_09336_));
 sg13g2_antennanp ANTENNA_2072 (.A(_09349_));
 sg13g2_antennanp ANTENNA_2073 (.A(_09349_));
 sg13g2_antennanp ANTENNA_2074 (.A(_09349_));
 sg13g2_antennanp ANTENNA_2075 (.A(_09349_));
 sg13g2_antennanp ANTENNA_2076 (.A(_09349_));
 sg13g2_antennanp ANTENNA_2077 (.A(_09349_));
 sg13g2_antennanp ANTENNA_2078 (.A(_09380_));
 sg13g2_antennanp ANTENNA_2079 (.A(_09380_));
 sg13g2_antennanp ANTENNA_2080 (.A(_09380_));
 sg13g2_antennanp ANTENNA_2081 (.A(_09380_));
 sg13g2_antennanp ANTENNA_2082 (.A(_09385_));
 sg13g2_antennanp ANTENNA_2083 (.A(_09385_));
 sg13g2_antennanp ANTENNA_2084 (.A(_09385_));
 sg13g2_antennanp ANTENNA_2085 (.A(_09385_));
 sg13g2_antennanp ANTENNA_2086 (.A(_09385_));
 sg13g2_antennanp ANTENNA_2087 (.A(_09385_));
 sg13g2_antennanp ANTENNA_2088 (.A(_09385_));
 sg13g2_antennanp ANTENNA_2089 (.A(_09385_));
 sg13g2_antennanp ANTENNA_2090 (.A(_09385_));
 sg13g2_antennanp ANTENNA_2091 (.A(_09386_));
 sg13g2_antennanp ANTENNA_2092 (.A(_09386_));
 sg13g2_antennanp ANTENNA_2093 (.A(_09386_));
 sg13g2_antennanp ANTENNA_2094 (.A(_09386_));
 sg13g2_antennanp ANTENNA_2095 (.A(_09386_));
 sg13g2_antennanp ANTENNA_2096 (.A(_09386_));
 sg13g2_antennanp ANTENNA_2097 (.A(_09386_));
 sg13g2_antennanp ANTENNA_2098 (.A(_09386_));
 sg13g2_antennanp ANTENNA_2099 (.A(_09388_));
 sg13g2_antennanp ANTENNA_2100 (.A(_09388_));
 sg13g2_antennanp ANTENNA_2101 (.A(_09388_));
 sg13g2_antennanp ANTENNA_2102 (.A(_09388_));
 sg13g2_antennanp ANTENNA_2103 (.A(_09389_));
 sg13g2_antennanp ANTENNA_2104 (.A(_09389_));
 sg13g2_antennanp ANTENNA_2105 (.A(_09389_));
 sg13g2_antennanp ANTENNA_2106 (.A(_09389_));
 sg13g2_antennanp ANTENNA_2107 (.A(_09389_));
 sg13g2_antennanp ANTENNA_2108 (.A(_09389_));
 sg13g2_antennanp ANTENNA_2109 (.A(_09389_));
 sg13g2_antennanp ANTENNA_2110 (.A(_09390_));
 sg13g2_antennanp ANTENNA_2111 (.A(_09390_));
 sg13g2_antennanp ANTENNA_2112 (.A(_09390_));
 sg13g2_antennanp ANTENNA_2113 (.A(_09444_));
 sg13g2_antennanp ANTENNA_2114 (.A(_09444_));
 sg13g2_antennanp ANTENNA_2115 (.A(_09444_));
 sg13g2_antennanp ANTENNA_2116 (.A(_09444_));
 sg13g2_antennanp ANTENNA_2117 (.A(_09444_));
 sg13g2_antennanp ANTENNA_2118 (.A(_09444_));
 sg13g2_antennanp ANTENNA_2119 (.A(_09445_));
 sg13g2_antennanp ANTENNA_2120 (.A(_09445_));
 sg13g2_antennanp ANTENNA_2121 (.A(_09445_));
 sg13g2_antennanp ANTENNA_2122 (.A(_09445_));
 sg13g2_antennanp ANTENNA_2123 (.A(_09554_));
 sg13g2_antennanp ANTENNA_2124 (.A(_09554_));
 sg13g2_antennanp ANTENNA_2125 (.A(_09587_));
 sg13g2_antennanp ANTENNA_2126 (.A(_09608_));
 sg13g2_antennanp ANTENNA_2127 (.A(_09665_));
 sg13g2_antennanp ANTENNA_2128 (.A(_09695_));
 sg13g2_antennanp ANTENNA_2129 (.A(_09721_));
 sg13g2_antennanp ANTENNA_2130 (.A(_09742_));
 sg13g2_antennanp ANTENNA_2131 (.A(_09765_));
 sg13g2_antennanp ANTENNA_2132 (.A(_09765_));
 sg13g2_antennanp ANTENNA_2133 (.A(_09794_));
 sg13g2_antennanp ANTENNA_2134 (.A(_09796_));
 sg13g2_antennanp ANTENNA_2135 (.A(_09912_));
 sg13g2_antennanp ANTENNA_2136 (.A(_09990_));
 sg13g2_antennanp ANTENNA_2137 (.A(_09990_));
 sg13g2_antennanp ANTENNA_2138 (.A(_09990_));
 sg13g2_antennanp ANTENNA_2139 (.A(_09990_));
 sg13g2_antennanp ANTENNA_2140 (.A(_09990_));
 sg13g2_antennanp ANTENNA_2141 (.A(_09990_));
 sg13g2_antennanp ANTENNA_2142 (.A(_09990_));
 sg13g2_antennanp ANTENNA_2143 (.A(_09990_));
 sg13g2_antennanp ANTENNA_2144 (.A(_09990_));
 sg13g2_antennanp ANTENNA_2145 (.A(_09990_));
 sg13g2_antennanp ANTENNA_2146 (.A(_10302_));
 sg13g2_antennanp ANTENNA_2147 (.A(_10302_));
 sg13g2_antennanp ANTENNA_2148 (.A(_10302_));
 sg13g2_antennanp ANTENNA_2149 (.A(_10302_));
 sg13g2_antennanp ANTENNA_2150 (.A(_10302_));
 sg13g2_antennanp ANTENNA_2151 (.A(_10302_));
 sg13g2_antennanp ANTENNA_2152 (.A(_10302_));
 sg13g2_antennanp ANTENNA_2153 (.A(_10302_));
 sg13g2_antennanp ANTENNA_2154 (.A(_10307_));
 sg13g2_antennanp ANTENNA_2155 (.A(_10307_));
 sg13g2_antennanp ANTENNA_2156 (.A(_10307_));
 sg13g2_antennanp ANTENNA_2157 (.A(_10307_));
 sg13g2_antennanp ANTENNA_2158 (.A(_10307_));
 sg13g2_antennanp ANTENNA_2159 (.A(_10307_));
 sg13g2_antennanp ANTENNA_2160 (.A(_10307_));
 sg13g2_antennanp ANTENNA_2161 (.A(_10307_));
 sg13g2_antennanp ANTENNA_2162 (.A(_10312_));
 sg13g2_antennanp ANTENNA_2163 (.A(_10312_));
 sg13g2_antennanp ANTENNA_2164 (.A(_10312_));
 sg13g2_antennanp ANTENNA_2165 (.A(_10312_));
 sg13g2_antennanp ANTENNA_2166 (.A(_10312_));
 sg13g2_antennanp ANTENNA_2167 (.A(_10312_));
 sg13g2_antennanp ANTENNA_2168 (.A(_10312_));
 sg13g2_antennanp ANTENNA_2169 (.A(_10312_));
 sg13g2_antennanp ANTENNA_2170 (.A(_10326_));
 sg13g2_antennanp ANTENNA_2171 (.A(_10326_));
 sg13g2_antennanp ANTENNA_2172 (.A(_10326_));
 sg13g2_antennanp ANTENNA_2173 (.A(_10326_));
 sg13g2_antennanp ANTENNA_2174 (.A(_10326_));
 sg13g2_antennanp ANTENNA_2175 (.A(_10326_));
 sg13g2_antennanp ANTENNA_2176 (.A(_10326_));
 sg13g2_antennanp ANTENNA_2177 (.A(_10326_));
 sg13g2_antennanp ANTENNA_2178 (.A(_10339_));
 sg13g2_antennanp ANTENNA_2179 (.A(_10339_));
 sg13g2_antennanp ANTENNA_2180 (.A(_10339_));
 sg13g2_antennanp ANTENNA_2181 (.A(_10339_));
 sg13g2_antennanp ANTENNA_2182 (.A(_10339_));
 sg13g2_antennanp ANTENNA_2183 (.A(_10339_));
 sg13g2_antennanp ANTENNA_2184 (.A(_10339_));
 sg13g2_antennanp ANTENNA_2185 (.A(_10344_));
 sg13g2_antennanp ANTENNA_2186 (.A(_10344_));
 sg13g2_antennanp ANTENNA_2187 (.A(_10344_));
 sg13g2_antennanp ANTENNA_2188 (.A(_10344_));
 sg13g2_antennanp ANTENNA_2189 (.A(_10344_));
 sg13g2_antennanp ANTENNA_2190 (.A(_10344_));
 sg13g2_antennanp ANTENNA_2191 (.A(_10344_));
 sg13g2_antennanp ANTENNA_2192 (.A(_10344_));
 sg13g2_antennanp ANTENNA_2193 (.A(_10645_));
 sg13g2_antennanp ANTENNA_2194 (.A(_10645_));
 sg13g2_antennanp ANTENNA_2195 (.A(_11129_));
 sg13g2_antennanp ANTENNA_2196 (.A(_12058_));
 sg13g2_antennanp ANTENNA_2197 (.A(_12058_));
 sg13g2_antennanp ANTENNA_2198 (.A(_12058_));
 sg13g2_antennanp ANTENNA_2199 (.A(_12058_));
 sg13g2_antennanp ANTENNA_2200 (.A(_12058_));
 sg13g2_antennanp ANTENNA_2201 (.A(_12058_));
 sg13g2_antennanp ANTENNA_2202 (.A(_12058_));
 sg13g2_antennanp ANTENNA_2203 (.A(_12058_));
 sg13g2_antennanp ANTENNA_2204 (.A(_12058_));
 sg13g2_antennanp ANTENNA_2205 (.A(_12127_));
 sg13g2_antennanp ANTENNA_2206 (.A(_12127_));
 sg13g2_antennanp ANTENNA_2207 (.A(_12127_));
 sg13g2_antennanp ANTENNA_2208 (.A(_12127_));
 sg13g2_antennanp ANTENNA_2209 (.A(_12127_));
 sg13g2_antennanp ANTENNA_2210 (.A(_12127_));
 sg13g2_antennanp ANTENNA_2211 (.A(_12127_));
 sg13g2_antennanp ANTENNA_2212 (.A(_12127_));
 sg13g2_antennanp ANTENNA_2213 (.A(_12127_));
 sg13g2_antennanp ANTENNA_2214 (.A(_12152_));
 sg13g2_antennanp ANTENNA_2215 (.A(_12152_));
 sg13g2_antennanp ANTENNA_2216 (.A(_12152_));
 sg13g2_antennanp ANTENNA_2217 (.A(_12152_));
 sg13g2_antennanp ANTENNA_2218 (.A(_12152_));
 sg13g2_antennanp ANTENNA_2219 (.A(_12152_));
 sg13g2_antennanp ANTENNA_2220 (.A(_12152_));
 sg13g2_antennanp ANTENNA_2221 (.A(_12152_));
 sg13g2_antennanp ANTENNA_2222 (.A(_12218_));
 sg13g2_antennanp ANTENNA_2223 (.A(_12218_));
 sg13g2_antennanp ANTENNA_2224 (.A(_12218_));
 sg13g2_antennanp ANTENNA_2225 (.A(_12218_));
 sg13g2_antennanp ANTENNA_2226 (.A(_12218_));
 sg13g2_antennanp ANTENNA_2227 (.A(_12218_));
 sg13g2_antennanp ANTENNA_2228 (.A(_12218_));
 sg13g2_antennanp ANTENNA_2229 (.A(_12218_));
 sg13g2_antennanp ANTENNA_2230 (.A(_12218_));
 sg13g2_antennanp ANTENNA_2231 (.A(_12223_));
 sg13g2_antennanp ANTENNA_2232 (.A(_12223_));
 sg13g2_antennanp ANTENNA_2233 (.A(_12223_));
 sg13g2_antennanp ANTENNA_2234 (.A(_12223_));
 sg13g2_antennanp ANTENNA_2235 (.A(_12223_));
 sg13g2_antennanp ANTENNA_2236 (.A(_12223_));
 sg13g2_antennanp ANTENNA_2237 (.A(_12223_));
 sg13g2_antennanp ANTENNA_2238 (.A(_12223_));
 sg13g2_antennanp ANTENNA_2239 (.A(_12223_));
 sg13g2_antennanp ANTENNA_2240 (.A(_12229_));
 sg13g2_antennanp ANTENNA_2241 (.A(_12229_));
 sg13g2_antennanp ANTENNA_2242 (.A(_12229_));
 sg13g2_antennanp ANTENNA_2243 (.A(_12229_));
 sg13g2_antennanp ANTENNA_2244 (.A(_12229_));
 sg13g2_antennanp ANTENNA_2245 (.A(_12229_));
 sg13g2_antennanp ANTENNA_2246 (.A(_12229_));
 sg13g2_antennanp ANTENNA_2247 (.A(_12229_));
 sg13g2_antennanp ANTENNA_2248 (.A(_12229_));
 sg13g2_antennanp ANTENNA_2249 (.A(_12558_));
 sg13g2_antennanp ANTENNA_2250 (.A(_12558_));
 sg13g2_antennanp ANTENNA_2251 (.A(_12558_));
 sg13g2_antennanp ANTENNA_2252 (.A(_12558_));
 sg13g2_antennanp ANTENNA_2253 (.A(_12558_));
 sg13g2_antennanp ANTENNA_2254 (.A(_12558_));
 sg13g2_antennanp ANTENNA_2255 (.A(_12558_));
 sg13g2_antennanp ANTENNA_2256 (.A(_12726_));
 sg13g2_antennanp ANTENNA_2257 (.A(_12726_));
 sg13g2_antennanp ANTENNA_2258 (.A(_12726_));
 sg13g2_antennanp ANTENNA_2259 (.A(_12726_));
 sg13g2_antennanp ANTENNA_2260 (.A(clk));
 sg13g2_antennanp ANTENNA_2261 (.A(clk));
 sg13g2_antennanp ANTENNA_2262 (.A(\cpu.ex.pc[3] ));
 sg13g2_antennanp ANTENNA_2263 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_2264 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_2265 (.A(net12));
 sg13g2_antennanp ANTENNA_2266 (.A(net12));
 sg13g2_antennanp ANTENNA_2267 (.A(net12));
 sg13g2_antennanp ANTENNA_2268 (.A(net13));
 sg13g2_antennanp ANTENNA_2269 (.A(net13));
 sg13g2_antennanp ANTENNA_2270 (.A(net13));
 sg13g2_antennanp ANTENNA_2271 (.A(net437));
 sg13g2_antennanp ANTENNA_2272 (.A(net437));
 sg13g2_antennanp ANTENNA_2273 (.A(net437));
 sg13g2_antennanp ANTENNA_2274 (.A(net437));
 sg13g2_antennanp ANTENNA_2275 (.A(net437));
 sg13g2_antennanp ANTENNA_2276 (.A(net437));
 sg13g2_antennanp ANTENNA_2277 (.A(net437));
 sg13g2_antennanp ANTENNA_2278 (.A(net437));
 sg13g2_antennanp ANTENNA_2279 (.A(net437));
 sg13g2_antennanp ANTENNA_2280 (.A(net524));
 sg13g2_antennanp ANTENNA_2281 (.A(net524));
 sg13g2_antennanp ANTENNA_2282 (.A(net524));
 sg13g2_antennanp ANTENNA_2283 (.A(net524));
 sg13g2_antennanp ANTENNA_2284 (.A(net524));
 sg13g2_antennanp ANTENNA_2285 (.A(net524));
 sg13g2_antennanp ANTENNA_2286 (.A(net524));
 sg13g2_antennanp ANTENNA_2287 (.A(net524));
 sg13g2_antennanp ANTENNA_2288 (.A(net524));
 sg13g2_antennanp ANTENNA_2289 (.A(net524));
 sg13g2_antennanp ANTENNA_2290 (.A(net524));
 sg13g2_antennanp ANTENNA_2291 (.A(net524));
 sg13g2_antennanp ANTENNA_2292 (.A(net524));
 sg13g2_antennanp ANTENNA_2293 (.A(net524));
 sg13g2_antennanp ANTENNA_2294 (.A(net524));
 sg13g2_antennanp ANTENNA_2295 (.A(net656));
 sg13g2_antennanp ANTENNA_2296 (.A(net656));
 sg13g2_antennanp ANTENNA_2297 (.A(net656));
 sg13g2_antennanp ANTENNA_2298 (.A(net656));
 sg13g2_antennanp ANTENNA_2299 (.A(net656));
 sg13g2_antennanp ANTENNA_2300 (.A(net656));
 sg13g2_antennanp ANTENNA_2301 (.A(net656));
 sg13g2_antennanp ANTENNA_2302 (.A(net656));
 sg13g2_antennanp ANTENNA_2303 (.A(net656));
 sg13g2_antennanp ANTENNA_2304 (.A(net685));
 sg13g2_antennanp ANTENNA_2305 (.A(net685));
 sg13g2_antennanp ANTENNA_2306 (.A(net685));
 sg13g2_antennanp ANTENNA_2307 (.A(net685));
 sg13g2_antennanp ANTENNA_2308 (.A(net685));
 sg13g2_antennanp ANTENNA_2309 (.A(net685));
 sg13g2_antennanp ANTENNA_2310 (.A(net685));
 sg13g2_antennanp ANTENNA_2311 (.A(net685));
 sg13g2_antennanp ANTENNA_2312 (.A(net685));
 sg13g2_antennanp ANTENNA_2313 (.A(net707));
 sg13g2_antennanp ANTENNA_2314 (.A(net707));
 sg13g2_antennanp ANTENNA_2315 (.A(net707));
 sg13g2_antennanp ANTENNA_2316 (.A(net707));
 sg13g2_antennanp ANTENNA_2317 (.A(net707));
 sg13g2_antennanp ANTENNA_2318 (.A(net707));
 sg13g2_antennanp ANTENNA_2319 (.A(net707));
 sg13g2_antennanp ANTENNA_2320 (.A(net707));
 sg13g2_antennanp ANTENNA_2321 (.A(net707));
 sg13g2_antennanp ANTENNA_2322 (.A(net803));
 sg13g2_antennanp ANTENNA_2323 (.A(net803));
 sg13g2_antennanp ANTENNA_2324 (.A(net803));
 sg13g2_antennanp ANTENNA_2325 (.A(net803));
 sg13g2_antennanp ANTENNA_2326 (.A(net803));
 sg13g2_antennanp ANTENNA_2327 (.A(net803));
 sg13g2_antennanp ANTENNA_2328 (.A(net803));
 sg13g2_antennanp ANTENNA_2329 (.A(net803));
 sg13g2_antennanp ANTENNA_2330 (.A(net803));
 sg13g2_antennanp ANTENNA_2331 (.A(net803));
 sg13g2_antennanp ANTENNA_2332 (.A(net803));
 sg13g2_antennanp ANTENNA_2333 (.A(net803));
 sg13g2_antennanp ANTENNA_2334 (.A(net803));
 sg13g2_antennanp ANTENNA_2335 (.A(net803));
 sg13g2_antennanp ANTENNA_2336 (.A(net888));
 sg13g2_antennanp ANTENNA_2337 (.A(net888));
 sg13g2_antennanp ANTENNA_2338 (.A(net888));
 sg13g2_antennanp ANTENNA_2339 (.A(net888));
 sg13g2_antennanp ANTENNA_2340 (.A(net888));
 sg13g2_antennanp ANTENNA_2341 (.A(net888));
 sg13g2_antennanp ANTENNA_2342 (.A(net888));
 sg13g2_antennanp ANTENNA_2343 (.A(net888));
 sg13g2_antennanp ANTENNA_2344 (.A(net928));
 sg13g2_antennanp ANTENNA_2345 (.A(net928));
 sg13g2_antennanp ANTENNA_2346 (.A(net928));
 sg13g2_antennanp ANTENNA_2347 (.A(net928));
 sg13g2_antennanp ANTENNA_2348 (.A(net928));
 sg13g2_antennanp ANTENNA_2349 (.A(net928));
 sg13g2_antennanp ANTENNA_2350 (.A(net928));
 sg13g2_antennanp ANTENNA_2351 (.A(net928));
 sg13g2_antennanp ANTENNA_2352 (.A(net928));
 sg13g2_antennanp ANTENNA_2353 (.A(net983));
 sg13g2_antennanp ANTENNA_2354 (.A(net983));
 sg13g2_antennanp ANTENNA_2355 (.A(net983));
 sg13g2_antennanp ANTENNA_2356 (.A(net983));
 sg13g2_antennanp ANTENNA_2357 (.A(net983));
 sg13g2_antennanp ANTENNA_2358 (.A(net983));
 sg13g2_antennanp ANTENNA_2359 (.A(net983));
 sg13g2_antennanp ANTENNA_2360 (.A(net983));
 sg13g2_antennanp ANTENNA_2361 (.A(net984));
 sg13g2_antennanp ANTENNA_2362 (.A(net984));
 sg13g2_antennanp ANTENNA_2363 (.A(net984));
 sg13g2_antennanp ANTENNA_2364 (.A(net984));
 sg13g2_antennanp ANTENNA_2365 (.A(net984));
 sg13g2_antennanp ANTENNA_2366 (.A(net984));
 sg13g2_antennanp ANTENNA_2367 (.A(net984));
 sg13g2_antennanp ANTENNA_2368 (.A(net984));
 sg13g2_antennanp ANTENNA_2369 (.A(net984));
 sg13g2_antennanp ANTENNA_2370 (.A(net984));
 sg13g2_antennanp ANTENNA_2371 (.A(net984));
 sg13g2_antennanp ANTENNA_2372 (.A(net984));
 sg13g2_antennanp ANTENNA_2373 (.A(net984));
 sg13g2_antennanp ANTENNA_2374 (.A(net984));
 sg13g2_antennanp ANTENNA_2375 (.A(net984));
 sg13g2_antennanp ANTENNA_2376 (.A(net984));
 sg13g2_antennanp ANTENNA_2377 (.A(net984));
 sg13g2_antennanp ANTENNA_2378 (.A(net984));
 sg13g2_antennanp ANTENNA_2379 (.A(net984));
 sg13g2_antennanp ANTENNA_2380 (.A(net984));
 sg13g2_antennanp ANTENNA_2381 (.A(net984));
 sg13g2_antennanp ANTENNA_2382 (.A(net984));
 sg13g2_antennanp ANTENNA_2383 (.A(net984));
 sg13g2_antennanp ANTENNA_2384 (.A(net984));
 sg13g2_antennanp ANTENNA_2385 (.A(net984));
 sg13g2_antennanp ANTENNA_2386 (.A(net984));
 sg13g2_antennanp ANTENNA_2387 (.A(net984));
 sg13g2_antennanp ANTENNA_2388 (.A(net984));
 sg13g2_antennanp ANTENNA_2389 (.A(net984));
 sg13g2_antennanp ANTENNA_2390 (.A(net984));
 sg13g2_antennanp ANTENNA_2391 (.A(_00190_));
 sg13g2_antennanp ANTENNA_2392 (.A(_00228_));
 sg13g2_antennanp ANTENNA_2393 (.A(_00228_));
 sg13g2_antennanp ANTENNA_2394 (.A(_00235_));
 sg13g2_antennanp ANTENNA_2395 (.A(_00235_));
 sg13g2_antennanp ANTENNA_2396 (.A(_01052_));
 sg13g2_antennanp ANTENNA_2397 (.A(_01052_));
 sg13g2_antennanp ANTENNA_2398 (.A(_02953_));
 sg13g2_antennanp ANTENNA_2399 (.A(_02953_));
 sg13g2_antennanp ANTENNA_2400 (.A(_02953_));
 sg13g2_antennanp ANTENNA_2401 (.A(_02953_));
 sg13g2_antennanp ANTENNA_2402 (.A(_02965_));
 sg13g2_antennanp ANTENNA_2403 (.A(_02965_));
 sg13g2_antennanp ANTENNA_2404 (.A(_02965_));
 sg13g2_antennanp ANTENNA_2405 (.A(_02965_));
 sg13g2_antennanp ANTENNA_2406 (.A(_02965_));
 sg13g2_antennanp ANTENNA_2407 (.A(_02965_));
 sg13g2_antennanp ANTENNA_2408 (.A(_02965_));
 sg13g2_antennanp ANTENNA_2409 (.A(_02965_));
 sg13g2_antennanp ANTENNA_2410 (.A(_02965_));
 sg13g2_antennanp ANTENNA_2411 (.A(_02965_));
 sg13g2_antennanp ANTENNA_2412 (.A(_03429_));
 sg13g2_antennanp ANTENNA_2413 (.A(_03429_));
 sg13g2_antennanp ANTENNA_2414 (.A(_03429_));
 sg13g2_antennanp ANTENNA_2415 (.A(_03429_));
 sg13g2_antennanp ANTENNA_2416 (.A(_03435_));
 sg13g2_antennanp ANTENNA_2417 (.A(_03435_));
 sg13g2_antennanp ANTENNA_2418 (.A(_03435_));
 sg13g2_antennanp ANTENNA_2419 (.A(_03435_));
 sg13g2_antennanp ANTENNA_2420 (.A(_03435_));
 sg13g2_antennanp ANTENNA_2421 (.A(_03435_));
 sg13g2_antennanp ANTENNA_2422 (.A(_03435_));
 sg13g2_antennanp ANTENNA_2423 (.A(_03435_));
 sg13g2_antennanp ANTENNA_2424 (.A(_03435_));
 sg13g2_antennanp ANTENNA_2425 (.A(_04742_));
 sg13g2_antennanp ANTENNA_2426 (.A(_04742_));
 sg13g2_antennanp ANTENNA_2427 (.A(_04742_));
 sg13g2_antennanp ANTENNA_2428 (.A(_04742_));
 sg13g2_antennanp ANTENNA_2429 (.A(_04887_));
 sg13g2_antennanp ANTENNA_2430 (.A(_04887_));
 sg13g2_antennanp ANTENNA_2431 (.A(_04887_));
 sg13g2_antennanp ANTENNA_2432 (.A(_04887_));
 sg13g2_antennanp ANTENNA_2433 (.A(_04894_));
 sg13g2_antennanp ANTENNA_2434 (.A(_05015_));
 sg13g2_antennanp ANTENNA_2435 (.A(_05169_));
 sg13g2_antennanp ANTENNA_2436 (.A(_05278_));
 sg13g2_antennanp ANTENNA_2437 (.A(_05280_));
 sg13g2_antennanp ANTENNA_2438 (.A(_05372_));
 sg13g2_antennanp ANTENNA_2439 (.A(_05432_));
 sg13g2_antennanp ANTENNA_2440 (.A(_05508_));
 sg13g2_antennanp ANTENNA_2441 (.A(_05646_));
 sg13g2_antennanp ANTENNA_2442 (.A(_05650_));
 sg13g2_antennanp ANTENNA_2443 (.A(_05654_));
 sg13g2_antennanp ANTENNA_2444 (.A(_05742_));
 sg13g2_antennanp ANTENNA_2445 (.A(_05763_));
 sg13g2_antennanp ANTENNA_2446 (.A(_05763_));
 sg13g2_antennanp ANTENNA_2447 (.A(_05763_));
 sg13g2_antennanp ANTENNA_2448 (.A(_05763_));
 sg13g2_antennanp ANTENNA_2449 (.A(_05763_));
 sg13g2_antennanp ANTENNA_2450 (.A(_05763_));
 sg13g2_antennanp ANTENNA_2451 (.A(_05763_));
 sg13g2_antennanp ANTENNA_2452 (.A(_05766_));
 sg13g2_antennanp ANTENNA_2453 (.A(_05766_));
 sg13g2_antennanp ANTENNA_2454 (.A(_05766_));
 sg13g2_antennanp ANTENNA_2455 (.A(_05770_));
 sg13g2_antennanp ANTENNA_2456 (.A(_05770_));
 sg13g2_antennanp ANTENNA_2457 (.A(_05770_));
 sg13g2_antennanp ANTENNA_2458 (.A(_05770_));
 sg13g2_antennanp ANTENNA_2459 (.A(_05770_));
 sg13g2_antennanp ANTENNA_2460 (.A(_05770_));
 sg13g2_antennanp ANTENNA_2461 (.A(_05770_));
 sg13g2_antennanp ANTENNA_2462 (.A(_05770_));
 sg13g2_antennanp ANTENNA_2463 (.A(_05775_));
 sg13g2_antennanp ANTENNA_2464 (.A(_05775_));
 sg13g2_antennanp ANTENNA_2465 (.A(_05775_));
 sg13g2_antennanp ANTENNA_2466 (.A(_05785_));
 sg13g2_antennanp ANTENNA_2467 (.A(_05785_));
 sg13g2_antennanp ANTENNA_2468 (.A(_05785_));
 sg13g2_antennanp ANTENNA_2469 (.A(_05785_));
 sg13g2_antennanp ANTENNA_2470 (.A(_05785_));
 sg13g2_antennanp ANTENNA_2471 (.A(_05835_));
 sg13g2_antennanp ANTENNA_2472 (.A(_05835_));
 sg13g2_antennanp ANTENNA_2473 (.A(_05835_));
 sg13g2_antennanp ANTENNA_2474 (.A(_05835_));
 sg13g2_antennanp ANTENNA_2475 (.A(_05835_));
 sg13g2_antennanp ANTENNA_2476 (.A(_06843_));
 sg13g2_antennanp ANTENNA_2477 (.A(_06843_));
 sg13g2_antennanp ANTENNA_2478 (.A(_06843_));
 sg13g2_antennanp ANTENNA_2479 (.A(_07398_));
 sg13g2_antennanp ANTENNA_2480 (.A(_07433_));
 sg13g2_antennanp ANTENNA_2481 (.A(_07434_));
 sg13g2_antennanp ANTENNA_2482 (.A(_08297_));
 sg13g2_antennanp ANTENNA_2483 (.A(_08297_));
 sg13g2_antennanp ANTENNA_2484 (.A(_08502_));
 sg13g2_antennanp ANTENNA_2485 (.A(_08502_));
 sg13g2_antennanp ANTENNA_2486 (.A(_08502_));
 sg13g2_antennanp ANTENNA_2487 (.A(_08502_));
 sg13g2_antennanp ANTENNA_2488 (.A(_08502_));
 sg13g2_antennanp ANTENNA_2489 (.A(_08502_));
 sg13g2_antennanp ANTENNA_2490 (.A(_08502_));
 sg13g2_antennanp ANTENNA_2491 (.A(_08533_));
 sg13g2_antennanp ANTENNA_2492 (.A(_08533_));
 sg13g2_antennanp ANTENNA_2493 (.A(_08533_));
 sg13g2_antennanp ANTENNA_2494 (.A(_08533_));
 sg13g2_antennanp ANTENNA_2495 (.A(_08533_));
 sg13g2_antennanp ANTENNA_2496 (.A(_08533_));
 sg13g2_antennanp ANTENNA_2497 (.A(_08558_));
 sg13g2_antennanp ANTENNA_2498 (.A(_08558_));
 sg13g2_antennanp ANTENNA_2499 (.A(_08558_));
 sg13g2_antennanp ANTENNA_2500 (.A(_08558_));
 sg13g2_antennanp ANTENNA_2501 (.A(_08558_));
 sg13g2_antennanp ANTENNA_2502 (.A(_08558_));
 sg13g2_antennanp ANTENNA_2503 (.A(_08558_));
 sg13g2_antennanp ANTENNA_2504 (.A(_08558_));
 sg13g2_antennanp ANTENNA_2505 (.A(_08558_));
 sg13g2_antennanp ANTENNA_2506 (.A(_08634_));
 sg13g2_antennanp ANTENNA_2507 (.A(_08634_));
 sg13g2_antennanp ANTENNA_2508 (.A(_08634_));
 sg13g2_antennanp ANTENNA_2509 (.A(_08634_));
 sg13g2_antennanp ANTENNA_2510 (.A(_08634_));
 sg13g2_antennanp ANTENNA_2511 (.A(_08634_));
 sg13g2_antennanp ANTENNA_2512 (.A(_08634_));
 sg13g2_antennanp ANTENNA_2513 (.A(_08634_));
 sg13g2_antennanp ANTENNA_2514 (.A(_08634_));
 sg13g2_antennanp ANTENNA_2515 (.A(_08679_));
 sg13g2_antennanp ANTENNA_2516 (.A(_08679_));
 sg13g2_antennanp ANTENNA_2517 (.A(_08679_));
 sg13g2_antennanp ANTENNA_2518 (.A(_08698_));
 sg13g2_antennanp ANTENNA_2519 (.A(_08698_));
 sg13g2_antennanp ANTENNA_2520 (.A(_08698_));
 sg13g2_antennanp ANTENNA_2521 (.A(_08728_));
 sg13g2_antennanp ANTENNA_2522 (.A(_08728_));
 sg13g2_antennanp ANTENNA_2523 (.A(_08728_));
 sg13g2_antennanp ANTENNA_2524 (.A(_08853_));
 sg13g2_antennanp ANTENNA_2525 (.A(_08918_));
 sg13g2_antennanp ANTENNA_2526 (.A(_08918_));
 sg13g2_antennanp ANTENNA_2527 (.A(_08918_));
 sg13g2_antennanp ANTENNA_2528 (.A(_08918_));
 sg13g2_antennanp ANTENNA_2529 (.A(_08918_));
 sg13g2_antennanp ANTENNA_2530 (.A(_08918_));
 sg13g2_antennanp ANTENNA_2531 (.A(_08918_));
 sg13g2_antennanp ANTENNA_2532 (.A(_08918_));
 sg13g2_antennanp ANTENNA_2533 (.A(_08918_));
 sg13g2_antennanp ANTENNA_2534 (.A(_08938_));
 sg13g2_antennanp ANTENNA_2535 (.A(_08959_));
 sg13g2_antennanp ANTENNA_2536 (.A(_08970_));
 sg13g2_antennanp ANTENNA_2537 (.A(_08970_));
 sg13g2_antennanp ANTENNA_2538 (.A(_08970_));
 sg13g2_antennanp ANTENNA_2539 (.A(_08970_));
 sg13g2_antennanp ANTENNA_2540 (.A(_09158_));
 sg13g2_antennanp ANTENNA_2541 (.A(_09158_));
 sg13g2_antennanp ANTENNA_2542 (.A(_09158_));
 sg13g2_antennanp ANTENNA_2543 (.A(_09158_));
 sg13g2_antennanp ANTENNA_2544 (.A(_09158_));
 sg13g2_antennanp ANTENNA_2545 (.A(_09158_));
 sg13g2_antennanp ANTENNA_2546 (.A(_09158_));
 sg13g2_antennanp ANTENNA_2547 (.A(_09158_));
 sg13g2_antennanp ANTENNA_2548 (.A(_09158_));
 sg13g2_antennanp ANTENNA_2549 (.A(_09167_));
 sg13g2_antennanp ANTENNA_2550 (.A(_09336_));
 sg13g2_antennanp ANTENNA_2551 (.A(_09336_));
 sg13g2_antennanp ANTENNA_2552 (.A(_09349_));
 sg13g2_antennanp ANTENNA_2553 (.A(_09349_));
 sg13g2_antennanp ANTENNA_2554 (.A(_09349_));
 sg13g2_antennanp ANTENNA_2555 (.A(_09349_));
 sg13g2_antennanp ANTENNA_2556 (.A(_09349_));
 sg13g2_antennanp ANTENNA_2557 (.A(_09349_));
 sg13g2_antennanp ANTENNA_2558 (.A(_09349_));
 sg13g2_antennanp ANTENNA_2559 (.A(_09349_));
 sg13g2_antennanp ANTENNA_2560 (.A(_09349_));
 sg13g2_antennanp ANTENNA_2561 (.A(_09349_));
 sg13g2_antennanp ANTENNA_2562 (.A(_09351_));
 sg13g2_antennanp ANTENNA_2563 (.A(_09351_));
 sg13g2_antennanp ANTENNA_2564 (.A(_09351_));
 sg13g2_antennanp ANTENNA_2565 (.A(_09351_));
 sg13g2_antennanp ANTENNA_2566 (.A(_09351_));
 sg13g2_antennanp ANTENNA_2567 (.A(_09351_));
 sg13g2_antennanp ANTENNA_2568 (.A(_09351_));
 sg13g2_antennanp ANTENNA_2569 (.A(_09351_));
 sg13g2_antennanp ANTENNA_2570 (.A(_09351_));
 sg13g2_antennanp ANTENNA_2571 (.A(_09380_));
 sg13g2_antennanp ANTENNA_2572 (.A(_09380_));
 sg13g2_antennanp ANTENNA_2573 (.A(_09380_));
 sg13g2_antennanp ANTENNA_2574 (.A(_09380_));
 sg13g2_antennanp ANTENNA_2575 (.A(_09386_));
 sg13g2_antennanp ANTENNA_2576 (.A(_09386_));
 sg13g2_antennanp ANTENNA_2577 (.A(_09386_));
 sg13g2_antennanp ANTENNA_2578 (.A(_09386_));
 sg13g2_antennanp ANTENNA_2579 (.A(_09386_));
 sg13g2_antennanp ANTENNA_2580 (.A(_09386_));
 sg13g2_antennanp ANTENNA_2581 (.A(_09386_));
 sg13g2_antennanp ANTENNA_2582 (.A(_09386_));
 sg13g2_antennanp ANTENNA_2583 (.A(_09388_));
 sg13g2_antennanp ANTENNA_2584 (.A(_09388_));
 sg13g2_antennanp ANTENNA_2585 (.A(_09388_));
 sg13g2_antennanp ANTENNA_2586 (.A(_09388_));
 sg13g2_antennanp ANTENNA_2587 (.A(_09389_));
 sg13g2_antennanp ANTENNA_2588 (.A(_09389_));
 sg13g2_antennanp ANTENNA_2589 (.A(_09389_));
 sg13g2_antennanp ANTENNA_2590 (.A(_09389_));
 sg13g2_antennanp ANTENNA_2591 (.A(_09389_));
 sg13g2_antennanp ANTENNA_2592 (.A(_09389_));
 sg13g2_antennanp ANTENNA_2593 (.A(_09389_));
 sg13g2_antennanp ANTENNA_2594 (.A(_09390_));
 sg13g2_antennanp ANTENNA_2595 (.A(_09390_));
 sg13g2_antennanp ANTENNA_2596 (.A(_09390_));
 sg13g2_antennanp ANTENNA_2597 (.A(_09390_));
 sg13g2_antennanp ANTENNA_2598 (.A(_09444_));
 sg13g2_antennanp ANTENNA_2599 (.A(_09444_));
 sg13g2_antennanp ANTENNA_2600 (.A(_09444_));
 sg13g2_antennanp ANTENNA_2601 (.A(_09444_));
 sg13g2_antennanp ANTENNA_2602 (.A(_09445_));
 sg13g2_antennanp ANTENNA_2603 (.A(_09445_));
 sg13g2_antennanp ANTENNA_2604 (.A(_09445_));
 sg13g2_antennanp ANTENNA_2605 (.A(_09445_));
 sg13g2_antennanp ANTENNA_2606 (.A(_09554_));
 sg13g2_antennanp ANTENNA_2607 (.A(_09554_));
 sg13g2_antennanp ANTENNA_2608 (.A(_09587_));
 sg13g2_antennanp ANTENNA_2609 (.A(_09608_));
 sg13g2_antennanp ANTENNA_2610 (.A(_09665_));
 sg13g2_antennanp ANTENNA_2611 (.A(_09695_));
 sg13g2_antennanp ANTENNA_2612 (.A(_09721_));
 sg13g2_antennanp ANTENNA_2613 (.A(_09742_));
 sg13g2_antennanp ANTENNA_2614 (.A(_09765_));
 sg13g2_antennanp ANTENNA_2615 (.A(_09765_));
 sg13g2_antennanp ANTENNA_2616 (.A(_09794_));
 sg13g2_antennanp ANTENNA_2617 (.A(_09796_));
 sg13g2_antennanp ANTENNA_2618 (.A(_09912_));
 sg13g2_antennanp ANTENNA_2619 (.A(_09990_));
 sg13g2_antennanp ANTENNA_2620 (.A(_09990_));
 sg13g2_antennanp ANTENNA_2621 (.A(_09990_));
 sg13g2_antennanp ANTENNA_2622 (.A(_09990_));
 sg13g2_antennanp ANTENNA_2623 (.A(_09990_));
 sg13g2_antennanp ANTENNA_2624 (.A(_09990_));
 sg13g2_antennanp ANTENNA_2625 (.A(_09990_));
 sg13g2_antennanp ANTENNA_2626 (.A(_09990_));
 sg13g2_antennanp ANTENNA_2627 (.A(_09990_));
 sg13g2_antennanp ANTENNA_2628 (.A(_09990_));
 sg13g2_antennanp ANTENNA_2629 (.A(_10246_));
 sg13g2_antennanp ANTENNA_2630 (.A(_10246_));
 sg13g2_antennanp ANTENNA_2631 (.A(_10246_));
 sg13g2_antennanp ANTENNA_2632 (.A(_10246_));
 sg13g2_antennanp ANTENNA_2633 (.A(_10246_));
 sg13g2_antennanp ANTENNA_2634 (.A(_10302_));
 sg13g2_antennanp ANTENNA_2635 (.A(_10302_));
 sg13g2_antennanp ANTENNA_2636 (.A(_10302_));
 sg13g2_antennanp ANTENNA_2637 (.A(_10302_));
 sg13g2_antennanp ANTENNA_2638 (.A(_10302_));
 sg13g2_antennanp ANTENNA_2639 (.A(_10302_));
 sg13g2_antennanp ANTENNA_2640 (.A(_10302_));
 sg13g2_antennanp ANTENNA_2641 (.A(_10302_));
 sg13g2_antennanp ANTENNA_2642 (.A(_10307_));
 sg13g2_antennanp ANTENNA_2643 (.A(_10307_));
 sg13g2_antennanp ANTENNA_2644 (.A(_10307_));
 sg13g2_antennanp ANTENNA_2645 (.A(_10307_));
 sg13g2_antennanp ANTENNA_2646 (.A(_10307_));
 sg13g2_antennanp ANTENNA_2647 (.A(_10307_));
 sg13g2_antennanp ANTENNA_2648 (.A(_10307_));
 sg13g2_antennanp ANTENNA_2649 (.A(_10307_));
 sg13g2_antennanp ANTENNA_2650 (.A(_10312_));
 sg13g2_antennanp ANTENNA_2651 (.A(_10312_));
 sg13g2_antennanp ANTENNA_2652 (.A(_10312_));
 sg13g2_antennanp ANTENNA_2653 (.A(_10312_));
 sg13g2_antennanp ANTENNA_2654 (.A(_10312_));
 sg13g2_antennanp ANTENNA_2655 (.A(_10312_));
 sg13g2_antennanp ANTENNA_2656 (.A(_10312_));
 sg13g2_antennanp ANTENNA_2657 (.A(_10312_));
 sg13g2_antennanp ANTENNA_2658 (.A(_10326_));
 sg13g2_antennanp ANTENNA_2659 (.A(_10326_));
 sg13g2_antennanp ANTENNA_2660 (.A(_10326_));
 sg13g2_antennanp ANTENNA_2661 (.A(_10326_));
 sg13g2_antennanp ANTENNA_2662 (.A(_10326_));
 sg13g2_antennanp ANTENNA_2663 (.A(_10326_));
 sg13g2_antennanp ANTENNA_2664 (.A(_10326_));
 sg13g2_antennanp ANTENNA_2665 (.A(_10326_));
 sg13g2_antennanp ANTENNA_2666 (.A(_10339_));
 sg13g2_antennanp ANTENNA_2667 (.A(_10339_));
 sg13g2_antennanp ANTENNA_2668 (.A(_10339_));
 sg13g2_antennanp ANTENNA_2669 (.A(_10339_));
 sg13g2_antennanp ANTENNA_2670 (.A(_10339_));
 sg13g2_antennanp ANTENNA_2671 (.A(_10339_));
 sg13g2_antennanp ANTENNA_2672 (.A(_10339_));
 sg13g2_antennanp ANTENNA_2673 (.A(_10344_));
 sg13g2_antennanp ANTENNA_2674 (.A(_10344_));
 sg13g2_antennanp ANTENNA_2675 (.A(_10344_));
 sg13g2_antennanp ANTENNA_2676 (.A(_10344_));
 sg13g2_antennanp ANTENNA_2677 (.A(_10344_));
 sg13g2_antennanp ANTENNA_2678 (.A(_10344_));
 sg13g2_antennanp ANTENNA_2679 (.A(_10344_));
 sg13g2_antennanp ANTENNA_2680 (.A(_10344_));
 sg13g2_antennanp ANTENNA_2681 (.A(_10645_));
 sg13g2_antennanp ANTENNA_2682 (.A(_10645_));
 sg13g2_antennanp ANTENNA_2683 (.A(_11129_));
 sg13g2_antennanp ANTENNA_2684 (.A(_12004_));
 sg13g2_antennanp ANTENNA_2685 (.A(_12004_));
 sg13g2_antennanp ANTENNA_2686 (.A(_12004_));
 sg13g2_antennanp ANTENNA_2687 (.A(_12004_));
 sg13g2_antennanp ANTENNA_2688 (.A(_12058_));
 sg13g2_antennanp ANTENNA_2689 (.A(_12058_));
 sg13g2_antennanp ANTENNA_2690 (.A(_12058_));
 sg13g2_antennanp ANTENNA_2691 (.A(_12058_));
 sg13g2_antennanp ANTENNA_2692 (.A(_12058_));
 sg13g2_antennanp ANTENNA_2693 (.A(_12058_));
 sg13g2_antennanp ANTENNA_2694 (.A(_12058_));
 sg13g2_antennanp ANTENNA_2695 (.A(_12058_));
 sg13g2_antennanp ANTENNA_2696 (.A(_12058_));
 sg13g2_antennanp ANTENNA_2697 (.A(_12127_));
 sg13g2_antennanp ANTENNA_2698 (.A(_12127_));
 sg13g2_antennanp ANTENNA_2699 (.A(_12127_));
 sg13g2_antennanp ANTENNA_2700 (.A(_12127_));
 sg13g2_antennanp ANTENNA_2701 (.A(_12127_));
 sg13g2_antennanp ANTENNA_2702 (.A(_12127_));
 sg13g2_antennanp ANTENNA_2703 (.A(_12127_));
 sg13g2_antennanp ANTENNA_2704 (.A(_12127_));
 sg13g2_antennanp ANTENNA_2705 (.A(_12127_));
 sg13g2_antennanp ANTENNA_2706 (.A(_12152_));
 sg13g2_antennanp ANTENNA_2707 (.A(_12152_));
 sg13g2_antennanp ANTENNA_2708 (.A(_12152_));
 sg13g2_antennanp ANTENNA_2709 (.A(_12152_));
 sg13g2_antennanp ANTENNA_2710 (.A(_12152_));
 sg13g2_antennanp ANTENNA_2711 (.A(_12152_));
 sg13g2_antennanp ANTENNA_2712 (.A(_12152_));
 sg13g2_antennanp ANTENNA_2713 (.A(_12152_));
 sg13g2_antennanp ANTENNA_2714 (.A(_12218_));
 sg13g2_antennanp ANTENNA_2715 (.A(_12218_));
 sg13g2_antennanp ANTENNA_2716 (.A(_12218_));
 sg13g2_antennanp ANTENNA_2717 (.A(_12218_));
 sg13g2_antennanp ANTENNA_2718 (.A(_12218_));
 sg13g2_antennanp ANTENNA_2719 (.A(_12218_));
 sg13g2_antennanp ANTENNA_2720 (.A(_12218_));
 sg13g2_antennanp ANTENNA_2721 (.A(_12218_));
 sg13g2_antennanp ANTENNA_2722 (.A(_12218_));
 sg13g2_antennanp ANTENNA_2723 (.A(_12223_));
 sg13g2_antennanp ANTENNA_2724 (.A(_12223_));
 sg13g2_antennanp ANTENNA_2725 (.A(_12223_));
 sg13g2_antennanp ANTENNA_2726 (.A(_12223_));
 sg13g2_antennanp ANTENNA_2727 (.A(_12223_));
 sg13g2_antennanp ANTENNA_2728 (.A(_12223_));
 sg13g2_antennanp ANTENNA_2729 (.A(_12223_));
 sg13g2_antennanp ANTENNA_2730 (.A(_12223_));
 sg13g2_antennanp ANTENNA_2731 (.A(_12223_));
 sg13g2_antennanp ANTENNA_2732 (.A(_12229_));
 sg13g2_antennanp ANTENNA_2733 (.A(_12229_));
 sg13g2_antennanp ANTENNA_2734 (.A(_12229_));
 sg13g2_antennanp ANTENNA_2735 (.A(_12229_));
 sg13g2_antennanp ANTENNA_2736 (.A(_12229_));
 sg13g2_antennanp ANTENNA_2737 (.A(_12229_));
 sg13g2_antennanp ANTENNA_2738 (.A(_12229_));
 sg13g2_antennanp ANTENNA_2739 (.A(_12229_));
 sg13g2_antennanp ANTENNA_2740 (.A(_12229_));
 sg13g2_antennanp ANTENNA_2741 (.A(_12558_));
 sg13g2_antennanp ANTENNA_2742 (.A(_12558_));
 sg13g2_antennanp ANTENNA_2743 (.A(_12558_));
 sg13g2_antennanp ANTENNA_2744 (.A(_12558_));
 sg13g2_antennanp ANTENNA_2745 (.A(_12558_));
 sg13g2_antennanp ANTENNA_2746 (.A(_12558_));
 sg13g2_antennanp ANTENNA_2747 (.A(_12558_));
 sg13g2_antennanp ANTENNA_2748 (.A(_12558_));
 sg13g2_antennanp ANTENNA_2749 (.A(_12558_));
 sg13g2_antennanp ANTENNA_2750 (.A(_12558_));
 sg13g2_antennanp ANTENNA_2751 (.A(_12726_));
 sg13g2_antennanp ANTENNA_2752 (.A(_12726_));
 sg13g2_antennanp ANTENNA_2753 (.A(_12726_));
 sg13g2_antennanp ANTENNA_2754 (.A(clk));
 sg13g2_antennanp ANTENNA_2755 (.A(clk));
 sg13g2_antennanp ANTENNA_2756 (.A(\cpu.ex.pc[3] ));
 sg13g2_antennanp ANTENNA_2757 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_2758 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_2759 (.A(net12));
 sg13g2_antennanp ANTENNA_2760 (.A(net12));
 sg13g2_antennanp ANTENNA_2761 (.A(net12));
 sg13g2_antennanp ANTENNA_2762 (.A(net437));
 sg13g2_antennanp ANTENNA_2763 (.A(net437));
 sg13g2_antennanp ANTENNA_2764 (.A(net437));
 sg13g2_antennanp ANTENNA_2765 (.A(net437));
 sg13g2_antennanp ANTENNA_2766 (.A(net437));
 sg13g2_antennanp ANTENNA_2767 (.A(net437));
 sg13g2_antennanp ANTENNA_2768 (.A(net437));
 sg13g2_antennanp ANTENNA_2769 (.A(net437));
 sg13g2_antennanp ANTENNA_2770 (.A(net437));
 sg13g2_antennanp ANTENNA_2771 (.A(net437));
 sg13g2_antennanp ANTENNA_2772 (.A(net437));
 sg13g2_antennanp ANTENNA_2773 (.A(net437));
 sg13g2_antennanp ANTENNA_2774 (.A(net437));
 sg13g2_antennanp ANTENNA_2775 (.A(net437));
 sg13g2_antennanp ANTENNA_2776 (.A(net437));
 sg13g2_antennanp ANTENNA_2777 (.A(net437));
 sg13g2_antennanp ANTENNA_2778 (.A(net437));
 sg13g2_antennanp ANTENNA_2779 (.A(net656));
 sg13g2_antennanp ANTENNA_2780 (.A(net656));
 sg13g2_antennanp ANTENNA_2781 (.A(net656));
 sg13g2_antennanp ANTENNA_2782 (.A(net656));
 sg13g2_antennanp ANTENNA_2783 (.A(net656));
 sg13g2_antennanp ANTENNA_2784 (.A(net656));
 sg13g2_antennanp ANTENNA_2785 (.A(net656));
 sg13g2_antennanp ANTENNA_2786 (.A(net656));
 sg13g2_antennanp ANTENNA_2787 (.A(net656));
 sg13g2_antennanp ANTENNA_2788 (.A(net656));
 sg13g2_antennanp ANTENNA_2789 (.A(net656));
 sg13g2_antennanp ANTENNA_2790 (.A(net656));
 sg13g2_antennanp ANTENNA_2791 (.A(net656));
 sg13g2_antennanp ANTENNA_2792 (.A(net656));
 sg13g2_antennanp ANTENNA_2793 (.A(net656));
 sg13g2_antennanp ANTENNA_2794 (.A(net656));
 sg13g2_antennanp ANTENNA_2795 (.A(net656));
 sg13g2_antennanp ANTENNA_2796 (.A(net685));
 sg13g2_antennanp ANTENNA_2797 (.A(net685));
 sg13g2_antennanp ANTENNA_2798 (.A(net685));
 sg13g2_antennanp ANTENNA_2799 (.A(net685));
 sg13g2_antennanp ANTENNA_2800 (.A(net685));
 sg13g2_antennanp ANTENNA_2801 (.A(net685));
 sg13g2_antennanp ANTENNA_2802 (.A(net685));
 sg13g2_antennanp ANTENNA_2803 (.A(net685));
 sg13g2_antennanp ANTENNA_2804 (.A(net685));
 sg13g2_antennanp ANTENNA_2805 (.A(net707));
 sg13g2_antennanp ANTENNA_2806 (.A(net707));
 sg13g2_antennanp ANTENNA_2807 (.A(net707));
 sg13g2_antennanp ANTENNA_2808 (.A(net707));
 sg13g2_antennanp ANTENNA_2809 (.A(net707));
 sg13g2_antennanp ANTENNA_2810 (.A(net707));
 sg13g2_antennanp ANTENNA_2811 (.A(net707));
 sg13g2_antennanp ANTENNA_2812 (.A(net707));
 sg13g2_antennanp ANTENNA_2813 (.A(net707));
 sg13g2_antennanp ANTENNA_2814 (.A(net803));
 sg13g2_antennanp ANTENNA_2815 (.A(net803));
 sg13g2_antennanp ANTENNA_2816 (.A(net803));
 sg13g2_antennanp ANTENNA_2817 (.A(net803));
 sg13g2_antennanp ANTENNA_2818 (.A(net803));
 sg13g2_antennanp ANTENNA_2819 (.A(net803));
 sg13g2_antennanp ANTENNA_2820 (.A(net803));
 sg13g2_antennanp ANTENNA_2821 (.A(net803));
 sg13g2_antennanp ANTENNA_2822 (.A(net803));
 sg13g2_antennanp ANTENNA_2823 (.A(net803));
 sg13g2_antennanp ANTENNA_2824 (.A(net803));
 sg13g2_antennanp ANTENNA_2825 (.A(net803));
 sg13g2_antennanp ANTENNA_2826 (.A(net803));
 sg13g2_antennanp ANTENNA_2827 (.A(net803));
 sg13g2_antennanp ANTENNA_2828 (.A(net888));
 sg13g2_antennanp ANTENNA_2829 (.A(net888));
 sg13g2_antennanp ANTENNA_2830 (.A(net888));
 sg13g2_antennanp ANTENNA_2831 (.A(net888));
 sg13g2_antennanp ANTENNA_2832 (.A(net888));
 sg13g2_antennanp ANTENNA_2833 (.A(net888));
 sg13g2_antennanp ANTENNA_2834 (.A(net888));
 sg13g2_antennanp ANTENNA_2835 (.A(net888));
 sg13g2_antennanp ANTENNA_2836 (.A(net888));
 sg13g2_antennanp ANTENNA_2837 (.A(net928));
 sg13g2_antennanp ANTENNA_2838 (.A(net928));
 sg13g2_antennanp ANTENNA_2839 (.A(net928));
 sg13g2_antennanp ANTENNA_2840 (.A(net928));
 sg13g2_antennanp ANTENNA_2841 (.A(net928));
 sg13g2_antennanp ANTENNA_2842 (.A(net928));
 sg13g2_antennanp ANTENNA_2843 (.A(net928));
 sg13g2_antennanp ANTENNA_2844 (.A(net928));
 sg13g2_antennanp ANTENNA_2845 (.A(net928));
 sg13g2_antennanp ANTENNA_2846 (.A(net984));
 sg13g2_antennanp ANTENNA_2847 (.A(net984));
 sg13g2_antennanp ANTENNA_2848 (.A(net984));
 sg13g2_antennanp ANTENNA_2849 (.A(net984));
 sg13g2_antennanp ANTENNA_2850 (.A(net984));
 sg13g2_antennanp ANTENNA_2851 (.A(net984));
 sg13g2_antennanp ANTENNA_2852 (.A(net984));
 sg13g2_antennanp ANTENNA_2853 (.A(net984));
 sg13g2_antennanp ANTENNA_2854 (.A(net984));
 sg13g2_antennanp ANTENNA_2855 (.A(net984));
 sg13g2_antennanp ANTENNA_2856 (.A(net984));
 sg13g2_antennanp ANTENNA_2857 (.A(net984));
 sg13g2_antennanp ANTENNA_2858 (.A(net984));
 sg13g2_antennanp ANTENNA_2859 (.A(net984));
 sg13g2_antennanp ANTENNA_2860 (.A(net984));
 sg13g2_antennanp ANTENNA_2861 (.A(net984));
 sg13g2_antennanp ANTENNA_2862 (.A(net984));
 sg13g2_antennanp ANTENNA_2863 (.A(net984));
 sg13g2_antennanp ANTENNA_2864 (.A(net984));
 sg13g2_antennanp ANTENNA_2865 (.A(net984));
 sg13g2_antennanp ANTENNA_2866 (.A(net984));
 sg13g2_antennanp ANTENNA_2867 (.A(net984));
 sg13g2_antennanp ANTENNA_2868 (.A(net984));
 sg13g2_antennanp ANTENNA_2869 (.A(net984));
 sg13g2_antennanp ANTENNA_2870 (.A(net984));
 sg13g2_antennanp ANTENNA_2871 (.A(net984));
 sg13g2_antennanp ANTENNA_2872 (.A(net984));
 sg13g2_antennanp ANTENNA_2873 (.A(net984));
 sg13g2_antennanp ANTENNA_2874 (.A(net984));
 sg13g2_antennanp ANTENNA_2875 (.A(net984));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_fill_2 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_96 ();
 sg13g2_decap_8 FILLER_0_103 ();
 sg13g2_decap_8 FILLER_0_110 ();
 sg13g2_decap_8 FILLER_0_117 ();
 sg13g2_decap_8 FILLER_0_124 ();
 sg13g2_decap_8 FILLER_0_131 ();
 sg13g2_decap_8 FILLER_0_138 ();
 sg13g2_decap_8 FILLER_0_145 ();
 sg13g2_decap_8 FILLER_0_152 ();
 sg13g2_decap_8 FILLER_0_159 ();
 sg13g2_decap_8 FILLER_0_166 ();
 sg13g2_decap_8 FILLER_0_173 ();
 sg13g2_decap_8 FILLER_0_180 ();
 sg13g2_decap_8 FILLER_0_187 ();
 sg13g2_decap_8 FILLER_0_194 ();
 sg13g2_decap_8 FILLER_0_201 ();
 sg13g2_decap_8 FILLER_0_208 ();
 sg13g2_decap_8 FILLER_0_256 ();
 sg13g2_decap_4 FILLER_0_263 ();
 sg13g2_fill_1 FILLER_0_267 ();
 sg13g2_fill_2 FILLER_0_330 ();
 sg13g2_fill_1 FILLER_0_339 ();
 sg13g2_fill_1 FILLER_0_355 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_438 ();
 sg13g2_decap_8 FILLER_0_445 ();
 sg13g2_fill_1 FILLER_0_452 ();
 sg13g2_fill_1 FILLER_0_457 ();
 sg13g2_decap_8 FILLER_0_475 ();
 sg13g2_decap_8 FILLER_0_482 ();
 sg13g2_decap_4 FILLER_0_489 ();
 sg13g2_fill_2 FILLER_0_493 ();
 sg13g2_decap_8 FILLER_0_499 ();
 sg13g2_decap_8 FILLER_0_506 ();
 sg13g2_decap_4 FILLER_0_513 ();
 sg13g2_fill_1 FILLER_0_517 ();
 sg13g2_decap_8 FILLER_0_544 ();
 sg13g2_decap_4 FILLER_0_551 ();
 sg13g2_fill_1 FILLER_0_555 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_fill_2 FILLER_0_567 ();
 sg13g2_fill_1 FILLER_0_569 ();
 sg13g2_decap_4 FILLER_0_609 ();
 sg13g2_fill_2 FILLER_0_613 ();
 sg13g2_decap_8 FILLER_0_619 ();
 sg13g2_decap_8 FILLER_0_626 ();
 sg13g2_decap_8 FILLER_0_633 ();
 sg13g2_decap_8 FILLER_0_640 ();
 sg13g2_decap_8 FILLER_0_647 ();
 sg13g2_decap_4 FILLER_0_654 ();
 sg13g2_decap_8 FILLER_0_662 ();
 sg13g2_decap_8 FILLER_0_669 ();
 sg13g2_decap_8 FILLER_0_676 ();
 sg13g2_decap_8 FILLER_0_683 ();
 sg13g2_fill_1 FILLER_0_690 ();
 sg13g2_decap_4 FILLER_0_695 ();
 sg13g2_fill_1 FILLER_0_699 ();
 sg13g2_decap_4 FILLER_0_708 ();
 sg13g2_fill_1 FILLER_0_712 ();
 sg13g2_decap_8 FILLER_0_717 ();
 sg13g2_fill_2 FILLER_0_724 ();
 sg13g2_fill_1 FILLER_0_726 ();
 sg13g2_decap_8 FILLER_0_731 ();
 sg13g2_decap_8 FILLER_0_738 ();
 sg13g2_decap_8 FILLER_0_745 ();
 sg13g2_decap_8 FILLER_0_752 ();
 sg13g2_decap_8 FILLER_0_759 ();
 sg13g2_decap_4 FILLER_0_766 ();
 sg13g2_fill_1 FILLER_0_770 ();
 sg13g2_fill_2 FILLER_0_780 ();
 sg13g2_decap_8 FILLER_0_786 ();
 sg13g2_decap_8 FILLER_0_793 ();
 sg13g2_decap_8 FILLER_0_800 ();
 sg13g2_decap_8 FILLER_0_807 ();
 sg13g2_decap_8 FILLER_0_814 ();
 sg13g2_decap_4 FILLER_0_821 ();
 sg13g2_fill_1 FILLER_0_825 ();
 sg13g2_decap_4 FILLER_0_830 ();
 sg13g2_fill_1 FILLER_0_834 ();
 sg13g2_decap_4 FILLER_0_840 ();
 sg13g2_fill_1 FILLER_0_844 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_decap_8 FILLER_0_861 ();
 sg13g2_fill_2 FILLER_0_868 ();
 sg13g2_fill_2 FILLER_0_896 ();
 sg13g2_decap_8 FILLER_0_919 ();
 sg13g2_decap_4 FILLER_0_926 ();
 sg13g2_fill_1 FILLER_0_930 ();
 sg13g2_decap_8 FILLER_0_935 ();
 sg13g2_decap_8 FILLER_0_942 ();
 sg13g2_fill_2 FILLER_0_949 ();
 sg13g2_fill_1 FILLER_0_951 ();
 sg13g2_decap_8 FILLER_0_982 ();
 sg13g2_decap_8 FILLER_0_989 ();
 sg13g2_decap_8 FILLER_0_996 ();
 sg13g2_decap_8 FILLER_0_1003 ();
 sg13g2_decap_8 FILLER_0_1010 ();
 sg13g2_decap_8 FILLER_0_1017 ();
 sg13g2_decap_8 FILLER_0_1024 ();
 sg13g2_decap_4 FILLER_0_1031 ();
 sg13g2_fill_2 FILLER_0_1035 ();
 sg13g2_fill_2 FILLER_0_1049 ();
 sg13g2_fill_1 FILLER_0_1051 ();
 sg13g2_fill_2 FILLER_0_1073 ();
 sg13g2_fill_1 FILLER_0_1075 ();
 sg13g2_fill_2 FILLER_0_1080 ();
 sg13g2_decap_8 FILLER_0_1090 ();
 sg13g2_decap_8 FILLER_0_1097 ();
 sg13g2_fill_1 FILLER_0_1104 ();
 sg13g2_decap_8 FILLER_0_1118 ();
 sg13g2_decap_8 FILLER_0_1125 ();
 sg13g2_fill_2 FILLER_0_1132 ();
 sg13g2_fill_1 FILLER_0_1134 ();
 sg13g2_decap_8 FILLER_0_1143 ();
 sg13g2_decap_8 FILLER_0_1150 ();
 sg13g2_decap_8 FILLER_0_1157 ();
 sg13g2_fill_2 FILLER_0_1164 ();
 sg13g2_decap_8 FILLER_0_1170 ();
 sg13g2_decap_8 FILLER_0_1177 ();
 sg13g2_fill_1 FILLER_0_1188 ();
 sg13g2_decap_8 FILLER_0_1193 ();
 sg13g2_decap_8 FILLER_0_1200 ();
 sg13g2_decap_8 FILLER_0_1207 ();
 sg13g2_decap_8 FILLER_0_1214 ();
 sg13g2_decap_8 FILLER_0_1221 ();
 sg13g2_decap_8 FILLER_0_1228 ();
 sg13g2_decap_8 FILLER_0_1235 ();
 sg13g2_fill_1 FILLER_0_1242 ();
 sg13g2_decap_8 FILLER_0_1269 ();
 sg13g2_decap_4 FILLER_0_1302 ();
 sg13g2_fill_2 FILLER_0_1306 ();
 sg13g2_decap_8 FILLER_0_1312 ();
 sg13g2_decap_8 FILLER_0_1319 ();
 sg13g2_decap_8 FILLER_0_1326 ();
 sg13g2_decap_8 FILLER_0_1333 ();
 sg13g2_decap_8 FILLER_0_1340 ();
 sg13g2_fill_2 FILLER_0_1347 ();
 sg13g2_fill_1 FILLER_0_1349 ();
 sg13g2_decap_8 FILLER_0_1376 ();
 sg13g2_decap_8 FILLER_0_1383 ();
 sg13g2_fill_2 FILLER_0_1390 ();
 sg13g2_fill_1 FILLER_0_1392 ();
 sg13g2_decap_8 FILLER_0_1397 ();
 sg13g2_decap_8 FILLER_0_1408 ();
 sg13g2_decap_8 FILLER_0_1415 ();
 sg13g2_decap_8 FILLER_0_1422 ();
 sg13g2_decap_8 FILLER_0_1429 ();
 sg13g2_decap_4 FILLER_0_1436 ();
 sg13g2_fill_1 FILLER_0_1440 ();
 sg13g2_decap_8 FILLER_0_1467 ();
 sg13g2_decap_8 FILLER_0_1474 ();
 sg13g2_decap_8 FILLER_0_1481 ();
 sg13g2_decap_4 FILLER_0_1488 ();
 sg13g2_fill_1 FILLER_0_1496 ();
 sg13g2_decap_8 FILLER_0_1501 ();
 sg13g2_decap_8 FILLER_0_1508 ();
 sg13g2_decap_8 FILLER_0_1515 ();
 sg13g2_decap_8 FILLER_0_1522 ();
 sg13g2_decap_8 FILLER_0_1529 ();
 sg13g2_decap_8 FILLER_0_1536 ();
 sg13g2_fill_1 FILLER_0_1551 ();
 sg13g2_decap_8 FILLER_0_1582 ();
 sg13g2_decap_8 FILLER_0_1589 ();
 sg13g2_decap_4 FILLER_0_1596 ();
 sg13g2_fill_1 FILLER_0_1600 ();
 sg13g2_decap_8 FILLER_0_1605 ();
 sg13g2_decap_8 FILLER_0_1612 ();
 sg13g2_decap_8 FILLER_0_1619 ();
 sg13g2_decap_8 FILLER_0_1626 ();
 sg13g2_decap_8 FILLER_0_1643 ();
 sg13g2_decap_8 FILLER_0_1650 ();
 sg13g2_decap_8 FILLER_0_1657 ();
 sg13g2_decap_8 FILLER_0_1664 ();
 sg13g2_fill_1 FILLER_0_1671 ();
 sg13g2_fill_1 FILLER_0_1676 ();
 sg13g2_decap_8 FILLER_0_1687 ();
 sg13g2_decap_8 FILLER_0_1694 ();
 sg13g2_decap_8 FILLER_0_1701 ();
 sg13g2_decap_8 FILLER_0_1708 ();
 sg13g2_decap_8 FILLER_0_1715 ();
 sg13g2_decap_8 FILLER_0_1722 ();
 sg13g2_decap_8 FILLER_0_1729 ();
 sg13g2_decap_8 FILLER_0_1736 ();
 sg13g2_decap_4 FILLER_0_1753 ();
 sg13g2_fill_2 FILLER_0_1757 ();
 sg13g2_decap_8 FILLER_0_1789 ();
 sg13g2_decap_8 FILLER_0_1796 ();
 sg13g2_decap_8 FILLER_0_1803 ();
 sg13g2_decap_8 FILLER_0_1810 ();
 sg13g2_decap_8 FILLER_0_1817 ();
 sg13g2_decap_8 FILLER_0_1824 ();
 sg13g2_decap_8 FILLER_0_1831 ();
 sg13g2_decap_8 FILLER_0_1838 ();
 sg13g2_decap_4 FILLER_0_1845 ();
 sg13g2_fill_2 FILLER_0_1849 ();
 sg13g2_fill_1 FILLER_0_1877 ();
 sg13g2_decap_8 FILLER_0_1899 ();
 sg13g2_decap_4 FILLER_0_1920 ();
 sg13g2_decap_8 FILLER_0_1928 ();
 sg13g2_decap_8 FILLER_0_1935 ();
 sg13g2_decap_8 FILLER_0_1942 ();
 sg13g2_decap_8 FILLER_0_1949 ();
 sg13g2_fill_2 FILLER_0_1956 ();
 sg13g2_fill_1 FILLER_0_1958 ();
 sg13g2_fill_1 FILLER_0_1963 ();
 sg13g2_decap_8 FILLER_0_1968 ();
 sg13g2_decap_8 FILLER_0_1975 ();
 sg13g2_decap_8 FILLER_0_1982 ();
 sg13g2_decap_4 FILLER_0_1989 ();
 sg13g2_fill_1 FILLER_0_1993 ();
 sg13g2_fill_2 FILLER_0_2008 ();
 sg13g2_decap_8 FILLER_0_2014 ();
 sg13g2_decap_8 FILLER_0_2021 ();
 sg13g2_decap_8 FILLER_0_2028 ();
 sg13g2_decap_8 FILLER_0_2035 ();
 sg13g2_decap_8 FILLER_0_2042 ();
 sg13g2_decap_8 FILLER_0_2049 ();
 sg13g2_decap_8 FILLER_0_2056 ();
 sg13g2_decap_8 FILLER_0_2063 ();
 sg13g2_fill_2 FILLER_0_2070 ();
 sg13g2_fill_1 FILLER_0_2072 ();
 sg13g2_decap_8 FILLER_0_2094 ();
 sg13g2_fill_2 FILLER_0_2101 ();
 sg13g2_decap_8 FILLER_0_2122 ();
 sg13g2_decap_8 FILLER_0_2129 ();
 sg13g2_decap_8 FILLER_0_2136 ();
 sg13g2_decap_8 FILLER_0_2143 ();
 sg13g2_decap_8 FILLER_0_2150 ();
 sg13g2_decap_8 FILLER_0_2157 ();
 sg13g2_decap_4 FILLER_0_2164 ();
 sg13g2_fill_1 FILLER_0_2168 ();
 sg13g2_decap_8 FILLER_0_2173 ();
 sg13g2_fill_2 FILLER_0_2180 ();
 sg13g2_fill_1 FILLER_0_2182 ();
 sg13g2_decap_8 FILLER_0_2197 ();
 sg13g2_decap_8 FILLER_0_2204 ();
 sg13g2_decap_8 FILLER_0_2211 ();
 sg13g2_decap_8 FILLER_0_2218 ();
 sg13g2_fill_2 FILLER_0_2225 ();
 sg13g2_fill_1 FILLER_0_2227 ();
 sg13g2_decap_8 FILLER_0_2232 ();
 sg13g2_decap_8 FILLER_0_2239 ();
 sg13g2_decap_8 FILLER_0_2246 ();
 sg13g2_decap_4 FILLER_0_2253 ();
 sg13g2_fill_2 FILLER_0_2257 ();
 sg13g2_fill_2 FILLER_0_2264 ();
 sg13g2_fill_1 FILLER_0_2266 ();
 sg13g2_decap_8 FILLER_0_2293 ();
 sg13g2_decap_8 FILLER_0_2300 ();
 sg13g2_decap_8 FILLER_0_2307 ();
 sg13g2_decap_8 FILLER_0_2314 ();
 sg13g2_decap_8 FILLER_0_2321 ();
 sg13g2_decap_8 FILLER_0_2328 ();
 sg13g2_fill_2 FILLER_0_2335 ();
 sg13g2_decap_8 FILLER_0_2373 ();
 sg13g2_decap_8 FILLER_0_2380 ();
 sg13g2_decap_8 FILLER_0_2387 ();
 sg13g2_decap_8 FILLER_0_2394 ();
 sg13g2_decap_8 FILLER_0_2401 ();
 sg13g2_decap_8 FILLER_0_2408 ();
 sg13g2_decap_8 FILLER_0_2415 ();
 sg13g2_decap_8 FILLER_0_2422 ();
 sg13g2_decap_8 FILLER_0_2429 ();
 sg13g2_decap_8 FILLER_0_2436 ();
 sg13g2_decap_8 FILLER_0_2443 ();
 sg13g2_decap_8 FILLER_0_2450 ();
 sg13g2_decap_8 FILLER_0_2457 ();
 sg13g2_decap_8 FILLER_0_2464 ();
 sg13g2_decap_8 FILLER_0_2471 ();
 sg13g2_decap_8 FILLER_0_2478 ();
 sg13g2_decap_8 FILLER_0_2485 ();
 sg13g2_decap_8 FILLER_0_2492 ();
 sg13g2_decap_8 FILLER_0_2499 ();
 sg13g2_decap_8 FILLER_0_2506 ();
 sg13g2_decap_8 FILLER_0_2513 ();
 sg13g2_decap_8 FILLER_0_2520 ();
 sg13g2_decap_8 FILLER_0_2527 ();
 sg13g2_decap_8 FILLER_0_2534 ();
 sg13g2_decap_8 FILLER_0_2541 ();
 sg13g2_decap_8 FILLER_0_2548 ();
 sg13g2_decap_8 FILLER_0_2555 ();
 sg13g2_decap_8 FILLER_0_2562 ();
 sg13g2_decap_8 FILLER_0_2569 ();
 sg13g2_decap_8 FILLER_0_2576 ();
 sg13g2_decap_8 FILLER_0_2583 ();
 sg13g2_decap_8 FILLER_0_2590 ();
 sg13g2_decap_8 FILLER_0_2597 ();
 sg13g2_decap_8 FILLER_0_2604 ();
 sg13g2_decap_8 FILLER_0_2611 ();
 sg13g2_decap_8 FILLER_0_2618 ();
 sg13g2_decap_8 FILLER_0_2625 ();
 sg13g2_decap_8 FILLER_0_2632 ();
 sg13g2_decap_8 FILLER_0_2639 ();
 sg13g2_decap_8 FILLER_0_2646 ();
 sg13g2_decap_8 FILLER_0_2653 ();
 sg13g2_decap_8 FILLER_0_2660 ();
 sg13g2_fill_2 FILLER_0_2667 ();
 sg13g2_fill_1 FILLER_0_2669 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_4 FILLER_1_15 ();
 sg13g2_fill_1 FILLER_1_19 ();
 sg13g2_decap_8 FILLER_1_24 ();
 sg13g2_fill_2 FILLER_1_31 ();
 sg13g2_fill_1 FILLER_1_33 ();
 sg13g2_fill_1 FILLER_1_72 ();
 sg13g2_decap_8 FILLER_1_107 ();
 sg13g2_fill_1 FILLER_1_114 ();
 sg13g2_decap_8 FILLER_1_145 ();
 sg13g2_decap_8 FILLER_1_152 ();
 sg13g2_decap_8 FILLER_1_159 ();
 sg13g2_decap_8 FILLER_1_166 ();
 sg13g2_decap_8 FILLER_1_173 ();
 sg13g2_decap_8 FILLER_1_180 ();
 sg13g2_decap_8 FILLER_1_187 ();
 sg13g2_decap_8 FILLER_1_194 ();
 sg13g2_decap_8 FILLER_1_201 ();
 sg13g2_fill_2 FILLER_1_208 ();
 sg13g2_fill_2 FILLER_1_274 ();
 sg13g2_fill_1 FILLER_1_282 ();
 sg13g2_fill_1 FILLER_1_315 ();
 sg13g2_fill_1 FILLER_1_319 ();
 sg13g2_fill_1 FILLER_1_355 ();
 sg13g2_decap_8 FILLER_1_366 ();
 sg13g2_decap_8 FILLER_1_373 ();
 sg13g2_decap_8 FILLER_1_380 ();
 sg13g2_fill_2 FILLER_1_439 ();
 sg13g2_decap_8 FILLER_1_472 ();
 sg13g2_decap_4 FILLER_1_479 ();
 sg13g2_fill_1 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_514 ();
 sg13g2_fill_1 FILLER_1_551 ();
 sg13g2_fill_2 FILLER_1_583 ();
 sg13g2_fill_2 FILLER_1_611 ();
 sg13g2_fill_1 FILLER_1_613 ();
 sg13g2_fill_2 FILLER_1_619 ();
 sg13g2_fill_1 FILLER_1_621 ();
 sg13g2_fill_2 FILLER_1_648 ();
 sg13g2_fill_1 FILLER_1_650 ();
 sg13g2_decap_8 FILLER_1_677 ();
 sg13g2_decap_4 FILLER_1_741 ();
 sg13g2_decap_8 FILLER_1_801 ();
 sg13g2_fill_1 FILLER_1_808 ();
 sg13g2_fill_1 FILLER_1_827 ();
 sg13g2_decap_8 FILLER_1_858 ();
 sg13g2_decap_4 FILLER_1_865 ();
 sg13g2_fill_1 FILLER_1_869 ();
 sg13g2_fill_1 FILLER_1_879 ();
 sg13g2_fill_2 FILLER_1_922 ();
 sg13g2_fill_1 FILLER_1_924 ();
 sg13g2_fill_2 FILLER_1_955 ();
 sg13g2_decap_4 FILLER_1_978 ();
 sg13g2_fill_2 FILLER_1_982 ();
 sg13g2_fill_2 FILLER_1_989 ();
 sg13g2_fill_1 FILLER_1_1029 ();
 sg13g2_decap_8 FILLER_1_1064 ();
 sg13g2_fill_2 FILLER_1_1097 ();
 sg13g2_fill_2 FILLER_1_1155 ();
 sg13g2_fill_1 FILLER_1_1157 ();
 sg13g2_fill_2 FILLER_1_1214 ();
 sg13g2_decap_4 FILLER_1_1226 ();
 sg13g2_fill_2 FILLER_1_1240 ();
 sg13g2_fill_1 FILLER_1_1242 ();
 sg13g2_decap_8 FILLER_1_1253 ();
 sg13g2_decap_8 FILLER_1_1260 ();
 sg13g2_decap_8 FILLER_1_1267 ();
 sg13g2_decap_8 FILLER_1_1284 ();
 sg13g2_fill_2 FILLER_1_1291 ();
 sg13g2_fill_1 FILLER_1_1293 ();
 sg13g2_fill_1 FILLER_1_1314 ();
 sg13g2_decap_4 FILLER_1_1341 ();
 sg13g2_fill_1 FILLER_1_1345 ();
 sg13g2_decap_8 FILLER_1_1376 ();
 sg13g2_decap_4 FILLER_1_1383 ();
 sg13g2_fill_1 FILLER_1_1387 ();
 sg13g2_decap_8 FILLER_1_1423 ();
 sg13g2_fill_2 FILLER_1_1430 ();
 sg13g2_fill_1 FILLER_1_1432 ();
 sg13g2_decap_8 FILLER_1_1458 ();
 sg13g2_fill_2 FILLER_1_1465 ();
 sg13g2_decap_8 FILLER_1_1471 ();
 sg13g2_fill_2 FILLER_1_1478 ();
 sg13g2_fill_1 FILLER_1_1480 ();
 sg13g2_fill_2 FILLER_1_1515 ();
 sg13g2_fill_2 FILLER_1_1553 ();
 sg13g2_fill_1 FILLER_1_1565 ();
 sg13g2_fill_2 FILLER_1_1592 ();
 sg13g2_decap_4 FILLER_1_1620 ();
 sg13g2_fill_1 FILLER_1_1624 ();
 sg13g2_fill_1 FILLER_1_1629 ();
 sg13g2_decap_4 FILLER_1_1656 ();
 sg13g2_fill_1 FILLER_1_1690 ();
 sg13g2_decap_8 FILLER_1_1727 ();
 sg13g2_fill_2 FILLER_1_1734 ();
 sg13g2_decap_8 FILLER_1_1797 ();
 sg13g2_decap_8 FILLER_1_1804 ();
 sg13g2_decap_8 FILLER_1_1811 ();
 sg13g2_fill_2 FILLER_1_1826 ();
 sg13g2_fill_1 FILLER_1_1828 ();
 sg13g2_fill_2 FILLER_1_1855 ();
 sg13g2_fill_1 FILLER_1_1857 ();
 sg13g2_decap_4 FILLER_1_1862 ();
 sg13g2_fill_2 FILLER_1_1912 ();
 sg13g2_fill_1 FILLER_1_1914 ();
 sg13g2_fill_2 FILLER_1_1941 ();
 sg13g2_fill_2 FILLER_1_1969 ();
 sg13g2_decap_4 FILLER_1_1991 ();
 sg13g2_decap_8 FILLER_1_2021 ();
 sg13g2_decap_4 FILLER_1_2028 ();
 sg13g2_fill_1 FILLER_1_2032 ();
 sg13g2_fill_1 FILLER_1_2059 ();
 sg13g2_fill_1 FILLER_1_2070 ();
 sg13g2_fill_2 FILLER_1_2081 ();
 sg13g2_fill_2 FILLER_1_2109 ();
 sg13g2_decap_8 FILLER_1_2151 ();
 sg13g2_fill_2 FILLER_1_2158 ();
 sg13g2_fill_1 FILLER_1_2170 ();
 sg13g2_decap_4 FILLER_1_2181 ();
 sg13g2_decap_8 FILLER_1_2211 ();
 sg13g2_fill_2 FILLER_1_2218 ();
 sg13g2_fill_1 FILLER_1_2220 ();
 sg13g2_decap_4 FILLER_1_2261 ();
 sg13g2_decap_4 FILLER_1_2337 ();
 sg13g2_fill_1 FILLER_1_2341 ();
 sg13g2_decap_8 FILLER_1_2352 ();
 sg13g2_decap_8 FILLER_1_2359 ();
 sg13g2_decap_8 FILLER_1_2366 ();
 sg13g2_decap_8 FILLER_1_2373 ();
 sg13g2_decap_8 FILLER_1_2380 ();
 sg13g2_decap_8 FILLER_1_2387 ();
 sg13g2_decap_8 FILLER_1_2394 ();
 sg13g2_decap_8 FILLER_1_2401 ();
 sg13g2_decap_8 FILLER_1_2408 ();
 sg13g2_decap_8 FILLER_1_2415 ();
 sg13g2_decap_8 FILLER_1_2422 ();
 sg13g2_decap_8 FILLER_1_2429 ();
 sg13g2_decap_8 FILLER_1_2436 ();
 sg13g2_decap_8 FILLER_1_2443 ();
 sg13g2_decap_8 FILLER_1_2450 ();
 sg13g2_decap_8 FILLER_1_2457 ();
 sg13g2_decap_8 FILLER_1_2464 ();
 sg13g2_decap_8 FILLER_1_2471 ();
 sg13g2_decap_8 FILLER_1_2478 ();
 sg13g2_decap_8 FILLER_1_2485 ();
 sg13g2_decap_8 FILLER_1_2492 ();
 sg13g2_decap_8 FILLER_1_2499 ();
 sg13g2_decap_8 FILLER_1_2506 ();
 sg13g2_decap_8 FILLER_1_2513 ();
 sg13g2_decap_8 FILLER_1_2520 ();
 sg13g2_decap_8 FILLER_1_2527 ();
 sg13g2_decap_8 FILLER_1_2534 ();
 sg13g2_decap_8 FILLER_1_2541 ();
 sg13g2_decap_8 FILLER_1_2548 ();
 sg13g2_decap_8 FILLER_1_2555 ();
 sg13g2_decap_8 FILLER_1_2562 ();
 sg13g2_decap_8 FILLER_1_2569 ();
 sg13g2_decap_8 FILLER_1_2576 ();
 sg13g2_decap_8 FILLER_1_2583 ();
 sg13g2_decap_8 FILLER_1_2590 ();
 sg13g2_decap_8 FILLER_1_2597 ();
 sg13g2_decap_8 FILLER_1_2604 ();
 sg13g2_decap_8 FILLER_1_2611 ();
 sg13g2_decap_8 FILLER_1_2618 ();
 sg13g2_decap_8 FILLER_1_2625 ();
 sg13g2_decap_8 FILLER_1_2632 ();
 sg13g2_decap_8 FILLER_1_2639 ();
 sg13g2_decap_8 FILLER_1_2646 ();
 sg13g2_decap_8 FILLER_1_2653 ();
 sg13g2_decap_8 FILLER_1_2660 ();
 sg13g2_fill_2 FILLER_1_2667 ();
 sg13g2_fill_1 FILLER_1_2669 ();
 sg13g2_fill_2 FILLER_2_0 ();
 sg13g2_fill_2 FILLER_2_48 ();
 sg13g2_fill_2 FILLER_2_81 ();
 sg13g2_fill_1 FILLER_2_83 ();
 sg13g2_fill_1 FILLER_2_89 ();
 sg13g2_fill_2 FILLER_2_95 ();
 sg13g2_fill_2 FILLER_2_101 ();
 sg13g2_fill_2 FILLER_2_107 ();
 sg13g2_fill_1 FILLER_2_109 ();
 sg13g2_decap_4 FILLER_2_136 ();
 sg13g2_fill_1 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_151 ();
 sg13g2_decap_8 FILLER_2_158 ();
 sg13g2_decap_8 FILLER_2_165 ();
 sg13g2_decap_8 FILLER_2_172 ();
 sg13g2_decap_8 FILLER_2_179 ();
 sg13g2_decap_8 FILLER_2_186 ();
 sg13g2_decap_4 FILLER_2_193 ();
 sg13g2_fill_1 FILLER_2_230 ();
 sg13g2_fill_1 FILLER_2_278 ();
 sg13g2_fill_1 FILLER_2_289 ();
 sg13g2_fill_1 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_366 ();
 sg13g2_decap_8 FILLER_2_373 ();
 sg13g2_fill_2 FILLER_2_413 ();
 sg13g2_fill_2 FILLER_2_445 ();
 sg13g2_fill_2 FILLER_2_478 ();
 sg13g2_fill_2 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_523 ();
 sg13g2_decap_4 FILLER_2_530 ();
 sg13g2_fill_1 FILLER_2_534 ();
 sg13g2_decap_4 FILLER_2_539 ();
 sg13g2_fill_1 FILLER_2_543 ();
 sg13g2_decap_4 FILLER_2_548 ();
 sg13g2_fill_1 FILLER_2_561 ();
 sg13g2_fill_1 FILLER_2_566 ();
 sg13g2_fill_1 FILLER_2_576 ();
 sg13g2_fill_2 FILLER_2_581 ();
 sg13g2_decap_4 FILLER_2_588 ();
 sg13g2_fill_1 FILLER_2_596 ();
 sg13g2_decap_4 FILLER_2_645 ();
 sg13g2_fill_2 FILLER_2_685 ();
 sg13g2_fill_2 FILLER_2_723 ();
 sg13g2_decap_4 FILLER_2_751 ();
 sg13g2_fill_1 FILLER_2_755 ();
 sg13g2_fill_2 FILLER_2_786 ();
 sg13g2_fill_1 FILLER_2_788 ();
 sg13g2_fill_1 FILLER_2_836 ();
 sg13g2_fill_1 FILLER_2_863 ();
 sg13g2_fill_1 FILLER_2_895 ();
 sg13g2_fill_1 FILLER_2_974 ();
 sg13g2_fill_1 FILLER_2_1001 ();
 sg13g2_fill_1 FILLER_2_1006 ();
 sg13g2_fill_1 FILLER_2_1033 ();
 sg13g2_fill_1 FILLER_2_1065 ();
 sg13g2_fill_1 FILLER_2_1139 ();
 sg13g2_fill_1 FILLER_2_1180 ();
 sg13g2_decap_8 FILLER_2_1211 ();
 sg13g2_fill_2 FILLER_2_1218 ();
 sg13g2_decap_4 FILLER_2_1343 ();
 sg13g2_fill_2 FILLER_2_1347 ();
 sg13g2_fill_2 FILLER_2_1385 ();
 sg13g2_fill_2 FILLER_2_1424 ();
 sg13g2_fill_2 FILLER_2_1432 ();
 sg13g2_fill_2 FILLER_2_1518 ();
 sg13g2_fill_1 FILLER_2_1520 ();
 sg13g2_fill_1 FILLER_2_1547 ();
 sg13g2_fill_1 FILLER_2_1587 ();
 sg13g2_decap_4 FILLER_2_1654 ();
 sg13g2_fill_2 FILLER_2_1705 ();
 sg13g2_fill_1 FILLER_2_1707 ();
 sg13g2_decap_8 FILLER_2_1734 ();
 sg13g2_fill_2 FILLER_2_1741 ();
 sg13g2_fill_2 FILLER_2_1812 ();
 sg13g2_decap_4 FILLER_2_1858 ();
 sg13g2_fill_2 FILLER_2_1862 ();
 sg13g2_decap_8 FILLER_2_1930 ();
 sg13g2_fill_2 FILLER_2_1937 ();
 sg13g2_fill_1 FILLER_2_1939 ();
 sg13g2_decap_8 FILLER_2_2013 ();
 sg13g2_decap_4 FILLER_2_2020 ();
 sg13g2_fill_1 FILLER_2_2024 ();
 sg13g2_fill_1 FILLER_2_2107 ();
 sg13g2_fill_2 FILLER_2_2134 ();
 sg13g2_fill_1 FILLER_2_2136 ();
 sg13g2_fill_1 FILLER_2_2215 ();
 sg13g2_decap_4 FILLER_2_2256 ();
 sg13g2_fill_2 FILLER_2_2277 ();
 sg13g2_decap_8 FILLER_2_2378 ();
 sg13g2_decap_8 FILLER_2_2385 ();
 sg13g2_decap_8 FILLER_2_2392 ();
 sg13g2_decap_8 FILLER_2_2399 ();
 sg13g2_decap_8 FILLER_2_2406 ();
 sg13g2_decap_8 FILLER_2_2413 ();
 sg13g2_decap_8 FILLER_2_2420 ();
 sg13g2_decap_8 FILLER_2_2427 ();
 sg13g2_decap_8 FILLER_2_2434 ();
 sg13g2_decap_8 FILLER_2_2441 ();
 sg13g2_decap_8 FILLER_2_2448 ();
 sg13g2_decap_8 FILLER_2_2455 ();
 sg13g2_decap_8 FILLER_2_2462 ();
 sg13g2_decap_8 FILLER_2_2469 ();
 sg13g2_decap_8 FILLER_2_2476 ();
 sg13g2_decap_8 FILLER_2_2483 ();
 sg13g2_decap_8 FILLER_2_2490 ();
 sg13g2_decap_8 FILLER_2_2497 ();
 sg13g2_decap_8 FILLER_2_2504 ();
 sg13g2_decap_8 FILLER_2_2511 ();
 sg13g2_decap_8 FILLER_2_2518 ();
 sg13g2_decap_8 FILLER_2_2525 ();
 sg13g2_decap_8 FILLER_2_2532 ();
 sg13g2_decap_8 FILLER_2_2539 ();
 sg13g2_decap_8 FILLER_2_2546 ();
 sg13g2_decap_8 FILLER_2_2553 ();
 sg13g2_decap_8 FILLER_2_2560 ();
 sg13g2_decap_8 FILLER_2_2567 ();
 sg13g2_decap_8 FILLER_2_2574 ();
 sg13g2_decap_8 FILLER_2_2581 ();
 sg13g2_decap_8 FILLER_2_2588 ();
 sg13g2_decap_8 FILLER_2_2595 ();
 sg13g2_decap_8 FILLER_2_2602 ();
 sg13g2_decap_8 FILLER_2_2609 ();
 sg13g2_decap_8 FILLER_2_2616 ();
 sg13g2_decap_8 FILLER_2_2623 ();
 sg13g2_decap_8 FILLER_2_2630 ();
 sg13g2_decap_8 FILLER_2_2637 ();
 sg13g2_decap_8 FILLER_2_2644 ();
 sg13g2_decap_8 FILLER_2_2651 ();
 sg13g2_decap_8 FILLER_2_2658 ();
 sg13g2_decap_4 FILLER_2_2665 ();
 sg13g2_fill_1 FILLER_2_2669 ();
 sg13g2_fill_2 FILLER_3_0 ();
 sg13g2_fill_2 FILLER_3_53 ();
 sg13g2_fill_1 FILLER_3_81 ();
 sg13g2_fill_2 FILLER_3_94 ();
 sg13g2_decap_4 FILLER_3_100 ();
 sg13g2_fill_2 FILLER_3_104 ();
 sg13g2_fill_1 FILLER_3_116 ();
 sg13g2_fill_1 FILLER_3_121 ();
 sg13g2_decap_8 FILLER_3_132 ();
 sg13g2_fill_2 FILLER_3_139 ();
 sg13g2_decap_8 FILLER_3_171 ();
 sg13g2_decap_8 FILLER_3_178 ();
 sg13g2_decap_8 FILLER_3_185 ();
 sg13g2_fill_2 FILLER_3_192 ();
 sg13g2_fill_2 FILLER_3_207 ();
 sg13g2_fill_1 FILLER_3_214 ();
 sg13g2_fill_1 FILLER_3_234 ();
 sg13g2_fill_2 FILLER_3_240 ();
 sg13g2_fill_2 FILLER_3_275 ();
 sg13g2_fill_1 FILLER_3_301 ();
 sg13g2_fill_1 FILLER_3_305 ();
 sg13g2_fill_2 FILLER_3_420 ();
 sg13g2_fill_1 FILLER_3_426 ();
 sg13g2_fill_2 FILLER_3_432 ();
 sg13g2_fill_2 FILLER_3_449 ();
 sg13g2_decap_4 FILLER_3_477 ();
 sg13g2_fill_1 FILLER_3_486 ();
 sg13g2_fill_2 FILLER_3_566 ();
 sg13g2_decap_4 FILLER_3_592 ();
 sg13g2_fill_2 FILLER_3_596 ();
 sg13g2_decap_4 FILLER_3_671 ();
 sg13g2_fill_2 FILLER_3_675 ();
 sg13g2_fill_2 FILLER_3_687 ();
 sg13g2_fill_1 FILLER_3_732 ();
 sg13g2_fill_1 FILLER_3_750 ();
 sg13g2_fill_1 FILLER_3_811 ();
 sg13g2_fill_1 FILLER_3_838 ();
 sg13g2_decap_8 FILLER_3_864 ();
 sg13g2_fill_2 FILLER_3_875 ();
 sg13g2_fill_2 FILLER_3_881 ();
 sg13g2_fill_1 FILLER_3_883 ();
 sg13g2_fill_1 FILLER_3_893 ();
 sg13g2_decap_8 FILLER_3_920 ();
 sg13g2_fill_1 FILLER_3_927 ();
 sg13g2_fill_1 FILLER_3_932 ();
 sg13g2_fill_1 FILLER_3_938 ();
 sg13g2_fill_2 FILLER_3_948 ();
 sg13g2_fill_1 FILLER_3_950 ();
 sg13g2_fill_1 FILLER_3_959 ();
 sg13g2_fill_1 FILLER_3_1037 ();
 sg13g2_fill_2 FILLER_3_1089 ();
 sg13g2_fill_2 FILLER_3_1127 ();
 sg13g2_fill_2 FILLER_3_1169 ();
 sg13g2_fill_1 FILLER_3_1171 ();
 sg13g2_fill_2 FILLER_3_1265 ();
 sg13g2_fill_1 FILLER_3_1271 ();
 sg13g2_fill_2 FILLER_3_1298 ();
 sg13g2_fill_1 FILLER_3_1326 ();
 sg13g2_fill_2 FILLER_3_1331 ();
 sg13g2_decap_8 FILLER_3_1337 ();
 sg13g2_decap_4 FILLER_3_1344 ();
 sg13g2_fill_2 FILLER_3_1348 ();
 sg13g2_fill_1 FILLER_3_1354 ();
 sg13g2_fill_1 FILLER_3_1363 ();
 sg13g2_fill_1 FILLER_3_1368 ();
 sg13g2_fill_2 FILLER_3_1374 ();
 sg13g2_fill_1 FILLER_3_1376 ();
 sg13g2_fill_1 FILLER_3_1434 ();
 sg13g2_fill_1 FILLER_3_1439 ();
 sg13g2_fill_2 FILLER_3_1450 ();
 sg13g2_fill_1 FILLER_3_1462 ();
 sg13g2_decap_8 FILLER_3_1473 ();
 sg13g2_fill_1 FILLER_3_1480 ();
 sg13g2_fill_2 FILLER_3_1487 ();
 sg13g2_fill_1 FILLER_3_1489 ();
 sg13g2_fill_2 FILLER_3_1496 ();
 sg13g2_fill_1 FILLER_3_1498 ();
 sg13g2_fill_1 FILLER_3_1576 ();
 sg13g2_decap_8 FILLER_3_1581 ();
 sg13g2_decap_8 FILLER_3_1588 ();
 sg13g2_fill_2 FILLER_3_1595 ();
 sg13g2_fill_1 FILLER_3_1597 ();
 sg13g2_decap_4 FILLER_3_1628 ();
 sg13g2_fill_2 FILLER_3_1708 ();
 sg13g2_fill_1 FILLER_3_1710 ();
 sg13g2_fill_1 FILLER_3_1737 ();
 sg13g2_fill_2 FILLER_3_1772 ();
 sg13g2_fill_1 FILLER_3_1774 ();
 sg13g2_fill_1 FILLER_3_1785 ();
 sg13g2_fill_1 FILLER_3_1812 ();
 sg13g2_fill_2 FILLER_3_1823 ();
 sg13g2_fill_1 FILLER_3_1833 ();
 sg13g2_decap_8 FILLER_3_1855 ();
 sg13g2_fill_1 FILLER_3_1909 ();
 sg13g2_fill_2 FILLER_3_1940 ();
 sg13g2_decap_4 FILLER_3_1982 ();
 sg13g2_fill_2 FILLER_3_1986 ();
 sg13g2_fill_1 FILLER_3_2024 ();
 sg13g2_fill_1 FILLER_3_2035 ();
 sg13g2_fill_2 FILLER_3_2040 ();
 sg13g2_fill_2 FILLER_3_2052 ();
 sg13g2_fill_1 FILLER_3_2107 ();
 sg13g2_decap_8 FILLER_3_2134 ();
 sg13g2_fill_2 FILLER_3_2141 ();
 sg13g2_fill_1 FILLER_3_2143 ();
 sg13g2_fill_1 FILLER_3_2154 ();
 sg13g2_fill_1 FILLER_3_2185 ();
 sg13g2_fill_2 FILLER_3_2216 ();
 sg13g2_fill_1 FILLER_3_2218 ();
 sg13g2_decap_8 FILLER_3_2249 ();
 sg13g2_fill_2 FILLER_3_2256 ();
 sg13g2_decap_4 FILLER_3_2268 ();
 sg13g2_fill_2 FILLER_3_2272 ();
 sg13g2_decap_8 FILLER_3_2278 ();
 sg13g2_fill_2 FILLER_3_2285 ();
 sg13g2_fill_1 FILLER_3_2287 ();
 sg13g2_decap_8 FILLER_3_2298 ();
 sg13g2_fill_1 FILLER_3_2305 ();
 sg13g2_fill_2 FILLER_3_2310 ();
 sg13g2_decap_8 FILLER_3_2316 ();
 sg13g2_decap_4 FILLER_3_2323 ();
 sg13g2_decap_8 FILLER_3_2378 ();
 sg13g2_decap_8 FILLER_3_2385 ();
 sg13g2_decap_8 FILLER_3_2392 ();
 sg13g2_decap_8 FILLER_3_2399 ();
 sg13g2_decap_8 FILLER_3_2406 ();
 sg13g2_decap_8 FILLER_3_2413 ();
 sg13g2_decap_8 FILLER_3_2420 ();
 sg13g2_decap_8 FILLER_3_2427 ();
 sg13g2_decap_8 FILLER_3_2434 ();
 sg13g2_decap_8 FILLER_3_2441 ();
 sg13g2_decap_8 FILLER_3_2448 ();
 sg13g2_decap_8 FILLER_3_2455 ();
 sg13g2_decap_8 FILLER_3_2462 ();
 sg13g2_decap_8 FILLER_3_2469 ();
 sg13g2_decap_8 FILLER_3_2476 ();
 sg13g2_decap_8 FILLER_3_2483 ();
 sg13g2_decap_8 FILLER_3_2490 ();
 sg13g2_decap_8 FILLER_3_2497 ();
 sg13g2_decap_8 FILLER_3_2504 ();
 sg13g2_decap_8 FILLER_3_2511 ();
 sg13g2_decap_8 FILLER_3_2518 ();
 sg13g2_decap_8 FILLER_3_2525 ();
 sg13g2_decap_8 FILLER_3_2532 ();
 sg13g2_decap_8 FILLER_3_2539 ();
 sg13g2_decap_8 FILLER_3_2546 ();
 sg13g2_decap_8 FILLER_3_2553 ();
 sg13g2_decap_8 FILLER_3_2560 ();
 sg13g2_decap_8 FILLER_3_2567 ();
 sg13g2_decap_8 FILLER_3_2574 ();
 sg13g2_decap_8 FILLER_3_2581 ();
 sg13g2_decap_8 FILLER_3_2588 ();
 sg13g2_decap_8 FILLER_3_2595 ();
 sg13g2_decap_8 FILLER_3_2602 ();
 sg13g2_decap_8 FILLER_3_2609 ();
 sg13g2_decap_8 FILLER_3_2616 ();
 sg13g2_decap_8 FILLER_3_2623 ();
 sg13g2_decap_8 FILLER_3_2630 ();
 sg13g2_decap_8 FILLER_3_2637 ();
 sg13g2_decap_8 FILLER_3_2644 ();
 sg13g2_decap_8 FILLER_3_2651 ();
 sg13g2_decap_8 FILLER_3_2658 ();
 sg13g2_decap_4 FILLER_3_2665 ();
 sg13g2_fill_1 FILLER_3_2669 ();
 sg13g2_fill_2 FILLER_4_0 ();
 sg13g2_fill_1 FILLER_4_6 ();
 sg13g2_fill_1 FILLER_4_17 ();
 sg13g2_fill_1 FILLER_4_44 ();
 sg13g2_fill_1 FILLER_4_81 ();
 sg13g2_fill_1 FILLER_4_112 ();
 sg13g2_fill_1 FILLER_4_139 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_fill_1 FILLER_4_182 ();
 sg13g2_fill_1 FILLER_4_209 ();
 sg13g2_fill_1 FILLER_4_225 ();
 sg13g2_decap_8 FILLER_4_348 ();
 sg13g2_decap_4 FILLER_4_355 ();
 sg13g2_fill_2 FILLER_4_359 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_4 FILLER_4_385 ();
 sg13g2_fill_1 FILLER_4_389 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_4_421 ();
 sg13g2_fill_2 FILLER_4_458 ();
 sg13g2_decap_8 FILLER_4_464 ();
 sg13g2_fill_1 FILLER_4_471 ();
 sg13g2_decap_4 FILLER_4_482 ();
 sg13g2_fill_2 FILLER_4_525 ();
 sg13g2_fill_1 FILLER_4_527 ();
 sg13g2_decap_4 FILLER_4_577 ();
 sg13g2_fill_2 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_587 ();
 sg13g2_decap_4 FILLER_4_594 ();
 sg13g2_fill_1 FILLER_4_598 ();
 sg13g2_fill_1 FILLER_4_620 ();
 sg13g2_decap_8 FILLER_4_641 ();
 sg13g2_fill_1 FILLER_4_688 ();
 sg13g2_fill_2 FILLER_4_703 ();
 sg13g2_fill_1 FILLER_4_713 ();
 sg13g2_fill_2 FILLER_4_719 ();
 sg13g2_fill_1 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_740 ();
 sg13g2_decap_8 FILLER_4_747 ();
 sg13g2_decap_4 FILLER_4_754 ();
 sg13g2_fill_2 FILLER_4_785 ();
 sg13g2_fill_1 FILLER_4_817 ();
 sg13g2_decap_4 FILLER_4_827 ();
 sg13g2_decap_4 FILLER_4_835 ();
 sg13g2_fill_2 FILLER_4_839 ();
 sg13g2_fill_1 FILLER_4_876 ();
 sg13g2_fill_1 FILLER_4_887 ();
 sg13g2_fill_1 FILLER_4_902 ();
 sg13g2_decap_8 FILLER_4_913 ();
 sg13g2_decap_8 FILLER_4_920 ();
 sg13g2_decap_8 FILLER_4_927 ();
 sg13g2_decap_8 FILLER_4_934 ();
 sg13g2_fill_2 FILLER_4_959 ();
 sg13g2_fill_2 FILLER_4_971 ();
 sg13g2_fill_1 FILLER_4_973 ();
 sg13g2_decap_4 FILLER_4_986 ();
 sg13g2_fill_1 FILLER_4_990 ();
 sg13g2_fill_2 FILLER_4_1005 ();
 sg13g2_fill_2 FILLER_4_1011 ();
 sg13g2_fill_2 FILLER_4_1022 ();
 sg13g2_fill_1 FILLER_4_1024 ();
 sg13g2_fill_2 FILLER_4_1046 ();
 sg13g2_fill_1 FILLER_4_1101 ();
 sg13g2_fill_2 FILLER_4_1110 ();
 sg13g2_fill_1 FILLER_4_1142 ();
 sg13g2_fill_1 FILLER_4_1148 ();
 sg13g2_fill_1 FILLER_4_1153 ();
 sg13g2_fill_1 FILLER_4_1158 ();
 sg13g2_fill_2 FILLER_4_1163 ();
 sg13g2_fill_1 FILLER_4_1165 ();
 sg13g2_fill_2 FILLER_4_1221 ();
 sg13g2_fill_2 FILLER_4_1227 ();
 sg13g2_fill_1 FILLER_4_1233 ();
 sg13g2_fill_2 FILLER_4_1238 ();
 sg13g2_decap_8 FILLER_4_1261 ();
 sg13g2_fill_1 FILLER_4_1268 ();
 sg13g2_decap_4 FILLER_4_1282 ();
 sg13g2_decap_8 FILLER_4_1322 ();
 sg13g2_decap_8 FILLER_4_1329 ();
 sg13g2_decap_8 FILLER_4_1336 ();
 sg13g2_decap_8 FILLER_4_1343 ();
 sg13g2_decap_4 FILLER_4_1350 ();
 sg13g2_decap_4 FILLER_4_1377 ();
 sg13g2_fill_2 FILLER_4_1428 ();
 sg13g2_fill_1 FILLER_4_1434 ();
 sg13g2_fill_1 FILLER_4_1461 ();
 sg13g2_fill_1 FILLER_4_1477 ();
 sg13g2_fill_1 FILLER_4_1487 ();
 sg13g2_fill_1 FILLER_4_1523 ();
 sg13g2_decap_8 FILLER_4_1536 ();
 sg13g2_decap_4 FILLER_4_1543 ();
 sg13g2_fill_1 FILLER_4_1547 ();
 sg13g2_decap_8 FILLER_4_1564 ();
 sg13g2_decap_8 FILLER_4_1571 ();
 sg13g2_decap_8 FILLER_4_1578 ();
 sg13g2_decap_8 FILLER_4_1585 ();
 sg13g2_decap_4 FILLER_4_1592 ();
 sg13g2_fill_2 FILLER_4_1600 ();
 sg13g2_fill_1 FILLER_4_1602 ();
 sg13g2_decap_4 FILLER_4_1607 ();
 sg13g2_fill_2 FILLER_4_1611 ();
 sg13g2_decap_4 FILLER_4_1655 ();
 sg13g2_fill_2 FILLER_4_1659 ();
 sg13g2_decap_4 FILLER_4_1671 ();
 sg13g2_fill_2 FILLER_4_1675 ();
 sg13g2_decap_8 FILLER_4_1681 ();
 sg13g2_decap_8 FILLER_4_1688 ();
 sg13g2_decap_8 FILLER_4_1695 ();
 sg13g2_decap_4 FILLER_4_1702 ();
 sg13g2_fill_2 FILLER_4_1716 ();
 sg13g2_fill_1 FILLER_4_1722 ();
 sg13g2_decap_8 FILLER_4_1727 ();
 sg13g2_decap_8 FILLER_4_1734 ();
 sg13g2_decap_4 FILLER_4_1741 ();
 sg13g2_fill_1 FILLER_4_1745 ();
 sg13g2_decap_8 FILLER_4_1760 ();
 sg13g2_fill_2 FILLER_4_1767 ();
 sg13g2_fill_1 FILLER_4_1769 ();
 sg13g2_fill_2 FILLER_4_1774 ();
 sg13g2_fill_1 FILLER_4_1776 ();
 sg13g2_fill_1 FILLER_4_1787 ();
 sg13g2_fill_1 FILLER_4_1792 ();
 sg13g2_fill_2 FILLER_4_1797 ();
 sg13g2_fill_1 FILLER_4_1817 ();
 sg13g2_fill_2 FILLER_4_1872 ();
 sg13g2_fill_1 FILLER_4_1874 ();
 sg13g2_fill_2 FILLER_4_1901 ();
 sg13g2_fill_1 FILLER_4_1903 ();
 sg13g2_fill_1 FILLER_4_2015 ();
 sg13g2_fill_1 FILLER_4_2029 ();
 sg13g2_fill_1 FILLER_4_2048 ();
 sg13g2_decap_8 FILLER_4_2057 ();
 sg13g2_decap_8 FILLER_4_2068 ();
 sg13g2_fill_2 FILLER_4_2085 ();
 sg13g2_fill_1 FILLER_4_2087 ();
 sg13g2_decap_8 FILLER_4_2129 ();
 sg13g2_fill_1 FILLER_4_2136 ();
 sg13g2_decap_4 FILLER_4_2147 ();
 sg13g2_fill_1 FILLER_4_2151 ();
 sg13g2_fill_1 FILLER_4_2209 ();
 sg13g2_decap_8 FILLER_4_2240 ();
 sg13g2_decap_4 FILLER_4_2247 ();
 sg13g2_fill_1 FILLER_4_2272 ();
 sg13g2_decap_8 FILLER_4_2309 ();
 sg13g2_decap_8 FILLER_4_2316 ();
 sg13g2_decap_8 FILLER_4_2323 ();
 sg13g2_decap_8 FILLER_4_2330 ();
 sg13g2_decap_8 FILLER_4_2337 ();
 sg13g2_fill_2 FILLER_4_2358 ();
 sg13g2_decap_8 FILLER_4_2368 ();
 sg13g2_decap_8 FILLER_4_2375 ();
 sg13g2_decap_8 FILLER_4_2382 ();
 sg13g2_decap_8 FILLER_4_2389 ();
 sg13g2_decap_8 FILLER_4_2396 ();
 sg13g2_decap_8 FILLER_4_2403 ();
 sg13g2_decap_8 FILLER_4_2410 ();
 sg13g2_decap_8 FILLER_4_2417 ();
 sg13g2_decap_8 FILLER_4_2424 ();
 sg13g2_decap_8 FILLER_4_2431 ();
 sg13g2_decap_8 FILLER_4_2438 ();
 sg13g2_decap_8 FILLER_4_2445 ();
 sg13g2_decap_8 FILLER_4_2452 ();
 sg13g2_decap_8 FILLER_4_2459 ();
 sg13g2_decap_8 FILLER_4_2466 ();
 sg13g2_decap_8 FILLER_4_2473 ();
 sg13g2_decap_8 FILLER_4_2480 ();
 sg13g2_decap_8 FILLER_4_2487 ();
 sg13g2_decap_8 FILLER_4_2494 ();
 sg13g2_decap_8 FILLER_4_2501 ();
 sg13g2_decap_8 FILLER_4_2508 ();
 sg13g2_decap_8 FILLER_4_2515 ();
 sg13g2_decap_8 FILLER_4_2522 ();
 sg13g2_decap_8 FILLER_4_2529 ();
 sg13g2_decap_8 FILLER_4_2536 ();
 sg13g2_decap_8 FILLER_4_2543 ();
 sg13g2_decap_8 FILLER_4_2550 ();
 sg13g2_decap_8 FILLER_4_2557 ();
 sg13g2_decap_8 FILLER_4_2564 ();
 sg13g2_decap_8 FILLER_4_2571 ();
 sg13g2_decap_8 FILLER_4_2578 ();
 sg13g2_decap_8 FILLER_4_2585 ();
 sg13g2_decap_8 FILLER_4_2592 ();
 sg13g2_decap_8 FILLER_4_2599 ();
 sg13g2_decap_8 FILLER_4_2606 ();
 sg13g2_decap_8 FILLER_4_2613 ();
 sg13g2_decap_8 FILLER_4_2620 ();
 sg13g2_decap_8 FILLER_4_2627 ();
 sg13g2_decap_8 FILLER_4_2634 ();
 sg13g2_decap_8 FILLER_4_2641 ();
 sg13g2_decap_8 FILLER_4_2648 ();
 sg13g2_decap_8 FILLER_4_2655 ();
 sg13g2_decap_8 FILLER_4_2662 ();
 sg13g2_fill_1 FILLER_4_2669 ();
 sg13g2_decap_4 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_4 ();
 sg13g2_decap_4 FILLER_5_12 ();
 sg13g2_fill_1 FILLER_5_24 ();
 sg13g2_fill_1 FILLER_5_29 ();
 sg13g2_fill_2 FILLER_5_46 ();
 sg13g2_fill_1 FILLER_5_48 ();
 sg13g2_fill_2 FILLER_5_60 ();
 sg13g2_fill_1 FILLER_5_62 ();
 sg13g2_decap_8 FILLER_5_97 ();
 sg13g2_fill_2 FILLER_5_104 ();
 sg13g2_fill_2 FILLER_5_116 ();
 sg13g2_decap_8 FILLER_5_122 ();
 sg13g2_fill_2 FILLER_5_129 ();
 sg13g2_fill_1 FILLER_5_131 ();
 sg13g2_fill_2 FILLER_5_168 ();
 sg13g2_fill_1 FILLER_5_232 ();
 sg13g2_fill_1 FILLER_5_240 ();
 sg13g2_fill_1 FILLER_5_277 ();
 sg13g2_fill_2 FILLER_5_304 ();
 sg13g2_fill_1 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_347 ();
 sg13g2_decap_4 FILLER_5_354 ();
 sg13g2_fill_2 FILLER_5_358 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_4 FILLER_5_468 ();
 sg13g2_fill_2 FILLER_5_472 ();
 sg13g2_decap_8 FILLER_5_484 ();
 sg13g2_decap_4 FILLER_5_491 ();
 sg13g2_fill_2 FILLER_5_495 ();
 sg13g2_fill_2 FILLER_5_510 ();
 sg13g2_fill_1 FILLER_5_512 ();
 sg13g2_decap_4 FILLER_5_533 ();
 sg13g2_fill_1 FILLER_5_537 ();
 sg13g2_decap_4 FILLER_5_542 ();
 sg13g2_fill_2 FILLER_5_574 ();
 sg13g2_fill_1 FILLER_5_576 ();
 sg13g2_fill_2 FILLER_5_603 ();
 sg13g2_fill_2 FILLER_5_628 ();
 sg13g2_fill_1 FILLER_5_630 ();
 sg13g2_decap_4 FILLER_5_641 ();
 sg13g2_fill_1 FILLER_5_655 ();
 sg13g2_fill_1 FILLER_5_661 ();
 sg13g2_fill_1 FILLER_5_692 ();
 sg13g2_fill_1 FILLER_5_698 ();
 sg13g2_fill_2 FILLER_5_709 ();
 sg13g2_decap_8 FILLER_5_751 ();
 sg13g2_fill_1 FILLER_5_758 ();
 sg13g2_fill_2 FILLER_5_789 ();
 sg13g2_decap_8 FILLER_5_821 ();
 sg13g2_decap_8 FILLER_5_828 ();
 sg13g2_decap_8 FILLER_5_835 ();
 sg13g2_decap_4 FILLER_5_842 ();
 sg13g2_fill_2 FILLER_5_855 ();
 sg13g2_decap_4 FILLER_5_862 ();
 sg13g2_fill_1 FILLER_5_870 ();
 sg13g2_fill_1 FILLER_5_881 ();
 sg13g2_fill_1 FILLER_5_908 ();
 sg13g2_fill_1 FILLER_5_935 ();
 sg13g2_fill_1 FILLER_5_941 ();
 sg13g2_fill_1 FILLER_5_946 ();
 sg13g2_fill_2 FILLER_5_956 ();
 sg13g2_decap_4 FILLER_5_984 ();
 sg13g2_decap_8 FILLER_5_992 ();
 sg13g2_decap_8 FILLER_5_999 ();
 sg13g2_decap_8 FILLER_5_1006 ();
 sg13g2_decap_8 FILLER_5_1013 ();
 sg13g2_decap_4 FILLER_5_1020 ();
 sg13g2_fill_2 FILLER_5_1024 ();
 sg13g2_fill_2 FILLER_5_1061 ();
 sg13g2_fill_2 FILLER_5_1102 ();
 sg13g2_fill_1 FILLER_5_1104 ();
 sg13g2_fill_2 FILLER_5_1109 ();
 sg13g2_fill_1 FILLER_5_1111 ();
 sg13g2_decap_4 FILLER_5_1117 ();
 sg13g2_fill_1 FILLER_5_1121 ();
 sg13g2_decap_8 FILLER_5_1130 ();
 sg13g2_decap_4 FILLER_5_1137 ();
 sg13g2_decap_4 FILLER_5_1145 ();
 sg13g2_fill_1 FILLER_5_1149 ();
 sg13g2_decap_8 FILLER_5_1223 ();
 sg13g2_decap_8 FILLER_5_1230 ();
 sg13g2_decap_8 FILLER_5_1237 ();
 sg13g2_decap_8 FILLER_5_1244 ();
 sg13g2_decap_8 FILLER_5_1251 ();
 sg13g2_decap_4 FILLER_5_1294 ();
 sg13g2_decap_8 FILLER_5_1334 ();
 sg13g2_decap_4 FILLER_5_1341 ();
 sg13g2_fill_2 FILLER_5_1345 ();
 sg13g2_fill_2 FILLER_5_1377 ();
 sg13g2_fill_1 FILLER_5_1379 ();
 sg13g2_fill_1 FILLER_5_1403 ();
 sg13g2_fill_1 FILLER_5_1423 ();
 sg13g2_fill_2 FILLER_5_1442 ();
 sg13g2_fill_1 FILLER_5_1444 ();
 sg13g2_decap_4 FILLER_5_1477 ();
 sg13g2_decap_4 FILLER_5_1486 ();
 sg13g2_fill_1 FILLER_5_1490 ();
 sg13g2_decap_8 FILLER_5_1495 ();
 sg13g2_decap_4 FILLER_5_1502 ();
 sg13g2_fill_1 FILLER_5_1506 ();
 sg13g2_fill_1 FILLER_5_1519 ();
 sg13g2_fill_2 FILLER_5_1525 ();
 sg13g2_fill_1 FILLER_5_1527 ();
 sg13g2_fill_1 FILLER_5_1548 ();
 sg13g2_fill_2 FILLER_5_1553 ();
 sg13g2_decap_8 FILLER_5_1585 ();
 sg13g2_fill_2 FILLER_5_1626 ();
 sg13g2_fill_1 FILLER_5_1628 ();
 sg13g2_decap_4 FILLER_5_1659 ();
 sg13g2_fill_2 FILLER_5_1663 ();
 sg13g2_decap_4 FILLER_5_1679 ();
 sg13g2_fill_1 FILLER_5_1683 ();
 sg13g2_fill_1 FILLER_5_1737 ();
 sg13g2_decap_8 FILLER_5_1760 ();
 sg13g2_decap_8 FILLER_5_1767 ();
 sg13g2_fill_1 FILLER_5_1774 ();
 sg13g2_decap_4 FILLER_5_1811 ();
 sg13g2_decap_4 FILLER_5_1861 ();
 sg13g2_fill_1 FILLER_5_1865 ();
 sg13g2_decap_8 FILLER_5_1874 ();
 sg13g2_fill_2 FILLER_5_1881 ();
 sg13g2_decap_8 FILLER_5_1897 ();
 sg13g2_fill_1 FILLER_5_1904 ();
 sg13g2_decap_8 FILLER_5_1935 ();
 sg13g2_fill_2 FILLER_5_1942 ();
 sg13g2_fill_1 FILLER_5_1944 ();
 sg13g2_decap_4 FILLER_5_1981 ();
 sg13g2_fill_2 FILLER_5_2011 ();
 sg13g2_fill_2 FILLER_5_2033 ();
 sg13g2_fill_1 FILLER_5_2035 ();
 sg13g2_fill_2 FILLER_5_2062 ();
 sg13g2_fill_1 FILLER_5_2064 ();
 sg13g2_fill_1 FILLER_5_2105 ();
 sg13g2_decap_8 FILLER_5_2127 ();
 sg13g2_decap_8 FILLER_5_2168 ();
 sg13g2_fill_2 FILLER_5_2175 ();
 sg13g2_decap_8 FILLER_5_2211 ();
 sg13g2_decap_8 FILLER_5_2218 ();
 sg13g2_decap_4 FILLER_5_2225 ();
 sg13g2_fill_1 FILLER_5_2229 ();
 sg13g2_decap_4 FILLER_5_2270 ();
 sg13g2_fill_1 FILLER_5_2274 ();
 sg13g2_fill_2 FILLER_5_2301 ();
 sg13g2_fill_1 FILLER_5_2303 ();
 sg13g2_fill_2 FILLER_5_2330 ();
 sg13g2_fill_1 FILLER_5_2332 ();
 sg13g2_decap_8 FILLER_5_2373 ();
 sg13g2_decap_8 FILLER_5_2380 ();
 sg13g2_decap_8 FILLER_5_2387 ();
 sg13g2_decap_8 FILLER_5_2394 ();
 sg13g2_decap_8 FILLER_5_2401 ();
 sg13g2_decap_8 FILLER_5_2408 ();
 sg13g2_decap_8 FILLER_5_2415 ();
 sg13g2_decap_8 FILLER_5_2422 ();
 sg13g2_decap_8 FILLER_5_2429 ();
 sg13g2_decap_8 FILLER_5_2436 ();
 sg13g2_decap_8 FILLER_5_2443 ();
 sg13g2_decap_8 FILLER_5_2450 ();
 sg13g2_decap_8 FILLER_5_2457 ();
 sg13g2_decap_8 FILLER_5_2464 ();
 sg13g2_decap_8 FILLER_5_2471 ();
 sg13g2_decap_8 FILLER_5_2478 ();
 sg13g2_decap_8 FILLER_5_2485 ();
 sg13g2_decap_8 FILLER_5_2492 ();
 sg13g2_decap_8 FILLER_5_2499 ();
 sg13g2_decap_8 FILLER_5_2506 ();
 sg13g2_decap_8 FILLER_5_2513 ();
 sg13g2_decap_8 FILLER_5_2520 ();
 sg13g2_decap_8 FILLER_5_2527 ();
 sg13g2_decap_8 FILLER_5_2534 ();
 sg13g2_decap_8 FILLER_5_2541 ();
 sg13g2_decap_8 FILLER_5_2548 ();
 sg13g2_decap_8 FILLER_5_2555 ();
 sg13g2_decap_8 FILLER_5_2562 ();
 sg13g2_decap_8 FILLER_5_2569 ();
 sg13g2_decap_8 FILLER_5_2576 ();
 sg13g2_decap_8 FILLER_5_2583 ();
 sg13g2_decap_8 FILLER_5_2590 ();
 sg13g2_decap_8 FILLER_5_2597 ();
 sg13g2_decap_8 FILLER_5_2604 ();
 sg13g2_decap_8 FILLER_5_2611 ();
 sg13g2_decap_8 FILLER_5_2618 ();
 sg13g2_decap_8 FILLER_5_2625 ();
 sg13g2_decap_8 FILLER_5_2632 ();
 sg13g2_decap_8 FILLER_5_2639 ();
 sg13g2_decap_8 FILLER_5_2646 ();
 sg13g2_decap_8 FILLER_5_2653 ();
 sg13g2_decap_8 FILLER_5_2660 ();
 sg13g2_fill_2 FILLER_5_2667 ();
 sg13g2_fill_1 FILLER_5_2669 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_fill_2 FILLER_6_35 ();
 sg13g2_fill_1 FILLER_6_46 ();
 sg13g2_decap_8 FILLER_6_57 ();
 sg13g2_decap_8 FILLER_6_73 ();
 sg13g2_decap_4 FILLER_6_80 ();
 sg13g2_fill_1 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_89 ();
 sg13g2_decap_8 FILLER_6_96 ();
 sg13g2_decap_8 FILLER_6_103 ();
 sg13g2_decap_8 FILLER_6_110 ();
 sg13g2_decap_8 FILLER_6_117 ();
 sg13g2_decap_8 FILLER_6_124 ();
 sg13g2_fill_2 FILLER_6_131 ();
 sg13g2_fill_1 FILLER_6_133 ();
 sg13g2_fill_2 FILLER_6_138 ();
 sg13g2_fill_2 FILLER_6_242 ();
 sg13g2_fill_1 FILLER_6_249 ();
 sg13g2_fill_1 FILLER_6_335 ();
 sg13g2_decap_8 FILLER_6_340 ();
 sg13g2_decap_8 FILLER_6_347 ();
 sg13g2_decap_8 FILLER_6_354 ();
 sg13g2_decap_8 FILLER_6_361 ();
 sg13g2_decap_8 FILLER_6_415 ();
 sg13g2_fill_1 FILLER_6_422 ();
 sg13g2_fill_2 FILLER_6_469 ();
 sg13g2_decap_4 FILLER_6_492 ();
 sg13g2_fill_1 FILLER_6_496 ();
 sg13g2_fill_1 FILLER_6_520 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_4 FILLER_6_539 ();
 sg13g2_fill_1 FILLER_6_543 ();
 sg13g2_fill_1 FILLER_6_558 ();
 sg13g2_fill_1 FILLER_6_565 ();
 sg13g2_fill_1 FILLER_6_576 ();
 sg13g2_fill_2 FILLER_6_582 ();
 sg13g2_fill_1 FILLER_6_610 ();
 sg13g2_fill_2 FILLER_6_617 ();
 sg13g2_fill_1 FILLER_6_619 ();
 sg13g2_fill_2 FILLER_6_646 ();
 sg13g2_fill_1 FILLER_6_648 ();
 sg13g2_fill_1 FILLER_6_653 ();
 sg13g2_decap_8 FILLER_6_664 ();
 sg13g2_fill_2 FILLER_6_671 ();
 sg13g2_fill_1 FILLER_6_673 ();
 sg13g2_fill_2 FILLER_6_678 ();
 sg13g2_decap_4 FILLER_6_706 ();
 sg13g2_fill_2 FILLER_6_723 ();
 sg13g2_fill_1 FILLER_6_725 ();
 sg13g2_decap_4 FILLER_6_752 ();
 sg13g2_fill_1 FILLER_6_756 ();
 sg13g2_fill_1 FILLER_6_783 ();
 sg13g2_fill_2 FILLER_6_841 ();
 sg13g2_fill_2 FILLER_6_847 ();
 sg13g2_fill_2 FILLER_6_857 ();
 sg13g2_fill_1 FILLER_6_859 ();
 sg13g2_fill_2 FILLER_6_886 ();
 sg13g2_fill_1 FILLER_6_888 ();
 sg13g2_fill_1 FILLER_6_936 ();
 sg13g2_decap_8 FILLER_6_971 ();
 sg13g2_fill_1 FILLER_6_978 ();
 sg13g2_decap_8 FILLER_6_1022 ();
 sg13g2_decap_8 FILLER_6_1059 ();
 sg13g2_decap_4 FILLER_6_1066 ();
 sg13g2_fill_1 FILLER_6_1070 ();
 sg13g2_decap_8 FILLER_6_1080 ();
 sg13g2_decap_8 FILLER_6_1087 ();
 sg13g2_decap_8 FILLER_6_1094 ();
 sg13g2_decap_4 FILLER_6_1101 ();
 sg13g2_fill_2 FILLER_6_1105 ();
 sg13g2_fill_2 FILLER_6_1155 ();
 sg13g2_fill_2 FILLER_6_1193 ();
 sg13g2_fill_2 FILLER_6_1199 ();
 sg13g2_fill_1 FILLER_6_1205 ();
 sg13g2_fill_2 FILLER_6_1227 ();
 sg13g2_fill_2 FILLER_6_1233 ();
 sg13g2_decap_4 FILLER_6_1239 ();
 sg13g2_decap_4 FILLER_6_1264 ();
 sg13g2_fill_2 FILLER_6_1272 ();
 sg13g2_decap_8 FILLER_6_1278 ();
 sg13g2_fill_1 FILLER_6_1306 ();
 sg13g2_decap_4 FILLER_6_1311 ();
 sg13g2_decap_8 FILLER_6_1319 ();
 sg13g2_decap_8 FILLER_6_1326 ();
 sg13g2_decap_8 FILLER_6_1333 ();
 sg13g2_decap_8 FILLER_6_1340 ();
 sg13g2_decap_4 FILLER_6_1347 ();
 sg13g2_fill_1 FILLER_6_1351 ();
 sg13g2_fill_1 FILLER_6_1356 ();
 sg13g2_fill_1 FILLER_6_1388 ();
 sg13g2_fill_1 FILLER_6_1420 ();
 sg13g2_fill_2 FILLER_6_1447 ();
 sg13g2_fill_1 FILLER_6_1449 ();
 sg13g2_fill_2 FILLER_6_1456 ();
 sg13g2_decap_8 FILLER_6_1463 ();
 sg13g2_fill_2 FILLER_6_1511 ();
 sg13g2_fill_1 FILLER_6_1527 ();
 sg13g2_fill_1 FILLER_6_1554 ();
 sg13g2_fill_2 FILLER_6_1560 ();
 sg13g2_fill_2 FILLER_6_1566 ();
 sg13g2_fill_2 FILLER_6_1573 ();
 sg13g2_decap_8 FILLER_6_1580 ();
 sg13g2_decap_8 FILLER_6_1587 ();
 sg13g2_decap_8 FILLER_6_1594 ();
 sg13g2_fill_1 FILLER_6_1605 ();
 sg13g2_fill_1 FILLER_6_1616 ();
 sg13g2_fill_1 FILLER_6_1637 ();
 sg13g2_decap_4 FILLER_6_1659 ();
 sg13g2_fill_1 FILLER_6_1663 ();
 sg13g2_fill_1 FILLER_6_1695 ();
 sg13g2_fill_1 FILLER_6_1706 ();
 sg13g2_decap_4 FILLER_6_1728 ();
 sg13g2_fill_1 FILLER_6_1732 ();
 sg13g2_decap_4 FILLER_6_1769 ();
 sg13g2_fill_2 FILLER_6_1773 ();
 sg13g2_decap_4 FILLER_6_1815 ();
 sg13g2_fill_2 FILLER_6_1819 ();
 sg13g2_decap_8 FILLER_6_1869 ();
 sg13g2_fill_1 FILLER_6_1876 ();
 sg13g2_decap_8 FILLER_6_1891 ();
 sg13g2_decap_8 FILLER_6_1898 ();
 sg13g2_decap_8 FILLER_6_1905 ();
 sg13g2_decap_4 FILLER_6_1912 ();
 sg13g2_fill_1 FILLER_6_1916 ();
 sg13g2_fill_2 FILLER_6_1932 ();
 sg13g2_fill_1 FILLER_6_1934 ();
 sg13g2_decap_8 FILLER_6_1948 ();
 sg13g2_decap_8 FILLER_6_1955 ();
 sg13g2_decap_8 FILLER_6_1962 ();
 sg13g2_decap_8 FILLER_6_1969 ();
 sg13g2_fill_2 FILLER_6_1976 ();
 sg13g2_decap_4 FILLER_6_1995 ();
 sg13g2_fill_2 FILLER_6_1999 ();
 sg13g2_fill_2 FILLER_6_2014 ();
 sg13g2_fill_1 FILLER_6_2016 ();
 sg13g2_decap_4 FILLER_6_2043 ();
 sg13g2_fill_2 FILLER_6_2047 ();
 sg13g2_decap_4 FILLER_6_2070 ();
 sg13g2_decap_8 FILLER_6_2100 ();
 sg13g2_fill_1 FILLER_6_2107 ();
 sg13g2_decap_8 FILLER_6_2134 ();
 sg13g2_decap_8 FILLER_6_2141 ();
 sg13g2_fill_1 FILLER_6_2148 ();
 sg13g2_fill_1 FILLER_6_2185 ();
 sg13g2_decap_8 FILLER_6_2190 ();
 sg13g2_fill_2 FILLER_6_2197 ();
 sg13g2_decap_8 FILLER_6_2203 ();
 sg13g2_decap_8 FILLER_6_2210 ();
 sg13g2_decap_4 FILLER_6_2217 ();
 sg13g2_decap_4 FILLER_6_2275 ();
 sg13g2_fill_2 FILLER_6_2296 ();
 sg13g2_fill_1 FILLER_6_2298 ();
 sg13g2_decap_4 FILLER_6_2317 ();
 sg13g2_fill_2 FILLER_6_2321 ();
 sg13g2_fill_2 FILLER_6_2327 ();
 sg13g2_fill_1 FILLER_6_2329 ();
 sg13g2_decap_8 FILLER_6_2366 ();
 sg13g2_decap_8 FILLER_6_2373 ();
 sg13g2_decap_4 FILLER_6_2380 ();
 sg13g2_fill_2 FILLER_6_2384 ();
 sg13g2_decap_8 FILLER_6_2399 ();
 sg13g2_decap_8 FILLER_6_2406 ();
 sg13g2_decap_8 FILLER_6_2413 ();
 sg13g2_decap_8 FILLER_6_2420 ();
 sg13g2_decap_8 FILLER_6_2427 ();
 sg13g2_decap_8 FILLER_6_2434 ();
 sg13g2_decap_8 FILLER_6_2441 ();
 sg13g2_decap_8 FILLER_6_2448 ();
 sg13g2_decap_8 FILLER_6_2455 ();
 sg13g2_decap_8 FILLER_6_2462 ();
 sg13g2_decap_8 FILLER_6_2469 ();
 sg13g2_decap_8 FILLER_6_2476 ();
 sg13g2_decap_8 FILLER_6_2483 ();
 sg13g2_decap_8 FILLER_6_2490 ();
 sg13g2_decap_8 FILLER_6_2497 ();
 sg13g2_decap_8 FILLER_6_2504 ();
 sg13g2_decap_8 FILLER_6_2511 ();
 sg13g2_decap_8 FILLER_6_2518 ();
 sg13g2_decap_8 FILLER_6_2525 ();
 sg13g2_decap_8 FILLER_6_2532 ();
 sg13g2_decap_8 FILLER_6_2539 ();
 sg13g2_decap_8 FILLER_6_2546 ();
 sg13g2_decap_8 FILLER_6_2553 ();
 sg13g2_decap_8 FILLER_6_2560 ();
 sg13g2_decap_8 FILLER_6_2567 ();
 sg13g2_decap_8 FILLER_6_2574 ();
 sg13g2_decap_8 FILLER_6_2581 ();
 sg13g2_decap_8 FILLER_6_2588 ();
 sg13g2_decap_8 FILLER_6_2595 ();
 sg13g2_decap_8 FILLER_6_2602 ();
 sg13g2_decap_8 FILLER_6_2609 ();
 sg13g2_decap_8 FILLER_6_2616 ();
 sg13g2_decap_8 FILLER_6_2623 ();
 sg13g2_decap_8 FILLER_6_2630 ();
 sg13g2_decap_8 FILLER_6_2637 ();
 sg13g2_decap_8 FILLER_6_2644 ();
 sg13g2_decap_8 FILLER_6_2651 ();
 sg13g2_decap_8 FILLER_6_2658 ();
 sg13g2_decap_4 FILLER_6_2665 ();
 sg13g2_fill_1 FILLER_6_2669 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_4 FILLER_7_35 ();
 sg13g2_decap_4 FILLER_7_75 ();
 sg13g2_fill_2 FILLER_7_79 ();
 sg13g2_decap_8 FILLER_7_104 ();
 sg13g2_fill_2 FILLER_7_111 ();
 sg13g2_decap_8 FILLER_7_117 ();
 sg13g2_fill_2 FILLER_7_124 ();
 sg13g2_fill_1 FILLER_7_126 ();
 sg13g2_fill_2 FILLER_7_165 ();
 sg13g2_fill_2 FILLER_7_223 ();
 sg13g2_fill_2 FILLER_7_233 ();
 sg13g2_fill_1 FILLER_7_252 ();
 sg13g2_fill_1 FILLER_7_283 ();
 sg13g2_fill_2 FILLER_7_389 ();
 sg13g2_fill_2 FILLER_7_398 ();
 sg13g2_decap_8 FILLER_7_412 ();
 sg13g2_fill_2 FILLER_7_419 ();
 sg13g2_fill_1 FILLER_7_421 ();
 sg13g2_fill_1 FILLER_7_448 ();
 sg13g2_fill_2 FILLER_7_558 ();
 sg13g2_fill_1 FILLER_7_560 ();
 sg13g2_fill_2 FILLER_7_566 ();
 sg13g2_fill_1 FILLER_7_573 ();
 sg13g2_fill_1 FILLER_7_608 ();
 sg13g2_fill_2 FILLER_7_624 ();
 sg13g2_fill_1 FILLER_7_626 ();
 sg13g2_decap_8 FILLER_7_631 ();
 sg13g2_fill_1 FILLER_7_638 ();
 sg13g2_fill_2 FILLER_7_649 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_fill_2 FILLER_7_672 ();
 sg13g2_fill_1 FILLER_7_674 ();
 sg13g2_decap_8 FILLER_7_681 ();
 sg13g2_decap_4 FILLER_7_692 ();
 sg13g2_fill_2 FILLER_7_696 ();
 sg13g2_fill_1 FILLER_7_713 ();
 sg13g2_decap_8 FILLER_7_744 ();
 sg13g2_decap_8 FILLER_7_751 ();
 sg13g2_decap_4 FILLER_7_758 ();
 sg13g2_fill_2 FILLER_7_762 ();
 sg13g2_fill_1 FILLER_7_777 ();
 sg13g2_fill_2 FILLER_7_787 ();
 sg13g2_fill_2 FILLER_7_806 ();
 sg13g2_fill_2 FILLER_7_826 ();
 sg13g2_fill_2 FILLER_7_833 ();
 sg13g2_decap_4 FILLER_7_861 ();
 sg13g2_fill_2 FILLER_7_901 ();
 sg13g2_fill_2 FILLER_7_913 ();
 sg13g2_fill_1 FILLER_7_915 ();
 sg13g2_decap_8 FILLER_7_924 ();
 sg13g2_fill_1 FILLER_7_931 ();
 sg13g2_fill_1 FILLER_7_936 ();
 sg13g2_decap_4 FILLER_7_977 ();
 sg13g2_fill_2 FILLER_7_981 ();
 sg13g2_fill_2 FILLER_7_987 ();
 sg13g2_decap_8 FILLER_7_1024 ();
 sg13g2_fill_1 FILLER_7_1031 ();
 sg13g2_fill_2 FILLER_7_1037 ();
 sg13g2_decap_8 FILLER_7_1043 ();
 sg13g2_decap_4 FILLER_7_1050 ();
 sg13g2_decap_8 FILLER_7_1058 ();
 sg13g2_decap_8 FILLER_7_1065 ();
 sg13g2_decap_4 FILLER_7_1072 ();
 sg13g2_fill_2 FILLER_7_1076 ();
 sg13g2_decap_8 FILLER_7_1112 ();
 sg13g2_fill_1 FILLER_7_1119 ();
 sg13g2_fill_2 FILLER_7_1129 ();
 sg13g2_decap_8 FILLER_7_1161 ();
 sg13g2_decap_8 FILLER_7_1168 ();
 sg13g2_fill_2 FILLER_7_1175 ();
 sg13g2_fill_1 FILLER_7_1177 ();
 sg13g2_fill_2 FILLER_7_1222 ();
 sg13g2_fill_1 FILLER_7_1224 ();
 sg13g2_fill_2 FILLER_7_1251 ();
 sg13g2_fill_1 FILLER_7_1253 ();
 sg13g2_fill_2 FILLER_7_1290 ();
 sg13g2_decap_4 FILLER_7_1302 ();
 sg13g2_fill_1 FILLER_7_1306 ();
 sg13g2_decap_8 FILLER_7_1311 ();
 sg13g2_decap_8 FILLER_7_1322 ();
 sg13g2_decap_4 FILLER_7_1329 ();
 sg13g2_fill_2 FILLER_7_1333 ();
 sg13g2_decap_8 FILLER_7_1339 ();
 sg13g2_decap_8 FILLER_7_1393 ();
 sg13g2_decap_4 FILLER_7_1400 ();
 sg13g2_fill_2 FILLER_7_1404 ();
 sg13g2_fill_2 FILLER_7_1410 ();
 sg13g2_fill_1 FILLER_7_1412 ();
 sg13g2_fill_2 FILLER_7_1417 ();
 sg13g2_decap_4 FILLER_7_1427 ();
 sg13g2_fill_1 FILLER_7_1431 ();
 sg13g2_fill_1 FILLER_7_1435 ();
 sg13g2_decap_4 FILLER_7_1442 ();
 sg13g2_fill_1 FILLER_7_1446 ();
 sg13g2_decap_8 FILLER_7_1462 ();
 sg13g2_fill_2 FILLER_7_1469 ();
 sg13g2_decap_8 FILLER_7_1563 ();
 sg13g2_decap_8 FILLER_7_1570 ();
 sg13g2_decap_8 FILLER_7_1577 ();
 sg13g2_decap_4 FILLER_7_1584 ();
 sg13g2_fill_1 FILLER_7_1588 ();
 sg13g2_decap_8 FILLER_7_1623 ();
 sg13g2_decap_4 FILLER_7_1630 ();
 sg13g2_decap_4 FILLER_7_1664 ();
 sg13g2_fill_2 FILLER_7_1698 ();
 sg13g2_fill_1 FILLER_7_1700 ();
 sg13g2_decap_8 FILLER_7_1722 ();
 sg13g2_decap_8 FILLER_7_1729 ();
 sg13g2_fill_2 FILLER_7_1736 ();
 sg13g2_fill_1 FILLER_7_1815 ();
 sg13g2_fill_2 FILLER_7_1911 ();
 sg13g2_fill_1 FILLER_7_1913 ();
 sg13g2_decap_8 FILLER_7_1954 ();
 sg13g2_decap_8 FILLER_7_1974 ();
 sg13g2_decap_8 FILLER_7_1981 ();
 sg13g2_fill_1 FILLER_7_1988 ();
 sg13g2_decap_4 FILLER_7_2002 ();
 sg13g2_decap_4 FILLER_7_2076 ();
 sg13g2_fill_1 FILLER_7_2080 ();
 sg13g2_fill_1 FILLER_7_2085 ();
 sg13g2_decap_8 FILLER_7_2090 ();
 sg13g2_decap_4 FILLER_7_2097 ();
 sg13g2_decap_4 FILLER_7_2111 ();
 sg13g2_fill_2 FILLER_7_2115 ();
 sg13g2_decap_4 FILLER_7_2129 ();
 sg13g2_fill_2 FILLER_7_2181 ();
 sg13g2_decap_4 FILLER_7_2255 ();
 sg13g2_decap_8 FILLER_7_2306 ();
 sg13g2_fill_2 FILLER_7_2313 ();
 sg13g2_decap_8 FILLER_7_2381 ();
 sg13g2_decap_8 FILLER_7_2388 ();
 sg13g2_decap_8 FILLER_7_2395 ();
 sg13g2_decap_8 FILLER_7_2402 ();
 sg13g2_decap_8 FILLER_7_2409 ();
 sg13g2_decap_8 FILLER_7_2416 ();
 sg13g2_decap_8 FILLER_7_2423 ();
 sg13g2_decap_8 FILLER_7_2430 ();
 sg13g2_decap_8 FILLER_7_2437 ();
 sg13g2_decap_8 FILLER_7_2444 ();
 sg13g2_decap_8 FILLER_7_2451 ();
 sg13g2_decap_8 FILLER_7_2458 ();
 sg13g2_decap_8 FILLER_7_2465 ();
 sg13g2_decap_8 FILLER_7_2472 ();
 sg13g2_decap_8 FILLER_7_2479 ();
 sg13g2_decap_8 FILLER_7_2486 ();
 sg13g2_decap_8 FILLER_7_2493 ();
 sg13g2_decap_8 FILLER_7_2500 ();
 sg13g2_decap_8 FILLER_7_2507 ();
 sg13g2_decap_8 FILLER_7_2514 ();
 sg13g2_decap_8 FILLER_7_2521 ();
 sg13g2_decap_8 FILLER_7_2528 ();
 sg13g2_decap_8 FILLER_7_2535 ();
 sg13g2_decap_8 FILLER_7_2542 ();
 sg13g2_decap_8 FILLER_7_2549 ();
 sg13g2_decap_8 FILLER_7_2556 ();
 sg13g2_decap_8 FILLER_7_2563 ();
 sg13g2_decap_8 FILLER_7_2570 ();
 sg13g2_decap_8 FILLER_7_2577 ();
 sg13g2_decap_8 FILLER_7_2584 ();
 sg13g2_decap_8 FILLER_7_2591 ();
 sg13g2_decap_8 FILLER_7_2598 ();
 sg13g2_decap_8 FILLER_7_2605 ();
 sg13g2_decap_8 FILLER_7_2612 ();
 sg13g2_decap_8 FILLER_7_2619 ();
 sg13g2_decap_8 FILLER_7_2626 ();
 sg13g2_decap_8 FILLER_7_2633 ();
 sg13g2_decap_8 FILLER_7_2640 ();
 sg13g2_decap_8 FILLER_7_2647 ();
 sg13g2_decap_8 FILLER_7_2654 ();
 sg13g2_decap_8 FILLER_7_2661 ();
 sg13g2_fill_2 FILLER_7_2668 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_fill_2 FILLER_8_21 ();
 sg13g2_fill_1 FILLER_8_23 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_4 FILLER_8_42 ();
 sg13g2_fill_1 FILLER_8_102 ();
 sg13g2_fill_2 FILLER_8_113 ();
 sg13g2_fill_2 FILLER_8_145 ();
 sg13g2_fill_2 FILLER_8_173 ();
 sg13g2_fill_1 FILLER_8_227 ();
 sg13g2_fill_2 FILLER_8_243 ();
 sg13g2_fill_1 FILLER_8_287 ();
 sg13g2_fill_2 FILLER_8_304 ();
 sg13g2_fill_2 FILLER_8_314 ();
 sg13g2_fill_1 FILLER_8_389 ();
 sg13g2_decap_8 FILLER_8_410 ();
 sg13g2_fill_2 FILLER_8_417 ();
 sg13g2_fill_2 FILLER_8_432 ();
 sg13g2_fill_2 FILLER_8_444 ();
 sg13g2_decap_8 FILLER_8_461 ();
 sg13g2_fill_1 FILLER_8_468 ();
 sg13g2_decap_8 FILLER_8_473 ();
 sg13g2_fill_1 FILLER_8_480 ();
 sg13g2_fill_2 FILLER_8_487 ();
 sg13g2_fill_2 FILLER_8_509 ();
 sg13g2_decap_4 FILLER_8_535 ();
 sg13g2_fill_1 FILLER_8_539 ();
 sg13g2_fill_1 FILLER_8_544 ();
 sg13g2_fill_1 FILLER_8_550 ();
 sg13g2_fill_1 FILLER_8_557 ();
 sg13g2_decap_4 FILLER_8_562 ();
 sg13g2_decap_8 FILLER_8_576 ();
 sg13g2_fill_1 FILLER_8_583 ();
 sg13g2_decap_4 FILLER_8_588 ();
 sg13g2_fill_1 FILLER_8_592 ();
 sg13g2_decap_8 FILLER_8_597 ();
 sg13g2_decap_8 FILLER_8_604 ();
 sg13g2_decap_8 FILLER_8_611 ();
 sg13g2_fill_1 FILLER_8_618 ();
 sg13g2_fill_2 FILLER_8_633 ();
 sg13g2_decap_8 FILLER_8_641 ();
 sg13g2_fill_1 FILLER_8_648 ();
 sg13g2_decap_8 FILLER_8_674 ();
 sg13g2_decap_8 FILLER_8_681 ();
 sg13g2_decap_8 FILLER_8_688 ();
 sg13g2_fill_1 FILLER_8_695 ();
 sg13g2_decap_8 FILLER_8_722 ();
 sg13g2_fill_2 FILLER_8_729 ();
 sg13g2_fill_1 FILLER_8_731 ();
 sg13g2_decap_8 FILLER_8_762 ();
 sg13g2_decap_8 FILLER_8_769 ();
 sg13g2_fill_2 FILLER_8_776 ();
 sg13g2_fill_1 FILLER_8_778 ();
 sg13g2_fill_1 FILLER_8_784 ();
 sg13g2_fill_1 FILLER_8_801 ();
 sg13g2_fill_2 FILLER_8_807 ();
 sg13g2_fill_1 FILLER_8_809 ();
 sg13g2_fill_2 FILLER_8_815 ();
 sg13g2_fill_1 FILLER_8_817 ();
 sg13g2_fill_2 FILLER_8_848 ();
 sg13g2_fill_1 FILLER_8_850 ();
 sg13g2_decap_4 FILLER_8_855 ();
 sg13g2_fill_1 FILLER_8_859 ();
 sg13g2_decap_8 FILLER_8_919 ();
 sg13g2_decap_4 FILLER_8_926 ();
 sg13g2_fill_1 FILLER_8_930 ();
 sg13g2_decap_4 FILLER_8_961 ();
 sg13g2_decap_4 FILLER_8_1034 ();
 sg13g2_fill_1 FILLER_8_1064 ();
 sg13g2_decap_4 FILLER_8_1069 ();
 sg13g2_fill_2 FILLER_8_1073 ();
 sg13g2_fill_2 FILLER_8_1088 ();
 sg13g2_fill_1 FILLER_8_1090 ();
 sg13g2_fill_2 FILLER_8_1126 ();
 sg13g2_fill_2 FILLER_8_1168 ();
 sg13g2_fill_1 FILLER_8_1219 ();
 sg13g2_decap_4 FILLER_8_1246 ();
 sg13g2_fill_1 FILLER_8_1250 ();
 sg13g2_fill_2 FILLER_8_1338 ();
 sg13g2_decap_4 FILLER_8_1348 ();
 sg13g2_fill_1 FILLER_8_1356 ();
 sg13g2_fill_2 FILLER_8_1369 ();
 sg13g2_decap_8 FILLER_8_1392 ();
 sg13g2_fill_2 FILLER_8_1399 ();
 sg13g2_fill_1 FILLER_8_1401 ();
 sg13g2_fill_1 FILLER_8_1419 ();
 sg13g2_fill_1 FILLER_8_1441 ();
 sg13g2_fill_1 FILLER_8_1503 ();
 sg13g2_fill_2 FILLER_8_1542 ();
 sg13g2_decap_8 FILLER_8_1576 ();
 sg13g2_fill_2 FILLER_8_1583 ();
 sg13g2_fill_1 FILLER_8_1585 ();
 sg13g2_fill_1 FILLER_8_1626 ();
 sg13g2_fill_2 FILLER_8_1676 ();
 sg13g2_fill_1 FILLER_8_1678 ();
 sg13g2_fill_2 FILLER_8_1683 ();
 sg13g2_fill_2 FILLER_8_1711 ();
 sg13g2_decap_8 FILLER_8_1734 ();
 sg13g2_fill_1 FILLER_8_1741 ();
 sg13g2_fill_1 FILLER_8_1793 ();
 sg13g2_decap_8 FILLER_8_1798 ();
 sg13g2_fill_2 FILLER_8_1805 ();
 sg13g2_fill_1 FILLER_8_1902 ();
 sg13g2_fill_2 FILLER_8_1950 ();
 sg13g2_decap_4 FILLER_8_1978 ();
 sg13g2_fill_2 FILLER_8_1982 ();
 sg13g2_decap_8 FILLER_8_2002 ();
 sg13g2_fill_2 FILLER_8_2009 ();
 sg13g2_fill_1 FILLER_8_2011 ();
 sg13g2_fill_1 FILLER_8_2029 ();
 sg13g2_decap_8 FILLER_8_2034 ();
 sg13g2_fill_2 FILLER_8_2041 ();
 sg13g2_decap_8 FILLER_8_2069 ();
 sg13g2_decap_8 FILLER_8_2076 ();
 sg13g2_decap_4 FILLER_8_2083 ();
 sg13g2_fill_2 FILLER_8_2095 ();
 sg13g2_decap_8 FILLER_8_2174 ();
 sg13g2_fill_1 FILLER_8_2207 ();
 sg13g2_fill_1 FILLER_8_2218 ();
 sg13g2_fill_1 FILLER_8_2233 ();
 sg13g2_fill_1 FILLER_8_2260 ();
 sg13g2_decap_8 FILLER_8_2282 ();
 sg13g2_decap_8 FILLER_8_2289 ();
 sg13g2_fill_2 FILLER_8_2296 ();
 sg13g2_fill_1 FILLER_8_2298 ();
 sg13g2_decap_4 FILLER_8_2356 ();
 sg13g2_decap_8 FILLER_8_2364 ();
 sg13g2_decap_8 FILLER_8_2371 ();
 sg13g2_decap_8 FILLER_8_2378 ();
 sg13g2_decap_8 FILLER_8_2385 ();
 sg13g2_decap_8 FILLER_8_2392 ();
 sg13g2_decap_8 FILLER_8_2399 ();
 sg13g2_decap_8 FILLER_8_2406 ();
 sg13g2_decap_8 FILLER_8_2413 ();
 sg13g2_decap_8 FILLER_8_2420 ();
 sg13g2_decap_8 FILLER_8_2427 ();
 sg13g2_decap_8 FILLER_8_2434 ();
 sg13g2_decap_8 FILLER_8_2441 ();
 sg13g2_decap_8 FILLER_8_2448 ();
 sg13g2_decap_8 FILLER_8_2455 ();
 sg13g2_decap_8 FILLER_8_2462 ();
 sg13g2_decap_8 FILLER_8_2469 ();
 sg13g2_decap_8 FILLER_8_2476 ();
 sg13g2_decap_8 FILLER_8_2483 ();
 sg13g2_decap_8 FILLER_8_2490 ();
 sg13g2_decap_8 FILLER_8_2497 ();
 sg13g2_decap_8 FILLER_8_2504 ();
 sg13g2_decap_8 FILLER_8_2511 ();
 sg13g2_decap_8 FILLER_8_2518 ();
 sg13g2_decap_8 FILLER_8_2525 ();
 sg13g2_decap_8 FILLER_8_2532 ();
 sg13g2_decap_8 FILLER_8_2539 ();
 sg13g2_decap_8 FILLER_8_2546 ();
 sg13g2_decap_8 FILLER_8_2553 ();
 sg13g2_decap_8 FILLER_8_2560 ();
 sg13g2_decap_8 FILLER_8_2567 ();
 sg13g2_decap_8 FILLER_8_2574 ();
 sg13g2_decap_8 FILLER_8_2581 ();
 sg13g2_decap_8 FILLER_8_2588 ();
 sg13g2_decap_8 FILLER_8_2595 ();
 sg13g2_decap_8 FILLER_8_2602 ();
 sg13g2_decap_8 FILLER_8_2609 ();
 sg13g2_decap_8 FILLER_8_2616 ();
 sg13g2_decap_8 FILLER_8_2623 ();
 sg13g2_decap_8 FILLER_8_2630 ();
 sg13g2_decap_8 FILLER_8_2637 ();
 sg13g2_decap_8 FILLER_8_2644 ();
 sg13g2_decap_8 FILLER_8_2651 ();
 sg13g2_decap_8 FILLER_8_2658 ();
 sg13g2_decap_4 FILLER_8_2665 ();
 sg13g2_fill_1 FILLER_8_2669 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_47 ();
 sg13g2_fill_1 FILLER_9_54 ();
 sg13g2_fill_2 FILLER_9_99 ();
 sg13g2_fill_1 FILLER_9_101 ();
 sg13g2_fill_2 FILLER_9_128 ();
 sg13g2_fill_1 FILLER_9_130 ();
 sg13g2_fill_1 FILLER_9_167 ();
 sg13g2_fill_1 FILLER_9_175 ();
 sg13g2_fill_1 FILLER_9_230 ();
 sg13g2_fill_1 FILLER_9_267 ();
 sg13g2_fill_1 FILLER_9_305 ();
 sg13g2_fill_2 FILLER_9_317 ();
 sg13g2_fill_2 FILLER_9_353 ();
 sg13g2_fill_1 FILLER_9_369 ();
 sg13g2_fill_1 FILLER_9_374 ();
 sg13g2_fill_1 FILLER_9_389 ();
 sg13g2_decap_8 FILLER_9_409 ();
 sg13g2_fill_2 FILLER_9_416 ();
 sg13g2_fill_1 FILLER_9_448 ();
 sg13g2_fill_2 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_fill_1 FILLER_9_490 ();
 sg13g2_fill_1 FILLER_9_556 ();
 sg13g2_decap_4 FILLER_9_561 ();
 sg13g2_fill_1 FILLER_9_565 ();
 sg13g2_fill_1 FILLER_9_570 ();
 sg13g2_fill_1 FILLER_9_580 ();
 sg13g2_decap_8 FILLER_9_585 ();
 sg13g2_fill_2 FILLER_9_592 ();
 sg13g2_decap_8 FILLER_9_599 ();
 sg13g2_decap_4 FILLER_9_606 ();
 sg13g2_fill_1 FILLER_9_610 ();
 sg13g2_fill_1 FILLER_9_615 ();
 sg13g2_fill_2 FILLER_9_625 ();
 sg13g2_decap_8 FILLER_9_677 ();
 sg13g2_decap_8 FILLER_9_684 ();
 sg13g2_decap_4 FILLER_9_691 ();
 sg13g2_decap_4 FILLER_9_703 ();
 sg13g2_fill_1 FILLER_9_712 ();
 sg13g2_fill_2 FILLER_9_717 ();
 sg13g2_fill_1 FILLER_9_734 ();
 sg13g2_decap_4 FILLER_9_739 ();
 sg13g2_decap_8 FILLER_9_747 ();
 sg13g2_decap_8 FILLER_9_754 ();
 sg13g2_decap_4 FILLER_9_761 ();
 sg13g2_fill_2 FILLER_9_765 ();
 sg13g2_fill_2 FILLER_9_845 ();
 sg13g2_fill_1 FILLER_9_847 ();
 sg13g2_fill_2 FILLER_9_853 ();
 sg13g2_decap_8 FILLER_9_902 ();
 sg13g2_decap_8 FILLER_9_943 ();
 sg13g2_decap_8 FILLER_9_950 ();
 sg13g2_fill_2 FILLER_9_957 ();
 sg13g2_fill_1 FILLER_9_959 ();
 sg13g2_fill_2 FILLER_9_986 ();
 sg13g2_fill_1 FILLER_9_988 ();
 sg13g2_fill_2 FILLER_9_1036 ();
 sg13g2_decap_8 FILLER_9_1077 ();
 sg13g2_fill_1 FILLER_9_1097 ();
 sg13g2_decap_4 FILLER_9_1129 ();
 sg13g2_fill_1 FILLER_9_1133 ();
 sg13g2_decap_4 FILLER_9_1138 ();
 sg13g2_fill_1 FILLER_9_1151 ();
 sg13g2_fill_1 FILLER_9_1178 ();
 sg13g2_fill_1 FILLER_9_1188 ();
 sg13g2_fill_1 FILLER_9_1193 ();
 sg13g2_decap_4 FILLER_9_1220 ();
 sg13g2_fill_1 FILLER_9_1224 ();
 sg13g2_fill_1 FILLER_9_1291 ();
 sg13g2_decap_4 FILLER_9_1328 ();
 sg13g2_fill_1 FILLER_9_1332 ();
 sg13g2_decap_8 FILLER_9_1346 ();
 sg13g2_decap_8 FILLER_9_1353 ();
 sg13g2_fill_2 FILLER_9_1360 ();
 sg13g2_fill_1 FILLER_9_1362 ();
 sg13g2_fill_2 FILLER_9_1367 ();
 sg13g2_decap_8 FILLER_9_1373 ();
 sg13g2_decap_8 FILLER_9_1380 ();
 sg13g2_decap_4 FILLER_9_1387 ();
 sg13g2_fill_2 FILLER_9_1399 ();
 sg13g2_fill_1 FILLER_9_1401 ();
 sg13g2_fill_1 FILLER_9_1406 ();
 sg13g2_decap_4 FILLER_9_1432 ();
 sg13g2_decap_4 FILLER_9_1469 ();
 sg13g2_fill_2 FILLER_9_1491 ();
 sg13g2_fill_1 FILLER_9_1549 ();
 sg13g2_decap_4 FILLER_9_1576 ();
 sg13g2_fill_1 FILLER_9_1580 ();
 sg13g2_fill_2 FILLER_9_1598 ();
 sg13g2_fill_1 FILLER_9_1600 ();
 sg13g2_fill_2 FILLER_9_1609 ();
 sg13g2_fill_1 FILLER_9_1621 ();
 sg13g2_decap_4 FILLER_9_1630 ();
 sg13g2_decap_8 FILLER_9_1648 ();
 sg13g2_decap_8 FILLER_9_1655 ();
 sg13g2_decap_4 FILLER_9_1662 ();
 sg13g2_fill_2 FILLER_9_1666 ();
 sg13g2_fill_1 FILLER_9_1678 ();
 sg13g2_decap_4 FILLER_9_1771 ();
 sg13g2_fill_1 FILLER_9_1775 ();
 sg13g2_decap_8 FILLER_9_1780 ();
 sg13g2_fill_2 FILLER_9_1787 ();
 sg13g2_decap_4 FILLER_9_1810 ();
 sg13g2_decap_8 FILLER_9_1892 ();
 sg13g2_fill_2 FILLER_9_1899 ();
 sg13g2_fill_1 FILLER_9_1916 ();
 sg13g2_decap_4 FILLER_9_1942 ();
 sg13g2_fill_1 FILLER_9_1946 ();
 sg13g2_decap_8 FILLER_9_1974 ();
 sg13g2_decap_4 FILLER_9_1981 ();
 sg13g2_fill_1 FILLER_9_1985 ();
 sg13g2_fill_2 FILLER_9_2033 ();
 sg13g2_fill_1 FILLER_9_2035 ();
 sg13g2_fill_2 FILLER_9_2051 ();
 sg13g2_fill_1 FILLER_9_2053 ();
 sg13g2_fill_2 FILLER_9_2063 ();
 sg13g2_fill_1 FILLER_9_2101 ();
 sg13g2_fill_1 FILLER_9_2125 ();
 sg13g2_decap_8 FILLER_9_2147 ();
 sg13g2_decap_4 FILLER_9_2158 ();
 sg13g2_fill_1 FILLER_9_2183 ();
 sg13g2_decap_4 FILLER_9_2193 ();
 sg13g2_fill_2 FILLER_9_2197 ();
 sg13g2_decap_4 FILLER_9_2203 ();
 sg13g2_fill_1 FILLER_9_2207 ();
 sg13g2_fill_2 FILLER_9_2239 ();
 sg13g2_decap_8 FILLER_9_2262 ();
 sg13g2_decap_8 FILLER_9_2269 ();
 sg13g2_decap_4 FILLER_9_2276 ();
 sg13g2_decap_4 FILLER_9_2320 ();
 sg13g2_fill_2 FILLER_9_2324 ();
 sg13g2_fill_1 FILLER_9_2336 ();
 sg13g2_fill_2 FILLER_9_2358 ();
 sg13g2_fill_1 FILLER_9_2360 ();
 sg13g2_decap_8 FILLER_9_2387 ();
 sg13g2_decap_8 FILLER_9_2394 ();
 sg13g2_decap_8 FILLER_9_2401 ();
 sg13g2_decap_8 FILLER_9_2408 ();
 sg13g2_decap_8 FILLER_9_2415 ();
 sg13g2_fill_1 FILLER_9_2422 ();
 sg13g2_decap_8 FILLER_9_2427 ();
 sg13g2_decap_8 FILLER_9_2434 ();
 sg13g2_decap_8 FILLER_9_2441 ();
 sg13g2_decap_8 FILLER_9_2448 ();
 sg13g2_decap_8 FILLER_9_2455 ();
 sg13g2_decap_8 FILLER_9_2462 ();
 sg13g2_decap_8 FILLER_9_2469 ();
 sg13g2_decap_8 FILLER_9_2476 ();
 sg13g2_decap_8 FILLER_9_2483 ();
 sg13g2_decap_8 FILLER_9_2490 ();
 sg13g2_decap_8 FILLER_9_2497 ();
 sg13g2_decap_8 FILLER_9_2504 ();
 sg13g2_decap_8 FILLER_9_2511 ();
 sg13g2_decap_8 FILLER_9_2518 ();
 sg13g2_decap_8 FILLER_9_2525 ();
 sg13g2_decap_8 FILLER_9_2532 ();
 sg13g2_decap_8 FILLER_9_2539 ();
 sg13g2_decap_8 FILLER_9_2546 ();
 sg13g2_decap_8 FILLER_9_2553 ();
 sg13g2_decap_8 FILLER_9_2560 ();
 sg13g2_decap_8 FILLER_9_2567 ();
 sg13g2_decap_8 FILLER_9_2574 ();
 sg13g2_decap_8 FILLER_9_2581 ();
 sg13g2_decap_8 FILLER_9_2588 ();
 sg13g2_decap_8 FILLER_9_2595 ();
 sg13g2_decap_8 FILLER_9_2602 ();
 sg13g2_decap_8 FILLER_9_2609 ();
 sg13g2_decap_8 FILLER_9_2616 ();
 sg13g2_decap_8 FILLER_9_2623 ();
 sg13g2_decap_8 FILLER_9_2630 ();
 sg13g2_decap_8 FILLER_9_2637 ();
 sg13g2_decap_8 FILLER_9_2644 ();
 sg13g2_decap_8 FILLER_9_2651 ();
 sg13g2_decap_8 FILLER_9_2658 ();
 sg13g2_decap_4 FILLER_9_2665 ();
 sg13g2_fill_1 FILLER_9_2669 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_4 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_34 ();
 sg13g2_decap_8 FILLER_10_41 ();
 sg13g2_decap_4 FILLER_10_48 ();
 sg13g2_fill_2 FILLER_10_52 ();
 sg13g2_fill_1 FILLER_10_118 ();
 sg13g2_fill_1 FILLER_10_192 ();
 sg13g2_fill_2 FILLER_10_280 ();
 sg13g2_fill_2 FILLER_10_293 ();
 sg13g2_fill_1 FILLER_10_354 ();
 sg13g2_fill_1 FILLER_10_361 ();
 sg13g2_fill_2 FILLER_10_368 ();
 sg13g2_fill_2 FILLER_10_396 ();
 sg13g2_decap_4 FILLER_10_424 ();
 sg13g2_fill_2 FILLER_10_463 ();
 sg13g2_fill_1 FILLER_10_465 ();
 sg13g2_decap_8 FILLER_10_502 ();
 sg13g2_decap_8 FILLER_10_509 ();
 sg13g2_decap_4 FILLER_10_516 ();
 sg13g2_decap_8 FILLER_10_524 ();
 sg13g2_decap_4 FILLER_10_531 ();
 sg13g2_decap_4 FILLER_10_541 ();
 sg13g2_fill_2 FILLER_10_545 ();
 sg13g2_fill_2 FILLER_10_604 ();
 sg13g2_fill_1 FILLER_10_616 ();
 sg13g2_fill_2 FILLER_10_643 ();
 sg13g2_fill_1 FILLER_10_713 ();
 sg13g2_fill_2 FILLER_10_753 ();
 sg13g2_decap_8 FILLER_10_759 ();
 sg13g2_decap_8 FILLER_10_766 ();
 sg13g2_fill_1 FILLER_10_825 ();
 sg13g2_decap_8 FILLER_10_830 ();
 sg13g2_fill_1 FILLER_10_837 ();
 sg13g2_fill_2 FILLER_10_859 ();
 sg13g2_fill_1 FILLER_10_861 ();
 sg13g2_decap_4 FILLER_10_880 ();
 sg13g2_decap_8 FILLER_10_888 ();
 sg13g2_decap_8 FILLER_10_895 ();
 sg13g2_decap_8 FILLER_10_902 ();
 sg13g2_fill_1 FILLER_10_923 ();
 sg13g2_decap_8 FILLER_10_950 ();
 sg13g2_decap_8 FILLER_10_957 ();
 sg13g2_fill_2 FILLER_10_964 ();
 sg13g2_decap_8 FILLER_10_979 ();
 sg13g2_decap_8 FILLER_10_986 ();
 sg13g2_decap_8 FILLER_10_993 ();
 sg13g2_fill_2 FILLER_10_1000 ();
 sg13g2_fill_1 FILLER_10_1006 ();
 sg13g2_fill_1 FILLER_10_1016 ();
 sg13g2_decap_8 FILLER_10_1030 ();
 sg13g2_fill_1 FILLER_10_1037 ();
 sg13g2_fill_1 FILLER_10_1082 ();
 sg13g2_decap_8 FILLER_10_1121 ();
 sg13g2_decap_8 FILLER_10_1128 ();
 sg13g2_decap_8 FILLER_10_1135 ();
 sg13g2_fill_2 FILLER_10_1156 ();
 sg13g2_fill_2 FILLER_10_1162 ();
 sg13g2_fill_2 FILLER_10_1185 ();
 sg13g2_fill_2 FILLER_10_1192 ();
 sg13g2_fill_1 FILLER_10_1194 ();
 sg13g2_fill_2 FILLER_10_1199 ();
 sg13g2_fill_1 FILLER_10_1201 ();
 sg13g2_fill_2 FILLER_10_1206 ();
 sg13g2_fill_1 FILLER_10_1208 ();
 sg13g2_decap_8 FILLER_10_1213 ();
 sg13g2_decap_4 FILLER_10_1220 ();
 sg13g2_fill_2 FILLER_10_1224 ();
 sg13g2_decap_8 FILLER_10_1236 ();
 sg13g2_decap_4 FILLER_10_1243 ();
 sg13g2_fill_1 FILLER_10_1261 ();
 sg13g2_decap_4 FILLER_10_1266 ();
 sg13g2_fill_1 FILLER_10_1270 ();
 sg13g2_fill_2 FILLER_10_1323 ();
 sg13g2_decap_8 FILLER_10_1329 ();
 sg13g2_decap_8 FILLER_10_1336 ();
 sg13g2_decap_8 FILLER_10_1343 ();
 sg13g2_fill_2 FILLER_10_1350 ();
 sg13g2_fill_1 FILLER_10_1382 ();
 sg13g2_decap_8 FILLER_10_1391 ();
 sg13g2_fill_2 FILLER_10_1402 ();
 sg13g2_fill_1 FILLER_10_1410 ();
 sg13g2_fill_1 FILLER_10_1416 ();
 sg13g2_fill_2 FILLER_10_1422 ();
 sg13g2_fill_2 FILLER_10_1429 ();
 sg13g2_fill_1 FILLER_10_1431 ();
 sg13g2_fill_1 FILLER_10_1455 ();
 sg13g2_fill_1 FILLER_10_1515 ();
 sg13g2_decap_4 FILLER_10_1529 ();
 sg13g2_decap_4 FILLER_10_1562 ();
 sg13g2_fill_1 FILLER_10_1566 ();
 sg13g2_fill_1 FILLER_10_1580 ();
 sg13g2_decap_4 FILLER_10_1586 ();
 sg13g2_fill_1 FILLER_10_1590 ();
 sg13g2_fill_2 FILLER_10_1595 ();
 sg13g2_fill_1 FILLER_10_1597 ();
 sg13g2_fill_2 FILLER_10_1607 ();
 sg13g2_decap_4 FILLER_10_1621 ();
 sg13g2_fill_2 FILLER_10_1635 ();
 sg13g2_fill_1 FILLER_10_1637 ();
 sg13g2_decap_8 FILLER_10_1648 ();
 sg13g2_decap_8 FILLER_10_1655 ();
 sg13g2_decap_8 FILLER_10_1662 ();
 sg13g2_decap_4 FILLER_10_1669 ();
 sg13g2_fill_1 FILLER_10_1673 ();
 sg13g2_decap_4 FILLER_10_1679 ();
 sg13g2_fill_1 FILLER_10_1683 ();
 sg13g2_fill_1 FILLER_10_1688 ();
 sg13g2_fill_2 FILLER_10_1697 ();
 sg13g2_decap_4 FILLER_10_1717 ();
 sg13g2_decap_8 FILLER_10_1725 ();
 sg13g2_decap_8 FILLER_10_1732 ();
 sg13g2_decap_8 FILLER_10_1739 ();
 sg13g2_decap_4 FILLER_10_1746 ();
 sg13g2_decap_8 FILLER_10_1754 ();
 sg13g2_decap_8 FILLER_10_1761 ();
 sg13g2_decap_8 FILLER_10_1768 ();
 sg13g2_decap_4 FILLER_10_1800 ();
 sg13g2_fill_1 FILLER_10_1804 ();
 sg13g2_decap_4 FILLER_10_1809 ();
 sg13g2_fill_2 FILLER_10_1813 ();
 sg13g2_fill_2 FILLER_10_1827 ();
 sg13g2_fill_1 FILLER_10_1865 ();
 sg13g2_decap_4 FILLER_10_1870 ();
 sg13g2_fill_2 FILLER_10_1955 ();
 sg13g2_fill_1 FILLER_10_1957 ();
 sg13g2_decap_8 FILLER_10_1966 ();
 sg13g2_decap_4 FILLER_10_1983 ();
 sg13g2_fill_1 FILLER_10_1987 ();
 sg13g2_fill_1 FILLER_10_2042 ();
 sg13g2_fill_1 FILLER_10_2047 ();
 sg13g2_fill_1 FILLER_10_2069 ();
 sg13g2_fill_1 FILLER_10_2096 ();
 sg13g2_decap_8 FILLER_10_2101 ();
 sg13g2_decap_4 FILLER_10_2160 ();
 sg13g2_decap_8 FILLER_10_2185 ();
 sg13g2_decap_4 FILLER_10_2192 ();
 sg13g2_fill_1 FILLER_10_2196 ();
 sg13g2_fill_2 FILLER_10_2233 ();
 sg13g2_fill_2 FILLER_10_2239 ();
 sg13g2_decap_8 FILLER_10_2251 ();
 sg13g2_decap_8 FILLER_10_2258 ();
 sg13g2_decap_8 FILLER_10_2265 ();
 sg13g2_decap_8 FILLER_10_2277 ();
 sg13g2_decap_8 FILLER_10_2284 ();
 sg13g2_decap_4 FILLER_10_2291 ();
 sg13g2_fill_1 FILLER_10_2295 ();
 sg13g2_decap_8 FILLER_10_2310 ();
 sg13g2_decap_8 FILLER_10_2317 ();
 sg13g2_decap_8 FILLER_10_2324 ();
 sg13g2_fill_2 FILLER_10_2331 ();
 sg13g2_decap_8 FILLER_10_2395 ();
 sg13g2_decap_8 FILLER_10_2402 ();
 sg13g2_decap_4 FILLER_10_2409 ();
 sg13g2_fill_1 FILLER_10_2413 ();
 sg13g2_decap_8 FILLER_10_2457 ();
 sg13g2_decap_4 FILLER_10_2464 ();
 sg13g2_decap_8 FILLER_10_2498 ();
 sg13g2_decap_8 FILLER_10_2505 ();
 sg13g2_decap_8 FILLER_10_2512 ();
 sg13g2_decap_8 FILLER_10_2519 ();
 sg13g2_decap_8 FILLER_10_2526 ();
 sg13g2_decap_8 FILLER_10_2533 ();
 sg13g2_decap_8 FILLER_10_2540 ();
 sg13g2_decap_8 FILLER_10_2547 ();
 sg13g2_decap_8 FILLER_10_2554 ();
 sg13g2_decap_8 FILLER_10_2561 ();
 sg13g2_decap_8 FILLER_10_2568 ();
 sg13g2_decap_8 FILLER_10_2575 ();
 sg13g2_decap_8 FILLER_10_2582 ();
 sg13g2_decap_8 FILLER_10_2589 ();
 sg13g2_decap_8 FILLER_10_2596 ();
 sg13g2_decap_8 FILLER_10_2603 ();
 sg13g2_decap_8 FILLER_10_2610 ();
 sg13g2_decap_8 FILLER_10_2617 ();
 sg13g2_decap_8 FILLER_10_2624 ();
 sg13g2_decap_8 FILLER_10_2631 ();
 sg13g2_decap_8 FILLER_10_2638 ();
 sg13g2_decap_8 FILLER_10_2645 ();
 sg13g2_decap_8 FILLER_10_2652 ();
 sg13g2_decap_8 FILLER_10_2659 ();
 sg13g2_decap_4 FILLER_10_2666 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_41 ();
 sg13g2_fill_1 FILLER_11_73 ();
 sg13g2_fill_2 FILLER_11_146 ();
 sg13g2_fill_1 FILLER_11_217 ();
 sg13g2_fill_1 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_fill_1 FILLER_11_287 ();
 sg13g2_fill_1 FILLER_11_304 ();
 sg13g2_fill_1 FILLER_11_313 ();
 sg13g2_fill_1 FILLER_11_328 ();
 sg13g2_fill_1 FILLER_11_382 ();
 sg13g2_fill_1 FILLER_11_390 ();
 sg13g2_fill_2 FILLER_11_395 ();
 sg13g2_fill_1 FILLER_11_403 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_fill_2 FILLER_11_443 ();
 sg13g2_fill_1 FILLER_11_458 ();
 sg13g2_fill_2 FILLER_11_482 ();
 sg13g2_decap_4 FILLER_11_510 ();
 sg13g2_fill_1 FILLER_11_514 ();
 sg13g2_fill_1 FILLER_11_547 ();
 sg13g2_fill_2 FILLER_11_586 ();
 sg13g2_fill_1 FILLER_11_619 ();
 sg13g2_fill_1 FILLER_11_624 ();
 sg13g2_fill_1 FILLER_11_641 ();
 sg13g2_fill_2 FILLER_11_656 ();
 sg13g2_fill_2 FILLER_11_672 ();
 sg13g2_fill_1 FILLER_11_678 ();
 sg13g2_fill_2 FILLER_11_683 ();
 sg13g2_fill_2 FILLER_11_726 ();
 sg13g2_fill_1 FILLER_11_728 ();
 sg13g2_fill_2 FILLER_11_734 ();
 sg13g2_decap_4 FILLER_11_762 ();
 sg13g2_decap_8 FILLER_11_826 ();
 sg13g2_decap_8 FILLER_11_833 ();
 sg13g2_decap_8 FILLER_11_840 ();
 sg13g2_decap_8 FILLER_11_847 ();
 sg13g2_fill_1 FILLER_11_858 ();
 sg13g2_fill_2 FILLER_11_869 ();
 sg13g2_decap_8 FILLER_11_875 ();
 sg13g2_decap_4 FILLER_11_882 ();
 sg13g2_decap_8 FILLER_11_901 ();
 sg13g2_fill_2 FILLER_11_908 ();
 sg13g2_decap_4 FILLER_11_960 ();
 sg13g2_decap_8 FILLER_11_968 ();
 sg13g2_decap_8 FILLER_11_975 ();
 sg13g2_decap_8 FILLER_11_982 ();
 sg13g2_fill_2 FILLER_11_1010 ();
 sg13g2_fill_1 FILLER_11_1042 ();
 sg13g2_fill_1 FILLER_11_1053 ();
 sg13g2_fill_1 FILLER_11_1062 ();
 sg13g2_decap_8 FILLER_11_1088 ();
 sg13g2_fill_2 FILLER_11_1095 ();
 sg13g2_fill_1 FILLER_11_1097 ();
 sg13g2_decap_8 FILLER_11_1124 ();
 sg13g2_decap_8 FILLER_11_1131 ();
 sg13g2_decap_4 FILLER_11_1138 ();
 sg13g2_decap_8 FILLER_11_1171 ();
 sg13g2_decap_8 FILLER_11_1178 ();
 sg13g2_decap_4 FILLER_11_1216 ();
 sg13g2_decap_4 FILLER_11_1225 ();
 sg13g2_fill_2 FILLER_11_1229 ();
 sg13g2_decap_4 FILLER_11_1241 ();
 sg13g2_fill_1 FILLER_11_1245 ();
 sg13g2_decap_4 FILLER_11_1272 ();
 sg13g2_fill_1 FILLER_11_1276 ();
 sg13g2_fill_1 FILLER_11_1318 ();
 sg13g2_fill_1 FILLER_11_1345 ();
 sg13g2_fill_1 FILLER_11_1372 ();
 sg13g2_fill_1 FILLER_11_1416 ();
 sg13g2_decap_8 FILLER_11_1426 ();
 sg13g2_fill_1 FILLER_11_1433 ();
 sg13g2_decap_4 FILLER_11_1439 ();
 sg13g2_fill_1 FILLER_11_1443 ();
 sg13g2_fill_2 FILLER_11_1481 ();
 sg13g2_fill_1 FILLER_11_1487 ();
 sg13g2_decap_8 FILLER_11_1515 ();
 sg13g2_decap_8 FILLER_11_1522 ();
 sg13g2_decap_8 FILLER_11_1529 ();
 sg13g2_fill_2 FILLER_11_1563 ();
 sg13g2_fill_2 FILLER_11_1570 ();
 sg13g2_fill_1 FILLER_11_1572 ();
 sg13g2_fill_1 FILLER_11_1592 ();
 sg13g2_fill_1 FILLER_11_1597 ();
 sg13g2_fill_2 FILLER_11_1658 ();
 sg13g2_decap_4 FILLER_11_1706 ();
 sg13g2_fill_1 FILLER_11_1720 ();
 sg13g2_decap_8 FILLER_11_1725 ();
 sg13g2_decap_8 FILLER_11_1732 ();
 sg13g2_decap_8 FILLER_11_1739 ();
 sg13g2_decap_8 FILLER_11_1746 ();
 sg13g2_decap_4 FILLER_11_1753 ();
 sg13g2_decap_4 FILLER_11_1793 ();
 sg13g2_fill_2 FILLER_11_1801 ();
 sg13g2_decap_4 FILLER_11_1811 ();
 sg13g2_fill_2 FILLER_11_1815 ();
 sg13g2_decap_8 FILLER_11_1821 ();
 sg13g2_decap_8 FILLER_11_1828 ();
 sg13g2_decap_4 FILLER_11_1843 ();
 sg13g2_fill_1 FILLER_11_1847 ();
 sg13g2_fill_2 FILLER_11_1856 ();
 sg13g2_fill_1 FILLER_11_1876 ();
 sg13g2_fill_2 FILLER_11_1887 ();
 sg13g2_fill_2 FILLER_11_1897 ();
 sg13g2_fill_1 FILLER_11_1907 ();
 sg13g2_decap_8 FILLER_11_1916 ();
 sg13g2_fill_2 FILLER_11_1923 ();
 sg13g2_fill_1 FILLER_11_1935 ();
 sg13g2_decap_4 FILLER_11_1940 ();
 sg13g2_fill_2 FILLER_11_1944 ();
 sg13g2_decap_4 FILLER_11_1956 ();
 sg13g2_fill_2 FILLER_11_1960 ();
 sg13g2_decap_4 FILLER_11_1987 ();
 sg13g2_fill_2 FILLER_11_1991 ();
 sg13g2_decap_8 FILLER_11_1997 ();
 sg13g2_fill_1 FILLER_11_2004 ();
 sg13g2_fill_2 FILLER_11_2031 ();
 sg13g2_fill_1 FILLER_11_2059 ();
 sg13g2_decap_8 FILLER_11_2145 ();
 sg13g2_fill_2 FILLER_11_2152 ();
 sg13g2_fill_1 FILLER_11_2154 ();
 sg13g2_decap_8 FILLER_11_2176 ();
 sg13g2_decap_8 FILLER_11_2183 ();
 sg13g2_fill_2 FILLER_11_2190 ();
 sg13g2_fill_1 FILLER_11_2192 ();
 sg13g2_fill_1 FILLER_11_2228 ();
 sg13g2_fill_2 FILLER_11_2269 ();
 sg13g2_fill_1 FILLER_11_2271 ();
 sg13g2_fill_1 FILLER_11_2298 ();
 sg13g2_fill_1 FILLER_11_2303 ();
 sg13g2_fill_2 FILLER_11_2334 ();
 sg13g2_fill_1 FILLER_11_2336 ();
 sg13g2_decap_8 FILLER_11_2361 ();
 sg13g2_decap_4 FILLER_11_2372 ();
 sg13g2_decap_8 FILLER_11_2380 ();
 sg13g2_fill_1 FILLER_11_2387 ();
 sg13g2_decap_8 FILLER_11_2448 ();
 sg13g2_fill_1 FILLER_11_2455 ();
 sg13g2_decap_8 FILLER_11_2486 ();
 sg13g2_decap_8 FILLER_11_2493 ();
 sg13g2_decap_4 FILLER_11_2500 ();
 sg13g2_decap_8 FILLER_11_2534 ();
 sg13g2_decap_8 FILLER_11_2541 ();
 sg13g2_decap_8 FILLER_11_2548 ();
 sg13g2_decap_8 FILLER_11_2555 ();
 sg13g2_decap_8 FILLER_11_2562 ();
 sg13g2_decap_8 FILLER_11_2569 ();
 sg13g2_decap_8 FILLER_11_2576 ();
 sg13g2_decap_8 FILLER_11_2583 ();
 sg13g2_decap_8 FILLER_11_2590 ();
 sg13g2_decap_8 FILLER_11_2597 ();
 sg13g2_decap_8 FILLER_11_2604 ();
 sg13g2_decap_8 FILLER_11_2611 ();
 sg13g2_decap_8 FILLER_11_2618 ();
 sg13g2_decap_8 FILLER_11_2625 ();
 sg13g2_decap_8 FILLER_11_2632 ();
 sg13g2_decap_8 FILLER_11_2639 ();
 sg13g2_decap_8 FILLER_11_2646 ();
 sg13g2_decap_8 FILLER_11_2653 ();
 sg13g2_decap_8 FILLER_11_2660 ();
 sg13g2_fill_2 FILLER_11_2667 ();
 sg13g2_fill_1 FILLER_11_2669 ();
 sg13g2_fill_1 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_5 ();
 sg13g2_fill_1 FILLER_12_32 ();
 sg13g2_decap_4 FILLER_12_38 ();
 sg13g2_fill_1 FILLER_12_63 ();
 sg13g2_fill_1 FILLER_12_94 ();
 sg13g2_fill_1 FILLER_12_99 ();
 sg13g2_fill_1 FILLER_12_122 ();
 sg13g2_fill_2 FILLER_12_128 ();
 sg13g2_fill_2 FILLER_12_135 ();
 sg13g2_fill_2 FILLER_12_141 ();
 sg13g2_fill_2 FILLER_12_148 ();
 sg13g2_fill_2 FILLER_12_168 ();
 sg13g2_fill_1 FILLER_12_223 ();
 sg13g2_fill_1 FILLER_12_296 ();
 sg13g2_fill_1 FILLER_12_305 ();
 sg13g2_fill_2 FILLER_12_320 ();
 sg13g2_fill_1 FILLER_12_361 ();
 sg13g2_fill_1 FILLER_12_367 ();
 sg13g2_fill_1 FILLER_12_377 ();
 sg13g2_fill_1 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_12_425 ();
 sg13g2_decap_8 FILLER_12_432 ();
 sg13g2_fill_1 FILLER_12_443 ();
 sg13g2_fill_1 FILLER_12_478 ();
 sg13g2_fill_2 FILLER_12_493 ();
 sg13g2_fill_1 FILLER_12_495 ();
 sg13g2_fill_1 FILLER_12_502 ();
 sg13g2_decap_4 FILLER_12_538 ();
 sg13g2_fill_2 FILLER_12_542 ();
 sg13g2_fill_1 FILLER_12_554 ();
 sg13g2_fill_1 FILLER_12_565 ();
 sg13g2_fill_1 FILLER_12_585 ();
 sg13g2_fill_1 FILLER_12_596 ();
 sg13g2_fill_1 FILLER_12_609 ();
 sg13g2_fill_1 FILLER_12_615 ();
 sg13g2_decap_4 FILLER_12_657 ();
 sg13g2_decap_8 FILLER_12_670 ();
 sg13g2_decap_8 FILLER_12_677 ();
 sg13g2_fill_2 FILLER_12_684 ();
 sg13g2_fill_1 FILLER_12_686 ();
 sg13g2_fill_1 FILLER_12_715 ();
 sg13g2_fill_2 FILLER_12_739 ();
 sg13g2_fill_1 FILLER_12_741 ();
 sg13g2_decap_8 FILLER_12_768 ();
 sg13g2_fill_2 FILLER_12_775 ();
 sg13g2_fill_1 FILLER_12_777 ();
 sg13g2_decap_4 FILLER_12_782 ();
 sg13g2_decap_8 FILLER_12_790 ();
 sg13g2_decap_8 FILLER_12_797 ();
 sg13g2_decap_4 FILLER_12_804 ();
 sg13g2_fill_1 FILLER_12_808 ();
 sg13g2_decap_8 FILLER_12_818 ();
 sg13g2_decap_8 FILLER_12_825 ();
 sg13g2_fill_2 FILLER_12_832 ();
 sg13g2_fill_1 FILLER_12_834 ();
 sg13g2_decap_8 FILLER_12_875 ();
 sg13g2_fill_2 FILLER_12_882 ();
 sg13g2_fill_2 FILLER_12_954 ();
 sg13g2_fill_1 FILLER_12_956 ();
 sg13g2_fill_2 FILLER_12_1039 ();
 sg13g2_decap_8 FILLER_12_1045 ();
 sg13g2_fill_1 FILLER_12_1052 ();
 sg13g2_fill_2 FILLER_12_1118 ();
 sg13g2_decap_4 FILLER_12_1124 ();
 sg13g2_fill_1 FILLER_12_1128 ();
 sg13g2_decap_8 FILLER_12_1164 ();
 sg13g2_decap_8 FILLER_12_1171 ();
 sg13g2_decap_4 FILLER_12_1178 ();
 sg13g2_fill_2 FILLER_12_1187 ();
 sg13g2_fill_2 FILLER_12_1194 ();
 sg13g2_fill_1 FILLER_12_1196 ();
 sg13g2_fill_1 FILLER_12_1201 ();
 sg13g2_decap_4 FILLER_12_1228 ();
 sg13g2_decap_4 FILLER_12_1281 ();
 sg13g2_fill_1 FILLER_12_1285 ();
 sg13g2_decap_8 FILLER_12_1290 ();
 sg13g2_decap_4 FILLER_12_1297 ();
 sg13g2_fill_1 FILLER_12_1312 ();
 sg13g2_decap_8 FILLER_12_1317 ();
 sg13g2_decap_8 FILLER_12_1324 ();
 sg13g2_decap_8 FILLER_12_1331 ();
 sg13g2_fill_2 FILLER_12_1338 ();
 sg13g2_fill_1 FILLER_12_1340 ();
 sg13g2_fill_1 FILLER_12_1371 ();
 sg13g2_decap_8 FILLER_12_1388 ();
 sg13g2_decap_8 FILLER_12_1395 ();
 sg13g2_fill_2 FILLER_12_1402 ();
 sg13g2_fill_2 FILLER_12_1414 ();
 sg13g2_decap_4 FILLER_12_1429 ();
 sg13g2_fill_2 FILLER_12_1433 ();
 sg13g2_fill_2 FILLER_12_1453 ();
 sg13g2_fill_1 FILLER_12_1455 ();
 sg13g2_fill_1 FILLER_12_1505 ();
 sg13g2_fill_2 FILLER_12_1520 ();
 sg13g2_fill_1 FILLER_12_1522 ();
 sg13g2_fill_2 FILLER_12_1527 ();
 sg13g2_fill_1 FILLER_12_1540 ();
 sg13g2_decap_4 FILLER_12_1567 ();
 sg13g2_fill_1 FILLER_12_1571 ();
 sg13g2_fill_2 FILLER_12_1576 ();
 sg13g2_decap_4 FILLER_12_1663 ();
 sg13g2_decap_4 FILLER_12_1740 ();
 sg13g2_fill_2 FILLER_12_1744 ();
 sg13g2_fill_2 FILLER_12_1822 ();
 sg13g2_fill_1 FILLER_12_1824 ();
 sg13g2_fill_2 FILLER_12_1835 ();
 sg13g2_fill_1 FILLER_12_1837 ();
 sg13g2_fill_1 FILLER_12_1864 ();
 sg13g2_decap_4 FILLER_12_1895 ();
 sg13g2_fill_1 FILLER_12_1899 ();
 sg13g2_fill_2 FILLER_12_1926 ();
 sg13g2_fill_1 FILLER_12_1971 ();
 sg13g2_fill_2 FILLER_12_1998 ();
 sg13g2_fill_1 FILLER_12_2000 ();
 sg13g2_fill_2 FILLER_12_2009 ();
 sg13g2_fill_2 FILLER_12_2054 ();
 sg13g2_fill_1 FILLER_12_2056 ();
 sg13g2_fill_2 FILLER_12_2074 ();
 sg13g2_decap_8 FILLER_12_2102 ();
 sg13g2_fill_1 FILLER_12_2109 ();
 sg13g2_decap_8 FILLER_12_2114 ();
 sg13g2_decap_4 FILLER_12_2134 ();
 sg13g2_fill_1 FILLER_12_2138 ();
 sg13g2_fill_2 FILLER_12_2165 ();
 sg13g2_fill_1 FILLER_12_2167 ();
 sg13g2_fill_2 FILLER_12_2172 ();
 sg13g2_fill_1 FILLER_12_2230 ();
 sg13g2_fill_2 FILLER_12_2241 ();
 sg13g2_fill_1 FILLER_12_2310 ();
 sg13g2_decap_4 FILLER_12_2319 ();
 sg13g2_decap_8 FILLER_12_2349 ();
 sg13g2_decap_8 FILLER_12_2356 ();
 sg13g2_decap_8 FILLER_12_2363 ();
 sg13g2_decap_8 FILLER_12_2370 ();
 sg13g2_decap_4 FILLER_12_2377 ();
 sg13g2_decap_8 FILLER_12_2407 ();
 sg13g2_fill_1 FILLER_12_2414 ();
 sg13g2_fill_2 FILLER_12_2487 ();
 sg13g2_fill_1 FILLER_12_2489 ();
 sg13g2_fill_2 FILLER_12_2520 ();
 sg13g2_fill_1 FILLER_12_2522 ();
 sg13g2_decap_8 FILLER_12_2549 ();
 sg13g2_decap_8 FILLER_12_2556 ();
 sg13g2_decap_8 FILLER_12_2563 ();
 sg13g2_decap_8 FILLER_12_2570 ();
 sg13g2_decap_8 FILLER_12_2577 ();
 sg13g2_decap_8 FILLER_12_2584 ();
 sg13g2_decap_8 FILLER_12_2591 ();
 sg13g2_decap_8 FILLER_12_2598 ();
 sg13g2_decap_8 FILLER_12_2605 ();
 sg13g2_decap_8 FILLER_12_2612 ();
 sg13g2_decap_8 FILLER_12_2619 ();
 sg13g2_decap_8 FILLER_12_2626 ();
 sg13g2_decap_8 FILLER_12_2633 ();
 sg13g2_decap_8 FILLER_12_2640 ();
 sg13g2_decap_8 FILLER_12_2647 ();
 sg13g2_decap_8 FILLER_12_2654 ();
 sg13g2_decap_8 FILLER_12_2661 ();
 sg13g2_fill_2 FILLER_12_2668 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_7 ();
 sg13g2_fill_1 FILLER_13_9 ();
 sg13g2_fill_1 FILLER_13_85 ();
 sg13g2_fill_2 FILLER_13_99 ();
 sg13g2_fill_1 FILLER_13_132 ();
 sg13g2_fill_1 FILLER_13_141 ();
 sg13g2_fill_2 FILLER_13_146 ();
 sg13g2_fill_2 FILLER_13_160 ();
 sg13g2_fill_1 FILLER_13_169 ();
 sg13g2_fill_2 FILLER_13_182 ();
 sg13g2_fill_1 FILLER_13_187 ();
 sg13g2_fill_2 FILLER_13_219 ();
 sg13g2_fill_1 FILLER_13_226 ();
 sg13g2_fill_2 FILLER_13_239 ();
 sg13g2_fill_1 FILLER_13_267 ();
 sg13g2_decap_4 FILLER_13_278 ();
 sg13g2_fill_1 FILLER_13_282 ();
 sg13g2_fill_1 FILLER_13_313 ();
 sg13g2_fill_2 FILLER_13_354 ();
 sg13g2_fill_2 FILLER_13_365 ();
 sg13g2_fill_1 FILLER_13_393 ();
 sg13g2_decap_8 FILLER_13_432 ();
 sg13g2_decap_4 FILLER_13_439 ();
 sg13g2_fill_2 FILLER_13_443 ();
 sg13g2_fill_1 FILLER_13_455 ();
 sg13g2_fill_1 FILLER_13_460 ();
 sg13g2_fill_1 FILLER_13_465 ();
 sg13g2_fill_2 FILLER_13_471 ();
 sg13g2_decap_8 FILLER_13_477 ();
 sg13g2_fill_2 FILLER_13_489 ();
 sg13g2_fill_1 FILLER_13_491 ();
 sg13g2_fill_2 FILLER_13_496 ();
 sg13g2_fill_2 FILLER_13_518 ();
 sg13g2_fill_2 FILLER_13_550 ();
 sg13g2_fill_2 FILLER_13_584 ();
 sg13g2_fill_2 FILLER_13_591 ();
 sg13g2_fill_1 FILLER_13_610 ();
 sg13g2_fill_2 FILLER_13_626 ();
 sg13g2_fill_1 FILLER_13_632 ();
 sg13g2_fill_2 FILLER_13_637 ();
 sg13g2_decap_4 FILLER_13_649 ();
 sg13g2_fill_2 FILLER_13_653 ();
 sg13g2_fill_2 FILLER_13_659 ();
 sg13g2_fill_1 FILLER_13_667 ();
 sg13g2_fill_1 FILLER_13_672 ();
 sg13g2_fill_1 FILLER_13_677 ();
 sg13g2_fill_1 FILLER_13_682 ();
 sg13g2_decap_8 FILLER_13_693 ();
 sg13g2_fill_2 FILLER_13_700 ();
 sg13g2_fill_2 FILLER_13_713 ();
 sg13g2_fill_1 FILLER_13_719 ();
 sg13g2_decap_4 FILLER_13_734 ();
 sg13g2_fill_1 FILLER_13_742 ();
 sg13g2_decap_8 FILLER_13_760 ();
 sg13g2_decap_8 FILLER_13_767 ();
 sg13g2_decap_8 FILLER_13_774 ();
 sg13g2_decap_8 FILLER_13_781 ();
 sg13g2_decap_4 FILLER_13_788 ();
 sg13g2_fill_2 FILLER_13_792 ();
 sg13g2_fill_1 FILLER_13_820 ();
 sg13g2_fill_1 FILLER_13_825 ();
 sg13g2_fill_2 FILLER_13_906 ();
 sg13g2_fill_2 FILLER_13_912 ();
 sg13g2_fill_1 FILLER_13_914 ();
 sg13g2_fill_1 FILLER_13_944 ();
 sg13g2_fill_2 FILLER_13_1003 ();
 sg13g2_decap_4 FILLER_13_1009 ();
 sg13g2_fill_1 FILLER_13_1013 ();
 sg13g2_decap_4 FILLER_13_1053 ();
 sg13g2_fill_1 FILLER_13_1057 ();
 sg13g2_fill_2 FILLER_13_1074 ();
 sg13g2_decap_8 FILLER_13_1080 ();
 sg13g2_fill_2 FILLER_13_1087 ();
 sg13g2_fill_2 FILLER_13_1093 ();
 sg13g2_fill_1 FILLER_13_1104 ();
 sg13g2_fill_1 FILLER_13_1131 ();
 sg13g2_fill_2 FILLER_13_1177 ();
 sg13g2_fill_1 FILLER_13_1183 ();
 sg13g2_fill_2 FILLER_13_1214 ();
 sg13g2_fill_1 FILLER_13_1216 ();
 sg13g2_fill_2 FILLER_13_1221 ();
 sg13g2_fill_2 FILLER_13_1249 ();
 sg13g2_fill_2 FILLER_13_1261 ();
 sg13g2_fill_1 FILLER_13_1263 ();
 sg13g2_decap_8 FILLER_13_1294 ();
 sg13g2_decap_8 FILLER_13_1322 ();
 sg13g2_decap_8 FILLER_13_1329 ();
 sg13g2_decap_8 FILLER_13_1336 ();
 sg13g2_decap_4 FILLER_13_1343 ();
 sg13g2_fill_2 FILLER_13_1347 ();
 sg13g2_fill_1 FILLER_13_1361 ();
 sg13g2_fill_2 FILLER_13_1366 ();
 sg13g2_decap_4 FILLER_13_1384 ();
 sg13g2_fill_1 FILLER_13_1393 ();
 sg13g2_fill_1 FILLER_13_1402 ();
 sg13g2_fill_2 FILLER_13_1443 ();
 sg13g2_fill_1 FILLER_13_1445 ();
 sg13g2_fill_2 FILLER_13_1451 ();
 sg13g2_fill_1 FILLER_13_1472 ();
 sg13g2_fill_1 FILLER_13_1476 ();
 sg13g2_decap_8 FILLER_13_1569 ();
 sg13g2_fill_2 FILLER_13_1576 ();
 sg13g2_decap_8 FILLER_13_1587 ();
 sg13g2_fill_2 FILLER_13_1594 ();
 sg13g2_fill_2 FILLER_13_1600 ();
 sg13g2_fill_1 FILLER_13_1606 ();
 sg13g2_fill_1 FILLER_13_1612 ();
 sg13g2_fill_2 FILLER_13_1633 ();
 sg13g2_fill_1 FILLER_13_1635 ();
 sg13g2_decap_8 FILLER_13_1649 ();
 sg13g2_decap_8 FILLER_13_1656 ();
 sg13g2_decap_8 FILLER_13_1663 ();
 sg13g2_decap_4 FILLER_13_1670 ();
 sg13g2_fill_1 FILLER_13_1674 ();
 sg13g2_fill_2 FILLER_13_1679 ();
 sg13g2_decap_8 FILLER_13_1721 ();
 sg13g2_fill_2 FILLER_13_1728 ();
 sg13g2_fill_1 FILLER_13_1730 ();
 sg13g2_fill_2 FILLER_13_1769 ();
 sg13g2_fill_2 FILLER_13_1788 ();
 sg13g2_fill_1 FILLER_13_1790 ();
 sg13g2_fill_2 FILLER_13_1817 ();
 sg13g2_fill_1 FILLER_13_1854 ();
 sg13g2_fill_1 FILLER_13_1865 ();
 sg13g2_fill_2 FILLER_13_1936 ();
 sg13g2_decap_8 FILLER_13_1943 ();
 sg13g2_decap_8 FILLER_13_1950 ();
 sg13g2_fill_2 FILLER_13_1957 ();
 sg13g2_fill_1 FILLER_13_1959 ();
 sg13g2_decap_4 FILLER_13_1970 ();
 sg13g2_fill_2 FILLER_13_1974 ();
 sg13g2_decap_8 FILLER_13_1997 ();
 sg13g2_fill_2 FILLER_13_2004 ();
 sg13g2_fill_1 FILLER_13_2006 ();
 sg13g2_decap_4 FILLER_13_2017 ();
 sg13g2_fill_1 FILLER_13_2021 ();
 sg13g2_fill_2 FILLER_13_2026 ();
 sg13g2_fill_1 FILLER_13_2028 ();
 sg13g2_fill_1 FILLER_13_2050 ();
 sg13g2_decap_8 FILLER_13_2077 ();
 sg13g2_fill_2 FILLER_13_2084 ();
 sg13g2_decap_8 FILLER_13_2090 ();
 sg13g2_decap_8 FILLER_13_2189 ();
 sg13g2_decap_4 FILLER_13_2235 ();
 sg13g2_fill_2 FILLER_13_2239 ();
 sg13g2_fill_1 FILLER_13_2267 ();
 sg13g2_fill_1 FILLER_13_2276 ();
 sg13g2_decap_4 FILLER_13_2298 ();
 sg13g2_fill_2 FILLER_13_2302 ();
 sg13g2_fill_2 FILLER_13_2327 ();
 sg13g2_fill_1 FILLER_13_2329 ();
 sg13g2_fill_2 FILLER_13_2423 ();
 sg13g2_fill_1 FILLER_13_2425 ();
 sg13g2_fill_2 FILLER_13_2446 ();
 sg13g2_decap_4 FILLER_13_2462 ();
 sg13g2_decap_4 FILLER_13_2506 ();
 sg13g2_fill_2 FILLER_13_2510 ();
 sg13g2_decap_8 FILLER_13_2516 ();
 sg13g2_decap_4 FILLER_13_2523 ();
 sg13g2_fill_1 FILLER_13_2527 ();
 sg13g2_fill_1 FILLER_13_2538 ();
 sg13g2_decap_8 FILLER_13_2552 ();
 sg13g2_fill_2 FILLER_13_2559 ();
 sg13g2_decap_8 FILLER_13_2597 ();
 sg13g2_decap_8 FILLER_13_2604 ();
 sg13g2_decap_8 FILLER_13_2611 ();
 sg13g2_decap_8 FILLER_13_2618 ();
 sg13g2_decap_8 FILLER_13_2625 ();
 sg13g2_decap_8 FILLER_13_2632 ();
 sg13g2_decap_8 FILLER_13_2639 ();
 sg13g2_decap_8 FILLER_13_2646 ();
 sg13g2_decap_8 FILLER_13_2653 ();
 sg13g2_decap_8 FILLER_13_2660 ();
 sg13g2_fill_2 FILLER_13_2667 ();
 sg13g2_fill_1 FILLER_13_2669 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_37 ();
 sg13g2_decap_8 FILLER_14_52 ();
 sg13g2_fill_2 FILLER_14_63 ();
 sg13g2_fill_1 FILLER_14_69 ();
 sg13g2_fill_1 FILLER_14_74 ();
 sg13g2_fill_2 FILLER_14_83 ();
 sg13g2_fill_2 FILLER_14_93 ();
 sg13g2_decap_8 FILLER_14_104 ();
 sg13g2_fill_2 FILLER_14_111 ();
 sg13g2_fill_1 FILLER_14_132 ();
 sg13g2_fill_2 FILLER_14_165 ();
 sg13g2_fill_2 FILLER_14_206 ();
 sg13g2_fill_1 FILLER_14_241 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_fill_1 FILLER_14_292 ();
 sg13g2_fill_1 FILLER_14_304 ();
 sg13g2_fill_2 FILLER_14_335 ();
 sg13g2_fill_2 FILLER_14_342 ();
 sg13g2_fill_2 FILLER_14_348 ();
 sg13g2_fill_1 FILLER_14_353 ();
 sg13g2_fill_2 FILLER_14_376 ();
 sg13g2_fill_1 FILLER_14_388 ();
 sg13g2_fill_1 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_449 ();
 sg13g2_fill_1 FILLER_14_454 ();
 sg13g2_fill_2 FILLER_14_487 ();
 sg13g2_decap_4 FILLER_14_505 ();
 sg13g2_fill_1 FILLER_14_509 ();
 sg13g2_fill_1 FILLER_14_527 ();
 sg13g2_decap_8 FILLER_14_532 ();
 sg13g2_decap_8 FILLER_14_539 ();
 sg13g2_decap_4 FILLER_14_546 ();
 sg13g2_fill_1 FILLER_14_550 ();
 sg13g2_decap_4 FILLER_14_556 ();
 sg13g2_fill_1 FILLER_14_560 ();
 sg13g2_fill_1 FILLER_14_567 ();
 sg13g2_decap_4 FILLER_14_620 ();
 sg13g2_fill_1 FILLER_14_624 ();
 sg13g2_decap_4 FILLER_14_630 ();
 sg13g2_fill_1 FILLER_14_634 ();
 sg13g2_fill_1 FILLER_14_652 ();
 sg13g2_fill_2 FILLER_14_663 ();
 sg13g2_fill_1 FILLER_14_670 ();
 sg13g2_fill_2 FILLER_14_697 ();
 sg13g2_fill_1 FILLER_14_703 ();
 sg13g2_decap_8 FILLER_14_714 ();
 sg13g2_decap_8 FILLER_14_721 ();
 sg13g2_fill_2 FILLER_14_728 ();
 sg13g2_fill_1 FILLER_14_730 ();
 sg13g2_fill_1 FILLER_14_757 ();
 sg13g2_fill_2 FILLER_14_784 ();
 sg13g2_fill_2 FILLER_14_796 ();
 sg13g2_fill_2 FILLER_14_808 ();
 sg13g2_decap_8 FILLER_14_836 ();
 sg13g2_decap_4 FILLER_14_843 ();
 sg13g2_fill_1 FILLER_14_847 ();
 sg13g2_fill_2 FILLER_14_878 ();
 sg13g2_fill_2 FILLER_14_898 ();
 sg13g2_fill_1 FILLER_14_900 ();
 sg13g2_decap_8 FILLER_14_911 ();
 sg13g2_decap_8 FILLER_14_918 ();
 sg13g2_decap_8 FILLER_14_925 ();
 sg13g2_decap_8 FILLER_14_932 ();
 sg13g2_decap_8 FILLER_14_939 ();
 sg13g2_decap_8 FILLER_14_946 ();
 sg13g2_fill_1 FILLER_14_953 ();
 sg13g2_decap_8 FILLER_14_993 ();
 sg13g2_decap_8 FILLER_14_1000 ();
 sg13g2_decap_8 FILLER_14_1007 ();
 sg13g2_fill_1 FILLER_14_1019 ();
 sg13g2_fill_1 FILLER_14_1050 ();
 sg13g2_fill_1 FILLER_14_1055 ();
 sg13g2_decap_8 FILLER_14_1087 ();
 sg13g2_fill_2 FILLER_14_1098 ();
 sg13g2_fill_1 FILLER_14_1100 ();
 sg13g2_fill_2 FILLER_14_1119 ();
 sg13g2_fill_1 FILLER_14_1121 ();
 sg13g2_decap_8 FILLER_14_1126 ();
 sg13g2_decap_8 FILLER_14_1133 ();
 sg13g2_fill_1 FILLER_14_1140 ();
 sg13g2_decap_4 FILLER_14_1145 ();
 sg13g2_fill_1 FILLER_14_1149 ();
 sg13g2_fill_2 FILLER_14_1154 ();
 sg13g2_decap_8 FILLER_14_1160 ();
 sg13g2_decap_8 FILLER_14_1167 ();
 sg13g2_fill_1 FILLER_14_1174 ();
 sg13g2_decap_4 FILLER_14_1185 ();
 sg13g2_fill_1 FILLER_14_1201 ();
 sg13g2_decap_4 FILLER_14_1223 ();
 sg13g2_fill_1 FILLER_14_1227 ();
 sg13g2_fill_2 FILLER_14_1242 ();
 sg13g2_fill_2 FILLER_14_1265 ();
 sg13g2_fill_1 FILLER_14_1267 ();
 sg13g2_decap_8 FILLER_14_1287 ();
 sg13g2_fill_1 FILLER_14_1294 ();
 sg13g2_fill_2 FILLER_14_1331 ();
 sg13g2_fill_2 FILLER_14_1376 ();
 sg13g2_fill_2 FILLER_14_1402 ();
 sg13g2_fill_1 FILLER_14_1404 ();
 sg13g2_fill_1 FILLER_14_1437 ();
 sg13g2_fill_1 FILLER_14_1486 ();
 sg13g2_fill_1 FILLER_14_1491 ();
 sg13g2_fill_2 FILLER_14_1544 ();
 sg13g2_fill_1 FILLER_14_1546 ();
 sg13g2_fill_1 FILLER_14_1554 ();
 sg13g2_fill_1 FILLER_14_1565 ();
 sg13g2_decap_8 FILLER_14_1569 ();
 sg13g2_decap_8 FILLER_14_1576 ();
 sg13g2_decap_8 FILLER_14_1583 ();
 sg13g2_decap_4 FILLER_14_1590 ();
 sg13g2_fill_1 FILLER_14_1594 ();
 sg13g2_fill_1 FILLER_14_1621 ();
 sg13g2_decap_8 FILLER_14_1642 ();
 sg13g2_decap_8 FILLER_14_1649 ();
 sg13g2_decap_8 FILLER_14_1656 ();
 sg13g2_decap_8 FILLER_14_1663 ();
 sg13g2_decap_8 FILLER_14_1670 ();
 sg13g2_fill_2 FILLER_14_1677 ();
 sg13g2_fill_1 FILLER_14_1703 ();
 sg13g2_fill_2 FILLER_14_1769 ();
 sg13g2_decap_8 FILLER_14_1800 ();
 sg13g2_decap_8 FILLER_14_1807 ();
 sg13g2_decap_4 FILLER_14_1814 ();
 sg13g2_fill_1 FILLER_14_1818 ();
 sg13g2_fill_1 FILLER_14_1849 ();
 sg13g2_fill_1 FILLER_14_1875 ();
 sg13g2_fill_1 FILLER_14_1884 ();
 sg13g2_fill_1 FILLER_14_1924 ();
 sg13g2_decap_4 FILLER_14_1961 ();
 sg13g2_fill_1 FILLER_14_1965 ();
 sg13g2_fill_1 FILLER_14_2006 ();
 sg13g2_decap_8 FILLER_14_2015 ();
 sg13g2_fill_2 FILLER_14_2048 ();
 sg13g2_decap_4 FILLER_14_2083 ();
 sg13g2_fill_2 FILLER_14_2087 ();
 sg13g2_decap_8 FILLER_14_2110 ();
 sg13g2_decap_8 FILLER_14_2117 ();
 sg13g2_decap_8 FILLER_14_2124 ();
 sg13g2_fill_1 FILLER_14_2131 ();
 sg13g2_decap_4 FILLER_14_2151 ();
 sg13g2_fill_2 FILLER_14_2155 ();
 sg13g2_fill_2 FILLER_14_2167 ();
 sg13g2_fill_1 FILLER_14_2169 ();
 sg13g2_decap_8 FILLER_14_2180 ();
 sg13g2_decap_8 FILLER_14_2187 ();
 sg13g2_decap_4 FILLER_14_2194 ();
 sg13g2_fill_1 FILLER_14_2198 ();
 sg13g2_decap_8 FILLER_14_2209 ();
 sg13g2_decap_8 FILLER_14_2220 ();
 sg13g2_decap_8 FILLER_14_2227 ();
 sg13g2_fill_1 FILLER_14_2234 ();
 sg13g2_fill_1 FILLER_14_2305 ();
 sg13g2_decap_4 FILLER_14_2332 ();
 sg13g2_fill_2 FILLER_14_2336 ();
 sg13g2_decap_4 FILLER_14_2348 ();
 sg13g2_fill_1 FILLER_14_2352 ();
 sg13g2_decap_8 FILLER_14_2379 ();
 sg13g2_fill_1 FILLER_14_2404 ();
 sg13g2_fill_1 FILLER_14_2411 ();
 sg13g2_fill_1 FILLER_14_2422 ();
 sg13g2_fill_2 FILLER_14_2429 ();
 sg13g2_fill_2 FILLER_14_2437 ();
 sg13g2_fill_1 FILLER_14_2439 ();
 sg13g2_decap_8 FILLER_14_2450 ();
 sg13g2_decap_4 FILLER_14_2457 ();
 sg13g2_fill_2 FILLER_14_2461 ();
 sg13g2_decap_4 FILLER_14_2473 ();
 sg13g2_decap_8 FILLER_14_2483 ();
 sg13g2_fill_1 FILLER_14_2490 ();
 sg13g2_fill_2 FILLER_14_2511 ();
 sg13g2_fill_2 FILLER_14_2525 ();
 sg13g2_fill_2 FILLER_14_2553 ();
 sg13g2_decap_8 FILLER_14_2607 ();
 sg13g2_decap_8 FILLER_14_2614 ();
 sg13g2_decap_8 FILLER_14_2621 ();
 sg13g2_decap_8 FILLER_14_2628 ();
 sg13g2_decap_8 FILLER_14_2635 ();
 sg13g2_decap_8 FILLER_14_2642 ();
 sg13g2_decap_8 FILLER_14_2649 ();
 sg13g2_decap_8 FILLER_14_2656 ();
 sg13g2_decap_8 FILLER_14_2663 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_7 ();
 sg13g2_fill_1 FILLER_15_9 ();
 sg13g2_fill_1 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_19 ();
 sg13g2_decap_8 FILLER_15_34 ();
 sg13g2_decap_8 FILLER_15_41 ();
 sg13g2_decap_8 FILLER_15_48 ();
 sg13g2_decap_4 FILLER_15_55 ();
 sg13g2_decap_8 FILLER_15_89 ();
 sg13g2_decap_4 FILLER_15_96 ();
 sg13g2_fill_2 FILLER_15_100 ();
 sg13g2_fill_1 FILLER_15_107 ();
 sg13g2_fill_1 FILLER_15_139 ();
 sg13g2_fill_1 FILLER_15_163 ();
 sg13g2_fill_1 FILLER_15_169 ();
 sg13g2_fill_2 FILLER_15_219 ();
 sg13g2_fill_1 FILLER_15_233 ();
 sg13g2_fill_2 FILLER_15_240 ();
 sg13g2_fill_2 FILLER_15_280 ();
 sg13g2_fill_1 FILLER_15_282 ();
 sg13g2_decap_4 FILLER_15_288 ();
 sg13g2_fill_2 FILLER_15_324 ();
 sg13g2_fill_1 FILLER_15_383 ();
 sg13g2_fill_1 FILLER_15_422 ();
 sg13g2_fill_1 FILLER_15_518 ();
 sg13g2_fill_1 FILLER_15_524 ();
 sg13g2_decap_4 FILLER_15_530 ();
 sg13g2_decap_8 FILLER_15_539 ();
 sg13g2_decap_8 FILLER_15_550 ();
 sg13g2_decap_4 FILLER_15_557 ();
 sg13g2_fill_2 FILLER_15_561 ();
 sg13g2_decap_4 FILLER_15_567 ();
 sg13g2_decap_8 FILLER_15_575 ();
 sg13g2_decap_8 FILLER_15_582 ();
 sg13g2_decap_8 FILLER_15_589 ();
 sg13g2_decap_4 FILLER_15_596 ();
 sg13g2_fill_2 FILLER_15_600 ();
 sg13g2_fill_2 FILLER_15_612 ();
 sg13g2_fill_1 FILLER_15_628 ();
 sg13g2_fill_1 FILLER_15_633 ();
 sg13g2_fill_1 FILLER_15_660 ();
 sg13g2_fill_2 FILLER_15_687 ();
 sg13g2_fill_1 FILLER_15_715 ();
 sg13g2_fill_2 FILLER_15_732 ();
 sg13g2_fill_1 FILLER_15_734 ();
 sg13g2_decap_8 FILLER_15_761 ();
 sg13g2_fill_2 FILLER_15_768 ();
 sg13g2_fill_1 FILLER_15_770 ();
 sg13g2_fill_2 FILLER_15_883 ();
 sg13g2_fill_1 FILLER_15_885 ();
 sg13g2_decap_8 FILLER_15_941 ();
 sg13g2_fill_2 FILLER_15_948 ();
 sg13g2_fill_1 FILLER_15_950 ();
 sg13g2_fill_1 FILLER_15_977 ();
 sg13g2_fill_1 FILLER_15_1008 ();
 sg13g2_decap_4 FILLER_15_1013 ();
 sg13g2_fill_2 FILLER_15_1017 ();
 sg13g2_decap_8 FILLER_15_1031 ();
 sg13g2_fill_1 FILLER_15_1038 ();
 sg13g2_decap_8 FILLER_15_1044 ();
 sg13g2_decap_8 FILLER_15_1051 ();
 sg13g2_fill_2 FILLER_15_1093 ();
 sg13g2_fill_2 FILLER_15_1100 ();
 sg13g2_fill_1 FILLER_15_1102 ();
 sg13g2_decap_8 FILLER_15_1132 ();
 sg13g2_decap_4 FILLER_15_1139 ();
 sg13g2_fill_2 FILLER_15_1174 ();
 sg13g2_fill_1 FILLER_15_1176 ();
 sg13g2_decap_8 FILLER_15_1217 ();
 sg13g2_decap_4 FILLER_15_1224 ();
 sg13g2_fill_1 FILLER_15_1228 ();
 sg13g2_decap_4 FILLER_15_1255 ();
 sg13g2_fill_2 FILLER_15_1259 ();
 sg13g2_fill_2 FILLER_15_1305 ();
 sg13g2_decap_4 FILLER_15_1333 ();
 sg13g2_fill_2 FILLER_15_1341 ();
 sg13g2_fill_1 FILLER_15_1343 ();
 sg13g2_fill_1 FILLER_15_1459 ();
 sg13g2_fill_2 FILLER_15_1465 ();
 sg13g2_fill_1 FILLER_15_1494 ();
 sg13g2_fill_2 FILLER_15_1504 ();
 sg13g2_decap_8 FILLER_15_1558 ();
 sg13g2_fill_1 FILLER_15_1565 ();
 sg13g2_fill_2 FILLER_15_1571 ();
 sg13g2_decap_4 FILLER_15_1582 ();
 sg13g2_fill_2 FILLER_15_1590 ();
 sg13g2_decap_8 FILLER_15_1661 ();
 sg13g2_decap_4 FILLER_15_1668 ();
 sg13g2_fill_2 FILLER_15_1682 ();
 sg13g2_fill_2 FILLER_15_1715 ();
 sg13g2_fill_1 FILLER_15_1721 ();
 sg13g2_decap_8 FILLER_15_1748 ();
 sg13g2_fill_1 FILLER_15_1817 ();
 sg13g2_decap_8 FILLER_15_1824 ();
 sg13g2_fill_2 FILLER_15_1831 ();
 sg13g2_fill_1 FILLER_15_1833 ();
 sg13g2_decap_4 FILLER_15_1838 ();
 sg13g2_fill_2 FILLER_15_1842 ();
 sg13g2_fill_2 FILLER_15_1866 ();
 sg13g2_fill_1 FILLER_15_1886 ();
 sg13g2_decap_8 FILLER_15_1896 ();
 sg13g2_decap_8 FILLER_15_1903 ();
 sg13g2_decap_8 FILLER_15_1910 ();
 sg13g2_decap_8 FILLER_15_1917 ();
 sg13g2_decap_4 FILLER_15_1934 ();
 sg13g2_fill_1 FILLER_15_1938 ();
 sg13g2_fill_1 FILLER_15_1943 ();
 sg13g2_fill_2 FILLER_15_1980 ();
 sg13g2_fill_1 FILLER_15_1982 ();
 sg13g2_fill_2 FILLER_15_2013 ();
 sg13g2_decap_4 FILLER_15_2025 ();
 sg13g2_decap_8 FILLER_15_2033 ();
 sg13g2_decap_8 FILLER_15_2040 ();
 sg13g2_decap_4 FILLER_15_2047 ();
 sg13g2_decap_8 FILLER_15_2055 ();
 sg13g2_decap_8 FILLER_15_2062 ();
 sg13g2_decap_8 FILLER_15_2069 ();
 sg13g2_decap_8 FILLER_15_2128 ();
 sg13g2_decap_4 FILLER_15_2135 ();
 sg13g2_fill_2 FILLER_15_2139 ();
 sg13g2_decap_8 FILLER_15_2145 ();
 sg13g2_fill_2 FILLER_15_2152 ();
 sg13g2_fill_1 FILLER_15_2154 ();
 sg13g2_decap_8 FILLER_15_2165 ();
 sg13g2_fill_1 FILLER_15_2172 ();
 sg13g2_fill_2 FILLER_15_2183 ();
 sg13g2_fill_1 FILLER_15_2185 ();
 sg13g2_decap_4 FILLER_15_2217 ();
 sg13g2_decap_4 FILLER_15_2231 ();
 sg13g2_decap_8 FILLER_15_2240 ();
 sg13g2_fill_2 FILLER_15_2251 ();
 sg13g2_decap_4 FILLER_15_2257 ();
 sg13g2_fill_2 FILLER_15_2274 ();
 sg13g2_decap_4 FILLER_15_2280 ();
 sg13g2_decap_8 FILLER_15_2310 ();
 sg13g2_decap_8 FILLER_15_2317 ();
 sg13g2_decap_4 FILLER_15_2324 ();
 sg13g2_fill_2 FILLER_15_2328 ();
 sg13g2_decap_4 FILLER_15_2340 ();
 sg13g2_fill_1 FILLER_15_2344 ();
 sg13g2_fill_1 FILLER_15_2355 ();
 sg13g2_decap_8 FILLER_15_2364 ();
 sg13g2_decap_8 FILLER_15_2371 ();
 sg13g2_decap_8 FILLER_15_2378 ();
 sg13g2_decap_8 FILLER_15_2385 ();
 sg13g2_decap_8 FILLER_15_2392 ();
 sg13g2_decap_4 FILLER_15_2399 ();
 sg13g2_fill_1 FILLER_15_2459 ();
 sg13g2_decap_8 FILLER_15_2466 ();
 sg13g2_decap_8 FILLER_15_2473 ();
 sg13g2_decap_8 FILLER_15_2480 ();
 sg13g2_fill_2 FILLER_15_2487 ();
 sg13g2_fill_2 FILLER_15_2515 ();
 sg13g2_fill_1 FILLER_15_2517 ();
 sg13g2_fill_1 FILLER_15_2574 ();
 sg13g2_fill_2 FILLER_15_2589 ();
 sg13g2_decap_4 FILLER_15_2595 ();
 sg13g2_fill_2 FILLER_15_2599 ();
 sg13g2_decap_8 FILLER_15_2624 ();
 sg13g2_decap_8 FILLER_15_2631 ();
 sg13g2_decap_8 FILLER_15_2638 ();
 sg13g2_decap_8 FILLER_15_2645 ();
 sg13g2_decap_8 FILLER_15_2652 ();
 sg13g2_decap_8 FILLER_15_2659 ();
 sg13g2_decap_4 FILLER_15_2666 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_13 ();
 sg13g2_fill_2 FILLER_16_20 ();
 sg13g2_decap_8 FILLER_16_27 ();
 sg13g2_decap_8 FILLER_16_38 ();
 sg13g2_decap_8 FILLER_16_45 ();
 sg13g2_fill_2 FILLER_16_52 ();
 sg13g2_fill_1 FILLER_16_67 ();
 sg13g2_fill_2 FILLER_16_94 ();
 sg13g2_fill_1 FILLER_16_96 ();
 sg13g2_fill_2 FILLER_16_133 ();
 sg13g2_fill_2 FILLER_16_183 ();
 sg13g2_fill_1 FILLER_16_224 ();
 sg13g2_fill_1 FILLER_16_238 ();
 sg13g2_fill_1 FILLER_16_317 ();
 sg13g2_fill_1 FILLER_16_396 ();
 sg13g2_fill_2 FILLER_16_441 ();
 sg13g2_fill_1 FILLER_16_443 ();
 sg13g2_fill_1 FILLER_16_454 ();
 sg13g2_decap_8 FILLER_16_472 ();
 sg13g2_fill_2 FILLER_16_479 ();
 sg13g2_fill_1 FILLER_16_481 ();
 sg13g2_fill_1 FILLER_16_492 ();
 sg13g2_fill_2 FILLER_16_498 ();
 sg13g2_decap_8 FILLER_16_513 ();
 sg13g2_decap_4 FILLER_16_524 ();
 sg13g2_decap_4 FILLER_16_560 ();
 sg13g2_fill_1 FILLER_16_564 ();
 sg13g2_fill_2 FILLER_16_573 ();
 sg13g2_decap_4 FILLER_16_580 ();
 sg13g2_fill_1 FILLER_16_584 ();
 sg13g2_fill_2 FILLER_16_589 ();
 sg13g2_decap_4 FILLER_16_596 ();
 sg13g2_fill_1 FILLER_16_600 ();
 sg13g2_fill_1 FILLER_16_612 ();
 sg13g2_fill_2 FILLER_16_649 ();
 sg13g2_fill_2 FILLER_16_656 ();
 sg13g2_decap_4 FILLER_16_664 ();
 sg13g2_fill_2 FILLER_16_672 ();
 sg13g2_fill_2 FILLER_16_684 ();
 sg13g2_fill_2 FILLER_16_698 ();
 sg13g2_fill_1 FILLER_16_700 ();
 sg13g2_fill_1 FILLER_16_731 ();
 sg13g2_fill_2 FILLER_16_737 ();
 sg13g2_fill_1 FILLER_16_743 ();
 sg13g2_fill_2 FILLER_16_748 ();
 sg13g2_decap_8 FILLER_16_754 ();
 sg13g2_fill_1 FILLER_16_761 ();
 sg13g2_fill_2 FILLER_16_813 ();
 sg13g2_fill_2 FILLER_16_825 ();
 sg13g2_fill_1 FILLER_16_827 ();
 sg13g2_fill_1 FILLER_16_854 ();
 sg13g2_fill_2 FILLER_16_865 ();
 sg13g2_fill_1 FILLER_16_867 ();
 sg13g2_decap_4 FILLER_16_878 ();
 sg13g2_fill_2 FILLER_16_882 ();
 sg13g2_fill_2 FILLER_16_960 ();
 sg13g2_fill_1 FILLER_16_962 ();
 sg13g2_fill_1 FILLER_16_1036 ();
 sg13g2_fill_2 FILLER_16_1041 ();
 sg13g2_fill_2 FILLER_16_1064 ();
 sg13g2_fill_1 FILLER_16_1070 ();
 sg13g2_fill_1 FILLER_16_1140 ();
 sg13g2_fill_2 FILLER_16_1146 ();
 sg13g2_fill_1 FILLER_16_1152 ();
 sg13g2_decap_8 FILLER_16_1174 ();
 sg13g2_decap_8 FILLER_16_1211 ();
 sg13g2_decap_8 FILLER_16_1218 ();
 sg13g2_decap_8 FILLER_16_1225 ();
 sg13g2_decap_4 FILLER_16_1232 ();
 sg13g2_fill_1 FILLER_16_1236 ();
 sg13g2_fill_2 FILLER_16_1328 ();
 sg13g2_fill_1 FILLER_16_1330 ();
 sg13g2_fill_2 FILLER_16_1357 ();
 sg13g2_fill_1 FILLER_16_1359 ();
 sg13g2_fill_2 FILLER_16_1425 ();
 sg13g2_fill_1 FILLER_16_1427 ();
 sg13g2_fill_2 FILLER_16_1432 ();
 sg13g2_fill_1 FILLER_16_1448 ();
 sg13g2_fill_2 FILLER_16_1467 ();
 sg13g2_fill_1 FILLER_16_1476 ();
 sg13g2_fill_1 FILLER_16_1481 ();
 sg13g2_fill_1 FILLER_16_1526 ();
 sg13g2_fill_1 FILLER_16_1532 ();
 sg13g2_fill_1 FILLER_16_1539 ();
 sg13g2_decap_8 FILLER_16_1544 ();
 sg13g2_decap_4 FILLER_16_1551 ();
 sg13g2_decap_8 FILLER_16_1566 ();
 sg13g2_decap_8 FILLER_16_1573 ();
 sg13g2_decap_8 FILLER_16_1580 ();
 sg13g2_decap_4 FILLER_16_1587 ();
 sg13g2_fill_1 FILLER_16_1591 ();
 sg13g2_fill_2 FILLER_16_1602 ();
 sg13g2_fill_2 FILLER_16_1608 ();
 sg13g2_fill_2 FILLER_16_1620 ();
 sg13g2_fill_1 FILLER_16_1622 ();
 sg13g2_fill_2 FILLER_16_1627 ();
 sg13g2_fill_1 FILLER_16_1629 ();
 sg13g2_decap_8 FILLER_16_1661 ();
 sg13g2_fill_2 FILLER_16_1668 ();
 sg13g2_fill_1 FILLER_16_1696 ();
 sg13g2_fill_1 FILLER_16_1701 ();
 sg13g2_decap_8 FILLER_16_1723 ();
 sg13g2_fill_2 FILLER_16_1730 ();
 sg13g2_fill_1 FILLER_16_1732 ();
 sg13g2_fill_2 FILLER_16_1747 ();
 sg13g2_fill_1 FILLER_16_1753 ();
 sg13g2_decap_8 FILLER_16_1780 ();
 sg13g2_fill_2 FILLER_16_1787 ();
 sg13g2_fill_1 FILLER_16_1822 ();
 sg13g2_fill_2 FILLER_16_1837 ();
 sg13g2_fill_1 FILLER_16_1839 ();
 sg13g2_fill_2 FILLER_16_1896 ();
 sg13g2_decap_8 FILLER_16_1933 ();
 sg13g2_decap_8 FILLER_16_1940 ();
 sg13g2_decap_8 FILLER_16_1947 ();
 sg13g2_decap_4 FILLER_16_1954 ();
 sg13g2_fill_2 FILLER_16_1958 ();
 sg13g2_fill_1 FILLER_16_1978 ();
 sg13g2_decap_8 FILLER_16_2020 ();
 sg13g2_decap_4 FILLER_16_2027 ();
 sg13g2_decap_4 FILLER_16_2071 ();
 sg13g2_fill_1 FILLER_16_2075 ();
 sg13g2_fill_2 FILLER_16_2100 ();
 sg13g2_fill_1 FILLER_16_2102 ();
 sg13g2_decap_8 FILLER_16_2132 ();
 sg13g2_decap_8 FILLER_16_2139 ();
 sg13g2_fill_2 FILLER_16_2146 ();
 sg13g2_decap_4 FILLER_16_2235 ();
 sg13g2_fill_2 FILLER_16_2239 ();
 sg13g2_fill_2 FILLER_16_2245 ();
 sg13g2_fill_1 FILLER_16_2247 ();
 sg13g2_decap_8 FILLER_16_2298 ();
 sg13g2_decap_8 FILLER_16_2367 ();
 sg13g2_decap_8 FILLER_16_2374 ();
 sg13g2_decap_8 FILLER_16_2381 ();
 sg13g2_decap_8 FILLER_16_2388 ();
 sg13g2_decap_8 FILLER_16_2395 ();
 sg13g2_decap_4 FILLER_16_2402 ();
 sg13g2_fill_1 FILLER_16_2419 ();
 sg13g2_fill_2 FILLER_16_2469 ();
 sg13g2_decap_8 FILLER_16_2476 ();
 sg13g2_fill_1 FILLER_16_2487 ();
 sg13g2_fill_2 FILLER_16_2538 ();
 sg13g2_fill_1 FILLER_16_2550 ();
 sg13g2_decap_8 FILLER_16_2555 ();
 sg13g2_decap_8 FILLER_16_2562 ();
 sg13g2_fill_2 FILLER_16_2569 ();
 sg13g2_fill_1 FILLER_16_2571 ();
 sg13g2_fill_1 FILLER_16_2612 ();
 sg13g2_decap_8 FILLER_16_2639 ();
 sg13g2_decap_8 FILLER_16_2646 ();
 sg13g2_decap_8 FILLER_16_2653 ();
 sg13g2_decap_8 FILLER_16_2660 ();
 sg13g2_fill_2 FILLER_16_2667 ();
 sg13g2_fill_1 FILLER_16_2669 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_decap_4 FILLER_17_97 ();
 sg13g2_decap_4 FILLER_17_131 ();
 sg13g2_fill_1 FILLER_17_135 ();
 sg13g2_fill_1 FILLER_17_141 ();
 sg13g2_fill_1 FILLER_17_152 ();
 sg13g2_fill_2 FILLER_17_186 ();
 sg13g2_fill_1 FILLER_17_188 ();
 sg13g2_fill_1 FILLER_17_262 ();
 sg13g2_fill_1 FILLER_17_266 ();
 sg13g2_fill_1 FILLER_17_312 ();
 sg13g2_fill_1 FILLER_17_324 ();
 sg13g2_fill_2 FILLER_17_344 ();
 sg13g2_fill_2 FILLER_17_377 ();
 sg13g2_fill_1 FILLER_17_379 ();
 sg13g2_fill_1 FILLER_17_384 ();
 sg13g2_fill_1 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_433 ();
 sg13g2_decap_4 FILLER_17_438 ();
 sg13g2_fill_1 FILLER_17_442 ();
 sg13g2_decap_8 FILLER_17_467 ();
 sg13g2_decap_4 FILLER_17_474 ();
 sg13g2_fill_1 FILLER_17_503 ();
 sg13g2_fill_2 FILLER_17_528 ();
 sg13g2_fill_1 FILLER_17_544 ();
 sg13g2_fill_1 FILLER_17_558 ();
 sg13g2_fill_1 FILLER_17_585 ();
 sg13g2_fill_1 FILLER_17_590 ();
 sg13g2_fill_1 FILLER_17_603 ();
 sg13g2_fill_2 FILLER_17_615 ();
 sg13g2_fill_1 FILLER_17_617 ();
 sg13g2_fill_2 FILLER_17_623 ();
 sg13g2_fill_1 FILLER_17_625 ();
 sg13g2_fill_1 FILLER_17_630 ();
 sg13g2_fill_1 FILLER_17_635 ();
 sg13g2_fill_1 FILLER_17_646 ();
 sg13g2_fill_2 FILLER_17_667 ();
 sg13g2_fill_1 FILLER_17_669 ();
 sg13g2_decap_4 FILLER_17_674 ();
 sg13g2_decap_4 FILLER_17_688 ();
 sg13g2_fill_2 FILLER_17_692 ();
 sg13g2_decap_4 FILLER_17_707 ();
 sg13g2_fill_1 FILLER_17_711 ();
 sg13g2_fill_1 FILLER_17_722 ();
 sg13g2_fill_2 FILLER_17_727 ();
 sg13g2_fill_1 FILLER_17_729 ();
 sg13g2_decap_8 FILLER_17_756 ();
 sg13g2_decap_8 FILLER_17_763 ();
 sg13g2_fill_1 FILLER_17_770 ();
 sg13g2_fill_2 FILLER_17_789 ();
 sg13g2_decap_8 FILLER_17_801 ();
 sg13g2_decap_8 FILLER_17_808 ();
 sg13g2_decap_4 FILLER_17_819 ();
 sg13g2_fill_1 FILLER_17_853 ();
 sg13g2_fill_2 FILLER_17_916 ();
 sg13g2_fill_2 FILLER_17_958 ();
 sg13g2_fill_2 FILLER_17_973 ();
 sg13g2_fill_1 FILLER_17_975 ();
 sg13g2_fill_1 FILLER_17_990 ();
 sg13g2_fill_2 FILLER_17_1022 ();
 sg13g2_fill_2 FILLER_17_1050 ();
 sg13g2_fill_1 FILLER_17_1057 ();
 sg13g2_decap_8 FILLER_17_1101 ();
 sg13g2_decap_4 FILLER_17_1108 ();
 sg13g2_decap_4 FILLER_17_1116 ();
 sg13g2_decap_4 FILLER_17_1141 ();
 sg13g2_fill_1 FILLER_17_1154 ();
 sg13g2_decap_8 FILLER_17_1215 ();
 sg13g2_decap_8 FILLER_17_1222 ();
 sg13g2_decap_4 FILLER_17_1229 ();
 sg13g2_decap_4 FILLER_17_1257 ();
 sg13g2_fill_2 FILLER_17_1265 ();
 sg13g2_fill_1 FILLER_17_1267 ();
 sg13g2_fill_1 FILLER_17_1280 ();
 sg13g2_fill_1 FILLER_17_1289 ();
 sg13g2_fill_2 FILLER_17_1300 ();
 sg13g2_fill_1 FILLER_17_1302 ();
 sg13g2_fill_1 FILLER_17_1317 ();
 sg13g2_decap_8 FILLER_17_1322 ();
 sg13g2_decap_4 FILLER_17_1329 ();
 sg13g2_fill_2 FILLER_17_1333 ();
 sg13g2_decap_8 FILLER_17_1339 ();
 sg13g2_decap_4 FILLER_17_1346 ();
 sg13g2_fill_2 FILLER_17_1350 ();
 sg13g2_fill_2 FILLER_17_1356 ();
 sg13g2_fill_1 FILLER_17_1358 ();
 sg13g2_fill_2 FILLER_17_1459 ();
 sg13g2_fill_2 FILLER_17_1472 ();
 sg13g2_decap_8 FILLER_17_1539 ();
 sg13g2_fill_2 FILLER_17_1546 ();
 sg13g2_fill_1 FILLER_17_1548 ();
 sg13g2_decap_4 FILLER_17_1575 ();
 sg13g2_fill_1 FILLER_17_1579 ();
 sg13g2_fill_1 FILLER_17_1610 ();
 sg13g2_decap_8 FILLER_17_1667 ();
 sg13g2_fill_2 FILLER_17_1674 ();
 sg13g2_fill_1 FILLER_17_1676 ();
 sg13g2_fill_2 FILLER_17_1711 ();
 sg13g2_fill_1 FILLER_17_1713 ();
 sg13g2_fill_2 FILLER_17_1722 ();
 sg13g2_decap_4 FILLER_17_1741 ();
 sg13g2_fill_1 FILLER_17_1745 ();
 sg13g2_fill_1 FILLER_17_1761 ();
 sg13g2_fill_2 FILLER_17_1815 ();
 sg13g2_fill_1 FILLER_17_1817 ();
 sg13g2_fill_1 FILLER_17_1907 ();
 sg13g2_decap_8 FILLER_17_1918 ();
 sg13g2_decap_8 FILLER_17_1925 ();
 sg13g2_decap_8 FILLER_17_1932 ();
 sg13g2_decap_8 FILLER_17_1962 ();
 sg13g2_decap_4 FILLER_17_1969 ();
 sg13g2_decap_4 FILLER_17_1983 ();
 sg13g2_fill_2 FILLER_17_1987 ();
 sg13g2_fill_2 FILLER_17_2001 ();
 sg13g2_fill_1 FILLER_17_2037 ();
 sg13g2_decap_8 FILLER_17_2044 ();
 sg13g2_fill_2 FILLER_17_2051 ();
 sg13g2_decap_4 FILLER_17_2087 ();
 sg13g2_fill_2 FILLER_17_2091 ();
 sg13g2_fill_1 FILLER_17_2125 ();
 sg13g2_fill_1 FILLER_17_2133 ();
 sg13g2_fill_1 FILLER_17_2144 ();
 sg13g2_fill_1 FILLER_17_2171 ();
 sg13g2_fill_1 FILLER_17_2208 ();
 sg13g2_decap_8 FILLER_17_2265 ();
 sg13g2_fill_2 FILLER_17_2272 ();
 sg13g2_fill_1 FILLER_17_2274 ();
 sg13g2_fill_1 FILLER_17_2292 ();
 sg13g2_fill_1 FILLER_17_2350 ();
 sg13g2_decap_4 FILLER_17_2355 ();
 sg13g2_decap_8 FILLER_17_2425 ();
 sg13g2_fill_2 FILLER_17_2432 ();
 sg13g2_fill_1 FILLER_17_2434 ();
 sg13g2_fill_1 FILLER_17_2453 ();
 sg13g2_fill_2 FILLER_17_2464 ();
 sg13g2_fill_1 FILLER_17_2492 ();
 sg13g2_decap_8 FILLER_17_2517 ();
 sg13g2_fill_2 FILLER_17_2524 ();
 sg13g2_fill_1 FILLER_17_2526 ();
 sg13g2_decap_4 FILLER_17_2531 ();
 sg13g2_fill_1 FILLER_17_2535 ();
 sg13g2_decap_4 FILLER_17_2540 ();
 sg13g2_fill_1 FILLER_17_2544 ();
 sg13g2_fill_1 FILLER_17_2627 ();
 sg13g2_decap_8 FILLER_17_2636 ();
 sg13g2_decap_4 FILLER_17_2643 ();
 sg13g2_decap_8 FILLER_17_2651 ();
 sg13g2_decap_8 FILLER_17_2658 ();
 sg13g2_decap_4 FILLER_17_2665 ();
 sg13g2_fill_1 FILLER_17_2669 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_33 ();
 sg13g2_fill_2 FILLER_18_49 ();
 sg13g2_fill_2 FILLER_18_55 ();
 sg13g2_fill_2 FILLER_18_61 ();
 sg13g2_fill_1 FILLER_18_63 ();
 sg13g2_fill_2 FILLER_18_68 ();
 sg13g2_fill_1 FILLER_18_70 ();
 sg13g2_fill_1 FILLER_18_89 ();
 sg13g2_fill_2 FILLER_18_111 ();
 sg13g2_fill_2 FILLER_18_127 ();
 sg13g2_fill_1 FILLER_18_129 ();
 sg13g2_fill_1 FILLER_18_134 ();
 sg13g2_decap_4 FILLER_18_180 ();
 sg13g2_fill_1 FILLER_18_184 ();
 sg13g2_fill_1 FILLER_18_223 ();
 sg13g2_fill_2 FILLER_18_248 ();
 sg13g2_fill_2 FILLER_18_261 ();
 sg13g2_fill_1 FILLER_18_269 ();
 sg13g2_decap_4 FILLER_18_307 ();
 sg13g2_fill_1 FILLER_18_311 ();
 sg13g2_fill_1 FILLER_18_327 ();
 sg13g2_decap_8 FILLER_18_352 ();
 sg13g2_fill_1 FILLER_18_359 ();
 sg13g2_fill_2 FILLER_18_365 ();
 sg13g2_decap_4 FILLER_18_370 ();
 sg13g2_fill_1 FILLER_18_374 ();
 sg13g2_fill_2 FILLER_18_419 ();
 sg13g2_fill_1 FILLER_18_421 ();
 sg13g2_fill_1 FILLER_18_426 ();
 sg13g2_fill_2 FILLER_18_458 ();
 sg13g2_fill_1 FILLER_18_460 ();
 sg13g2_fill_2 FILLER_18_513 ();
 sg13g2_fill_1 FILLER_18_521 ();
 sg13g2_fill_2 FILLER_18_526 ();
 sg13g2_fill_2 FILLER_18_542 ();
 sg13g2_fill_2 FILLER_18_606 ();
 sg13g2_fill_1 FILLER_18_608 ();
 sg13g2_fill_1 FILLER_18_614 ();
 sg13g2_fill_1 FILLER_18_626 ();
 sg13g2_decap_8 FILLER_18_647 ();
 sg13g2_fill_1 FILLER_18_654 ();
 sg13g2_fill_2 FILLER_18_669 ();
 sg13g2_decap_8 FILLER_18_687 ();
 sg13g2_decap_4 FILLER_18_694 ();
 sg13g2_decap_4 FILLER_18_702 ();
 sg13g2_fill_2 FILLER_18_734 ();
 sg13g2_decap_8 FILLER_18_740 ();
 sg13g2_decap_8 FILLER_18_747 ();
 sg13g2_decap_8 FILLER_18_754 ();
 sg13g2_decap_8 FILLER_18_761 ();
 sg13g2_decap_8 FILLER_18_772 ();
 sg13g2_decap_8 FILLER_18_779 ();
 sg13g2_decap_8 FILLER_18_786 ();
 sg13g2_decap_8 FILLER_18_793 ();
 sg13g2_decap_8 FILLER_18_800 ();
 sg13g2_decap_8 FILLER_18_807 ();
 sg13g2_decap_8 FILLER_18_814 ();
 sg13g2_decap_8 FILLER_18_821 ();
 sg13g2_decap_8 FILLER_18_842 ();
 sg13g2_decap_8 FILLER_18_849 ();
 sg13g2_decap_8 FILLER_18_856 ();
 sg13g2_decap_8 FILLER_18_867 ();
 sg13g2_decap_8 FILLER_18_874 ();
 sg13g2_decap_8 FILLER_18_881 ();
 sg13g2_fill_1 FILLER_18_888 ();
 sg13g2_fill_2 FILLER_18_893 ();
 sg13g2_fill_1 FILLER_18_895 ();
 sg13g2_decap_4 FILLER_18_926 ();
 sg13g2_decap_8 FILLER_18_951 ();
 sg13g2_decap_8 FILLER_18_958 ();
 sg13g2_fill_2 FILLER_18_965 ();
 sg13g2_fill_1 FILLER_18_967 ();
 sg13g2_fill_2 FILLER_18_1008 ();
 sg13g2_fill_2 FILLER_18_1015 ();
 sg13g2_fill_1 FILLER_18_1017 ();
 sg13g2_decap_8 FILLER_18_1121 ();
 sg13g2_decap_8 FILLER_18_1128 ();
 sg13g2_decap_8 FILLER_18_1135 ();
 sg13g2_decap_8 FILLER_18_1142 ();
 sg13g2_decap_4 FILLER_18_1149 ();
 sg13g2_decap_8 FILLER_18_1162 ();
 sg13g2_decap_8 FILLER_18_1169 ();
 sg13g2_decap_4 FILLER_18_1176 ();
 sg13g2_fill_2 FILLER_18_1180 ();
 sg13g2_fill_1 FILLER_18_1186 ();
 sg13g2_decap_8 FILLER_18_1217 ();
 sg13g2_decap_8 FILLER_18_1254 ();
 sg13g2_decap_8 FILLER_18_1261 ();
 sg13g2_fill_2 FILLER_18_1268 ();
 sg13g2_fill_1 FILLER_18_1270 ();
 sg13g2_fill_2 FILLER_18_1275 ();
 sg13g2_fill_2 FILLER_18_1293 ();
 sg13g2_decap_4 FILLER_18_1304 ();
 sg13g2_fill_2 FILLER_18_1308 ();
 sg13g2_decap_8 FILLER_18_1314 ();
 sg13g2_decap_8 FILLER_18_1325 ();
 sg13g2_decap_8 FILLER_18_1332 ();
 sg13g2_decap_8 FILLER_18_1339 ();
 sg13g2_fill_2 FILLER_18_1382 ();
 sg13g2_fill_1 FILLER_18_1430 ();
 sg13g2_fill_1 FILLER_18_1444 ();
 sg13g2_fill_2 FILLER_18_1457 ();
 sg13g2_fill_2 FILLER_18_1555 ();
 sg13g2_fill_2 FILLER_18_1560 ();
 sg13g2_fill_1 FILLER_18_1571 ();
 sg13g2_decap_4 FILLER_18_1585 ();
 sg13g2_decap_4 FILLER_18_1593 ();
 sg13g2_fill_2 FILLER_18_1597 ();
 sg13g2_decap_8 FILLER_18_1604 ();
 sg13g2_decap_8 FILLER_18_1611 ();
 sg13g2_fill_2 FILLER_18_1618 ();
 sg13g2_fill_1 FILLER_18_1620 ();
 sg13g2_fill_1 FILLER_18_1625 ();
 sg13g2_decap_8 FILLER_18_1662 ();
 sg13g2_decap_4 FILLER_18_1669 ();
 sg13g2_fill_2 FILLER_18_1673 ();
 sg13g2_decap_4 FILLER_18_1685 ();
 sg13g2_fill_1 FILLER_18_1689 ();
 sg13g2_decap_4 FILLER_18_1700 ();
 sg13g2_fill_1 FILLER_18_1704 ();
 sg13g2_fill_1 FILLER_18_1744 ();
 sg13g2_fill_1 FILLER_18_1758 ();
 sg13g2_fill_2 FILLER_18_1799 ();
 sg13g2_fill_1 FILLER_18_1801 ();
 sg13g2_decap_8 FILLER_18_1922 ();
 sg13g2_decap_4 FILLER_18_1929 ();
 sg13g2_fill_1 FILLER_18_1933 ();
 sg13g2_fill_2 FILLER_18_1990 ();
 sg13g2_fill_1 FILLER_18_2040 ();
 sg13g2_decap_8 FILLER_18_2077 ();
 sg13g2_decap_8 FILLER_18_2084 ();
 sg13g2_fill_2 FILLER_18_2091 ();
 sg13g2_decap_8 FILLER_18_2119 ();
 sg13g2_decap_4 FILLER_18_2126 ();
 sg13g2_fill_1 FILLER_18_2169 ();
 sg13g2_fill_2 FILLER_18_2199 ();
 sg13g2_fill_1 FILLER_18_2253 ();
 sg13g2_decap_8 FILLER_18_2264 ();
 sg13g2_decap_8 FILLER_18_2271 ();
 sg13g2_decap_4 FILLER_18_2278 ();
 sg13g2_decap_8 FILLER_18_2303 ();
 sg13g2_fill_2 FILLER_18_2310 ();
 sg13g2_fill_1 FILLER_18_2312 ();
 sg13g2_decap_8 FILLER_18_2347 ();
 sg13g2_decap_8 FILLER_18_2354 ();
 sg13g2_decap_4 FILLER_18_2361 ();
 sg13g2_fill_2 FILLER_18_2365 ();
 sg13g2_fill_2 FILLER_18_2377 ();
 sg13g2_decap_8 FILLER_18_2433 ();
 sg13g2_fill_1 FILLER_18_2466 ();
 sg13g2_fill_1 FILLER_18_2473 ();
 sg13g2_fill_1 FILLER_18_2478 ();
 sg13g2_fill_1 FILLER_18_2487 ();
 sg13g2_decap_4 FILLER_18_2498 ();
 sg13g2_fill_2 FILLER_18_2538 ();
 sg13g2_fill_1 FILLER_18_2586 ();
 sg13g2_fill_1 FILLER_18_2591 ();
 sg13g2_fill_1 FILLER_18_2602 ();
 sg13g2_fill_1 FILLER_18_2629 ();
 sg13g2_decap_4 FILLER_18_2666 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_7 ();
 sg13g2_fill_1 FILLER_19_52 ();
 sg13g2_fill_1 FILLER_19_57 ();
 sg13g2_fill_2 FILLER_19_62 ();
 sg13g2_fill_2 FILLER_19_68 ();
 sg13g2_fill_2 FILLER_19_74 ();
 sg13g2_fill_2 FILLER_19_102 ();
 sg13g2_decap_4 FILLER_19_131 ();
 sg13g2_fill_2 FILLER_19_135 ();
 sg13g2_decap_8 FILLER_19_141 ();
 sg13g2_fill_1 FILLER_19_148 ();
 sg13g2_fill_2 FILLER_19_153 ();
 sg13g2_decap_8 FILLER_19_159 ();
 sg13g2_decap_8 FILLER_19_166 ();
 sg13g2_decap_4 FILLER_19_173 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_fill_2 FILLER_19_196 ();
 sg13g2_fill_1 FILLER_19_198 ();
 sg13g2_decap_4 FILLER_19_219 ();
 sg13g2_fill_1 FILLER_19_223 ();
 sg13g2_fill_2 FILLER_19_229 ();
 sg13g2_fill_2 FILLER_19_254 ();
 sg13g2_fill_2 FILLER_19_286 ();
 sg13g2_decap_8 FILLER_19_304 ();
 sg13g2_decap_8 FILLER_19_311 ();
 sg13g2_fill_2 FILLER_19_318 ();
 sg13g2_decap_4 FILLER_19_326 ();
 sg13g2_decap_4 FILLER_19_344 ();
 sg13g2_fill_1 FILLER_19_348 ();
 sg13g2_decap_8 FILLER_19_359 ();
 sg13g2_fill_2 FILLER_19_366 ();
 sg13g2_fill_1 FILLER_19_368 ();
 sg13g2_decap_8 FILLER_19_375 ();
 sg13g2_decap_8 FILLER_19_386 ();
 sg13g2_decap_4 FILLER_19_393 ();
 sg13g2_fill_1 FILLER_19_397 ();
 sg13g2_decap_4 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_410 ();
 sg13g2_decap_4 FILLER_19_456 ();
 sg13g2_fill_1 FILLER_19_460 ();
 sg13g2_decap_8 FILLER_19_544 ();
 sg13g2_fill_2 FILLER_19_551 ();
 sg13g2_fill_1 FILLER_19_553 ();
 sg13g2_fill_1 FILLER_19_558 ();
 sg13g2_decap_4 FILLER_19_563 ();
 sg13g2_fill_2 FILLER_19_581 ();
 sg13g2_fill_1 FILLER_19_593 ();
 sg13g2_fill_2 FILLER_19_598 ();
 sg13g2_fill_1 FILLER_19_600 ();
 sg13g2_fill_2 FILLER_19_611 ();
 sg13g2_fill_1 FILLER_19_613 ();
 sg13g2_fill_1 FILLER_19_640 ();
 sg13g2_fill_2 FILLER_19_645 ();
 sg13g2_fill_1 FILLER_19_647 ();
 sg13g2_fill_1 FILLER_19_663 ();
 sg13g2_fill_1 FILLER_19_690 ();
 sg13g2_decap_4 FILLER_19_757 ();
 sg13g2_decap_8 FILLER_19_787 ();
 sg13g2_fill_2 FILLER_19_794 ();
 sg13g2_decap_4 FILLER_19_822 ();
 sg13g2_fill_1 FILLER_19_826 ();
 sg13g2_decap_8 FILLER_19_848 ();
 sg13g2_decap_8 FILLER_19_855 ();
 sg13g2_decap_8 FILLER_19_862 ();
 sg13g2_decap_4 FILLER_19_872 ();
 sg13g2_fill_1 FILLER_19_876 ();
 sg13g2_fill_2 FILLER_19_887 ();
 sg13g2_fill_1 FILLER_19_889 ();
 sg13g2_fill_2 FILLER_19_918 ();
 sg13g2_decap_8 FILLER_19_956 ();
 sg13g2_decap_4 FILLER_19_963 ();
 sg13g2_fill_1 FILLER_19_967 ();
 sg13g2_fill_2 FILLER_19_977 ();
 sg13g2_decap_8 FILLER_19_1005 ();
 sg13g2_fill_2 FILLER_19_1016 ();
 sg13g2_fill_1 FILLER_19_1018 ();
 sg13g2_decap_4 FILLER_19_1027 ();
 sg13g2_decap_8 FILLER_19_1044 ();
 sg13g2_fill_1 FILLER_19_1051 ();
 sg13g2_fill_2 FILLER_19_1109 ();
 sg13g2_decap_8 FILLER_19_1115 ();
 sg13g2_decap_4 FILLER_19_1122 ();
 sg13g2_fill_1 FILLER_19_1126 ();
 sg13g2_fill_1 FILLER_19_1158 ();
 sg13g2_fill_1 FILLER_19_1173 ();
 sg13g2_fill_2 FILLER_19_1209 ();
 sg13g2_fill_1 FILLER_19_1211 ();
 sg13g2_decap_8 FILLER_19_1242 ();
 sg13g2_decap_8 FILLER_19_1249 ();
 sg13g2_fill_2 FILLER_19_1260 ();
 sg13g2_fill_2 FILLER_19_1275 ();
 sg13g2_fill_2 FILLER_19_1293 ();
 sg13g2_fill_1 FILLER_19_1309 ();
 sg13g2_fill_2 FILLER_19_1315 ();
 sg13g2_fill_1 FILLER_19_1321 ();
 sg13g2_decap_4 FILLER_19_1326 ();
 sg13g2_fill_2 FILLER_19_1339 ();
 sg13g2_fill_2 FILLER_19_1409 ();
 sg13g2_fill_1 FILLER_19_1411 ();
 sg13g2_fill_1 FILLER_19_1415 ();
 sg13g2_fill_2 FILLER_19_1471 ();
 sg13g2_fill_2 FILLER_19_1477 ();
 sg13g2_fill_1 FILLER_19_1494 ();
 sg13g2_fill_2 FILLER_19_1521 ();
 sg13g2_fill_1 FILLER_19_1574 ();
 sg13g2_fill_1 FILLER_19_1583 ();
 sg13g2_fill_2 FILLER_19_1596 ();
 sg13g2_fill_1 FILLER_19_1598 ();
 sg13g2_fill_1 FILLER_19_1629 ();
 sg13g2_fill_2 FILLER_19_1645 ();
 sg13g2_fill_2 FILLER_19_1651 ();
 sg13g2_decap_4 FILLER_19_1657 ();
 sg13g2_fill_2 FILLER_19_1661 ();
 sg13g2_decap_8 FILLER_19_1668 ();
 sg13g2_fill_1 FILLER_19_1675 ();
 sg13g2_fill_2 FILLER_19_1680 ();
 sg13g2_fill_1 FILLER_19_1682 ();
 sg13g2_fill_1 FILLER_19_1733 ();
 sg13g2_decap_8 FILLER_19_1738 ();
 sg13g2_fill_2 FILLER_19_1745 ();
 sg13g2_fill_1 FILLER_19_1747 ();
 sg13g2_decap_4 FILLER_19_1754 ();
 sg13g2_fill_1 FILLER_19_1758 ();
 sg13g2_decap_8 FILLER_19_1789 ();
 sg13g2_decap_8 FILLER_19_1796 ();
 sg13g2_decap_4 FILLER_19_1803 ();
 sg13g2_fill_2 FILLER_19_1807 ();
 sg13g2_decap_8 FILLER_19_1812 ();
 sg13g2_fill_1 FILLER_19_1860 ();
 sg13g2_fill_1 FILLER_19_1869 ();
 sg13g2_decap_4 FILLER_19_1901 ();
 sg13g2_fill_2 FILLER_19_1905 ();
 sg13g2_decap_4 FILLER_19_1945 ();
 sg13g2_fill_1 FILLER_19_1949 ();
 sg13g2_fill_1 FILLER_19_1964 ();
 sg13g2_decap_4 FILLER_19_1995 ();
 sg13g2_fill_1 FILLER_19_2034 ();
 sg13g2_fill_1 FILLER_19_2081 ();
 sg13g2_decap_4 FILLER_19_2096 ();
 sg13g2_fill_2 FILLER_19_2125 ();
 sg13g2_fill_2 FILLER_19_2134 ();
 sg13g2_decap_8 FILLER_19_2140 ();
 sg13g2_decap_8 FILLER_19_2147 ();
 sg13g2_fill_2 FILLER_19_2154 ();
 sg13g2_fill_1 FILLER_19_2156 ();
 sg13g2_decap_8 FILLER_19_2193 ();
 sg13g2_decap_8 FILLER_19_2200 ();
 sg13g2_decap_4 FILLER_19_2207 ();
 sg13g2_fill_2 FILLER_19_2275 ();
 sg13g2_decap_8 FILLER_19_2298 ();
 sg13g2_decap_8 FILLER_19_2305 ();
 sg13g2_decap_8 FILLER_19_2312 ();
 sg13g2_fill_2 FILLER_19_2319 ();
 sg13g2_fill_1 FILLER_19_2321 ();
 sg13g2_decap_8 FILLER_19_2336 ();
 sg13g2_decap_8 FILLER_19_2343 ();
 sg13g2_decap_8 FILLER_19_2350 ();
 sg13g2_decap_4 FILLER_19_2357 ();
 sg13g2_fill_1 FILLER_19_2361 ();
 sg13g2_fill_2 FILLER_19_2388 ();
 sg13g2_fill_1 FILLER_19_2390 ();
 sg13g2_decap_8 FILLER_19_2404 ();
 sg13g2_decap_8 FILLER_19_2425 ();
 sg13g2_decap_8 FILLER_19_2432 ();
 sg13g2_fill_2 FILLER_19_2445 ();
 sg13g2_decap_8 FILLER_19_2451 ();
 sg13g2_decap_4 FILLER_19_2458 ();
 sg13g2_decap_4 FILLER_19_2472 ();
 sg13g2_fill_2 FILLER_19_2476 ();
 sg13g2_fill_1 FILLER_19_2482 ();
 sg13g2_fill_2 FILLER_19_2532 ();
 sg13g2_decap_8 FILLER_19_2564 ();
 sg13g2_decap_4 FILLER_19_2571 ();
 sg13g2_fill_2 FILLER_19_2575 ();
 sg13g2_decap_8 FILLER_19_2581 ();
 sg13g2_decap_8 FILLER_19_2588 ();
 sg13g2_decap_8 FILLER_19_2595 ();
 sg13g2_decap_8 FILLER_19_2602 ();
 sg13g2_fill_2 FILLER_19_2609 ();
 sg13g2_fill_1 FILLER_19_2611 ();
 sg13g2_fill_1 FILLER_19_2616 ();
 sg13g2_decap_8 FILLER_19_2622 ();
 sg13g2_decap_8 FILLER_19_2629 ();
 sg13g2_decap_8 FILLER_19_2636 ();
 sg13g2_decap_8 FILLER_19_2643 ();
 sg13g2_decap_8 FILLER_19_2650 ();
 sg13g2_decap_8 FILLER_19_2657 ();
 sg13g2_decap_4 FILLER_19_2664 ();
 sg13g2_fill_2 FILLER_19_2668 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_28 ();
 sg13g2_fill_1 FILLER_20_55 ();
 sg13g2_fill_2 FILLER_20_61 ();
 sg13g2_fill_1 FILLER_20_63 ();
 sg13g2_decap_4 FILLER_20_68 ();
 sg13g2_fill_1 FILLER_20_72 ();
 sg13g2_decap_8 FILLER_20_130 ();
 sg13g2_decap_8 FILLER_20_137 ();
 sg13g2_fill_1 FILLER_20_181 ();
 sg13g2_fill_2 FILLER_20_208 ();
 sg13g2_fill_1 FILLER_20_214 ();
 sg13g2_fill_2 FILLER_20_222 ();
 sg13g2_fill_2 FILLER_20_229 ();
 sg13g2_fill_1 FILLER_20_231 ();
 sg13g2_fill_1 FILLER_20_266 ();
 sg13g2_fill_2 FILLER_20_271 ();
 sg13g2_fill_2 FILLER_20_277 ();
 sg13g2_decap_8 FILLER_20_283 ();
 sg13g2_fill_2 FILLER_20_290 ();
 sg13g2_decap_4 FILLER_20_324 ();
 sg13g2_fill_1 FILLER_20_328 ();
 sg13g2_fill_1 FILLER_20_339 ();
 sg13g2_fill_2 FILLER_20_366 ();
 sg13g2_fill_1 FILLER_20_368 ();
 sg13g2_decap_8 FILLER_20_373 ();
 sg13g2_decap_8 FILLER_20_380 ();
 sg13g2_decap_8 FILLER_20_387 ();
 sg13g2_fill_1 FILLER_20_394 ();
 sg13g2_decap_4 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_403 ();
 sg13g2_fill_2 FILLER_20_409 ();
 sg13g2_fill_1 FILLER_20_427 ();
 sg13g2_fill_2 FILLER_20_443 ();
 sg13g2_fill_1 FILLER_20_450 ();
 sg13g2_fill_1 FILLER_20_461 ();
 sg13g2_fill_1 FILLER_20_467 ();
 sg13g2_fill_1 FILLER_20_472 ();
 sg13g2_fill_2 FILLER_20_478 ();
 sg13g2_fill_1 FILLER_20_480 ();
 sg13g2_fill_2 FILLER_20_548 ();
 sg13g2_fill_2 FILLER_20_555 ();
 sg13g2_fill_1 FILLER_20_562 ();
 sg13g2_fill_1 FILLER_20_569 ();
 sg13g2_fill_2 FILLER_20_580 ();
 sg13g2_fill_1 FILLER_20_582 ();
 sg13g2_decap_8 FILLER_20_603 ();
 sg13g2_decap_8 FILLER_20_610 ();
 sg13g2_decap_4 FILLER_20_617 ();
 sg13g2_fill_2 FILLER_20_625 ();
 sg13g2_fill_1 FILLER_20_627 ();
 sg13g2_decap_4 FILLER_20_636 ();
 sg13g2_fill_1 FILLER_20_651 ();
 sg13g2_decap_4 FILLER_20_662 ();
 sg13g2_fill_2 FILLER_20_670 ();
 sg13g2_fill_1 FILLER_20_692 ();
 sg13g2_decap_8 FILLER_20_697 ();
 sg13g2_decap_4 FILLER_20_709 ();
 sg13g2_fill_2 FILLER_20_713 ();
 sg13g2_decap_4 FILLER_20_849 ();
 sg13g2_fill_2 FILLER_20_853 ();
 sg13g2_fill_1 FILLER_20_885 ();
 sg13g2_fill_1 FILLER_20_890 ();
 sg13g2_fill_1 FILLER_20_901 ();
 sg13g2_fill_2 FILLER_20_906 ();
 sg13g2_decap_4 FILLER_20_933 ();
 sg13g2_fill_1 FILLER_20_937 ();
 sg13g2_decap_8 FILLER_20_942 ();
 sg13g2_fill_2 FILLER_20_949 ();
 sg13g2_fill_1 FILLER_20_951 ();
 sg13g2_fill_1 FILLER_20_978 ();
 sg13g2_fill_2 FILLER_20_983 ();
 sg13g2_fill_2 FILLER_20_989 ();
 sg13g2_fill_2 FILLER_20_995 ();
 sg13g2_fill_2 FILLER_20_1028 ();
 sg13g2_fill_1 FILLER_20_1030 ();
 sg13g2_fill_1 FILLER_20_1036 ();
 sg13g2_fill_2 FILLER_20_1097 ();
 sg13g2_fill_1 FILLER_20_1099 ();
 sg13g2_fill_2 FILLER_20_1131 ();
 sg13g2_fill_1 FILLER_20_1173 ();
 sg13g2_fill_2 FILLER_20_1218 ();
 sg13g2_fill_2 FILLER_20_1256 ();
 sg13g2_fill_2 FILLER_20_1289 ();
 sg13g2_fill_1 FILLER_20_1291 ();
 sg13g2_fill_1 FILLER_20_1308 ();
 sg13g2_decap_8 FILLER_20_1314 ();
 sg13g2_decap_8 FILLER_20_1321 ();
 sg13g2_decap_8 FILLER_20_1328 ();
 sg13g2_decap_4 FILLER_20_1335 ();
 sg13g2_fill_2 FILLER_20_1345 ();
 sg13g2_fill_2 FILLER_20_1351 ();
 sg13g2_decap_8 FILLER_20_1357 ();
 sg13g2_fill_1 FILLER_20_1364 ();
 sg13g2_decap_8 FILLER_20_1369 ();
 sg13g2_fill_2 FILLER_20_1376 ();
 sg13g2_fill_1 FILLER_20_1378 ();
 sg13g2_fill_2 FILLER_20_1389 ();
 sg13g2_fill_2 FILLER_20_1409 ();
 sg13g2_fill_2 FILLER_20_1424 ();
 sg13g2_fill_2 FILLER_20_1432 ();
 sg13g2_fill_2 FILLER_20_1438 ();
 sg13g2_fill_2 FILLER_20_1481 ();
 sg13g2_fill_1 FILLER_20_1512 ();
 sg13g2_fill_2 FILLER_20_1518 ();
 sg13g2_fill_1 FILLER_20_1524 ();
 sg13g2_fill_2 FILLER_20_1542 ();
 sg13g2_fill_1 FILLER_20_1548 ();
 sg13g2_fill_2 FILLER_20_1559 ();
 sg13g2_decap_8 FILLER_20_1568 ();
 sg13g2_fill_2 FILLER_20_1575 ();
 sg13g2_fill_2 FILLER_20_1586 ();
 sg13g2_fill_1 FILLER_20_1588 ();
 sg13g2_fill_2 FILLER_20_1598 ();
 sg13g2_fill_2 FILLER_20_1605 ();
 sg13g2_fill_1 FILLER_20_1607 ();
 sg13g2_fill_2 FILLER_20_1634 ();
 sg13g2_fill_1 FILLER_20_1636 ();
 sg13g2_fill_2 FILLER_20_1647 ();
 sg13g2_decap_8 FILLER_20_1653 ();
 sg13g2_decap_8 FILLER_20_1660 ();
 sg13g2_decap_8 FILLER_20_1667 ();
 sg13g2_decap_8 FILLER_20_1674 ();
 sg13g2_fill_1 FILLER_20_1681 ();
 sg13g2_decap_4 FILLER_20_1703 ();
 sg13g2_fill_1 FILLER_20_1707 ();
 sg13g2_decap_8 FILLER_20_1744 ();
 sg13g2_decap_8 FILLER_20_1751 ();
 sg13g2_fill_2 FILLER_20_1758 ();
 sg13g2_fill_1 FILLER_20_1760 ();
 sg13g2_fill_1 FILLER_20_1775 ();
 sg13g2_fill_1 FILLER_20_1786 ();
 sg13g2_fill_1 FILLER_20_1791 ();
 sg13g2_decap_8 FILLER_20_1818 ();
 sg13g2_decap_4 FILLER_20_1825 ();
 sg13g2_fill_2 FILLER_20_1829 ();
 sg13g2_fill_2 FILLER_20_1843 ();
 sg13g2_fill_1 FILLER_20_1853 ();
 sg13g2_fill_2 FILLER_20_1864 ();
 sg13g2_fill_2 FILLER_20_1870 ();
 sg13g2_fill_1 FILLER_20_1872 ();
 sg13g2_fill_1 FILLER_20_1899 ();
 sg13g2_fill_2 FILLER_20_1926 ();
 sg13g2_fill_1 FILLER_20_1928 ();
 sg13g2_fill_2 FILLER_20_2005 ();
 sg13g2_fill_1 FILLER_20_2017 ();
 sg13g2_fill_2 FILLER_20_2073 ();
 sg13g2_decap_4 FILLER_20_2134 ();
 sg13g2_fill_1 FILLER_20_2138 ();
 sg13g2_decap_8 FILLER_20_2153 ();
 sg13g2_fill_2 FILLER_20_2160 ();
 sg13g2_fill_1 FILLER_20_2162 ();
 sg13g2_decap_8 FILLER_20_2167 ();
 sg13g2_fill_2 FILLER_20_2199 ();
 sg13g2_fill_1 FILLER_20_2201 ();
 sg13g2_decap_8 FILLER_20_2226 ();
 sg13g2_decap_4 FILLER_20_2269 ();
 sg13g2_fill_2 FILLER_20_2273 ();
 sg13g2_decap_8 FILLER_20_2305 ();
 sg13g2_decap_8 FILLER_20_2312 ();
 sg13g2_decap_8 FILLER_20_2319 ();
 sg13g2_decap_8 FILLER_20_2326 ();
 sg13g2_decap_4 FILLER_20_2395 ();
 sg13g2_fill_2 FILLER_20_2399 ();
 sg13g2_decap_8 FILLER_20_2437 ();
 sg13g2_decap_8 FILLER_20_2444 ();
 sg13g2_decap_8 FILLER_20_2451 ();
 sg13g2_fill_1 FILLER_20_2458 ();
 sg13g2_fill_2 FILLER_20_2499 ();
 sg13g2_fill_1 FILLER_20_2501 ();
 sg13g2_fill_2 FILLER_20_2512 ();
 sg13g2_fill_1 FILLER_20_2524 ();
 sg13g2_fill_1 FILLER_20_2543 ();
 sg13g2_decap_8 FILLER_20_2554 ();
 sg13g2_fill_2 FILLER_20_2561 ();
 sg13g2_fill_1 FILLER_20_2563 ();
 sg13g2_fill_2 FILLER_20_2615 ();
 sg13g2_decap_8 FILLER_20_2657 ();
 sg13g2_decap_4 FILLER_20_2664 ();
 sg13g2_fill_2 FILLER_20_2668 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_7 ();
 sg13g2_fill_1 FILLER_21_43 ();
 sg13g2_fill_2 FILLER_21_63 ();
 sg13g2_fill_2 FILLER_21_69 ();
 sg13g2_fill_1 FILLER_21_71 ();
 sg13g2_fill_1 FILLER_21_85 ();
 sg13g2_fill_1 FILLER_21_96 ();
 sg13g2_fill_1 FILLER_21_103 ();
 sg13g2_fill_1 FILLER_21_108 ();
 sg13g2_fill_1 FILLER_21_135 ();
 sg13g2_fill_2 FILLER_21_142 ();
 sg13g2_fill_1 FILLER_21_144 ();
 sg13g2_fill_1 FILLER_21_158 ();
 sg13g2_decap_8 FILLER_21_179 ();
 sg13g2_fill_1 FILLER_21_186 ();
 sg13g2_fill_2 FILLER_21_191 ();
 sg13g2_fill_1 FILLER_21_193 ();
 sg13g2_fill_1 FILLER_21_199 ();
 sg13g2_fill_2 FILLER_21_205 ();
 sg13g2_fill_2 FILLER_21_212 ();
 sg13g2_fill_1 FILLER_21_250 ();
 sg13g2_decap_4 FILLER_21_268 ();
 sg13g2_decap_8 FILLER_21_276 ();
 sg13g2_fill_2 FILLER_21_283 ();
 sg13g2_fill_1 FILLER_21_285 ();
 sg13g2_decap_4 FILLER_21_306 ();
 sg13g2_decap_4 FILLER_21_334 ();
 sg13g2_decap_4 FILLER_21_342 ();
 sg13g2_fill_2 FILLER_21_356 ();
 sg13g2_fill_2 FILLER_21_384 ();
 sg13g2_fill_2 FILLER_21_412 ();
 sg13g2_fill_2 FILLER_21_427 ();
 sg13g2_decap_8 FILLER_21_469 ();
 sg13g2_fill_2 FILLER_21_476 ();
 sg13g2_decap_4 FILLER_21_482 ();
 sg13g2_fill_2 FILLER_21_490 ();
 sg13g2_fill_1 FILLER_21_504 ();
 sg13g2_fill_1 FILLER_21_537 ();
 sg13g2_fill_2 FILLER_21_552 ();
 sg13g2_decap_4 FILLER_21_558 ();
 sg13g2_decap_4 FILLER_21_567 ();
 sg13g2_fill_2 FILLER_21_576 ();
 sg13g2_decap_4 FILLER_21_608 ();
 sg13g2_decap_8 FILLER_21_617 ();
 sg13g2_decap_4 FILLER_21_624 ();
 sg13g2_fill_1 FILLER_21_628 ();
 sg13g2_fill_2 FILLER_21_633 ();
 sg13g2_fill_2 FILLER_21_644 ();
 sg13g2_fill_1 FILLER_21_646 ();
 sg13g2_decap_4 FILLER_21_651 ();
 sg13g2_fill_2 FILLER_21_666 ();
 sg13g2_fill_2 FILLER_21_677 ();
 sg13g2_fill_1 FILLER_21_679 ();
 sg13g2_fill_2 FILLER_21_710 ();
 sg13g2_fill_1 FILLER_21_712 ();
 sg13g2_fill_2 FILLER_21_718 ();
 sg13g2_fill_2 FILLER_21_724 ();
 sg13g2_fill_1 FILLER_21_731 ();
 sg13g2_fill_2 FILLER_21_736 ();
 sg13g2_fill_2 FILLER_21_742 ();
 sg13g2_fill_2 FILLER_21_748 ();
 sg13g2_fill_1 FILLER_21_750 ();
 sg13g2_fill_2 FILLER_21_755 ();
 sg13g2_fill_1 FILLER_21_757 ();
 sg13g2_fill_2 FILLER_21_827 ();
 sg13g2_fill_1 FILLER_21_855 ();
 sg13g2_fill_1 FILLER_21_860 ();
 sg13g2_fill_1 FILLER_21_887 ();
 sg13g2_fill_2 FILLER_21_914 ();
 sg13g2_decap_8 FILLER_21_990 ();
 sg13g2_fill_2 FILLER_21_997 ();
 sg13g2_fill_1 FILLER_21_999 ();
 sg13g2_decap_4 FILLER_21_1009 ();
 sg13g2_decap_4 FILLER_21_1039 ();
 sg13g2_fill_1 FILLER_21_1043 ();
 sg13g2_decap_4 FILLER_21_1048 ();
 sg13g2_fill_1 FILLER_21_1065 ();
 sg13g2_fill_2 FILLER_21_1071 ();
 sg13g2_fill_1 FILLER_21_1073 ();
 sg13g2_fill_1 FILLER_21_1110 ();
 sg13g2_fill_1 FILLER_21_1201 ();
 sg13g2_fill_2 FILLER_21_1215 ();
 sg13g2_decap_8 FILLER_21_1263 ();
 sg13g2_fill_2 FILLER_21_1270 ();
 sg13g2_fill_1 FILLER_21_1272 ();
 sg13g2_decap_8 FILLER_21_1317 ();
 sg13g2_fill_2 FILLER_21_1324 ();
 sg13g2_fill_1 FILLER_21_1326 ();
 sg13g2_fill_1 FILLER_21_1336 ();
 sg13g2_decap_8 FILLER_21_1343 ();
 sg13g2_decap_4 FILLER_21_1350 ();
 sg13g2_fill_2 FILLER_21_1362 ();
 sg13g2_fill_2 FILLER_21_1374 ();
 sg13g2_fill_1 FILLER_21_1376 ();
 sg13g2_fill_2 FILLER_21_1433 ();
 sg13g2_fill_1 FILLER_21_1465 ();
 sg13g2_fill_1 FILLER_21_1508 ();
 sg13g2_fill_2 FILLER_21_1524 ();
 sg13g2_fill_1 FILLER_21_1551 ();
 sg13g2_fill_1 FILLER_21_1556 ();
 sg13g2_fill_2 FILLER_21_1561 ();
 sg13g2_fill_1 FILLER_21_1563 ();
 sg13g2_fill_2 FILLER_21_1568 ();
 sg13g2_fill_1 FILLER_21_1570 ();
 sg13g2_fill_2 FILLER_21_1576 ();
 sg13g2_fill_2 FILLER_21_1630 ();
 sg13g2_fill_2 FILLER_21_1751 ();
 sg13g2_fill_1 FILLER_21_1763 ();
 sg13g2_decap_4 FILLER_21_1819 ();
 sg13g2_fill_1 FILLER_21_1831 ();
 sg13g2_decap_4 FILLER_21_1842 ();
 sg13g2_fill_1 FILLER_21_1856 ();
 sg13g2_decap_4 FILLER_21_1889 ();
 sg13g2_fill_2 FILLER_21_1893 ();
 sg13g2_fill_2 FILLER_21_1905 ();
 sg13g2_decap_8 FILLER_21_1947 ();
 sg13g2_decap_4 FILLER_21_1954 ();
 sg13g2_fill_1 FILLER_21_1958 ();
 sg13g2_fill_2 FILLER_21_1973 ();
 sg13g2_fill_1 FILLER_21_1975 ();
 sg13g2_fill_2 FILLER_21_2020 ();
 sg13g2_fill_1 FILLER_21_2022 ();
 sg13g2_fill_2 FILLER_21_2058 ();
 sg13g2_decap_4 FILLER_21_2064 ();
 sg13g2_fill_2 FILLER_21_2068 ();
 sg13g2_decap_4 FILLER_21_2080 ();
 sg13g2_fill_2 FILLER_21_2127 ();
 sg13g2_fill_1 FILLER_21_2129 ();
 sg13g2_decap_8 FILLER_21_2147 ();
 sg13g2_fill_2 FILLER_21_2210 ();
 sg13g2_fill_1 FILLER_21_2212 ();
 sg13g2_decap_8 FILLER_21_2226 ();
 sg13g2_decap_8 FILLER_21_2233 ();
 sg13g2_decap_8 FILLER_21_2240 ();
 sg13g2_decap_4 FILLER_21_2247 ();
 sg13g2_fill_1 FILLER_21_2255 ();
 sg13g2_decap_4 FILLER_21_2260 ();
 sg13g2_fill_1 FILLER_21_2300 ();
 sg13g2_fill_2 FILLER_21_2311 ();
 sg13g2_fill_1 FILLER_21_2313 ();
 sg13g2_decap_8 FILLER_21_2324 ();
 sg13g2_decap_8 FILLER_21_2331 ();
 sg13g2_fill_2 FILLER_21_2356 ();
 sg13g2_fill_1 FILLER_21_2362 ();
 sg13g2_fill_2 FILLER_21_2373 ();
 sg13g2_fill_1 FILLER_21_2379 ();
 sg13g2_fill_2 FILLER_21_2384 ();
 sg13g2_fill_2 FILLER_21_2390 ();
 sg13g2_fill_2 FILLER_21_2397 ();
 sg13g2_fill_2 FILLER_21_2403 ();
 sg13g2_fill_2 FILLER_21_2411 ();
 sg13g2_fill_1 FILLER_21_2413 ();
 sg13g2_decap_8 FILLER_21_2423 ();
 sg13g2_fill_2 FILLER_21_2430 ();
 sg13g2_decap_8 FILLER_21_2458 ();
 sg13g2_decap_8 FILLER_21_2465 ();
 sg13g2_decap_8 FILLER_21_2472 ();
 sg13g2_fill_2 FILLER_21_2479 ();
 sg13g2_fill_1 FILLER_21_2481 ();
 sg13g2_fill_2 FILLER_21_2492 ();
 sg13g2_decap_4 FILLER_21_2498 ();
 sg13g2_fill_2 FILLER_21_2502 ();
 sg13g2_decap_4 FILLER_21_2510 ();
 sg13g2_fill_1 FILLER_21_2514 ();
 sg13g2_decap_8 FILLER_21_2541 ();
 sg13g2_decap_4 FILLER_21_2548 ();
 sg13g2_fill_1 FILLER_21_2552 ();
 sg13g2_fill_1 FILLER_21_2563 ();
 sg13g2_fill_2 FILLER_21_2568 ();
 sg13g2_decap_8 FILLER_21_2610 ();
 sg13g2_fill_1 FILLER_21_2617 ();
 sg13g2_decap_8 FILLER_21_2662 ();
 sg13g2_fill_1 FILLER_21_2669 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_fill_1 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_73 ();
 sg13g2_decap_8 FILLER_22_80 ();
 sg13g2_decap_8 FILLER_22_87 ();
 sg13g2_decap_8 FILLER_22_94 ();
 sg13g2_decap_4 FILLER_22_101 ();
 sg13g2_fill_2 FILLER_22_105 ();
 sg13g2_fill_1 FILLER_22_120 ();
 sg13g2_fill_2 FILLER_22_135 ();
 sg13g2_fill_1 FILLER_22_163 ();
 sg13g2_fill_2 FILLER_22_169 ();
 sg13g2_fill_1 FILLER_22_171 ();
 sg13g2_decap_8 FILLER_22_177 ();
 sg13g2_decap_8 FILLER_22_184 ();
 sg13g2_fill_1 FILLER_22_191 ();
 sg13g2_fill_1 FILLER_22_200 ();
 sg13g2_fill_2 FILLER_22_206 ();
 sg13g2_fill_1 FILLER_22_212 ();
 sg13g2_fill_2 FILLER_22_221 ();
 sg13g2_fill_2 FILLER_22_227 ();
 sg13g2_fill_2 FILLER_22_238 ();
 sg13g2_fill_1 FILLER_22_252 ();
 sg13g2_fill_2 FILLER_22_262 ();
 sg13g2_decap_8 FILLER_22_295 ();
 sg13g2_decap_8 FILLER_22_302 ();
 sg13g2_decap_4 FILLER_22_309 ();
 sg13g2_decap_4 FILLER_22_344 ();
 sg13g2_fill_1 FILLER_22_348 ();
 sg13g2_decap_8 FILLER_22_359 ();
 sg13g2_decap_8 FILLER_22_366 ();
 sg13g2_decap_8 FILLER_22_373 ();
 sg13g2_fill_2 FILLER_22_398 ();
 sg13g2_fill_2 FILLER_22_426 ();
 sg13g2_fill_2 FILLER_22_431 ();
 sg13g2_fill_1 FILLER_22_456 ();
 sg13g2_fill_2 FILLER_22_461 ();
 sg13g2_decap_8 FILLER_22_473 ();
 sg13g2_decap_8 FILLER_22_480 ();
 sg13g2_decap_8 FILLER_22_506 ();
 sg13g2_decap_4 FILLER_22_516 ();
 sg13g2_fill_1 FILLER_22_525 ();
 sg13g2_fill_2 FILLER_22_563 ();
 sg13g2_fill_1 FILLER_22_565 ();
 sg13g2_fill_2 FILLER_22_576 ();
 sg13g2_fill_2 FILLER_22_604 ();
 sg13g2_fill_1 FILLER_22_606 ();
 sg13g2_fill_1 FILLER_22_633 ();
 sg13g2_fill_2 FILLER_22_660 ();
 sg13g2_fill_1 FILLER_22_662 ();
 sg13g2_fill_2 FILLER_22_667 ();
 sg13g2_decap_8 FILLER_22_678 ();
 sg13g2_decap_8 FILLER_22_685 ();
 sg13g2_decap_4 FILLER_22_692 ();
 sg13g2_fill_2 FILLER_22_696 ();
 sg13g2_decap_4 FILLER_22_722 ();
 sg13g2_decap_8 FILLER_22_730 ();
 sg13g2_decap_8 FILLER_22_737 ();
 sg13g2_fill_2 FILLER_22_744 ();
 sg13g2_fill_1 FILLER_22_746 ();
 sg13g2_decap_8 FILLER_22_757 ();
 sg13g2_fill_2 FILLER_22_764 ();
 sg13g2_fill_1 FILLER_22_766 ();
 sg13g2_fill_2 FILLER_22_771 ();
 sg13g2_fill_2 FILLER_22_840 ();
 sg13g2_fill_1 FILLER_22_842 ();
 sg13g2_fill_2 FILLER_22_872 ();
 sg13g2_fill_2 FILLER_22_895 ();
 sg13g2_decap_8 FILLER_22_953 ();
 sg13g2_fill_1 FILLER_22_964 ();
 sg13g2_decap_8 FILLER_22_969 ();
 sg13g2_decap_4 FILLER_22_976 ();
 sg13g2_fill_1 FILLER_22_980 ();
 sg13g2_fill_1 FILLER_22_1016 ();
 sg13g2_decap_8 FILLER_22_1021 ();
 sg13g2_decap_8 FILLER_22_1028 ();
 sg13g2_fill_2 FILLER_22_1035 ();
 sg13g2_fill_1 FILLER_22_1037 ();
 sg13g2_decap_4 FILLER_22_1042 ();
 sg13g2_fill_1 FILLER_22_1050 ();
 sg13g2_fill_2 FILLER_22_1056 ();
 sg13g2_fill_1 FILLER_22_1058 ();
 sg13g2_fill_2 FILLER_22_1123 ();
 sg13g2_fill_1 FILLER_22_1125 ();
 sg13g2_fill_1 FILLER_22_1131 ();
 sg13g2_fill_1 FILLER_22_1184 ();
 sg13g2_decap_4 FILLER_22_1232 ();
 sg13g2_decap_8 FILLER_22_1257 ();
 sg13g2_fill_2 FILLER_22_1264 ();
 sg13g2_fill_1 FILLER_22_1266 ();
 sg13g2_decap_8 FILLER_22_1276 ();
 sg13g2_decap_8 FILLER_22_1283 ();
 sg13g2_fill_2 FILLER_22_1290 ();
 sg13g2_decap_4 FILLER_22_1318 ();
 sg13g2_fill_2 FILLER_22_1322 ();
 sg13g2_fill_2 FILLER_22_1334 ();
 sg13g2_decap_4 FILLER_22_1340 ();
 sg13g2_fill_1 FILLER_22_1361 ();
 sg13g2_fill_2 FILLER_22_1370 ();
 sg13g2_fill_1 FILLER_22_1372 ();
 sg13g2_fill_1 FILLER_22_1427 ();
 sg13g2_fill_2 FILLER_22_1486 ();
 sg13g2_fill_2 FILLER_22_1504 ();
 sg13g2_fill_1 FILLER_22_1562 ();
 sg13g2_fill_1 FILLER_22_1612 ();
 sg13g2_fill_1 FILLER_22_1617 ();
 sg13g2_decap_8 FILLER_22_1689 ();
 sg13g2_decap_8 FILLER_22_1696 ();
 sg13g2_decap_8 FILLER_22_1703 ();
 sg13g2_decap_8 FILLER_22_1710 ();
 sg13g2_fill_1 FILLER_22_1717 ();
 sg13g2_decap_8 FILLER_22_1739 ();
 sg13g2_decap_4 FILLER_22_1746 ();
 sg13g2_fill_1 FILLER_22_1784 ();
 sg13g2_fill_1 FILLER_22_1795 ();
 sg13g2_fill_1 FILLER_22_1800 ();
 sg13g2_decap_4 FILLER_22_1805 ();
 sg13g2_fill_2 FILLER_22_1809 ();
 sg13g2_fill_2 FILLER_22_1825 ();
 sg13g2_fill_2 FILLER_22_1853 ();
 sg13g2_fill_2 FILLER_22_1896 ();
 sg13g2_fill_1 FILLER_22_1898 ();
 sg13g2_decap_8 FILLER_22_1923 ();
 sg13g2_decap_8 FILLER_22_1930 ();
 sg13g2_fill_1 FILLER_22_1937 ();
 sg13g2_decap_4 FILLER_22_1942 ();
 sg13g2_decap_8 FILLER_22_1949 ();
 sg13g2_decap_8 FILLER_22_1956 ();
 sg13g2_fill_2 FILLER_22_1963 ();
 sg13g2_fill_1 FILLER_22_1965 ();
 sg13g2_decap_8 FILLER_22_1974 ();
 sg13g2_fill_1 FILLER_22_1981 ();
 sg13g2_fill_1 FILLER_22_2010 ();
 sg13g2_decap_8 FILLER_22_2037 ();
 sg13g2_decap_4 FILLER_22_2044 ();
 sg13g2_fill_2 FILLER_22_2048 ();
 sg13g2_decap_8 FILLER_22_2054 ();
 sg13g2_fill_1 FILLER_22_2061 ();
 sg13g2_fill_2 FILLER_22_2072 ();
 sg13g2_decap_8 FILLER_22_2078 ();
 sg13g2_fill_1 FILLER_22_2085 ();
 sg13g2_fill_1 FILLER_22_2096 ();
 sg13g2_fill_2 FILLER_22_2107 ();
 sg13g2_decap_8 FILLER_22_2113 ();
 sg13g2_fill_1 FILLER_22_2146 ();
 sg13g2_fill_2 FILLER_22_2173 ();
 sg13g2_fill_2 FILLER_22_2196 ();
 sg13g2_fill_2 FILLER_22_2202 ();
 sg13g2_decap_8 FILLER_22_2244 ();
 sg13g2_decap_8 FILLER_22_2251 ();
 sg13g2_decap_8 FILLER_22_2258 ();
 sg13g2_decap_4 FILLER_22_2265 ();
 sg13g2_fill_1 FILLER_22_2269 ();
 sg13g2_decap_8 FILLER_22_2274 ();
 sg13g2_decap_4 FILLER_22_2281 ();
 sg13g2_fill_2 FILLER_22_2285 ();
 sg13g2_fill_1 FILLER_22_2297 ();
 sg13g2_decap_8 FILLER_22_2329 ();
 sg13g2_decap_4 FILLER_22_2336 ();
 sg13g2_decap_4 FILLER_22_2376 ();
 sg13g2_fill_1 FILLER_22_2380 ();
 sg13g2_fill_1 FILLER_22_2441 ();
 sg13g2_decap_8 FILLER_22_2472 ();
 sg13g2_fill_1 FILLER_22_2479 ();
 sg13g2_fill_1 FILLER_22_2484 ();
 sg13g2_decap_8 FILLER_22_2509 ();
 sg13g2_decap_4 FILLER_22_2516 ();
 sg13g2_fill_2 FILLER_22_2524 ();
 sg13g2_fill_1 FILLER_22_2526 ();
 sg13g2_fill_2 FILLER_22_2551 ();
 sg13g2_fill_2 FILLER_22_2589 ();
 sg13g2_decap_4 FILLER_22_2601 ();
 sg13g2_decap_4 FILLER_22_2621 ();
 sg13g2_fill_1 FILLER_22_2625 ();
 sg13g2_fill_2 FILLER_22_2636 ();
 sg13g2_fill_1 FILLER_22_2638 ();
 sg13g2_fill_1 FILLER_22_2669 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_fill_1 FILLER_23_14 ();
 sg13g2_decap_4 FILLER_23_19 ();
 sg13g2_fill_2 FILLER_23_70 ();
 sg13g2_fill_2 FILLER_23_76 ();
 sg13g2_decap_8 FILLER_23_82 ();
 sg13g2_decap_8 FILLER_23_89 ();
 sg13g2_fill_2 FILLER_23_96 ();
 sg13g2_decap_8 FILLER_23_103 ();
 sg13g2_fill_1 FILLER_23_114 ();
 sg13g2_decap_8 FILLER_23_124 ();
 sg13g2_decap_4 FILLER_23_131 ();
 sg13g2_decap_4 FILLER_23_139 ();
 sg13g2_fill_2 FILLER_23_143 ();
 sg13g2_fill_2 FILLER_23_149 ();
 sg13g2_fill_2 FILLER_23_160 ();
 sg13g2_fill_2 FILLER_23_165 ();
 sg13g2_fill_1 FILLER_23_167 ();
 sg13g2_decap_8 FILLER_23_174 ();
 sg13g2_fill_2 FILLER_23_181 ();
 sg13g2_fill_1 FILLER_23_183 ();
 sg13g2_fill_2 FILLER_23_188 ();
 sg13g2_fill_2 FILLER_23_236 ();
 sg13g2_fill_1 FILLER_23_249 ();
 sg13g2_fill_1 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_291 ();
 sg13g2_decap_8 FILLER_23_298 ();
 sg13g2_decap_8 FILLER_23_305 ();
 sg13g2_decap_8 FILLER_23_312 ();
 sg13g2_fill_2 FILLER_23_385 ();
 sg13g2_fill_1 FILLER_23_420 ();
 sg13g2_fill_1 FILLER_23_427 ();
 sg13g2_decap_8 FILLER_23_502 ();
 sg13g2_fill_2 FILLER_23_509 ();
 sg13g2_fill_1 FILLER_23_515 ();
 sg13g2_fill_2 FILLER_23_573 ();
 sg13g2_decap_4 FILLER_23_579 ();
 sg13g2_fill_2 FILLER_23_588 ();
 sg13g2_fill_1 FILLER_23_590 ();
 sg13g2_decap_8 FILLER_23_595 ();
 sg13g2_decap_4 FILLER_23_602 ();
 sg13g2_decap_4 FILLER_23_628 ();
 sg13g2_fill_2 FILLER_23_632 ();
 sg13g2_fill_2 FILLER_23_643 ();
 sg13g2_fill_1 FILLER_23_654 ();
 sg13g2_fill_1 FILLER_23_681 ();
 sg13g2_decap_4 FILLER_23_692 ();
 sg13g2_fill_1 FILLER_23_696 ();
 sg13g2_decap_4 FILLER_23_738 ();
 sg13g2_fill_1 FILLER_23_742 ();
 sg13g2_decap_4 FILLER_23_760 ();
 sg13g2_fill_2 FILLER_23_764 ();
 sg13g2_decap_4 FILLER_23_792 ();
 sg13g2_fill_2 FILLER_23_796 ();
 sg13g2_decap_8 FILLER_23_806 ();
 sg13g2_decap_8 FILLER_23_813 ();
 sg13g2_fill_2 FILLER_23_833 ();
 sg13g2_fill_1 FILLER_23_835 ();
 sg13g2_fill_2 FILLER_23_846 ();
 sg13g2_fill_1 FILLER_23_858 ();
 sg13g2_fill_2 FILLER_23_864 ();
 sg13g2_fill_1 FILLER_23_883 ();
 sg13g2_fill_2 FILLER_23_917 ();
 sg13g2_fill_1 FILLER_23_919 ();
 sg13g2_decap_8 FILLER_23_941 ();
 sg13g2_decap_8 FILLER_23_948 ();
 sg13g2_fill_2 FILLER_23_955 ();
 sg13g2_fill_1 FILLER_23_966 ();
 sg13g2_decap_4 FILLER_23_971 ();
 sg13g2_fill_1 FILLER_23_979 ();
 sg13g2_fill_2 FILLER_23_1024 ();
 sg13g2_fill_1 FILLER_23_1052 ();
 sg13g2_fill_1 FILLER_23_1079 ();
 sg13g2_fill_2 FILLER_23_1089 ();
 sg13g2_decap_4 FILLER_23_1099 ();
 sg13g2_fill_2 FILLER_23_1103 ();
 sg13g2_fill_2 FILLER_23_1135 ();
 sg13g2_fill_1 FILLER_23_1137 ();
 sg13g2_fill_1 FILLER_23_1143 ();
 sg13g2_fill_1 FILLER_23_1148 ();
 sg13g2_decap_4 FILLER_23_1162 ();
 sg13g2_fill_1 FILLER_23_1166 ();
 sg13g2_fill_2 FILLER_23_1171 ();
 sg13g2_fill_1 FILLER_23_1173 ();
 sg13g2_decap_4 FILLER_23_1200 ();
 sg13g2_fill_2 FILLER_23_1214 ();
 sg13g2_fill_1 FILLER_23_1216 ();
 sg13g2_decap_4 FILLER_23_1221 ();
 sg13g2_decap_4 FILLER_23_1233 ();
 sg13g2_decap_8 FILLER_23_1241 ();
 sg13g2_decap_8 FILLER_23_1248 ();
 sg13g2_fill_1 FILLER_23_1255 ();
 sg13g2_fill_2 FILLER_23_1269 ();
 sg13g2_fill_1 FILLER_23_1271 ();
 sg13g2_decap_8 FILLER_23_1292 ();
 sg13g2_decap_4 FILLER_23_1299 ();
 sg13g2_fill_1 FILLER_23_1303 ();
 sg13g2_decap_8 FILLER_23_1307 ();
 sg13g2_decap_4 FILLER_23_1314 ();
 sg13g2_decap_8 FILLER_23_1323 ();
 sg13g2_decap_8 FILLER_23_1330 ();
 sg13g2_fill_1 FILLER_23_1337 ();
 sg13g2_fill_2 FILLER_23_1342 ();
 sg13g2_fill_1 FILLER_23_1359 ();
 sg13g2_fill_1 FILLER_23_1392 ();
 sg13g2_fill_2 FILLER_23_1428 ();
 sg13g2_fill_2 FILLER_23_1466 ();
 sg13g2_fill_2 FILLER_23_1525 ();
 sg13g2_fill_2 FILLER_23_1559 ();
 sg13g2_fill_2 FILLER_23_1580 ();
 sg13g2_fill_2 FILLER_23_1586 ();
 sg13g2_fill_1 FILLER_23_1588 ();
 sg13g2_fill_2 FILLER_23_1617 ();
 sg13g2_fill_2 FILLER_23_1623 ();
 sg13g2_fill_1 FILLER_23_1660 ();
 sg13g2_decap_8 FILLER_23_1695 ();
 sg13g2_decap_4 FILLER_23_1702 ();
 sg13g2_decap_4 FILLER_23_1727 ();
 sg13g2_fill_2 FILLER_23_1735 ();
 sg13g2_fill_2 FILLER_23_1741 ();
 sg13g2_fill_1 FILLER_23_1769 ();
 sg13g2_fill_2 FILLER_23_1808 ();
 sg13g2_fill_1 FILLER_23_1810 ();
 sg13g2_fill_1 FILLER_23_1837 ();
 sg13g2_fill_1 FILLER_23_1842 ();
 sg13g2_fill_1 FILLER_23_1869 ();
 sg13g2_fill_1 FILLER_23_1900 ();
 sg13g2_decap_8 FILLER_23_1931 ();
 sg13g2_decap_4 FILLER_23_1938 ();
 sg13g2_fill_1 FILLER_23_1942 ();
 sg13g2_fill_2 FILLER_23_2046 ();
 sg13g2_decap_8 FILLER_23_2084 ();
 sg13g2_decap_8 FILLER_23_2091 ();
 sg13g2_decap_8 FILLER_23_2098 ();
 sg13g2_decap_8 FILLER_23_2105 ();
 sg13g2_fill_1 FILLER_23_2112 ();
 sg13g2_fill_2 FILLER_23_2239 ();
 sg13g2_decap_8 FILLER_23_2267 ();
 sg13g2_fill_2 FILLER_23_2274 ();
 sg13g2_fill_2 FILLER_23_2306 ();
 sg13g2_decap_8 FILLER_23_2312 ();
 sg13g2_fill_1 FILLER_23_2319 ();
 sg13g2_decap_4 FILLER_23_2346 ();
 sg13g2_decap_4 FILLER_23_2355 ();
 sg13g2_fill_1 FILLER_23_2377 ();
 sg13g2_decap_8 FILLER_23_2388 ();
 sg13g2_decap_8 FILLER_23_2395 ();
 sg13g2_decap_4 FILLER_23_2402 ();
 sg13g2_decap_4 FILLER_23_2432 ();
 sg13g2_fill_2 FILLER_23_2454 ();
 sg13g2_fill_1 FILLER_23_2456 ();
 sg13g2_decap_4 FILLER_23_2565 ();
 sg13g2_decap_8 FILLER_23_2579 ();
 sg13g2_decap_4 FILLER_23_2612 ();
 sg13g2_fill_1 FILLER_23_2616 ();
 sg13g2_fill_2 FILLER_23_2637 ();
 sg13g2_fill_1 FILLER_23_2669 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_fill_2 FILLER_24_14 ();
 sg13g2_fill_2 FILLER_24_58 ();
 sg13g2_fill_1 FILLER_24_75 ();
 sg13g2_decap_4 FILLER_24_81 ();
 sg13g2_fill_1 FILLER_24_85 ();
 sg13g2_fill_1 FILLER_24_117 ();
 sg13g2_decap_4 FILLER_24_123 ();
 sg13g2_fill_2 FILLER_24_132 ();
 sg13g2_fill_1 FILLER_24_134 ();
 sg13g2_decap_4 FILLER_24_153 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_fill_2 FILLER_24_168 ();
 sg13g2_fill_1 FILLER_24_170 ();
 sg13g2_fill_1 FILLER_24_182 ();
 sg13g2_fill_1 FILLER_24_214 ();
 sg13g2_fill_1 FILLER_24_223 ();
 sg13g2_decap_8 FILLER_24_275 ();
 sg13g2_decap_8 FILLER_24_282 ();
 sg13g2_fill_1 FILLER_24_289 ();
 sg13g2_fill_2 FILLER_24_296 ();
 sg13g2_fill_1 FILLER_24_298 ();
 sg13g2_fill_2 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_335 ();
 sg13g2_decap_4 FILLER_24_352 ();
 sg13g2_fill_2 FILLER_24_356 ();
 sg13g2_fill_1 FILLER_24_417 ();
 sg13g2_decap_8 FILLER_24_468 ();
 sg13g2_fill_1 FILLER_24_475 ();
 sg13g2_fill_1 FILLER_24_512 ();
 sg13g2_decap_4 FILLER_24_518 ();
 sg13g2_fill_1 FILLER_24_522 ();
 sg13g2_decap_4 FILLER_24_527 ();
 sg13g2_fill_1 FILLER_24_531 ();
 sg13g2_fill_2 FILLER_24_538 ();
 sg13g2_fill_1 FILLER_24_540 ();
 sg13g2_fill_1 FILLER_24_545 ();
 sg13g2_fill_2 FILLER_24_551 ();
 sg13g2_fill_1 FILLER_24_553 ();
 sg13g2_fill_1 FILLER_24_600 ();
 sg13g2_fill_1 FILLER_24_654 ();
 sg13g2_fill_1 FILLER_24_665 ();
 sg13g2_fill_1 FILLER_24_676 ();
 sg13g2_fill_1 FILLER_24_703 ();
 sg13g2_fill_1 FILLER_24_730 ();
 sg13g2_fill_1 FILLER_24_735 ();
 sg13g2_fill_1 FILLER_24_762 ();
 sg13g2_fill_1 FILLER_24_815 ();
 sg13g2_decap_4 FILLER_24_837 ();
 sg13g2_fill_2 FILLER_24_845 ();
 sg13g2_fill_1 FILLER_24_847 ();
 sg13g2_fill_1 FILLER_24_853 ();
 sg13g2_fill_1 FILLER_24_869 ();
 sg13g2_decap_8 FILLER_24_934 ();
 sg13g2_decap_4 FILLER_24_941 ();
 sg13g2_fill_1 FILLER_24_945 ();
 sg13g2_decap_4 FILLER_24_954 ();
 sg13g2_fill_1 FILLER_24_958 ();
 sg13g2_fill_1 FILLER_24_989 ();
 sg13g2_fill_2 FILLER_24_994 ();
 sg13g2_fill_2 FILLER_24_1000 ();
 sg13g2_fill_2 FILLER_24_1023 ();
 sg13g2_fill_2 FILLER_24_1066 ();
 sg13g2_fill_1 FILLER_24_1068 ();
 sg13g2_decap_4 FILLER_24_1086 ();
 sg13g2_fill_2 FILLER_24_1090 ();
 sg13g2_fill_2 FILLER_24_1101 ();
 sg13g2_fill_2 FILLER_24_1108 ();
 sg13g2_fill_2 FILLER_24_1140 ();
 sg13g2_fill_2 FILLER_24_1146 ();
 sg13g2_fill_2 FILLER_24_1196 ();
 sg13g2_fill_1 FILLER_24_1198 ();
 sg13g2_fill_2 FILLER_24_1236 ();
 sg13g2_fill_1 FILLER_24_1238 ();
 sg13g2_fill_2 FILLER_24_1308 ();
 sg13g2_fill_1 FILLER_24_1340 ();
 sg13g2_fill_1 FILLER_24_1346 ();
 sg13g2_fill_1 FILLER_24_1351 ();
 sg13g2_fill_1 FILLER_24_1356 ();
 sg13g2_fill_1 FILLER_24_1365 ();
 sg13g2_fill_2 FILLER_24_1396 ();
 sg13g2_fill_1 FILLER_24_1409 ();
 sg13g2_fill_2 FILLER_24_1474 ();
 sg13g2_fill_2 FILLER_24_1483 ();
 sg13g2_decap_8 FILLER_24_1519 ();
 sg13g2_decap_8 FILLER_24_1526 ();
 sg13g2_fill_2 FILLER_24_1533 ();
 sg13g2_fill_2 FILLER_24_1565 ();
 sg13g2_fill_2 FILLER_24_1587 ();
 sg13g2_fill_2 FILLER_24_1593 ();
 sg13g2_decap_8 FILLER_24_1605 ();
 sg13g2_fill_2 FILLER_24_1612 ();
 sg13g2_fill_2 FILLER_24_1619 ();
 sg13g2_fill_2 FILLER_24_1626 ();
 sg13g2_decap_8 FILLER_24_1645 ();
 sg13g2_decap_4 FILLER_24_1652 ();
 sg13g2_decap_8 FILLER_24_1660 ();
 sg13g2_decap_8 FILLER_24_1667 ();
 sg13g2_fill_1 FILLER_24_1674 ();
 sg13g2_fill_1 FILLER_24_1679 ();
 sg13g2_decap_4 FILLER_24_1690 ();
 sg13g2_decap_8 FILLER_24_1735 ();
 sg13g2_decap_4 FILLER_24_1742 ();
 sg13g2_fill_2 FILLER_24_1746 ();
 sg13g2_fill_2 FILLER_24_1758 ();
 sg13g2_fill_2 FILLER_24_1789 ();
 sg13g2_fill_1 FILLER_24_1791 ();
 sg13g2_decap_4 FILLER_24_1796 ();
 sg13g2_decap_8 FILLER_24_1804 ();
 sg13g2_fill_2 FILLER_24_1811 ();
 sg13g2_fill_1 FILLER_24_1813 ();
 sg13g2_decap_4 FILLER_24_1833 ();
 sg13g2_fill_1 FILLER_24_1837 ();
 sg13g2_fill_2 FILLER_24_1866 ();
 sg13g2_fill_2 FILLER_24_1906 ();
 sg13g2_fill_1 FILLER_24_1908 ();
 sg13g2_decap_8 FILLER_24_1935 ();
 sg13g2_fill_1 FILLER_24_1942 ();
 sg13g2_fill_1 FILLER_24_1947 ();
 sg13g2_decap_4 FILLER_24_1982 ();
 sg13g2_fill_2 FILLER_24_1996 ();
 sg13g2_fill_1 FILLER_24_2009 ();
 sg13g2_decap_8 FILLER_24_2075 ();
 sg13g2_decap_8 FILLER_24_2108 ();
 sg13g2_decap_4 FILLER_24_2115 ();
 sg13g2_fill_1 FILLER_24_2119 ();
 sg13g2_fill_2 FILLER_24_2125 ();
 sg13g2_fill_2 FILLER_24_2131 ();
 sg13g2_decap_8 FILLER_24_2154 ();
 sg13g2_decap_8 FILLER_24_2161 ();
 sg13g2_decap_8 FILLER_24_2168 ();
 sg13g2_decap_8 FILLER_24_2175 ();
 sg13g2_fill_2 FILLER_24_2182 ();
 sg13g2_fill_1 FILLER_24_2188 ();
 sg13g2_fill_2 FILLER_24_2193 ();
 sg13g2_fill_1 FILLER_24_2195 ();
 sg13g2_decap_4 FILLER_24_2204 ();
 sg13g2_decap_8 FILLER_24_2233 ();
 sg13g2_decap_8 FILLER_24_2240 ();
 sg13g2_decap_4 FILLER_24_2247 ();
 sg13g2_decap_8 FILLER_24_2255 ();
 sg13g2_fill_2 FILLER_24_2262 ();
 sg13g2_decap_4 FILLER_24_2296 ();
 sg13g2_fill_1 FILLER_24_2300 ();
 sg13g2_decap_4 FILLER_24_2310 ();
 sg13g2_fill_1 FILLER_24_2314 ();
 sg13g2_decap_8 FILLER_24_2319 ();
 sg13g2_decap_8 FILLER_24_2330 ();
 sg13g2_decap_4 FILLER_24_2337 ();
 sg13g2_decap_8 FILLER_24_2391 ();
 sg13g2_decap_8 FILLER_24_2398 ();
 sg13g2_decap_8 FILLER_24_2405 ();
 sg13g2_decap_8 FILLER_24_2429 ();
 sg13g2_decap_4 FILLER_24_2436 ();
 sg13g2_fill_1 FILLER_24_2440 ();
 sg13g2_fill_2 FILLER_24_2473 ();
 sg13g2_fill_2 FILLER_24_2481 ();
 sg13g2_fill_1 FILLER_24_2489 ();
 sg13g2_fill_2 FILLER_24_2496 ();
 sg13g2_fill_2 FILLER_24_2510 ();
 sg13g2_decap_4 FILLER_24_2566 ();
 sg13g2_fill_1 FILLER_24_2570 ();
 sg13g2_fill_1 FILLER_24_2623 ();
 sg13g2_decap_4 FILLER_24_2634 ();
 sg13g2_fill_2 FILLER_24_2638 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_28 ();
 sg13g2_fill_1 FILLER_25_34 ();
 sg13g2_fill_1 FILLER_25_62 ();
 sg13g2_fill_2 FILLER_25_103 ();
 sg13g2_fill_2 FILLER_25_109 ();
 sg13g2_fill_2 FILLER_25_119 ();
 sg13g2_decap_4 FILLER_25_126 ();
 sg13g2_fill_2 FILLER_25_186 ();
 sg13g2_fill_1 FILLER_25_188 ();
 sg13g2_fill_1 FILLER_25_200 ();
 sg13g2_fill_1 FILLER_25_206 ();
 sg13g2_fill_2 FILLER_25_211 ();
 sg13g2_fill_2 FILLER_25_218 ();
 sg13g2_fill_2 FILLER_25_225 ();
 sg13g2_fill_1 FILLER_25_227 ();
 sg13g2_fill_2 FILLER_25_272 ();
 sg13g2_fill_1 FILLER_25_310 ();
 sg13g2_decap_8 FILLER_25_329 ();
 sg13g2_decap_8 FILLER_25_344 ();
 sg13g2_decap_4 FILLER_25_351 ();
 sg13g2_decap_8 FILLER_25_359 ();
 sg13g2_fill_1 FILLER_25_366 ();
 sg13g2_fill_1 FILLER_25_381 ();
 sg13g2_fill_1 FILLER_25_387 ();
 sg13g2_fill_1 FILLER_25_418 ();
 sg13g2_fill_1 FILLER_25_447 ();
 sg13g2_decap_4 FILLER_25_474 ();
 sg13g2_fill_2 FILLER_25_478 ();
 sg13g2_decap_4 FILLER_25_497 ();
 sg13g2_fill_1 FILLER_25_501 ();
 sg13g2_decap_4 FILLER_25_518 ();
 sg13g2_fill_1 FILLER_25_522 ();
 sg13g2_decap_8 FILLER_25_527 ();
 sg13g2_decap_4 FILLER_25_534 ();
 sg13g2_decap_4 FILLER_25_544 ();
 sg13g2_fill_1 FILLER_25_548 ();
 sg13g2_fill_2 FILLER_25_553 ();
 sg13g2_fill_1 FILLER_25_580 ();
 sg13g2_fill_2 FILLER_25_585 ();
 sg13g2_fill_1 FILLER_25_587 ();
 sg13g2_fill_1 FILLER_25_601 ();
 sg13g2_fill_2 FILLER_25_612 ();
 sg13g2_fill_2 FILLER_25_628 ();
 sg13g2_fill_2 FILLER_25_634 ();
 sg13g2_fill_2 FILLER_25_641 ();
 sg13g2_fill_1 FILLER_25_647 ();
 sg13g2_fill_1 FILLER_25_662 ();
 sg13g2_fill_1 FILLER_25_680 ();
 sg13g2_fill_2 FILLER_25_689 ();
 sg13g2_fill_1 FILLER_25_691 ();
 sg13g2_fill_1 FILLER_25_700 ();
 sg13g2_fill_2 FILLER_25_715 ();
 sg13g2_fill_2 FILLER_25_736 ();
 sg13g2_decap_8 FILLER_25_818 ();
 sg13g2_decap_8 FILLER_25_825 ();
 sg13g2_fill_2 FILLER_25_832 ();
 sg13g2_fill_1 FILLER_25_834 ();
 sg13g2_fill_2 FILLER_25_861 ();
 sg13g2_fill_2 FILLER_25_867 ();
 sg13g2_fill_2 FILLER_25_895 ();
 sg13g2_decap_8 FILLER_25_995 ();
 sg13g2_decap_8 FILLER_25_1002 ();
 sg13g2_fill_2 FILLER_25_1091 ();
 sg13g2_decap_8 FILLER_25_1123 ();
 sg13g2_fill_1 FILLER_25_1156 ();
 sg13g2_fill_2 FILLER_25_1242 ();
 sg13g2_fill_2 FILLER_25_1267 ();
 sg13g2_fill_1 FILLER_25_1286 ();
 sg13g2_fill_2 FILLER_25_1309 ();
 sg13g2_decap_4 FILLER_25_1315 ();
 sg13g2_fill_2 FILLER_25_1323 ();
 sg13g2_fill_2 FILLER_25_1342 ();
 sg13g2_fill_1 FILLER_25_1344 ();
 sg13g2_fill_1 FILLER_25_1353 ();
 sg13g2_fill_2 FILLER_25_1408 ();
 sg13g2_fill_1 FILLER_25_1415 ();
 sg13g2_fill_1 FILLER_25_1481 ();
 sg13g2_decap_8 FILLER_25_1495 ();
 sg13g2_decap_8 FILLER_25_1502 ();
 sg13g2_fill_2 FILLER_25_1518 ();
 sg13g2_fill_1 FILLER_25_1520 ();
 sg13g2_fill_2 FILLER_25_1526 ();
 sg13g2_fill_1 FILLER_25_1528 ();
 sg13g2_fill_2 FILLER_25_1556 ();
 sg13g2_fill_2 FILLER_25_1575 ();
 sg13g2_fill_1 FILLER_25_1628 ();
 sg13g2_decap_4 FILLER_25_1652 ();
 sg13g2_fill_1 FILLER_25_1656 ();
 sg13g2_fill_2 FILLER_25_1670 ();
 sg13g2_fill_1 FILLER_25_1672 ();
 sg13g2_decap_4 FILLER_25_1733 ();
 sg13g2_fill_2 FILLER_25_1737 ();
 sg13g2_fill_2 FILLER_25_1794 ();
 sg13g2_fill_1 FILLER_25_1796 ();
 sg13g2_decap_8 FILLER_25_1801 ();
 sg13g2_decap_8 FILLER_25_1832 ();
 sg13g2_fill_1 FILLER_25_1843 ();
 sg13g2_fill_1 FILLER_25_1854 ();
 sg13g2_fill_1 FILLER_25_1904 ();
 sg13g2_fill_2 FILLER_25_1930 ();
 sg13g2_fill_1 FILLER_25_1945 ();
 sg13g2_fill_2 FILLER_25_1956 ();
 sg13g2_decap_4 FILLER_25_1968 ();
 sg13g2_fill_2 FILLER_25_1993 ();
 sg13g2_fill_2 FILLER_25_2007 ();
 sg13g2_fill_1 FILLER_25_2020 ();
 sg13g2_decap_4 FILLER_25_2051 ();
 sg13g2_decap_4 FILLER_25_2094 ();
 sg13g2_fill_1 FILLER_25_2098 ();
 sg13g2_fill_1 FILLER_25_2135 ();
 sg13g2_fill_2 FILLER_25_2181 ();
 sg13g2_decap_8 FILLER_25_2191 ();
 sg13g2_decap_8 FILLER_25_2198 ();
 sg13g2_decap_8 FILLER_25_2205 ();
 sg13g2_decap_8 FILLER_25_2212 ();
 sg13g2_fill_1 FILLER_25_2219 ();
 sg13g2_fill_2 FILLER_25_2230 ();
 sg13g2_fill_1 FILLER_25_2232 ();
 sg13g2_decap_8 FILLER_25_2290 ();
 sg13g2_fill_1 FILLER_25_2297 ();
 sg13g2_decap_4 FILLER_25_2303 ();
 sg13g2_fill_1 FILLER_25_2307 ();
 sg13g2_fill_2 FILLER_25_2344 ();
 sg13g2_fill_1 FILLER_25_2346 ();
 sg13g2_decap_4 FILLER_25_2353 ();
 sg13g2_fill_1 FILLER_25_2357 ();
 sg13g2_fill_2 FILLER_25_2368 ();
 sg13g2_fill_1 FILLER_25_2400 ();
 sg13g2_fill_2 FILLER_25_2411 ();
 sg13g2_fill_1 FILLER_25_2413 ();
 sg13g2_decap_4 FILLER_25_2429 ();
 sg13g2_fill_2 FILLER_25_2463 ();
 sg13g2_fill_1 FILLER_25_2481 ();
 sg13g2_fill_2 FILLER_25_2490 ();
 sg13g2_fill_2 FILLER_25_2496 ();
 sg13g2_fill_2 FILLER_25_2506 ();
 sg13g2_fill_1 FILLER_25_2508 ();
 sg13g2_fill_1 FILLER_25_2514 ();
 sg13g2_decap_4 FILLER_25_2640 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_27 ();
 sg13g2_fill_1 FILLER_26_32 ();
 sg13g2_fill_1 FILLER_26_38 ();
 sg13g2_decap_8 FILLER_26_45 ();
 sg13g2_decap_4 FILLER_26_52 ();
 sg13g2_fill_2 FILLER_26_64 ();
 sg13g2_decap_4 FILLER_26_76 ();
 sg13g2_fill_2 FILLER_26_80 ();
 sg13g2_fill_2 FILLER_26_87 ();
 sg13g2_fill_1 FILLER_26_119 ();
 sg13g2_fill_1 FILLER_26_131 ();
 sg13g2_fill_1 FILLER_26_136 ();
 sg13g2_fill_2 FILLER_26_141 ();
 sg13g2_decap_8 FILLER_26_170 ();
 sg13g2_fill_2 FILLER_26_187 ();
 sg13g2_fill_2 FILLER_26_194 ();
 sg13g2_fill_2 FILLER_26_201 ();
 sg13g2_fill_1 FILLER_26_203 ();
 sg13g2_fill_1 FILLER_26_212 ();
 sg13g2_fill_2 FILLER_26_217 ();
 sg13g2_fill_1 FILLER_26_219 ();
 sg13g2_decap_8 FILLER_26_228 ();
 sg13g2_decap_8 FILLER_26_235 ();
 sg13g2_fill_1 FILLER_26_242 ();
 sg13g2_fill_1 FILLER_26_257 ();
 sg13g2_decap_8 FILLER_26_288 ();
 sg13g2_fill_1 FILLER_26_295 ();
 sg13g2_decap_8 FILLER_26_374 ();
 sg13g2_fill_1 FILLER_26_389 ();
 sg13g2_fill_2 FILLER_26_427 ();
 sg13g2_fill_1 FILLER_26_435 ();
 sg13g2_decap_4 FILLER_26_477 ();
 sg13g2_fill_2 FILLER_26_485 ();
 sg13g2_fill_2 FILLER_26_492 ();
 sg13g2_fill_1 FILLER_26_494 ();
 sg13g2_fill_2 FILLER_26_499 ();
 sg13g2_fill_1 FILLER_26_562 ();
 sg13g2_fill_1 FILLER_26_568 ();
 sg13g2_fill_1 FILLER_26_595 ();
 sg13g2_fill_1 FILLER_26_673 ();
 sg13g2_fill_1 FILLER_26_680 ();
 sg13g2_fill_1 FILLER_26_709 ();
 sg13g2_fill_2 FILLER_26_721 ();
 sg13g2_fill_1 FILLER_26_739 ();
 sg13g2_fill_1 FILLER_26_749 ();
 sg13g2_decap_8 FILLER_26_763 ();
 sg13g2_decap_4 FILLER_26_770 ();
 sg13g2_fill_1 FILLER_26_774 ();
 sg13g2_decap_4 FILLER_26_779 ();
 sg13g2_fill_1 FILLER_26_783 ();
 sg13g2_fill_2 FILLER_26_834 ();
 sg13g2_fill_1 FILLER_26_895 ();
 sg13g2_fill_1 FILLER_26_923 ();
 sg13g2_fill_2 FILLER_26_954 ();
 sg13g2_fill_1 FILLER_26_956 ();
 sg13g2_fill_2 FILLER_26_962 ();
 sg13g2_fill_2 FILLER_26_990 ();
 sg13g2_decap_4 FILLER_26_1013 ();
 sg13g2_fill_2 FILLER_26_1017 ();
 sg13g2_fill_2 FILLER_26_1023 ();
 sg13g2_fill_1 FILLER_26_1025 ();
 sg13g2_fill_2 FILLER_26_1030 ();
 sg13g2_fill_1 FILLER_26_1032 ();
 sg13g2_fill_2 FILLER_26_1037 ();
 sg13g2_fill_2 FILLER_26_1044 ();
 sg13g2_decap_8 FILLER_26_1054 ();
 sg13g2_fill_1 FILLER_26_1061 ();
 sg13g2_decap_4 FILLER_26_1070 ();
 sg13g2_fill_2 FILLER_26_1074 ();
 sg13g2_fill_2 FILLER_26_1101 ();
 sg13g2_fill_2 FILLER_26_1107 ();
 sg13g2_fill_1 FILLER_26_1109 ();
 sg13g2_fill_1 FILLER_26_1178 ();
 sg13g2_fill_2 FILLER_26_1184 ();
 sg13g2_fill_1 FILLER_26_1186 ();
 sg13g2_fill_2 FILLER_26_1191 ();
 sg13g2_fill_2 FILLER_26_1282 ();
 sg13g2_fill_1 FILLER_26_1284 ();
 sg13g2_decap_8 FILLER_26_1289 ();
 sg13g2_fill_1 FILLER_26_1296 ();
 sg13g2_decap_8 FILLER_26_1313 ();
 sg13g2_decap_8 FILLER_26_1320 ();
 sg13g2_fill_2 FILLER_26_1327 ();
 sg13g2_decap_8 FILLER_26_1333 ();
 sg13g2_decap_8 FILLER_26_1340 ();
 sg13g2_decap_4 FILLER_26_1347 ();
 sg13g2_fill_1 FILLER_26_1351 ();
 sg13g2_fill_2 FILLER_26_1360 ();
 sg13g2_fill_1 FILLER_26_1362 ();
 sg13g2_fill_2 FILLER_26_1401 ();
 sg13g2_fill_2 FILLER_26_1454 ();
 sg13g2_fill_1 FILLER_26_1474 ();
 sg13g2_decap_8 FILLER_26_1493 ();
 sg13g2_decap_4 FILLER_26_1500 ();
 sg13g2_fill_2 FILLER_26_1504 ();
 sg13g2_fill_2 FILLER_26_1526 ();
 sg13g2_fill_1 FILLER_26_1554 ();
 sg13g2_fill_2 FILLER_26_1565 ();
 sg13g2_fill_2 FILLER_26_1577 ();
 sg13g2_fill_2 FILLER_26_1583 ();
 sg13g2_fill_2 FILLER_26_1589 ();
 sg13g2_decap_4 FILLER_26_1612 ();
 sg13g2_fill_2 FILLER_26_1620 ();
 sg13g2_fill_1 FILLER_26_1682 ();
 sg13g2_fill_1 FILLER_26_1729 ();
 sg13g2_fill_1 FILLER_26_1796 ();
 sg13g2_decap_8 FILLER_26_1805 ();
 sg13g2_fill_2 FILLER_26_1812 ();
 sg13g2_fill_2 FILLER_26_1839 ();
 sg13g2_fill_1 FILLER_26_1841 ();
 sg13g2_fill_1 FILLER_26_1880 ();
 sg13g2_decap_4 FILLER_26_1936 ();
 sg13g2_fill_2 FILLER_26_1940 ();
 sg13g2_fill_2 FILLER_26_1968 ();
 sg13g2_fill_1 FILLER_26_1970 ();
 sg13g2_decap_8 FILLER_26_1975 ();
 sg13g2_decap_4 FILLER_26_1982 ();
 sg13g2_fill_2 FILLER_26_2048 ();
 sg13g2_fill_1 FILLER_26_2056 ();
 sg13g2_decap_4 FILLER_26_2135 ();
 sg13g2_fill_2 FILLER_26_2139 ();
 sg13g2_decap_8 FILLER_26_2197 ();
 sg13g2_fill_1 FILLER_26_2204 ();
 sg13g2_decap_4 FILLER_26_2225 ();
 sg13g2_decap_8 FILLER_26_2255 ();
 sg13g2_decap_4 FILLER_26_2262 ();
 sg13g2_fill_1 FILLER_26_2266 ();
 sg13g2_decap_4 FILLER_26_2293 ();
 sg13g2_fill_1 FILLER_26_2327 ();
 sg13g2_fill_2 FILLER_26_2354 ();
 sg13g2_fill_2 FILLER_26_2362 ();
 sg13g2_fill_2 FILLER_26_2368 ();
 sg13g2_fill_1 FILLER_26_2432 ();
 sg13g2_decap_4 FILLER_26_2459 ();
 sg13g2_fill_2 FILLER_26_2495 ();
 sg13g2_fill_1 FILLER_26_2497 ();
 sg13g2_fill_2 FILLER_26_2535 ();
 sg13g2_fill_1 FILLER_26_2543 ();
 sg13g2_fill_2 FILLER_26_2555 ();
 sg13g2_fill_1 FILLER_26_2557 ();
 sg13g2_decap_4 FILLER_26_2568 ();
 sg13g2_fill_1 FILLER_26_2572 ();
 sg13g2_fill_2 FILLER_26_2577 ();
 sg13g2_fill_1 FILLER_26_2579 ();
 sg13g2_decap_4 FILLER_26_2584 ();
 sg13g2_fill_1 FILLER_26_2588 ();
 sg13g2_decap_4 FILLER_26_2599 ();
 sg13g2_fill_1 FILLER_26_2603 ();
 sg13g2_fill_2 FILLER_26_2608 ();
 sg13g2_fill_1 FILLER_26_2610 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_15 ();
 sg13g2_decap_8 FILLER_27_34 ();
 sg13g2_decap_8 FILLER_27_41 ();
 sg13g2_decap_8 FILLER_27_48 ();
 sg13g2_decap_8 FILLER_27_55 ();
 sg13g2_decap_8 FILLER_27_62 ();
 sg13g2_fill_2 FILLER_27_69 ();
 sg13g2_decap_8 FILLER_27_75 ();
 sg13g2_decap_4 FILLER_27_82 ();
 sg13g2_fill_1 FILLER_27_86 ();
 sg13g2_fill_2 FILLER_27_91 ();
 sg13g2_fill_2 FILLER_27_97 ();
 sg13g2_fill_1 FILLER_27_99 ();
 sg13g2_fill_1 FILLER_27_126 ();
 sg13g2_fill_2 FILLER_27_145 ();
 sg13g2_fill_1 FILLER_27_164 ();
 sg13g2_fill_2 FILLER_27_170 ();
 sg13g2_fill_1 FILLER_27_172 ();
 sg13g2_fill_1 FILLER_27_187 ();
 sg13g2_fill_1 FILLER_27_211 ();
 sg13g2_decap_4 FILLER_27_219 ();
 sg13g2_fill_2 FILLER_27_223 ();
 sg13g2_fill_2 FILLER_27_230 ();
 sg13g2_fill_1 FILLER_27_232 ();
 sg13g2_decap_8 FILLER_27_272 ();
 sg13g2_decap_8 FILLER_27_279 ();
 sg13g2_decap_8 FILLER_27_286 ();
 sg13g2_fill_1 FILLER_27_293 ();
 sg13g2_decap_4 FILLER_27_302 ();
 sg13g2_fill_1 FILLER_27_306 ();
 sg13g2_fill_2 FILLER_27_321 ();
 sg13g2_fill_1 FILLER_27_323 ();
 sg13g2_decap_8 FILLER_27_329 ();
 sg13g2_fill_1 FILLER_27_336 ();
 sg13g2_fill_1 FILLER_27_341 ();
 sg13g2_fill_1 FILLER_27_346 ();
 sg13g2_decap_8 FILLER_27_360 ();
 sg13g2_fill_2 FILLER_27_367 ();
 sg13g2_fill_1 FILLER_27_369 ();
 sg13g2_fill_1 FILLER_27_374 ();
 sg13g2_fill_1 FILLER_27_428 ();
 sg13g2_fill_1 FILLER_27_447 ();
 sg13g2_fill_1 FILLER_27_458 ();
 sg13g2_fill_2 FILLER_27_480 ();
 sg13g2_fill_1 FILLER_27_482 ();
 sg13g2_fill_1 FILLER_27_554 ();
 sg13g2_fill_1 FILLER_27_560 ();
 sg13g2_fill_2 FILLER_27_581 ();
 sg13g2_fill_2 FILLER_27_644 ();
 sg13g2_fill_1 FILLER_27_662 ();
 sg13g2_fill_2 FILLER_27_697 ();
 sg13g2_fill_2 FILLER_27_733 ();
 sg13g2_fill_1 FILLER_27_750 ();
 sg13g2_fill_1 FILLER_27_759 ();
 sg13g2_decap_8 FILLER_27_770 ();
 sg13g2_decap_8 FILLER_27_777 ();
 sg13g2_decap_8 FILLER_27_784 ();
 sg13g2_decap_4 FILLER_27_791 ();
 sg13g2_decap_8 FILLER_27_811 ();
 sg13g2_fill_2 FILLER_27_818 ();
 sg13g2_decap_8 FILLER_27_829 ();
 sg13g2_fill_1 FILLER_27_836 ();
 sg13g2_fill_1 FILLER_27_888 ();
 sg13g2_fill_2 FILLER_27_902 ();
 sg13g2_fill_1 FILLER_27_925 ();
 sg13g2_decap_8 FILLER_27_1022 ();
 sg13g2_decap_8 FILLER_27_1029 ();
 sg13g2_fill_1 FILLER_27_1036 ();
 sg13g2_decap_8 FILLER_27_1045 ();
 sg13g2_decap_8 FILLER_27_1056 ();
 sg13g2_decap_8 FILLER_27_1098 ();
 sg13g2_decap_8 FILLER_27_1105 ();
 sg13g2_fill_2 FILLER_27_1112 ();
 sg13g2_decap_8 FILLER_27_1118 ();
 sg13g2_decap_8 FILLER_27_1125 ();
 sg13g2_fill_1 FILLER_27_1177 ();
 sg13g2_fill_2 FILLER_27_1207 ();
 sg13g2_fill_2 FILLER_27_1220 ();
 sg13g2_fill_1 FILLER_27_1248 ();
 sg13g2_decap_8 FILLER_27_1296 ();
 sg13g2_decap_8 FILLER_27_1303 ();
 sg13g2_decap_8 FILLER_27_1310 ();
 sg13g2_decap_8 FILLER_27_1321 ();
 sg13g2_fill_2 FILLER_27_1328 ();
 sg13g2_decap_8 FILLER_27_1356 ();
 sg13g2_fill_1 FILLER_27_1363 ();
 sg13g2_fill_1 FILLER_27_1368 ();
 sg13g2_fill_2 FILLER_27_1389 ();
 sg13g2_fill_2 FILLER_27_1426 ();
 sg13g2_fill_1 FILLER_27_1483 ();
 sg13g2_fill_1 FILLER_27_1489 ();
 sg13g2_fill_1 FILLER_27_1494 ();
 sg13g2_fill_2 FILLER_27_1517 ();
 sg13g2_fill_2 FILLER_27_1523 ();
 sg13g2_fill_1 FILLER_27_1560 ();
 sg13g2_decap_4 FILLER_27_1669 ();
 sg13g2_fill_1 FILLER_27_1673 ();
 sg13g2_fill_1 FILLER_27_1680 ();
 sg13g2_fill_1 FILLER_27_1691 ();
 sg13g2_fill_2 FILLER_27_1696 ();
 sg13g2_fill_1 FILLER_27_1698 ();
 sg13g2_fill_1 FILLER_27_1703 ();
 sg13g2_decap_8 FILLER_27_1712 ();
 sg13g2_decap_8 FILLER_27_1719 ();
 sg13g2_fill_2 FILLER_27_1726 ();
 sg13g2_fill_2 FILLER_27_1749 ();
 sg13g2_fill_1 FILLER_27_1777 ();
 sg13g2_fill_2 FILLER_27_1782 ();
 sg13g2_fill_1 FILLER_27_1784 ();
 sg13g2_decap_4 FILLER_27_1811 ();
 sg13g2_fill_2 FILLER_27_1815 ();
 sg13g2_fill_2 FILLER_27_1820 ();
 sg13g2_fill_1 FILLER_27_1848 ();
 sg13g2_fill_2 FILLER_27_1854 ();
 sg13g2_fill_1 FILLER_27_1877 ();
 sg13g2_fill_2 FILLER_27_1897 ();
 sg13g2_decap_8 FILLER_27_1979 ();
 sg13g2_decap_8 FILLER_27_1986 ();
 sg13g2_decap_8 FILLER_27_1993 ();
 sg13g2_decap_8 FILLER_27_2000 ();
 sg13g2_decap_8 FILLER_27_2007 ();
 sg13g2_fill_2 FILLER_27_2028 ();
 sg13g2_fill_2 FILLER_27_2061 ();
 sg13g2_decap_8 FILLER_27_2085 ();
 sg13g2_fill_2 FILLER_27_2092 ();
 sg13g2_fill_2 FILLER_27_2097 ();
 sg13g2_decap_4 FILLER_27_2120 ();
 sg13g2_decap_4 FILLER_27_2134 ();
 sg13g2_decap_4 FILLER_27_2174 ();
 sg13g2_fill_2 FILLER_27_2188 ();
 sg13g2_fill_1 FILLER_27_2190 ();
 sg13g2_decap_8 FILLER_27_2248 ();
 sg13g2_fill_2 FILLER_27_2255 ();
 sg13g2_fill_2 FILLER_27_2269 ();
 sg13g2_fill_1 FILLER_27_2271 ();
 sg13g2_fill_2 FILLER_27_2276 ();
 sg13g2_fill_1 FILLER_27_2278 ();
 sg13g2_fill_1 FILLER_27_2289 ();
 sg13g2_decap_8 FILLER_27_2316 ();
 sg13g2_fill_1 FILLER_27_2323 ();
 sg13g2_decap_4 FILLER_27_2386 ();
 sg13g2_fill_2 FILLER_27_2418 ();
 sg13g2_decap_8 FILLER_27_2424 ();
 sg13g2_fill_2 FILLER_27_2431 ();
 sg13g2_decap_4 FILLER_27_2465 ();
 sg13g2_fill_2 FILLER_27_2469 ();
 sg13g2_fill_2 FILLER_27_2481 ();
 sg13g2_fill_1 FILLER_27_2483 ();
 sg13g2_fill_2 FILLER_27_2488 ();
 sg13g2_fill_2 FILLER_27_2532 ();
 sg13g2_decap_8 FILLER_27_2570 ();
 sg13g2_decap_8 FILLER_27_2577 ();
 sg13g2_decap_8 FILLER_27_2584 ();
 sg13g2_decap_8 FILLER_27_2591 ();
 sg13g2_decap_8 FILLER_27_2598 ();
 sg13g2_decap_8 FILLER_27_2605 ();
 sg13g2_fill_2 FILLER_27_2612 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_7 ();
 sg13g2_fill_2 FILLER_28_11 ();
 sg13g2_fill_2 FILLER_28_31 ();
 sg13g2_fill_1 FILLER_28_33 ();
 sg13g2_decap_4 FILLER_28_38 ();
 sg13g2_fill_2 FILLER_28_42 ();
 sg13g2_fill_2 FILLER_28_48 ();
 sg13g2_fill_1 FILLER_28_50 ();
 sg13g2_decap_8 FILLER_28_55 ();
 sg13g2_decap_8 FILLER_28_62 ();
 sg13g2_fill_1 FILLER_28_69 ();
 sg13g2_fill_2 FILLER_28_74 ();
 sg13g2_fill_2 FILLER_28_80 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_fill_1 FILLER_28_119 ();
 sg13g2_fill_1 FILLER_28_161 ();
 sg13g2_fill_2 FILLER_28_201 ();
 sg13g2_fill_1 FILLER_28_229 ();
 sg13g2_fill_1 FILLER_28_256 ();
 sg13g2_decap_8 FILLER_28_261 ();
 sg13g2_decap_8 FILLER_28_268 ();
 sg13g2_fill_1 FILLER_28_275 ();
 sg13g2_fill_2 FILLER_28_298 ();
 sg13g2_decap_4 FILLER_28_328 ();
 sg13g2_decap_8 FILLER_28_358 ();
 sg13g2_fill_1 FILLER_28_365 ();
 sg13g2_decap_8 FILLER_28_371 ();
 sg13g2_fill_2 FILLER_28_378 ();
 sg13g2_fill_1 FILLER_28_380 ();
 sg13g2_decap_8 FILLER_28_389 ();
 sg13g2_fill_1 FILLER_28_396 ();
 sg13g2_fill_1 FILLER_28_417 ();
 sg13g2_fill_2 FILLER_28_433 ();
 sg13g2_decap_4 FILLER_28_481 ();
 sg13g2_fill_2 FILLER_28_485 ();
 sg13g2_fill_1 FILLER_28_513 ();
 sg13g2_fill_2 FILLER_28_518 ();
 sg13g2_fill_2 FILLER_28_525 ();
 sg13g2_fill_1 FILLER_28_531 ();
 sg13g2_fill_1 FILLER_28_548 ();
 sg13g2_decap_4 FILLER_28_558 ();
 sg13g2_fill_2 FILLER_28_562 ();
 sg13g2_fill_2 FILLER_28_585 ();
 sg13g2_fill_1 FILLER_28_614 ();
 sg13g2_fill_1 FILLER_28_630 ();
 sg13g2_fill_2 FILLER_28_641 ();
 sg13g2_fill_1 FILLER_28_648 ();
 sg13g2_fill_2 FILLER_28_659 ();
 sg13g2_fill_2 FILLER_28_701 ();
 sg13g2_fill_2 FILLER_28_708 ();
 sg13g2_fill_1 FILLER_28_720 ();
 sg13g2_fill_2 FILLER_28_738 ();
 sg13g2_fill_2 FILLER_28_744 ();
 sg13g2_decap_8 FILLER_28_780 ();
 sg13g2_decap_8 FILLER_28_787 ();
 sg13g2_decap_8 FILLER_28_794 ();
 sg13g2_fill_1 FILLER_28_801 ();
 sg13g2_decap_4 FILLER_28_853 ();
 sg13g2_fill_1 FILLER_28_857 ();
 sg13g2_decap_8 FILLER_28_871 ();
 sg13g2_fill_2 FILLER_28_878 ();
 sg13g2_fill_1 FILLER_28_884 ();
 sg13g2_fill_2 FILLER_28_917 ();
 sg13g2_fill_2 FILLER_28_933 ();
 sg13g2_fill_2 FILLER_28_939 ();
 sg13g2_fill_1 FILLER_28_941 ();
 sg13g2_fill_2 FILLER_28_967 ();
 sg13g2_fill_1 FILLER_28_969 ();
 sg13g2_fill_1 FILLER_28_974 ();
 sg13g2_decap_4 FILLER_28_1023 ();
 sg13g2_decap_4 FILLER_28_1031 ();
 sg13g2_decap_4 FILLER_28_1100 ();
 sg13g2_fill_2 FILLER_28_1104 ();
 sg13g2_decap_8 FILLER_28_1110 ();
 sg13g2_decap_8 FILLER_28_1117 ();
 sg13g2_fill_1 FILLER_28_1146 ();
 sg13g2_decap_8 FILLER_28_1152 ();
 sg13g2_fill_1 FILLER_28_1159 ();
 sg13g2_fill_2 FILLER_28_1191 ();
 sg13g2_fill_1 FILLER_28_1193 ();
 sg13g2_fill_2 FILLER_28_1198 ();
 sg13g2_fill_2 FILLER_28_1219 ();
 sg13g2_fill_1 FILLER_28_1233 ();
 sg13g2_fill_1 FILLER_28_1255 ();
 sg13g2_decap_8 FILLER_28_1292 ();
 sg13g2_fill_1 FILLER_28_1334 ();
 sg13g2_decap_8 FILLER_28_1339 ();
 sg13g2_fill_1 FILLER_28_1378 ();
 sg13g2_fill_1 FILLER_28_1388 ();
 sg13g2_fill_1 FILLER_28_1399 ();
 sg13g2_fill_2 FILLER_28_1408 ();
 sg13g2_fill_1 FILLER_28_1424 ();
 sg13g2_fill_1 FILLER_28_1468 ();
 sg13g2_fill_1 FILLER_28_1495 ();
 sg13g2_fill_1 FILLER_28_1501 ();
 sg13g2_fill_1 FILLER_28_1545 ();
 sg13g2_fill_1 FILLER_28_1557 ();
 sg13g2_fill_1 FILLER_28_1562 ();
 sg13g2_fill_2 FILLER_28_1585 ();
 sg13g2_decap_4 FILLER_28_1597 ();
 sg13g2_decap_8 FILLER_28_1605 ();
 sg13g2_fill_2 FILLER_28_1612 ();
 sg13g2_decap_8 FILLER_28_1617 ();
 sg13g2_decap_4 FILLER_28_1624 ();
 sg13g2_fill_1 FILLER_28_1628 ();
 sg13g2_fill_2 FILLER_28_1640 ();
 sg13g2_fill_2 FILLER_28_1650 ();
 sg13g2_decap_8 FILLER_28_1657 ();
 sg13g2_decap_8 FILLER_28_1664 ();
 sg13g2_fill_2 FILLER_28_1671 ();
 sg13g2_fill_1 FILLER_28_1673 ();
 sg13g2_decap_8 FILLER_28_1684 ();
 sg13g2_decap_8 FILLER_28_1717 ();
 sg13g2_decap_8 FILLER_28_1724 ();
 sg13g2_decap_8 FILLER_28_1731 ();
 sg13g2_decap_4 FILLER_28_1820 ();
 sg13g2_fill_2 FILLER_28_1824 ();
 sg13g2_fill_1 FILLER_28_1852 ();
 sg13g2_decap_4 FILLER_28_1887 ();
 sg13g2_fill_1 FILLER_28_1895 ();
 sg13g2_fill_2 FILLER_28_1935 ();
 sg13g2_decap_4 FILLER_28_1954 ();
 sg13g2_fill_2 FILLER_28_1958 ();
 sg13g2_fill_2 FILLER_28_1986 ();
 sg13g2_fill_2 FILLER_28_1993 ();
 sg13g2_fill_1 FILLER_28_2024 ();
 sg13g2_fill_1 FILLER_28_2107 ();
 sg13g2_fill_2 FILLER_28_2180 ();
 sg13g2_decap_4 FILLER_28_2218 ();
 sg13g2_fill_2 FILLER_28_2222 ();
 sg13g2_fill_1 FILLER_28_2228 ();
 sg13g2_decap_4 FILLER_28_2255 ();
 sg13g2_fill_2 FILLER_28_2259 ();
 sg13g2_decap_8 FILLER_28_2265 ();
 sg13g2_decap_8 FILLER_28_2272 ();
 sg13g2_decap_8 FILLER_28_2279 ();
 sg13g2_decap_4 FILLER_28_2286 ();
 sg13g2_fill_2 FILLER_28_2290 ();
 sg13g2_fill_1 FILLER_28_2316 ();
 sg13g2_fill_1 FILLER_28_2331 ();
 sg13g2_fill_1 FILLER_28_2346 ();
 sg13g2_fill_1 FILLER_28_2388 ();
 sg13g2_decap_8 FILLER_28_2399 ();
 sg13g2_fill_1 FILLER_28_2406 ();
 sg13g2_decap_8 FILLER_28_2426 ();
 sg13g2_decap_4 FILLER_28_2433 ();
 sg13g2_fill_2 FILLER_28_2437 ();
 sg13g2_decap_8 FILLER_28_2447 ();
 sg13g2_decap_8 FILLER_28_2454 ();
 sg13g2_decap_8 FILLER_28_2461 ();
 sg13g2_decap_8 FILLER_28_2468 ();
 sg13g2_fill_2 FILLER_28_2475 ();
 sg13g2_fill_1 FILLER_28_2495 ();
 sg13g2_fill_1 FILLER_28_2506 ();
 sg13g2_decap_8 FILLER_28_2542 ();
 sg13g2_decap_4 FILLER_28_2549 ();
 sg13g2_fill_2 FILLER_28_2553 ();
 sg13g2_decap_8 FILLER_28_2559 ();
 sg13g2_decap_8 FILLER_28_2566 ();
 sg13g2_fill_2 FILLER_28_2601 ();
 sg13g2_fill_1 FILLER_28_2603 ();
 sg13g2_fill_2 FILLER_28_2614 ();
 sg13g2_fill_2 FILLER_28_2662 ();
 sg13g2_fill_2 FILLER_28_2667 ();
 sg13g2_fill_1 FILLER_28_2669 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_fill_1 FILLER_29_28 ();
 sg13g2_fill_2 FILLER_29_68 ();
 sg13g2_fill_1 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_113 ();
 sg13g2_fill_2 FILLER_29_120 ();
 sg13g2_fill_2 FILLER_29_157 ();
 sg13g2_fill_1 FILLER_29_159 ();
 sg13g2_decap_4 FILLER_29_218 ();
 sg13g2_decap_8 FILLER_29_227 ();
 sg13g2_fill_2 FILLER_29_234 ();
 sg13g2_fill_1 FILLER_29_236 ();
 sg13g2_decap_4 FILLER_29_272 ();
 sg13g2_fill_1 FILLER_29_276 ();
 sg13g2_fill_2 FILLER_29_303 ();
 sg13g2_fill_2 FILLER_29_313 ();
 sg13g2_fill_2 FILLER_29_341 ();
 sg13g2_decap_4 FILLER_29_369 ();
 sg13g2_fill_2 FILLER_29_435 ();
 sg13g2_fill_1 FILLER_29_468 ();
 sg13g2_fill_2 FILLER_29_505 ();
 sg13g2_decap_4 FILLER_29_511 ();
 sg13g2_fill_2 FILLER_29_515 ();
 sg13g2_decap_8 FILLER_29_532 ();
 sg13g2_decap_4 FILLER_29_539 ();
 sg13g2_fill_2 FILLER_29_547 ();
 sg13g2_fill_1 FILLER_29_549 ();
 sg13g2_fill_1 FILLER_29_554 ();
 sg13g2_fill_1 FILLER_29_559 ();
 sg13g2_fill_2 FILLER_29_592 ();
 sg13g2_fill_1 FILLER_29_598 ();
 sg13g2_fill_1 FILLER_29_685 ();
 sg13g2_fill_2 FILLER_29_784 ();
 sg13g2_fill_1 FILLER_29_786 ();
 sg13g2_decap_4 FILLER_29_881 ();
 sg13g2_fill_1 FILLER_29_888 ();
 sg13g2_fill_1 FILLER_29_915 ();
 sg13g2_decap_4 FILLER_29_942 ();
 sg13g2_fill_2 FILLER_29_946 ();
 sg13g2_decap_8 FILLER_29_952 ();
 sg13g2_fill_2 FILLER_29_959 ();
 sg13g2_fill_1 FILLER_29_961 ();
 sg13g2_decap_8 FILLER_29_965 ();
 sg13g2_decap_8 FILLER_29_972 ();
 sg13g2_decap_8 FILLER_29_979 ();
 sg13g2_decap_4 FILLER_29_986 ();
 sg13g2_fill_1 FILLER_29_990 ();
 sg13g2_fill_1 FILLER_29_995 ();
 sg13g2_fill_1 FILLER_29_1007 ();
 sg13g2_fill_1 FILLER_29_1014 ();
 sg13g2_fill_1 FILLER_29_1029 ();
 sg13g2_fill_2 FILLER_29_1034 ();
 sg13g2_fill_2 FILLER_29_1062 ();
 sg13g2_fill_1 FILLER_29_1064 ();
 sg13g2_fill_1 FILLER_29_1078 ();
 sg13g2_decap_4 FILLER_29_1088 ();
 sg13g2_fill_2 FILLER_29_1123 ();
 sg13g2_fill_1 FILLER_29_1146 ();
 sg13g2_fill_1 FILLER_29_1160 ();
 sg13g2_decap_8 FILLER_29_1167 ();
 sg13g2_decap_4 FILLER_29_1174 ();
 sg13g2_fill_1 FILLER_29_1178 ();
 sg13g2_decap_4 FILLER_29_1183 ();
 sg13g2_fill_1 FILLER_29_1187 ();
 sg13g2_fill_1 FILLER_29_1214 ();
 sg13g2_fill_1 FILLER_29_1224 ();
 sg13g2_decap_4 FILLER_29_1234 ();
 sg13g2_fill_2 FILLER_29_1238 ();
 sg13g2_fill_2 FILLER_29_1250 ();
 sg13g2_decap_4 FILLER_29_1262 ();
 sg13g2_decap_8 FILLER_29_1333 ();
 sg13g2_decap_8 FILLER_29_1340 ();
 sg13g2_fill_2 FILLER_29_1347 ();
 sg13g2_fill_1 FILLER_29_1349 ();
 sg13g2_decap_8 FILLER_29_1358 ();
 sg13g2_fill_1 FILLER_29_1365 ();
 sg13g2_fill_2 FILLER_29_1370 ();
 sg13g2_fill_1 FILLER_29_1426 ();
 sg13g2_fill_1 FILLER_29_1435 ();
 sg13g2_fill_1 FILLER_29_1449 ();
 sg13g2_fill_1 FILLER_29_1469 ();
 sg13g2_fill_2 FILLER_29_1492 ();
 sg13g2_fill_2 FILLER_29_1509 ();
 sg13g2_fill_2 FILLER_29_1530 ();
 sg13g2_decap_4 FILLER_29_1570 ();
 sg13g2_decap_8 FILLER_29_1588 ();
 sg13g2_decap_8 FILLER_29_1595 ();
 sg13g2_decap_8 FILLER_29_1602 ();
 sg13g2_decap_8 FILLER_29_1609 ();
 sg13g2_fill_2 FILLER_29_1616 ();
 sg13g2_fill_1 FILLER_29_1618 ();
 sg13g2_decap_4 FILLER_29_1628 ();
 sg13g2_fill_1 FILLER_29_1632 ();
 sg13g2_decap_8 FILLER_29_1642 ();
 sg13g2_decap_4 FILLER_29_1659 ();
 sg13g2_fill_2 FILLER_29_1663 ();
 sg13g2_decap_8 FILLER_29_1669 ();
 sg13g2_fill_1 FILLER_29_1676 ();
 sg13g2_decap_8 FILLER_29_1680 ();
 sg13g2_decap_8 FILLER_29_1687 ();
 sg13g2_fill_2 FILLER_29_1694 ();
 sg13g2_fill_1 FILLER_29_1696 ();
 sg13g2_decap_8 FILLER_29_1714 ();
 sg13g2_decap_8 FILLER_29_1721 ();
 sg13g2_decap_8 FILLER_29_1728 ();
 sg13g2_decap_8 FILLER_29_1735 ();
 sg13g2_decap_8 FILLER_29_1742 ();
 sg13g2_decap_4 FILLER_29_1749 ();
 sg13g2_decap_4 FILLER_29_1776 ();
 sg13g2_fill_1 FILLER_29_1786 ();
 sg13g2_fill_2 FILLER_29_1831 ();
 sg13g2_fill_2 FILLER_29_1854 ();
 sg13g2_decap_4 FILLER_29_1868 ();
 sg13g2_fill_2 FILLER_29_1876 ();
 sg13g2_fill_1 FILLER_29_1878 ();
 sg13g2_decap_8 FILLER_29_1884 ();
 sg13g2_decap_8 FILLER_29_1891 ();
 sg13g2_decap_8 FILLER_29_1898 ();
 sg13g2_decap_8 FILLER_29_1905 ();
 sg13g2_decap_8 FILLER_29_1916 ();
 sg13g2_decap_8 FILLER_29_1927 ();
 sg13g2_decap_8 FILLER_29_1934 ();
 sg13g2_fill_2 FILLER_29_1941 ();
 sg13g2_fill_1 FILLER_29_1947 ();
 sg13g2_decap_8 FILLER_29_1961 ();
 sg13g2_decap_4 FILLER_29_1968 ();
 sg13g2_fill_1 FILLER_29_1998 ();
 sg13g2_fill_2 FILLER_29_2003 ();
 sg13g2_fill_1 FILLER_29_2005 ();
 sg13g2_fill_1 FILLER_29_2062 ();
 sg13g2_fill_1 FILLER_29_2092 ();
 sg13g2_fill_1 FILLER_29_2103 ();
 sg13g2_decap_8 FILLER_29_2137 ();
 sg13g2_decap_8 FILLER_29_2144 ();
 sg13g2_fill_1 FILLER_29_2151 ();
 sg13g2_decap_8 FILLER_29_2173 ();
 sg13g2_decap_8 FILLER_29_2180 ();
 sg13g2_fill_2 FILLER_29_2187 ();
 sg13g2_fill_1 FILLER_29_2189 ();
 sg13g2_decap_8 FILLER_29_2202 ();
 sg13g2_decap_8 FILLER_29_2209 ();
 sg13g2_fill_2 FILLER_29_2216 ();
 sg13g2_fill_1 FILLER_29_2218 ();
 sg13g2_decap_4 FILLER_29_2229 ();
 sg13g2_decap_8 FILLER_29_2241 ();
 sg13g2_decap_8 FILLER_29_2261 ();
 sg13g2_fill_2 FILLER_29_2268 ();
 sg13g2_fill_1 FILLER_29_2270 ();
 sg13g2_decap_8 FILLER_29_2275 ();
 sg13g2_fill_2 FILLER_29_2282 ();
 sg13g2_fill_1 FILLER_29_2299 ();
 sg13g2_decap_4 FILLER_29_2304 ();
 sg13g2_decap_8 FILLER_29_2318 ();
 sg13g2_decap_4 FILLER_29_2330 ();
 sg13g2_decap_8 FILLER_29_2347 ();
 sg13g2_fill_2 FILLER_29_2418 ();
 sg13g2_fill_1 FILLER_29_2420 ();
 sg13g2_decap_8 FILLER_29_2457 ();
 sg13g2_decap_8 FILLER_29_2464 ();
 sg13g2_fill_2 FILLER_29_2471 ();
 sg13g2_fill_1 FILLER_29_2473 ();
 sg13g2_fill_1 FILLER_29_2504 ();
 sg13g2_decap_4 FILLER_29_2518 ();
 sg13g2_decap_8 FILLER_29_2526 ();
 sg13g2_decap_4 FILLER_29_2533 ();
 sg13g2_fill_1 FILLER_29_2573 ();
 sg13g2_decap_8 FILLER_29_2604 ();
 sg13g2_fill_2 FILLER_29_2611 ();
 sg13g2_fill_1 FILLER_29_2661 ();
 sg13g2_fill_1 FILLER_29_2669 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_98 ();
 sg13g2_decap_4 FILLER_30_129 ();
 sg13g2_decap_8 FILLER_30_137 ();
 sg13g2_decap_4 FILLER_30_149 ();
 sg13g2_fill_2 FILLER_30_163 ();
 sg13g2_decap_8 FILLER_30_236 ();
 sg13g2_decap_8 FILLER_30_243 ();
 sg13g2_decap_4 FILLER_30_250 ();
 sg13g2_fill_2 FILLER_30_258 ();
 sg13g2_fill_2 FILLER_30_270 ();
 sg13g2_fill_1 FILLER_30_280 ();
 sg13g2_fill_1 FILLER_30_289 ();
 sg13g2_fill_1 FILLER_30_300 ();
 sg13g2_fill_1 FILLER_30_327 ();
 sg13g2_fill_1 FILLER_30_332 ();
 sg13g2_fill_1 FILLER_30_352 ();
 sg13g2_fill_1 FILLER_30_410 ();
 sg13g2_fill_2 FILLER_30_428 ();
 sg13g2_fill_2 FILLER_30_433 ();
 sg13g2_fill_2 FILLER_30_454 ();
 sg13g2_fill_1 FILLER_30_456 ();
 sg13g2_decap_8 FILLER_30_480 ();
 sg13g2_decap_8 FILLER_30_487 ();
 sg13g2_fill_2 FILLER_30_494 ();
 sg13g2_decap_4 FILLER_30_500 ();
 sg13g2_decap_8 FILLER_30_527 ();
 sg13g2_decap_4 FILLER_30_534 ();
 sg13g2_fill_1 FILLER_30_601 ();
 sg13g2_fill_1 FILLER_30_689 ();
 sg13g2_fill_2 FILLER_30_734 ();
 sg13g2_fill_1 FILLER_30_749 ();
 sg13g2_fill_1 FILLER_30_770 ();
 sg13g2_fill_1 FILLER_30_816 ();
 sg13g2_fill_1 FILLER_30_833 ();
 sg13g2_fill_1 FILLER_30_860 ();
 sg13g2_fill_1 FILLER_30_961 ();
 sg13g2_decap_8 FILLER_30_977 ();
 sg13g2_decap_8 FILLER_30_984 ();
 sg13g2_decap_8 FILLER_30_996 ();
 sg13g2_fill_1 FILLER_30_1003 ();
 sg13g2_fill_2 FILLER_30_1023 ();
 sg13g2_fill_2 FILLER_30_1060 ();
 sg13g2_fill_2 FILLER_30_1071 ();
 sg13g2_fill_1 FILLER_30_1073 ();
 sg13g2_decap_4 FILLER_30_1078 ();
 sg13g2_fill_2 FILLER_30_1086 ();
 sg13g2_fill_1 FILLER_30_1088 ();
 sg13g2_fill_2 FILLER_30_1093 ();
 sg13g2_fill_2 FILLER_30_1216 ();
 sg13g2_fill_1 FILLER_30_1221 ();
 sg13g2_decap_8 FILLER_30_1243 ();
 sg13g2_decap_4 FILLER_30_1250 ();
 sg13g2_decap_4 FILLER_30_1264 ();
 sg13g2_fill_2 FILLER_30_1268 ();
 sg13g2_fill_1 FILLER_30_1274 ();
 sg13g2_decap_8 FILLER_30_1285 ();
 sg13g2_fill_1 FILLER_30_1292 ();
 sg13g2_fill_2 FILLER_30_1314 ();
 sg13g2_fill_1 FILLER_30_1334 ();
 sg13g2_decap_8 FILLER_30_1342 ();
 sg13g2_decap_8 FILLER_30_1349 ();
 sg13g2_decap_8 FILLER_30_1356 ();
 sg13g2_decap_4 FILLER_30_1363 ();
 sg13g2_fill_1 FILLER_30_1367 ();
 sg13g2_decap_8 FILLER_30_1372 ();
 sg13g2_fill_2 FILLER_30_1379 ();
 sg13g2_fill_1 FILLER_30_1381 ();
 sg13g2_fill_1 FILLER_30_1409 ();
 sg13g2_fill_2 FILLER_30_1432 ();
 sg13g2_fill_2 FILLER_30_1440 ();
 sg13g2_fill_2 FILLER_30_1490 ();
 sg13g2_fill_1 FILLER_30_1504 ();
 sg13g2_fill_2 FILLER_30_1516 ();
 sg13g2_fill_2 FILLER_30_1538 ();
 sg13g2_fill_1 FILLER_30_1576 ();
 sg13g2_decap_8 FILLER_30_1603 ();
 sg13g2_decap_8 FILLER_30_1610 ();
 sg13g2_decap_8 FILLER_30_1617 ();
 sg13g2_decap_8 FILLER_30_1628 ();
 sg13g2_decap_4 FILLER_30_1635 ();
 sg13g2_fill_1 FILLER_30_1639 ();
 sg13g2_decap_4 FILLER_30_1653 ();
 sg13g2_fill_2 FILLER_30_1657 ();
 sg13g2_fill_2 FILLER_30_1702 ();
 sg13g2_fill_1 FILLER_30_1704 ();
 sg13g2_decap_8 FILLER_30_1748 ();
 sg13g2_decap_4 FILLER_30_1755 ();
 sg13g2_fill_1 FILLER_30_1759 ();
 sg13g2_fill_2 FILLER_30_1798 ();
 sg13g2_decap_4 FILLER_30_1821 ();
 sg13g2_fill_2 FILLER_30_1825 ();
 sg13g2_fill_2 FILLER_30_1835 ();
 sg13g2_fill_2 FILLER_30_1842 ();
 sg13g2_fill_1 FILLER_30_1844 ();
 sg13g2_decap_4 FILLER_30_1857 ();
 sg13g2_fill_1 FILLER_30_1861 ();
 sg13g2_fill_1 FILLER_30_1871 ();
 sg13g2_fill_2 FILLER_30_1877 ();
 sg13g2_fill_1 FILLER_30_1895 ();
 sg13g2_fill_1 FILLER_30_1908 ();
 sg13g2_decap_4 FILLER_30_1938 ();
 sg13g2_fill_2 FILLER_30_1942 ();
 sg13g2_decap_8 FILLER_30_1956 ();
 sg13g2_fill_1 FILLER_30_1963 ();
 sg13g2_decap_8 FILLER_30_1974 ();
 sg13g2_fill_2 FILLER_30_1985 ();
 sg13g2_fill_2 FILLER_30_2013 ();
 sg13g2_fill_1 FILLER_30_2045 ();
 sg13g2_fill_1 FILLER_30_2056 ();
 sg13g2_fill_1 FILLER_30_2133 ();
 sg13g2_decap_8 FILLER_30_2170 ();
 sg13g2_decap_8 FILLER_30_2189 ();
 sg13g2_fill_1 FILLER_30_2196 ();
 sg13g2_fill_1 FILLER_30_2207 ();
 sg13g2_fill_1 FILLER_30_2229 ();
 sg13g2_decap_8 FILLER_30_2256 ();
 sg13g2_fill_1 FILLER_30_2263 ();
 sg13g2_fill_2 FILLER_30_2290 ();
 sg13g2_fill_1 FILLER_30_2292 ();
 sg13g2_decap_4 FILLER_30_2319 ();
 sg13g2_fill_2 FILLER_30_2323 ();
 sg13g2_decap_8 FILLER_30_2350 ();
 sg13g2_decap_8 FILLER_30_2357 ();
 sg13g2_fill_2 FILLER_30_2364 ();
 sg13g2_fill_1 FILLER_30_2366 ();
 sg13g2_fill_1 FILLER_30_2377 ();
 sg13g2_fill_2 FILLER_30_2383 ();
 sg13g2_fill_1 FILLER_30_2385 ();
 sg13g2_fill_2 FILLER_30_2426 ();
 sg13g2_fill_1 FILLER_30_2428 ();
 sg13g2_fill_2 FILLER_30_2526 ();
 sg13g2_decap_8 FILLER_30_2564 ();
 sg13g2_decap_8 FILLER_30_2571 ();
 sg13g2_decap_4 FILLER_30_2578 ();
 sg13g2_fill_2 FILLER_30_2582 ();
 sg13g2_fill_2 FILLER_30_2668 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_32 ();
 sg13g2_fill_2 FILLER_31_48 ();
 sg13g2_fill_1 FILLER_31_50 ();
 sg13g2_fill_2 FILLER_31_77 ();
 sg13g2_fill_1 FILLER_31_79 ();
 sg13g2_fill_2 FILLER_31_93 ();
 sg13g2_fill_1 FILLER_31_108 ();
 sg13g2_fill_2 FILLER_31_113 ();
 sg13g2_fill_2 FILLER_31_119 ();
 sg13g2_fill_2 FILLER_31_125 ();
 sg13g2_decap_8 FILLER_31_153 ();
 sg13g2_decap_8 FILLER_31_160 ();
 sg13g2_decap_8 FILLER_31_167 ();
 sg13g2_fill_2 FILLER_31_174 ();
 sg13g2_fill_2 FILLER_31_180 ();
 sg13g2_fill_1 FILLER_31_182 ();
 sg13g2_decap_4 FILLER_31_187 ();
 sg13g2_fill_2 FILLER_31_191 ();
 sg13g2_decap_8 FILLER_31_200 ();
 sg13g2_decap_4 FILLER_31_207 ();
 sg13g2_fill_1 FILLER_31_211 ();
 sg13g2_fill_2 FILLER_31_224 ();
 sg13g2_fill_1 FILLER_31_226 ();
 sg13g2_decap_4 FILLER_31_236 ();
 sg13g2_fill_1 FILLER_31_244 ();
 sg13g2_fill_2 FILLER_31_271 ();
 sg13g2_fill_2 FILLER_31_299 ();
 sg13g2_fill_2 FILLER_31_311 ();
 sg13g2_fill_1 FILLER_31_313 ();
 sg13g2_fill_2 FILLER_31_322 ();
 sg13g2_fill_1 FILLER_31_324 ();
 sg13g2_decap_4 FILLER_31_345 ();
 sg13g2_fill_1 FILLER_31_353 ();
 sg13g2_decap_4 FILLER_31_390 ();
 sg13g2_fill_2 FILLER_31_399 ();
 sg13g2_fill_2 FILLER_31_414 ();
 sg13g2_fill_1 FILLER_31_416 ();
 sg13g2_decap_8 FILLER_31_443 ();
 sg13g2_fill_2 FILLER_31_450 ();
 sg13g2_fill_1 FILLER_31_452 ();
 sg13g2_decap_8 FILLER_31_457 ();
 sg13g2_decap_4 FILLER_31_464 ();
 sg13g2_decap_8 FILLER_31_472 ();
 sg13g2_fill_2 FILLER_31_479 ();
 sg13g2_fill_1 FILLER_31_481 ();
 sg13g2_decap_8 FILLER_31_508 ();
 sg13g2_decap_4 FILLER_31_525 ();
 sg13g2_fill_2 FILLER_31_533 ();
 sg13g2_fill_2 FILLER_31_569 ();
 sg13g2_fill_2 FILLER_31_621 ();
 sg13g2_fill_1 FILLER_31_643 ();
 sg13g2_fill_1 FILLER_31_653 ();
 sg13g2_fill_2 FILLER_31_678 ();
 sg13g2_fill_2 FILLER_31_699 ();
 sg13g2_fill_1 FILLER_31_711 ();
 sg13g2_fill_1 FILLER_31_730 ();
 sg13g2_fill_1 FILLER_31_741 ();
 sg13g2_fill_1 FILLER_31_745 ();
 sg13g2_decap_4 FILLER_31_784 ();
 sg13g2_fill_1 FILLER_31_788 ();
 sg13g2_decap_4 FILLER_31_825 ();
 sg13g2_fill_1 FILLER_31_829 ();
 sg13g2_fill_2 FILLER_31_834 ();
 sg13g2_fill_1 FILLER_31_836 ();
 sg13g2_fill_1 FILLER_31_847 ();
 sg13g2_decap_8 FILLER_31_852 ();
 sg13g2_decap_8 FILLER_31_859 ();
 sg13g2_decap_8 FILLER_31_866 ();
 sg13g2_decap_4 FILLER_31_883 ();
 sg13g2_fill_1 FILLER_31_887 ();
 sg13g2_fill_2 FILLER_31_927 ();
 sg13g2_fill_2 FILLER_31_972 ();
 sg13g2_decap_4 FILLER_31_978 ();
 sg13g2_fill_2 FILLER_31_982 ();
 sg13g2_decap_8 FILLER_31_992 ();
 sg13g2_fill_1 FILLER_31_1004 ();
 sg13g2_fill_2 FILLER_31_1027 ();
 sg13g2_fill_2 FILLER_31_1047 ();
 sg13g2_fill_1 FILLER_31_1067 ();
 sg13g2_fill_1 FILLER_31_1072 ();
 sg13g2_fill_1 FILLER_31_1104 ();
 sg13g2_fill_1 FILLER_31_1139 ();
 sg13g2_fill_2 FILLER_31_1148 ();
 sg13g2_fill_1 FILLER_31_1150 ();
 sg13g2_fill_1 FILLER_31_1279 ();
 sg13g2_fill_2 FILLER_31_1321 ();
 sg13g2_fill_1 FILLER_31_1394 ();
 sg13g2_fill_1 FILLER_31_1462 ();
 sg13g2_fill_1 FILLER_31_1550 ();
 sg13g2_fill_2 FILLER_31_1602 ();
 sg13g2_fill_2 FILLER_31_1630 ();
 sg13g2_decap_8 FILLER_31_1662 ();
 sg13g2_fill_2 FILLER_31_1682 ();
 sg13g2_decap_8 FILLER_31_1710 ();
 sg13g2_decap_8 FILLER_31_1717 ();
 sg13g2_fill_1 FILLER_31_1724 ();
 sg13g2_fill_1 FILLER_31_1729 ();
 sg13g2_decap_8 FILLER_31_1764 ();
 sg13g2_decap_8 FILLER_31_1809 ();
 sg13g2_fill_1 FILLER_31_1835 ();
 sg13g2_fill_1 FILLER_31_1841 ();
 sg13g2_fill_1 FILLER_31_1847 ();
 sg13g2_fill_2 FILLER_31_1892 ();
 sg13g2_fill_1 FILLER_31_1920 ();
 sg13g2_fill_2 FILLER_31_1931 ();
 sg13g2_fill_1 FILLER_31_1950 ();
 sg13g2_decap_8 FILLER_31_1955 ();
 sg13g2_decap_8 FILLER_31_1962 ();
 sg13g2_decap_8 FILLER_31_1969 ();
 sg13g2_decap_4 FILLER_31_1976 ();
 sg13g2_decap_8 FILLER_31_1990 ();
 sg13g2_fill_2 FILLER_31_1997 ();
 sg13g2_fill_1 FILLER_31_1999 ();
 sg13g2_decap_4 FILLER_31_2020 ();
 sg13g2_fill_2 FILLER_31_2024 ();
 sg13g2_decap_4 FILLER_31_2030 ();
 sg13g2_fill_2 FILLER_31_2034 ();
 sg13g2_decap_4 FILLER_31_2102 ();
 sg13g2_fill_1 FILLER_31_2106 ();
 sg13g2_fill_2 FILLER_31_2163 ();
 sg13g2_fill_1 FILLER_31_2165 ();
 sg13g2_fill_2 FILLER_31_2187 ();
 sg13g2_fill_1 FILLER_31_2189 ();
 sg13g2_decap_4 FILLER_31_2250 ();
 sg13g2_fill_1 FILLER_31_2266 ();
 sg13g2_decap_8 FILLER_31_2293 ();
 sg13g2_fill_2 FILLER_31_2300 ();
 sg13g2_decap_8 FILLER_31_2307 ();
 sg13g2_fill_2 FILLER_31_2314 ();
 sg13g2_fill_1 FILLER_31_2321 ();
 sg13g2_fill_1 FILLER_31_2327 ();
 sg13g2_fill_1 FILLER_31_2358 ();
 sg13g2_fill_2 FILLER_31_2373 ();
 sg13g2_fill_1 FILLER_31_2375 ();
 sg13g2_decap_8 FILLER_31_2380 ();
 sg13g2_decap_8 FILLER_31_2387 ();
 sg13g2_fill_1 FILLER_31_2394 ();
 sg13g2_decap_8 FILLER_31_2399 ();
 sg13g2_decap_4 FILLER_31_2406 ();
 sg13g2_fill_2 FILLER_31_2410 ();
 sg13g2_decap_8 FILLER_31_2418 ();
 sg13g2_fill_2 FILLER_31_2425 ();
 sg13g2_decap_4 FILLER_31_2460 ();
 sg13g2_decap_4 FILLER_31_2504 ();
 sg13g2_fill_1 FILLER_31_2508 ();
 sg13g2_fill_1 FILLER_31_2549 ();
 sg13g2_fill_2 FILLER_31_2586 ();
 sg13g2_fill_2 FILLER_31_2627 ();
 sg13g2_fill_2 FILLER_31_2668 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_38 ();
 sg13g2_decap_4 FILLER_32_45 ();
 sg13g2_fill_2 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_55 ();
 sg13g2_decap_8 FILLER_32_62 ();
 sg13g2_decap_8 FILLER_32_69 ();
 sg13g2_fill_2 FILLER_32_76 ();
 sg13g2_decap_8 FILLER_32_82 ();
 sg13g2_fill_2 FILLER_32_93 ();
 sg13g2_decap_8 FILLER_32_99 ();
 sg13g2_fill_2 FILLER_32_111 ();
 sg13g2_decap_8 FILLER_32_124 ();
 sg13g2_fill_2 FILLER_32_131 ();
 sg13g2_fill_2 FILLER_32_163 ();
 sg13g2_decap_8 FILLER_32_173 ();
 sg13g2_decap_8 FILLER_32_180 ();
 sg13g2_decap_8 FILLER_32_187 ();
 sg13g2_fill_2 FILLER_32_194 ();
 sg13g2_fill_1 FILLER_32_196 ();
 sg13g2_decap_4 FILLER_32_205 ();
 sg13g2_fill_1 FILLER_32_235 ();
 sg13g2_decap_8 FILLER_32_244 ();
 sg13g2_decap_8 FILLER_32_251 ();
 sg13g2_decap_8 FILLER_32_258 ();
 sg13g2_decap_8 FILLER_32_265 ();
 sg13g2_decap_4 FILLER_32_272 ();
 sg13g2_fill_1 FILLER_32_276 ();
 sg13g2_decap_8 FILLER_32_286 ();
 sg13g2_fill_2 FILLER_32_345 ();
 sg13g2_fill_2 FILLER_32_360 ();
 sg13g2_fill_1 FILLER_32_395 ();
 sg13g2_fill_1 FILLER_32_406 ();
 sg13g2_decap_8 FILLER_32_447 ();
 sg13g2_decap_4 FILLER_32_454 ();
 sg13g2_fill_1 FILLER_32_458 ();
 sg13g2_decap_8 FILLER_32_463 ();
 sg13g2_decap_8 FILLER_32_470 ();
 sg13g2_decap_8 FILLER_32_477 ();
 sg13g2_fill_2 FILLER_32_488 ();
 sg13g2_decap_4 FILLER_32_494 ();
 sg13g2_fill_1 FILLER_32_498 ();
 sg13g2_fill_2 FILLER_32_539 ();
 sg13g2_fill_2 FILLER_32_583 ();
 sg13g2_fill_1 FILLER_32_585 ();
 sg13g2_fill_2 FILLER_32_596 ();
 sg13g2_fill_1 FILLER_32_642 ();
 sg13g2_fill_2 FILLER_32_654 ();
 sg13g2_fill_1 FILLER_32_694 ();
 sg13g2_fill_2 FILLER_32_704 ();
 sg13g2_fill_1 FILLER_32_750 ();
 sg13g2_fill_2 FILLER_32_774 ();
 sg13g2_decap_8 FILLER_32_785 ();
 sg13g2_decap_4 FILLER_32_792 ();
 sg13g2_decap_4 FILLER_32_800 ();
 sg13g2_fill_2 FILLER_32_851 ();
 sg13g2_decap_8 FILLER_32_857 ();
 sg13g2_decap_8 FILLER_32_864 ();
 sg13g2_decap_8 FILLER_32_871 ();
 sg13g2_fill_2 FILLER_32_878 ();
 sg13g2_fill_1 FILLER_32_880 ();
 sg13g2_decap_4 FILLER_32_902 ();
 sg13g2_decap_4 FILLER_32_927 ();
 sg13g2_fill_1 FILLER_32_931 ();
 sg13g2_fill_2 FILLER_32_974 ();
 sg13g2_fill_2 FILLER_32_985 ();
 sg13g2_fill_1 FILLER_32_987 ();
 sg13g2_decap_8 FILLER_32_1094 ();
 sg13g2_decap_4 FILLER_32_1101 ();
 sg13g2_fill_2 FILLER_32_1105 ();
 sg13g2_fill_2 FILLER_32_1120 ();
 sg13g2_fill_1 FILLER_32_1122 ();
 sg13g2_decap_8 FILLER_32_1136 ();
 sg13g2_fill_2 FILLER_32_1148 ();
 sg13g2_fill_1 FILLER_32_1155 ();
 sg13g2_fill_1 FILLER_32_1176 ();
 sg13g2_fill_2 FILLER_32_1203 ();
 sg13g2_fill_2 FILLER_32_1209 ();
 sg13g2_fill_2 FILLER_32_1279 ();
 sg13g2_fill_1 FILLER_32_1281 ();
 sg13g2_fill_1 FILLER_32_1292 ();
 sg13g2_fill_1 FILLER_32_1316 ();
 sg13g2_decap_4 FILLER_32_1335 ();
 sg13g2_decap_4 FILLER_32_1375 ();
 sg13g2_fill_1 FILLER_32_1379 ();
 sg13g2_fill_2 FILLER_32_1393 ();
 sg13g2_fill_2 FILLER_32_1428 ();
 sg13g2_fill_2 FILLER_32_1458 ();
 sg13g2_fill_1 FILLER_32_1463 ();
 sg13g2_fill_2 FILLER_32_1528 ();
 sg13g2_fill_1 FILLER_32_1545 ();
 sg13g2_fill_2 FILLER_32_1551 ();
 sg13g2_fill_2 FILLER_32_1558 ();
 sg13g2_fill_2 FILLER_32_1586 ();
 sg13g2_fill_1 FILLER_32_1588 ();
 sg13g2_decap_8 FILLER_32_1619 ();
 sg13g2_fill_2 FILLER_32_1626 ();
 sg13g2_fill_1 FILLER_32_1628 ();
 sg13g2_fill_2 FILLER_32_1638 ();
 sg13g2_fill_2 FILLER_32_1666 ();
 sg13g2_fill_2 FILLER_32_1672 ();
 sg13g2_fill_1 FILLER_32_1674 ();
 sg13g2_decap_8 FILLER_32_1701 ();
 sg13g2_decap_8 FILLER_32_1708 ();
 sg13g2_decap_4 FILLER_32_1729 ();
 sg13g2_fill_2 FILLER_32_1733 ();
 sg13g2_fill_1 FILLER_32_1743 ();
 sg13g2_fill_2 FILLER_32_1748 ();
 sg13g2_fill_2 FILLER_32_1789 ();
 sg13g2_decap_8 FILLER_32_1795 ();
 sg13g2_fill_1 FILLER_32_1802 ();
 sg13g2_fill_2 FILLER_32_1880 ();
 sg13g2_fill_1 FILLER_32_1882 ();
 sg13g2_fill_1 FILLER_32_1897 ();
 sg13g2_fill_2 FILLER_32_1913 ();
 sg13g2_fill_1 FILLER_32_1920 ();
 sg13g2_fill_2 FILLER_32_1926 ();
 sg13g2_fill_2 FILLER_32_1965 ();
 sg13g2_decap_4 FILLER_32_1971 ();
 sg13g2_decap_4 FILLER_32_2001 ();
 sg13g2_fill_2 FILLER_32_2005 ();
 sg13g2_fill_2 FILLER_32_2011 ();
 sg13g2_fill_1 FILLER_32_2013 ();
 sg13g2_decap_8 FILLER_32_2024 ();
 sg13g2_fill_2 FILLER_32_2031 ();
 sg13g2_decap_4 FILLER_32_2038 ();
 sg13g2_fill_2 FILLER_32_2042 ();
 sg13g2_fill_1 FILLER_32_2069 ();
 sg13g2_decap_8 FILLER_32_2094 ();
 sg13g2_fill_1 FILLER_32_2101 ();
 sg13g2_fill_2 FILLER_32_2138 ();
 sg13g2_decap_4 FILLER_32_2161 ();
 sg13g2_fill_1 FILLER_32_2195 ();
 sg13g2_decap_8 FILLER_32_2204 ();
 sg13g2_fill_1 FILLER_32_2211 ();
 sg13g2_decap_4 FILLER_32_2222 ();
 sg13g2_decap_4 FILLER_32_2256 ();
 sg13g2_fill_2 FILLER_32_2260 ();
 sg13g2_fill_2 FILLER_32_2272 ();
 sg13g2_fill_1 FILLER_32_2274 ();
 sg13g2_decap_4 FILLER_32_2279 ();
 sg13g2_decap_8 FILLER_32_2288 ();
 sg13g2_fill_2 FILLER_32_2295 ();
 sg13g2_fill_1 FILLER_32_2301 ();
 sg13g2_decap_8 FILLER_32_2307 ();
 sg13g2_fill_1 FILLER_32_2314 ();
 sg13g2_decap_4 FILLER_32_2351 ();
 sg13g2_fill_2 FILLER_32_2395 ();
 sg13g2_fill_1 FILLER_32_2443 ();
 sg13g2_fill_1 FILLER_32_2454 ();
 sg13g2_fill_2 FILLER_32_2481 ();
 sg13g2_fill_1 FILLER_32_2504 ();
 sg13g2_fill_1 FILLER_32_2539 ();
 sg13g2_decap_4 FILLER_32_2564 ();
 sg13g2_fill_2 FILLER_32_2568 ();
 sg13g2_decap_8 FILLER_32_2574 ();
 sg13g2_fill_2 FILLER_32_2605 ();
 sg13g2_fill_1 FILLER_32_2607 ();
 sg13g2_decap_4 FILLER_32_2664 ();
 sg13g2_fill_2 FILLER_32_2668 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_41 ();
 sg13g2_fill_1 FILLER_33_43 ();
 sg13g2_decap_4 FILLER_33_57 ();
 sg13g2_fill_2 FILLER_33_61 ();
 sg13g2_fill_1 FILLER_33_81 ();
 sg13g2_fill_1 FILLER_33_86 ();
 sg13g2_fill_2 FILLER_33_95 ();
 sg13g2_fill_2 FILLER_33_189 ();
 sg13g2_fill_2 FILLER_33_197 ();
 sg13g2_fill_1 FILLER_33_199 ();
 sg13g2_fill_1 FILLER_33_205 ();
 sg13g2_fill_2 FILLER_33_214 ();
 sg13g2_decap_4 FILLER_33_247 ();
 sg13g2_fill_2 FILLER_33_251 ();
 sg13g2_decap_4 FILLER_33_262 ();
 sg13g2_fill_1 FILLER_33_266 ();
 sg13g2_decap_8 FILLER_33_280 ();
 sg13g2_decap_8 FILLER_33_287 ();
 sg13g2_fill_1 FILLER_33_312 ();
 sg13g2_fill_1 FILLER_33_319 ();
 sg13g2_fill_1 FILLER_33_330 ();
 sg13g2_fill_2 FILLER_33_367 ();
 sg13g2_fill_1 FILLER_33_369 ();
 sg13g2_fill_1 FILLER_33_376 ();
 sg13g2_fill_2 FILLER_33_441 ();
 sg13g2_fill_2 FILLER_33_447 ();
 sg13g2_fill_2 FILLER_33_483 ();
 sg13g2_fill_1 FILLER_33_485 ();
 sg13g2_fill_2 FILLER_33_494 ();
 sg13g2_fill_2 FILLER_33_525 ();
 sg13g2_fill_2 FILLER_33_557 ();
 sg13g2_fill_2 FILLER_33_657 ();
 sg13g2_fill_2 FILLER_33_663 ();
 sg13g2_fill_1 FILLER_33_706 ();
 sg13g2_fill_1 FILLER_33_730 ();
 sg13g2_fill_1 FILLER_33_745 ();
 sg13g2_fill_2 FILLER_33_766 ();
 sg13g2_fill_1 FILLER_33_779 ();
 sg13g2_fill_1 FILLER_33_790 ();
 sg13g2_decap_8 FILLER_33_795 ();
 sg13g2_decap_4 FILLER_33_868 ();
 sg13g2_decap_8 FILLER_33_876 ();
 sg13g2_decap_8 FILLER_33_893 ();
 sg13g2_decap_8 FILLER_33_900 ();
 sg13g2_decap_8 FILLER_33_907 ();
 sg13g2_decap_8 FILLER_33_914 ();
 sg13g2_decap_8 FILLER_33_921 ();
 sg13g2_decap_8 FILLER_33_928 ();
 sg13g2_fill_1 FILLER_33_935 ();
 sg13g2_fill_1 FILLER_33_981 ();
 sg13g2_fill_2 FILLER_33_1013 ();
 sg13g2_fill_2 FILLER_33_1019 ();
 sg13g2_fill_2 FILLER_33_1086 ();
 sg13g2_fill_2 FILLER_33_1092 ();
 sg13g2_decap_8 FILLER_33_1154 ();
 sg13g2_decap_8 FILLER_33_1165 ();
 sg13g2_fill_2 FILLER_33_1172 ();
 sg13g2_decap_4 FILLER_33_1191 ();
 sg13g2_fill_1 FILLER_33_1195 ();
 sg13g2_decap_4 FILLER_33_1201 ();
 sg13g2_fill_1 FILLER_33_1205 ();
 sg13g2_fill_2 FILLER_33_1237 ();
 sg13g2_fill_1 FILLER_33_1239 ();
 sg13g2_fill_1 FILLER_33_1266 ();
 sg13g2_fill_1 FILLER_33_1298 ();
 sg13g2_fill_1 FILLER_33_1313 ();
 sg13g2_decap_4 FILLER_33_1340 ();
 sg13g2_decap_4 FILLER_33_1384 ();
 sg13g2_fill_2 FILLER_33_1388 ();
 sg13g2_fill_1 FILLER_33_1405 ();
 sg13g2_decap_8 FILLER_33_1410 ();
 sg13g2_fill_1 FILLER_33_1417 ();
 sg13g2_fill_1 FILLER_33_1442 ();
 sg13g2_fill_2 FILLER_33_1450 ();
 sg13g2_fill_1 FILLER_33_1489 ();
 sg13g2_fill_1 FILLER_33_1503 ();
 sg13g2_fill_2 FILLER_33_1523 ();
 sg13g2_fill_1 FILLER_33_1542 ();
 sg13g2_fill_1 FILLER_33_1569 ();
 sg13g2_fill_1 FILLER_33_1575 ();
 sg13g2_fill_1 FILLER_33_1580 ();
 sg13g2_decap_8 FILLER_33_1597 ();
 sg13g2_decap_4 FILLER_33_1604 ();
 sg13g2_fill_2 FILLER_33_1634 ();
 sg13g2_fill_1 FILLER_33_1636 ();
 sg13g2_fill_2 FILLER_33_1695 ();
 sg13g2_fill_1 FILLER_33_1707 ();
 sg13g2_fill_1 FILLER_33_1734 ();
 sg13g2_decap_4 FILLER_33_1739 ();
 sg13g2_fill_2 FILLER_33_1743 ();
 sg13g2_fill_1 FILLER_33_1749 ();
 sg13g2_fill_1 FILLER_33_1755 ();
 sg13g2_fill_2 FILLER_33_1760 ();
 sg13g2_fill_1 FILLER_33_1762 ();
 sg13g2_fill_1 FILLER_33_1768 ();
 sg13g2_fill_1 FILLER_33_1773 ();
 sg13g2_decap_8 FILLER_33_1800 ();
 sg13g2_fill_1 FILLER_33_1822 ();
 sg13g2_fill_1 FILLER_33_1843 ();
 sg13g2_fill_1 FILLER_33_1849 ();
 sg13g2_fill_2 FILLER_33_1860 ();
 sg13g2_fill_1 FILLER_33_1862 ();
 sg13g2_fill_1 FILLER_33_1935 ();
 sg13g2_fill_1 FILLER_33_1942 ();
 sg13g2_fill_2 FILLER_33_1965 ();
 sg13g2_fill_2 FILLER_33_2005 ();
 sg13g2_fill_2 FILLER_33_2012 ();
 sg13g2_fill_2 FILLER_33_2018 ();
 sg13g2_fill_2 FILLER_33_2046 ();
 sg13g2_decap_8 FILLER_33_2077 ();
 sg13g2_decap_4 FILLER_33_2084 ();
 sg13g2_decap_8 FILLER_33_2122 ();
 sg13g2_fill_2 FILLER_33_2129 ();
 sg13g2_decap_8 FILLER_33_2156 ();
 sg13g2_fill_2 FILLER_33_2163 ();
 sg13g2_fill_1 FILLER_33_2165 ();
 sg13g2_fill_2 FILLER_33_2176 ();
 sg13g2_decap_8 FILLER_33_2203 ();
 sg13g2_decap_8 FILLER_33_2210 ();
 sg13g2_fill_2 FILLER_33_2217 ();
 sg13g2_fill_1 FILLER_33_2219 ();
 sg13g2_decap_8 FILLER_33_2230 ();
 sg13g2_fill_1 FILLER_33_2237 ();
 sg13g2_fill_1 FILLER_33_2249 ();
 sg13g2_decap_8 FILLER_33_2264 ();
 sg13g2_fill_2 FILLER_33_2271 ();
 sg13g2_decap_8 FILLER_33_2283 ();
 sg13g2_decap_8 FILLER_33_2290 ();
 sg13g2_decap_4 FILLER_33_2297 ();
 sg13g2_fill_1 FILLER_33_2301 ();
 sg13g2_fill_1 FILLER_33_2336 ();
 sg13g2_fill_1 FILLER_33_2409 ();
 sg13g2_decap_8 FILLER_33_2424 ();
 sg13g2_fill_2 FILLER_33_2431 ();
 sg13g2_fill_1 FILLER_33_2449 ();
 sg13g2_fill_2 FILLER_33_2468 ();
 sg13g2_decap_8 FILLER_33_2506 ();
 sg13g2_fill_1 FILLER_33_2513 ();
 sg13g2_decap_4 FILLER_33_2530 ();
 sg13g2_fill_2 FILLER_33_2534 ();
 sg13g2_fill_2 FILLER_33_2549 ();
 sg13g2_fill_2 FILLER_33_2582 ();
 sg13g2_fill_1 FILLER_33_2594 ();
 sg13g2_fill_2 FILLER_33_2633 ();
 sg13g2_fill_1 FILLER_33_2652 ();
 sg13g2_decap_8 FILLER_33_2663 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_4 FILLER_34_66 ();
 sg13g2_fill_2 FILLER_34_105 ();
 sg13g2_fill_1 FILLER_34_107 ();
 sg13g2_fill_1 FILLER_34_134 ();
 sg13g2_fill_2 FILLER_34_140 ();
 sg13g2_fill_2 FILLER_34_167 ();
 sg13g2_fill_2 FILLER_34_233 ();
 sg13g2_fill_2 FILLER_34_266 ();
 sg13g2_fill_2 FILLER_34_273 ();
 sg13g2_fill_2 FILLER_34_281 ();
 sg13g2_fill_1 FILLER_34_297 ();
 sg13g2_decap_4 FILLER_34_313 ();
 sg13g2_fill_1 FILLER_34_317 ();
 sg13g2_fill_2 FILLER_34_324 ();
 sg13g2_decap_8 FILLER_34_340 ();
 sg13g2_fill_2 FILLER_34_351 ();
 sg13g2_fill_1 FILLER_34_353 ();
 sg13g2_decap_4 FILLER_34_364 ();
 sg13g2_fill_2 FILLER_34_368 ();
 sg13g2_fill_1 FILLER_34_376 ();
 sg13g2_fill_2 FILLER_34_396 ();
 sg13g2_fill_1 FILLER_34_398 ();
 sg13g2_fill_2 FILLER_34_422 ();
 sg13g2_fill_1 FILLER_34_447 ();
 sg13g2_fill_2 FILLER_34_453 ();
 sg13g2_fill_2 FILLER_34_474 ();
 sg13g2_fill_1 FILLER_34_476 ();
 sg13g2_fill_2 FILLER_34_519 ();
 sg13g2_fill_1 FILLER_34_521 ();
 sg13g2_decap_8 FILLER_34_532 ();
 sg13g2_fill_1 FILLER_34_539 ();
 sg13g2_decap_8 FILLER_34_566 ();
 sg13g2_fill_1 FILLER_34_573 ();
 sg13g2_fill_2 FILLER_34_584 ();
 sg13g2_fill_1 FILLER_34_586 ();
 sg13g2_fill_2 FILLER_34_614 ();
 sg13g2_fill_2 FILLER_34_624 ();
 sg13g2_fill_2 FILLER_34_634 ();
 sg13g2_fill_2 FILLER_34_725 ();
 sg13g2_fill_1 FILLER_34_732 ();
 sg13g2_fill_1 FILLER_34_742 ();
 sg13g2_fill_1 FILLER_34_752 ();
 sg13g2_fill_1 FILLER_34_756 ();
 sg13g2_fill_1 FILLER_34_762 ();
 sg13g2_fill_1 FILLER_34_775 ();
 sg13g2_fill_2 FILLER_34_784 ();
 sg13g2_decap_4 FILLER_34_808 ();
 sg13g2_decap_8 FILLER_34_853 ();
 sg13g2_decap_4 FILLER_34_860 ();
 sg13g2_fill_1 FILLER_34_864 ();
 sg13g2_decap_4 FILLER_34_891 ();
 sg13g2_fill_2 FILLER_34_895 ();
 sg13g2_fill_2 FILLER_34_918 ();
 sg13g2_fill_1 FILLER_34_920 ();
 sg13g2_fill_2 FILLER_34_937 ();
 sg13g2_fill_2 FILLER_34_981 ();
 sg13g2_fill_1 FILLER_34_983 ();
 sg13g2_fill_2 FILLER_34_997 ();
 sg13g2_fill_2 FILLER_34_1003 ();
 sg13g2_fill_1 FILLER_34_1031 ();
 sg13g2_fill_2 FILLER_34_1063 ();
 sg13g2_fill_1 FILLER_34_1065 ();
 sg13g2_fill_2 FILLER_34_1070 ();
 sg13g2_fill_1 FILLER_34_1072 ();
 sg13g2_fill_2 FILLER_34_1077 ();
 sg13g2_fill_1 FILLER_34_1079 ();
 sg13g2_decap_8 FILLER_34_1111 ();
 sg13g2_fill_2 FILLER_34_1118 ();
 sg13g2_fill_1 FILLER_34_1120 ();
 sg13g2_fill_1 FILLER_34_1152 ();
 sg13g2_fill_1 FILLER_34_1179 ();
 sg13g2_fill_1 FILLER_34_1201 ();
 sg13g2_fill_1 FILLER_34_1207 ();
 sg13g2_fill_2 FILLER_34_1222 ();
 sg13g2_fill_1 FILLER_34_1254 ();
 sg13g2_fill_1 FILLER_34_1259 ();
 sg13g2_fill_1 FILLER_34_1265 ();
 sg13g2_fill_2 FILLER_34_1276 ();
 sg13g2_fill_2 FILLER_34_1304 ();
 sg13g2_fill_2 FILLER_34_1316 ();
 sg13g2_decap_8 FILLER_34_1344 ();
 sg13g2_decap_8 FILLER_34_1355 ();
 sg13g2_fill_2 FILLER_34_1362 ();
 sg13g2_fill_1 FILLER_34_1364 ();
 sg13g2_fill_1 FILLER_34_1368 ();
 sg13g2_fill_2 FILLER_34_1374 ();
 sg13g2_fill_1 FILLER_34_1376 ();
 sg13g2_decap_4 FILLER_34_1417 ();
 sg13g2_fill_1 FILLER_34_1421 ();
 sg13g2_fill_2 FILLER_34_1425 ();
 sg13g2_fill_1 FILLER_34_1453 ();
 sg13g2_fill_1 FILLER_34_1465 ();
 sg13g2_fill_1 FILLER_34_1472 ();
 sg13g2_fill_2 FILLER_34_1481 ();
 sg13g2_fill_1 FILLER_34_1493 ();
 sg13g2_fill_2 FILLER_34_1505 ();
 sg13g2_fill_2 FILLER_34_1536 ();
 sg13g2_fill_1 FILLER_34_1562 ();
 sg13g2_fill_2 FILLER_34_1568 ();
 sg13g2_decap_8 FILLER_34_1615 ();
 sg13g2_fill_2 FILLER_34_1622 ();
 sg13g2_decap_8 FILLER_34_1629 ();
 sg13g2_decap_4 FILLER_34_1636 ();
 sg13g2_fill_2 FILLER_34_1640 ();
 sg13g2_decap_4 FILLER_34_1646 ();
 sg13g2_fill_1 FILLER_34_1685 ();
 sg13g2_fill_1 FILLER_34_1693 ();
 sg13g2_fill_1 FILLER_34_1768 ();
 sg13g2_fill_1 FILLER_34_1778 ();
 sg13g2_fill_1 FILLER_34_1783 ();
 sg13g2_decap_8 FILLER_34_1803 ();
 sg13g2_fill_1 FILLER_34_1810 ();
 sg13g2_fill_2 FILLER_34_1854 ();
 sg13g2_fill_1 FILLER_34_1856 ();
 sg13g2_fill_2 FILLER_34_1890 ();
 sg13g2_fill_1 FILLER_34_1902 ();
 sg13g2_fill_1 FILLER_34_1913 ();
 sg13g2_fill_1 FILLER_34_1919 ();
 sg13g2_fill_2 FILLER_34_1994 ();
 sg13g2_fill_2 FILLER_34_2000 ();
 sg13g2_fill_1 FILLER_34_2002 ();
 sg13g2_fill_2 FILLER_34_2013 ();
 sg13g2_fill_1 FILLER_34_2015 ();
 sg13g2_decap_8 FILLER_34_2021 ();
 sg13g2_fill_1 FILLER_34_2028 ();
 sg13g2_decap_4 FILLER_34_2033 ();
 sg13g2_decap_8 FILLER_34_2077 ();
 sg13g2_decap_8 FILLER_34_2084 ();
 sg13g2_fill_1 FILLER_34_2091 ();
 sg13g2_decap_8 FILLER_34_2118 ();
 sg13g2_decap_8 FILLER_34_2125 ();
 sg13g2_fill_2 FILLER_34_2159 ();
 sg13g2_fill_2 FILLER_34_2177 ();
 sg13g2_fill_1 FILLER_34_2179 ();
 sg13g2_decap_8 FILLER_34_2216 ();
 sg13g2_decap_4 FILLER_34_2223 ();
 sg13g2_decap_8 FILLER_34_2311 ();
 sg13g2_decap_4 FILLER_34_2318 ();
 sg13g2_fill_1 FILLER_34_2322 ();
 sg13g2_fill_2 FILLER_34_2327 ();
 sg13g2_decap_8 FILLER_34_2339 ();
 sg13g2_fill_1 FILLER_34_2346 ();
 sg13g2_fill_2 FILLER_34_2357 ();
 sg13g2_fill_2 FILLER_34_2365 ();
 sg13g2_fill_2 FILLER_34_2399 ();
 sg13g2_fill_1 FILLER_34_2401 ();
 sg13g2_fill_1 FILLER_34_2428 ();
 sg13g2_fill_1 FILLER_34_2434 ();
 sg13g2_fill_1 FILLER_34_2439 ();
 sg13g2_fill_2 FILLER_34_2470 ();
 sg13g2_fill_1 FILLER_34_2482 ();
 sg13g2_fill_2 FILLER_34_2493 ();
 sg13g2_fill_2 FILLER_34_2499 ();
 sg13g2_fill_2 FILLER_34_2507 ();
 sg13g2_decap_4 FILLER_34_2515 ();
 sg13g2_fill_1 FILLER_34_2538 ();
 sg13g2_fill_1 FILLER_34_2580 ();
 sg13g2_fill_1 FILLER_34_2620 ();
 sg13g2_fill_2 FILLER_34_2664 ();
 sg13g2_fill_1 FILLER_34_2669 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_12 ();
 sg13g2_decap_8 FILLER_35_55 ();
 sg13g2_fill_2 FILLER_35_66 ();
 sg13g2_decap_4 FILLER_35_77 ();
 sg13g2_fill_2 FILLER_35_81 ();
 sg13g2_decap_8 FILLER_35_87 ();
 sg13g2_fill_1 FILLER_35_94 ();
 sg13g2_fill_1 FILLER_35_99 ();
 sg13g2_fill_1 FILLER_35_131 ();
 sg13g2_fill_1 FILLER_35_146 ();
 sg13g2_fill_1 FILLER_35_162 ();
 sg13g2_fill_1 FILLER_35_167 ();
 sg13g2_fill_1 FILLER_35_173 ();
 sg13g2_fill_1 FILLER_35_179 ();
 sg13g2_decap_4 FILLER_35_184 ();
 sg13g2_fill_1 FILLER_35_188 ();
 sg13g2_fill_2 FILLER_35_303 ();
 sg13g2_fill_2 FILLER_35_323 ();
 sg13g2_fill_1 FILLER_35_331 ();
 sg13g2_decap_8 FILLER_35_337 ();
 sg13g2_fill_1 FILLER_35_344 ();
 sg13g2_fill_1 FILLER_35_350 ();
 sg13g2_fill_1 FILLER_35_385 ();
 sg13g2_decap_8 FILLER_35_412 ();
 sg13g2_fill_2 FILLER_35_419 ();
 sg13g2_fill_1 FILLER_35_421 ();
 sg13g2_fill_1 FILLER_35_426 ();
 sg13g2_fill_1 FILLER_35_469 ();
 sg13g2_fill_1 FILLER_35_475 ();
 sg13g2_decap_8 FILLER_35_521 ();
 sg13g2_decap_4 FILLER_35_528 ();
 sg13g2_fill_2 FILLER_35_532 ();
 sg13g2_fill_1 FILLER_35_597 ();
 sg13g2_fill_1 FILLER_35_617 ();
 sg13g2_fill_2 FILLER_35_671 ();
 sg13g2_fill_2 FILLER_35_698 ();
 sg13g2_fill_1 FILLER_35_720 ();
 sg13g2_fill_1 FILLER_35_726 ();
 sg13g2_fill_2 FILLER_35_751 ();
 sg13g2_fill_1 FILLER_35_758 ();
 sg13g2_fill_1 FILLER_35_772 ();
 sg13g2_fill_2 FILLER_35_788 ();
 sg13g2_fill_2 FILLER_35_802 ();
 sg13g2_decap_8 FILLER_35_808 ();
 sg13g2_fill_2 FILLER_35_815 ();
 sg13g2_decap_4 FILLER_35_853 ();
 sg13g2_decap_4 FILLER_35_887 ();
 sg13g2_fill_2 FILLER_35_891 ();
 sg13g2_fill_2 FILLER_35_947 ();
 sg13g2_fill_2 FILLER_35_953 ();
 sg13g2_fill_1 FILLER_35_960 ();
 sg13g2_fill_2 FILLER_35_965 ();
 sg13g2_fill_1 FILLER_35_1003 ();
 sg13g2_fill_2 FILLER_35_1009 ();
 sg13g2_fill_2 FILLER_35_1015 ();
 sg13g2_fill_2 FILLER_35_1021 ();
 sg13g2_fill_1 FILLER_35_1041 ();
 sg13g2_decap_8 FILLER_35_1046 ();
 sg13g2_fill_2 FILLER_35_1053 ();
 sg13g2_fill_1 FILLER_35_1055 ();
 sg13g2_fill_1 FILLER_35_1065 ();
 sg13g2_fill_2 FILLER_35_1122 ();
 sg13g2_fill_2 FILLER_35_1129 ();
 sg13g2_fill_1 FILLER_35_1131 ();
 sg13g2_fill_2 FILLER_35_1140 ();
 sg13g2_fill_1 FILLER_35_1142 ();
 sg13g2_fill_1 FILLER_35_1147 ();
 sg13g2_decap_4 FILLER_35_1169 ();
 sg13g2_fill_2 FILLER_35_1173 ();
 sg13g2_decap_8 FILLER_35_1216 ();
 sg13g2_decap_8 FILLER_35_1223 ();
 sg13g2_fill_2 FILLER_35_1240 ();
 sg13g2_fill_1 FILLER_35_1242 ();
 sg13g2_decap_4 FILLER_35_1258 ();
 sg13g2_fill_2 FILLER_35_1262 ();
 sg13g2_fill_2 FILLER_35_1281 ();
 sg13g2_fill_1 FILLER_35_1327 ();
 sg13g2_decap_8 FILLER_35_1336 ();
 sg13g2_fill_2 FILLER_35_1343 ();
 sg13g2_fill_1 FILLER_35_1345 ();
 sg13g2_decap_8 FILLER_35_1382 ();
 sg13g2_fill_2 FILLER_35_1398 ();
 sg13g2_fill_1 FILLER_35_1400 ();
 sg13g2_fill_2 FILLER_35_1427 ();
 sg13g2_fill_1 FILLER_35_1429 ();
 sg13g2_fill_2 FILLER_35_1479 ();
 sg13g2_fill_1 FILLER_35_1525 ();
 sg13g2_fill_1 FILLER_35_1543 ();
 sg13g2_fill_2 FILLER_35_1564 ();
 sg13g2_fill_1 FILLER_35_1587 ();
 sg13g2_fill_2 FILLER_35_1591 ();
 sg13g2_decap_8 FILLER_35_1636 ();
 sg13g2_fill_2 FILLER_35_1643 ();
 sg13g2_fill_1 FILLER_35_1645 ();
 sg13g2_fill_1 FILLER_35_1682 ();
 sg13g2_fill_1 FILLER_35_1691 ();
 sg13g2_fill_2 FILLER_35_1722 ();
 sg13g2_fill_2 FILLER_35_1734 ();
 sg13g2_fill_1 FILLER_35_1740 ();
 sg13g2_fill_2 FILLER_35_1767 ();
 sg13g2_decap_8 FILLER_35_1804 ();
 sg13g2_decap_8 FILLER_35_1811 ();
 sg13g2_decap_4 FILLER_35_1818 ();
 sg13g2_fill_1 FILLER_35_1845 ();
 sg13g2_fill_1 FILLER_35_1851 ();
 sg13g2_fill_1 FILLER_35_1857 ();
 sg13g2_fill_2 FILLER_35_1865 ();
 sg13g2_fill_2 FILLER_35_1876 ();
 sg13g2_fill_2 FILLER_35_1909 ();
 sg13g2_fill_1 FILLER_35_1911 ();
 sg13g2_fill_2 FILLER_35_1961 ();
 sg13g2_fill_1 FILLER_35_1984 ();
 sg13g2_fill_1 FILLER_35_1996 ();
 sg13g2_fill_2 FILLER_35_2018 ();
 sg13g2_fill_1 FILLER_35_2024 ();
 sg13g2_fill_2 FILLER_35_2029 ();
 sg13g2_fill_1 FILLER_35_2035 ();
 sg13g2_fill_1 FILLER_35_2040 ();
 sg13g2_fill_1 FILLER_35_2051 ();
 sg13g2_fill_2 FILLER_35_2083 ();
 sg13g2_fill_1 FILLER_35_2116 ();
 sg13g2_decap_4 FILLER_35_2218 ();
 sg13g2_fill_1 FILLER_35_2222 ();
 sg13g2_fill_2 FILLER_35_2271 ();
 sg13g2_fill_1 FILLER_35_2277 ();
 sg13g2_fill_1 FILLER_35_2288 ();
 sg13g2_fill_2 FILLER_35_2294 ();
 sg13g2_decap_8 FILLER_35_2338 ();
 sg13g2_decap_8 FILLER_35_2345 ();
 sg13g2_decap_4 FILLER_35_2352 ();
 sg13g2_fill_1 FILLER_35_2356 ();
 sg13g2_fill_1 FILLER_35_2373 ();
 sg13g2_fill_1 FILLER_35_2422 ();
 sg13g2_decap_8 FILLER_35_2463 ();
 sg13g2_fill_2 FILLER_35_2470 ();
 sg13g2_fill_2 FILLER_35_2478 ();
 sg13g2_fill_2 FILLER_35_2486 ();
 sg13g2_fill_2 FILLER_35_2525 ();
 sg13g2_fill_1 FILLER_35_2557 ();
 sg13g2_fill_1 FILLER_35_2603 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_32 ();
 sg13g2_fill_1 FILLER_36_42 ();
 sg13g2_fill_2 FILLER_36_48 ();
 sg13g2_fill_2 FILLER_36_54 ();
 sg13g2_fill_2 FILLER_36_82 ();
 sg13g2_decap_4 FILLER_36_88 ();
 sg13g2_fill_2 FILLER_36_92 ();
 sg13g2_fill_1 FILLER_36_147 ();
 sg13g2_fill_2 FILLER_36_165 ();
 sg13g2_fill_1 FILLER_36_167 ();
 sg13g2_fill_2 FILLER_36_207 ();
 sg13g2_fill_2 FILLER_36_214 ();
 sg13g2_fill_1 FILLER_36_241 ();
 sg13g2_fill_2 FILLER_36_293 ();
 sg13g2_fill_1 FILLER_36_329 ();
 sg13g2_fill_2 FILLER_36_335 ();
 sg13g2_fill_1 FILLER_36_337 ();
 sg13g2_fill_2 FILLER_36_359 ();
 sg13g2_fill_1 FILLER_36_361 ();
 sg13g2_fill_2 FILLER_36_382 ();
 sg13g2_fill_1 FILLER_36_384 ();
 sg13g2_decap_4 FILLER_36_417 ();
 sg13g2_fill_2 FILLER_36_421 ();
 sg13g2_decap_4 FILLER_36_430 ();
 sg13g2_fill_1 FILLER_36_434 ();
 sg13g2_fill_2 FILLER_36_473 ();
 sg13g2_fill_2 FILLER_36_484 ();
 sg13g2_fill_1 FILLER_36_510 ();
 sg13g2_decap_8 FILLER_36_525 ();
 sg13g2_decap_4 FILLER_36_532 ();
 sg13g2_fill_2 FILLER_36_572 ();
 sg13g2_fill_1 FILLER_36_574 ();
 sg13g2_fill_2 FILLER_36_579 ();
 sg13g2_fill_2 FILLER_36_616 ();
 sg13g2_fill_2 FILLER_36_622 ();
 sg13g2_fill_2 FILLER_36_638 ();
 sg13g2_fill_1 FILLER_36_645 ();
 sg13g2_fill_1 FILLER_36_685 ();
 sg13g2_fill_1 FILLER_36_703 ();
 sg13g2_fill_2 FILLER_36_797 ();
 sg13g2_decap_4 FILLER_36_809 ();
 sg13g2_fill_2 FILLER_36_813 ();
 sg13g2_decap_8 FILLER_36_851 ();
 sg13g2_fill_1 FILLER_36_894 ();
 sg13g2_fill_1 FILLER_36_942 ();
 sg13g2_fill_2 FILLER_36_973 ();
 sg13g2_fill_1 FILLER_36_975 ();
 sg13g2_decap_4 FILLER_36_981 ();
 sg13g2_decap_4 FILLER_36_1010 ();
 sg13g2_fill_2 FILLER_36_1014 ();
 sg13g2_fill_1 FILLER_36_1021 ();
 sg13g2_decap_8 FILLER_36_1048 ();
 sg13g2_fill_1 FILLER_36_1055 ();
 sg13g2_fill_1 FILLER_36_1066 ();
 sg13g2_fill_2 FILLER_36_1084 ();
 sg13g2_fill_1 FILLER_36_1091 ();
 sg13g2_fill_1 FILLER_36_1101 ();
 sg13g2_decap_4 FILLER_36_1158 ();
 sg13g2_decap_4 FILLER_36_1166 ();
 sg13g2_fill_1 FILLER_36_1196 ();
 sg13g2_fill_1 FILLER_36_1205 ();
 sg13g2_decap_8 FILLER_36_1210 ();
 sg13g2_decap_4 FILLER_36_1222 ();
 sg13g2_decap_8 FILLER_36_1262 ();
 sg13g2_decap_8 FILLER_36_1269 ();
 sg13g2_fill_1 FILLER_36_1276 ();
 sg13g2_fill_1 FILLER_36_1313 ();
 sg13g2_fill_2 FILLER_36_1326 ();
 sg13g2_decap_8 FILLER_36_1343 ();
 sg13g2_fill_2 FILLER_36_1350 ();
 sg13g2_fill_2 FILLER_36_1378 ();
 sg13g2_fill_1 FILLER_36_1380 ();
 sg13g2_fill_2 FILLER_36_1407 ();
 sg13g2_fill_1 FILLER_36_1409 ();
 sg13g2_fill_1 FILLER_36_1414 ();
 sg13g2_fill_1 FILLER_36_1432 ();
 sg13g2_fill_2 FILLER_36_1438 ();
 sg13g2_fill_1 FILLER_36_1440 ();
 sg13g2_fill_1 FILLER_36_1472 ();
 sg13g2_fill_1 FILLER_36_1484 ();
 sg13g2_fill_2 FILLER_36_1497 ();
 sg13g2_fill_2 FILLER_36_1554 ();
 sg13g2_fill_2 FILLER_36_1630 ();
 sg13g2_fill_1 FILLER_36_1632 ();
 sg13g2_fill_1 FILLER_36_1667 ();
 sg13g2_fill_1 FILLER_36_1687 ();
 sg13g2_fill_2 FILLER_36_1728 ();
 sg13g2_fill_2 FILLER_36_1743 ();
 sg13g2_fill_1 FILLER_36_1771 ();
 sg13g2_fill_2 FILLER_36_1784 ();
 sg13g2_decap_8 FILLER_36_1794 ();
 sg13g2_decap_4 FILLER_36_1801 ();
 sg13g2_fill_1 FILLER_36_1805 ();
 sg13g2_fill_1 FILLER_36_1811 ();
 sg13g2_fill_1 FILLER_36_1816 ();
 sg13g2_decap_4 FILLER_36_1840 ();
 sg13g2_fill_2 FILLER_36_1844 ();
 sg13g2_decap_4 FILLER_36_1851 ();
 sg13g2_fill_1 FILLER_36_1855 ();
 sg13g2_fill_2 FILLER_36_1910 ();
 sg13g2_fill_2 FILLER_36_1917 ();
 sg13g2_fill_1 FILLER_36_1919 ();
 sg13g2_fill_1 FILLER_36_1925 ();
 sg13g2_fill_2 FILLER_36_1954 ();
 sg13g2_fill_1 FILLER_36_1974 ();
 sg13g2_fill_1 FILLER_36_1990 ();
 sg13g2_fill_1 FILLER_36_2006 ();
 sg13g2_fill_1 FILLER_36_2021 ();
 sg13g2_fill_2 FILLER_36_2034 ();
 sg13g2_fill_2 FILLER_36_2040 ();
 sg13g2_fill_1 FILLER_36_2042 ();
 sg13g2_fill_1 FILLER_36_2052 ();
 sg13g2_fill_1 FILLER_36_2057 ();
 sg13g2_fill_1 FILLER_36_2062 ();
 sg13g2_fill_1 FILLER_36_2068 ();
 sg13g2_fill_2 FILLER_36_2095 ();
 sg13g2_fill_1 FILLER_36_2097 ();
 sg13g2_fill_2 FILLER_36_2111 ();
 sg13g2_fill_1 FILLER_36_2139 ();
 sg13g2_fill_1 FILLER_36_2144 ();
 sg13g2_fill_2 FILLER_36_2198 ();
 sg13g2_fill_1 FILLER_36_2230 ();
 sg13g2_fill_2 FILLER_36_2243 ();
 sg13g2_fill_2 FILLER_36_2302 ();
 sg13g2_fill_1 FILLER_36_2384 ();
 sg13g2_fill_1 FILLER_36_2411 ();
 sg13g2_decap_4 FILLER_36_2444 ();
 sg13g2_fill_1 FILLER_36_2448 ();
 sg13g2_decap_8 FILLER_36_2499 ();
 sg13g2_decap_4 FILLER_36_2506 ();
 sg13g2_fill_1 FILLER_36_2510 ();
 sg13g2_fill_1 FILLER_36_2541 ();
 sg13g2_fill_1 FILLER_36_2614 ();
 sg13g2_decap_4 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_4 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_fill_1 FILLER_37_21 ();
 sg13g2_decap_4 FILLER_37_30 ();
 sg13g2_fill_2 FILLER_37_34 ();
 sg13g2_fill_2 FILLER_37_63 ();
 sg13g2_fill_1 FILLER_37_73 ();
 sg13g2_fill_2 FILLER_37_82 ();
 sg13g2_fill_2 FILLER_37_98 ();
 sg13g2_fill_1 FILLER_37_105 ();
 sg13g2_fill_1 FILLER_37_135 ();
 sg13g2_decap_4 FILLER_37_166 ();
 sg13g2_fill_2 FILLER_37_170 ();
 sg13g2_fill_2 FILLER_37_185 ();
 sg13g2_decap_8 FILLER_37_192 ();
 sg13g2_fill_1 FILLER_37_199 ();
 sg13g2_decap_8 FILLER_37_204 ();
 sg13g2_decap_8 FILLER_37_211 ();
 sg13g2_decap_8 FILLER_37_218 ();
 sg13g2_fill_2 FILLER_37_225 ();
 sg13g2_fill_2 FILLER_37_231 ();
 sg13g2_fill_1 FILLER_37_264 ();
 sg13g2_fill_1 FILLER_37_269 ();
 sg13g2_fill_1 FILLER_37_274 ();
 sg13g2_fill_1 FILLER_37_290 ();
 sg13g2_fill_2 FILLER_37_305 ();
 sg13g2_fill_1 FILLER_37_315 ();
 sg13g2_fill_1 FILLER_37_336 ();
 sg13g2_decap_8 FILLER_37_342 ();
 sg13g2_fill_2 FILLER_37_349 ();
 sg13g2_decap_4 FILLER_37_355 ();
 sg13g2_fill_2 FILLER_37_363 ();
 sg13g2_fill_1 FILLER_37_365 ();
 sg13g2_fill_1 FILLER_37_370 ();
 sg13g2_fill_1 FILLER_37_375 ();
 sg13g2_fill_2 FILLER_37_402 ();
 sg13g2_fill_2 FILLER_37_430 ();
 sg13g2_fill_2 FILLER_37_477 ();
 sg13g2_fill_1 FILLER_37_479 ();
 sg13g2_fill_1 FILLER_37_485 ();
 sg13g2_decap_4 FILLER_37_525 ();
 sg13g2_fill_1 FILLER_37_535 ();
 sg13g2_fill_1 FILLER_37_540 ();
 sg13g2_fill_1 FILLER_37_545 ();
 sg13g2_decap_4 FILLER_37_556 ();
 sg13g2_fill_1 FILLER_37_560 ();
 sg13g2_fill_2 FILLER_37_570 ();
 sg13g2_fill_1 FILLER_37_572 ();
 sg13g2_decap_4 FILLER_37_579 ();
 sg13g2_fill_1 FILLER_37_599 ();
 sg13g2_fill_1 FILLER_37_615 ();
 sg13g2_fill_1 FILLER_37_653 ();
 sg13g2_fill_1 FILLER_37_669 ();
 sg13g2_fill_1 FILLER_37_685 ();
 sg13g2_fill_1 FILLER_37_691 ();
 sg13g2_fill_2 FILLER_37_701 ();
 sg13g2_fill_2 FILLER_37_748 ();
 sg13g2_fill_2 FILLER_37_770 ();
 sg13g2_fill_2 FILLER_37_834 ();
 sg13g2_fill_1 FILLER_37_836 ();
 sg13g2_fill_2 FILLER_37_863 ();
 sg13g2_fill_1 FILLER_37_865 ();
 sg13g2_fill_2 FILLER_37_870 ();
 sg13g2_fill_1 FILLER_37_882 ();
 sg13g2_fill_1 FILLER_37_893 ();
 sg13g2_decap_8 FILLER_37_924 ();
 sg13g2_decap_4 FILLER_37_931 ();
 sg13g2_fill_1 FILLER_37_935 ();
 sg13g2_decap_8 FILLER_37_971 ();
 sg13g2_decap_4 FILLER_37_978 ();
 sg13g2_fill_1 FILLER_37_994 ();
 sg13g2_decap_4 FILLER_37_1020 ();
 sg13g2_fill_2 FILLER_37_1024 ();
 sg13g2_decap_4 FILLER_37_1034 ();
 sg13g2_fill_1 FILLER_37_1038 ();
 sg13g2_decap_8 FILLER_37_1044 ();
 sg13g2_decap_8 FILLER_37_1051 ();
 sg13g2_fill_1 FILLER_37_1058 ();
 sg13g2_decap_8 FILLER_37_1085 ();
 sg13g2_decap_8 FILLER_37_1170 ();
 sg13g2_fill_2 FILLER_37_1177 ();
 sg13g2_fill_1 FILLER_37_1179 ();
 sg13g2_decap_4 FILLER_37_1238 ();
 sg13g2_decap_8 FILLER_37_1246 ();
 sg13g2_decap_8 FILLER_37_1253 ();
 sg13g2_decap_4 FILLER_37_1260 ();
 sg13g2_fill_2 FILLER_37_1264 ();
 sg13g2_fill_2 FILLER_37_1295 ();
 sg13g2_fill_2 FILLER_37_1394 ();
 sg13g2_fill_2 FILLER_37_1406 ();
 sg13g2_decap_4 FILLER_37_1444 ();
 sg13g2_fill_1 FILLER_37_1448 ();
 sg13g2_fill_2 FILLER_37_1453 ();
 sg13g2_fill_1 FILLER_37_1479 ();
 sg13g2_fill_1 FILLER_37_1485 ();
 sg13g2_fill_2 FILLER_37_1509 ();
 sg13g2_fill_1 FILLER_37_1553 ();
 sg13g2_fill_2 FILLER_37_1571 ();
 sg13g2_fill_1 FILLER_37_1573 ();
 sg13g2_fill_2 FILLER_37_1583 ();
 sg13g2_fill_2 FILLER_37_1595 ();
 sg13g2_fill_2 FILLER_37_1601 ();
 sg13g2_fill_1 FILLER_37_1631 ();
 sg13g2_decap_8 FILLER_37_1645 ();
 sg13g2_decap_4 FILLER_37_1652 ();
 sg13g2_fill_2 FILLER_37_1656 ();
 sg13g2_decap_8 FILLER_37_1666 ();
 sg13g2_fill_2 FILLER_37_1683 ();
 sg13g2_decap_4 FILLER_37_1689 ();
 sg13g2_fill_2 FILLER_37_1693 ();
 sg13g2_decap_8 FILLER_37_1710 ();
 sg13g2_decap_8 FILLER_37_1717 ();
 sg13g2_fill_1 FILLER_37_1724 ();
 sg13g2_decap_8 FILLER_37_1729 ();
 sg13g2_decap_4 FILLER_37_1736 ();
 sg13g2_fill_2 FILLER_37_1745 ();
 sg13g2_fill_1 FILLER_37_1771 ();
 sg13g2_decap_4 FILLER_37_1798 ();
 sg13g2_fill_2 FILLER_37_1826 ();
 sg13g2_fill_2 FILLER_37_1833 ();
 sg13g2_fill_1 FILLER_37_1835 ();
 sg13g2_fill_1 FILLER_37_1841 ();
 sg13g2_fill_1 FILLER_37_1864 ();
 sg13g2_fill_1 FILLER_37_1923 ();
 sg13g2_fill_1 FILLER_37_1937 ();
 sg13g2_fill_1 FILLER_37_1942 ();
 sg13g2_decap_8 FILLER_37_1951 ();
 sg13g2_fill_2 FILLER_37_1958 ();
 sg13g2_fill_1 FILLER_37_1960 ();
 sg13g2_fill_1 FILLER_37_1966 ();
 sg13g2_fill_1 FILLER_37_1972 ();
 sg13g2_fill_2 FILLER_37_2011 ();
 sg13g2_fill_1 FILLER_37_2013 ();
 sg13g2_fill_1 FILLER_37_2019 ();
 sg13g2_fill_1 FILLER_37_2025 ();
 sg13g2_fill_1 FILLER_37_2030 ();
 sg13g2_decap_8 FILLER_37_2035 ();
 sg13g2_fill_2 FILLER_37_2042 ();
 sg13g2_fill_1 FILLER_37_2044 ();
 sg13g2_fill_1 FILLER_37_2052 ();
 sg13g2_fill_2 FILLER_37_2056 ();
 sg13g2_fill_2 FILLER_37_2077 ();
 sg13g2_fill_1 FILLER_37_2164 ();
 sg13g2_fill_1 FILLER_37_2185 ();
 sg13g2_fill_2 FILLER_37_2203 ();
 sg13g2_decap_8 FILLER_37_2231 ();
 sg13g2_decap_4 FILLER_37_2238 ();
 sg13g2_fill_2 FILLER_37_2242 ();
 sg13g2_decap_4 FILLER_37_2249 ();
 sg13g2_fill_2 FILLER_37_2253 ();
 sg13g2_decap_4 FILLER_37_2264 ();
 sg13g2_fill_1 FILLER_37_2268 ();
 sg13g2_fill_2 FILLER_37_2279 ();
 sg13g2_fill_1 FILLER_37_2281 ();
 sg13g2_decap_8 FILLER_37_2286 ();
 sg13g2_decap_8 FILLER_37_2293 ();
 sg13g2_decap_8 FILLER_37_2300 ();
 sg13g2_fill_1 FILLER_37_2307 ();
 sg13g2_fill_1 FILLER_37_2332 ();
 sg13g2_fill_2 FILLER_37_2383 ();
 sg13g2_fill_2 FILLER_37_2390 ();
 sg13g2_decap_4 FILLER_37_2396 ();
 sg13g2_decap_4 FILLER_37_2413 ();
 sg13g2_fill_1 FILLER_37_2417 ();
 sg13g2_decap_4 FILLER_37_2422 ();
 sg13g2_fill_2 FILLER_37_2432 ();
 sg13g2_fill_1 FILLER_37_2434 ();
 sg13g2_fill_2 FILLER_37_2441 ();
 sg13g2_fill_1 FILLER_37_2443 ();
 sg13g2_fill_2 FILLER_37_2448 ();
 sg13g2_fill_1 FILLER_37_2450 ();
 sg13g2_fill_2 FILLER_37_2477 ();
 sg13g2_fill_1 FILLER_37_2479 ();
 sg13g2_decap_8 FILLER_37_2492 ();
 sg13g2_decap_8 FILLER_37_2499 ();
 sg13g2_fill_1 FILLER_37_2523 ();
 sg13g2_fill_1 FILLER_37_2539 ();
 sg13g2_fill_1 FILLER_37_2572 ();
 sg13g2_fill_1 FILLER_37_2583 ();
 sg13g2_fill_2 FILLER_37_2604 ();
 sg13g2_fill_1 FILLER_37_2622 ();
 sg13g2_fill_1 FILLER_37_2669 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_fill_1 FILLER_38_22 ();
 sg13g2_fill_2 FILLER_38_60 ();
 sg13g2_fill_1 FILLER_38_62 ();
 sg13g2_fill_1 FILLER_38_104 ();
 sg13g2_fill_1 FILLER_38_113 ();
 sg13g2_decap_4 FILLER_38_174 ();
 sg13g2_fill_2 FILLER_38_178 ();
 sg13g2_decap_4 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_218 ();
 sg13g2_decap_8 FILLER_38_225 ();
 sg13g2_decap_4 FILLER_38_232 ();
 sg13g2_fill_2 FILLER_38_236 ();
 sg13g2_fill_2 FILLER_38_243 ();
 sg13g2_fill_1 FILLER_38_245 ();
 sg13g2_fill_2 FILLER_38_254 ();
 sg13g2_decap_4 FILLER_38_295 ();
 sg13g2_fill_1 FILLER_38_308 ();
 sg13g2_fill_2 FILLER_38_328 ();
 sg13g2_fill_1 FILLER_38_330 ();
 sg13g2_fill_1 FILLER_38_380 ();
 sg13g2_fill_1 FILLER_38_386 ();
 sg13g2_fill_2 FILLER_38_396 ();
 sg13g2_fill_1 FILLER_38_446 ();
 sg13g2_decap_8 FILLER_38_487 ();
 sg13g2_decap_8 FILLER_38_494 ();
 sg13g2_decap_8 FILLER_38_527 ();
 sg13g2_decap_4 FILLER_38_534 ();
 sg13g2_decap_4 FILLER_38_573 ();
 sg13g2_fill_1 FILLER_38_577 ();
 sg13g2_fill_2 FILLER_38_655 ();
 sg13g2_fill_1 FILLER_38_761 ();
 sg13g2_fill_2 FILLER_38_770 ();
 sg13g2_fill_2 FILLER_38_777 ();
 sg13g2_fill_2 FILLER_38_784 ();
 sg13g2_fill_1 FILLER_38_797 ();
 sg13g2_fill_1 FILLER_38_817 ();
 sg13g2_fill_1 FILLER_38_848 ();
 sg13g2_fill_2 FILLER_38_870 ();
 sg13g2_decap_4 FILLER_38_923 ();
 sg13g2_decap_4 FILLER_38_1001 ();
 sg13g2_fill_2 FILLER_38_1051 ();
 sg13g2_decap_8 FILLER_38_1092 ();
 sg13g2_decap_4 FILLER_38_1099 ();
 sg13g2_fill_1 FILLER_38_1103 ();
 sg13g2_decap_4 FILLER_38_1113 ();
 sg13g2_fill_1 FILLER_38_1117 ();
 sg13g2_fill_2 FILLER_38_1122 ();
 sg13g2_decap_8 FILLER_38_1129 ();
 sg13g2_decap_4 FILLER_38_1136 ();
 sg13g2_fill_2 FILLER_38_1145 ();
 sg13g2_fill_1 FILLER_38_1165 ();
 sg13g2_fill_1 FILLER_38_1195 ();
 sg13g2_fill_1 FILLER_38_1222 ();
 sg13g2_fill_1 FILLER_38_1228 ();
 sg13g2_fill_2 FILLER_38_1240 ();
 sg13g2_decap_8 FILLER_38_1253 ();
 sg13g2_decap_8 FILLER_38_1260 ();
 sg13g2_decap_8 FILLER_38_1267 ();
 sg13g2_fill_1 FILLER_38_1274 ();
 sg13g2_fill_2 FILLER_38_1335 ();
 sg13g2_fill_2 FILLER_38_1381 ();
 sg13g2_fill_1 FILLER_38_1383 ();
 sg13g2_decap_8 FILLER_38_1410 ();
 sg13g2_decap_8 FILLER_38_1417 ();
 sg13g2_decap_8 FILLER_38_1424 ();
 sg13g2_decap_8 FILLER_38_1431 ();
 sg13g2_decap_8 FILLER_38_1438 ();
 sg13g2_decap_4 FILLER_38_1445 ();
 sg13g2_fill_1 FILLER_38_1449 ();
 sg13g2_fill_1 FILLER_38_1499 ();
 sg13g2_fill_1 FILLER_38_1534 ();
 sg13g2_decap_4 FILLER_38_1578 ();
 sg13g2_fill_2 FILLER_38_1582 ();
 sg13g2_decap_4 FILLER_38_1644 ();
 sg13g2_fill_1 FILLER_38_1648 ();
 sg13g2_fill_1 FILLER_38_1656 ();
 sg13g2_decap_8 FILLER_38_1699 ();
 sg13g2_decap_4 FILLER_38_1709 ();
 sg13g2_fill_1 FILLER_38_1762 ();
 sg13g2_fill_2 FILLER_38_1778 ();
 sg13g2_fill_1 FILLER_38_1784 ();
 sg13g2_fill_2 FILLER_38_1789 ();
 sg13g2_fill_2 FILLER_38_1796 ();
 sg13g2_fill_1 FILLER_38_1803 ();
 sg13g2_fill_2 FILLER_38_1808 ();
 sg13g2_fill_1 FILLER_38_1819 ();
 sg13g2_fill_1 FILLER_38_1828 ();
 sg13g2_fill_1 FILLER_38_1833 ();
 sg13g2_decap_4 FILLER_38_1844 ();
 sg13g2_fill_1 FILLER_38_1848 ();
 sg13g2_fill_2 FILLER_38_1854 ();
 sg13g2_fill_1 FILLER_38_1856 ();
 sg13g2_fill_2 FILLER_38_1862 ();
 sg13g2_fill_1 FILLER_38_1916 ();
 sg13g2_decap_4 FILLER_38_1922 ();
 sg13g2_fill_1 FILLER_38_1926 ();
 sg13g2_fill_1 FILLER_38_1932 ();
 sg13g2_fill_2 FILLER_38_1947 ();
 sg13g2_fill_1 FILLER_38_1949 ();
 sg13g2_fill_1 FILLER_38_1999 ();
 sg13g2_fill_1 FILLER_38_2032 ();
 sg13g2_decap_8 FILLER_38_2036 ();
 sg13g2_decap_4 FILLER_38_2043 ();
 sg13g2_fill_1 FILLER_38_2047 ();
 sg13g2_fill_1 FILLER_38_2052 ();
 sg13g2_fill_2 FILLER_38_2063 ();
 sg13g2_fill_1 FILLER_38_2091 ();
 sg13g2_fill_2 FILLER_38_2100 ();
 sg13g2_fill_1 FILLER_38_2102 ();
 sg13g2_decap_8 FILLER_38_2119 ();
 sg13g2_fill_2 FILLER_38_2126 ();
 sg13g2_fill_1 FILLER_38_2128 ();
 sg13g2_decap_4 FILLER_38_2137 ();
 sg13g2_fill_2 FILLER_38_2164 ();
 sg13g2_fill_1 FILLER_38_2192 ();
 sg13g2_fill_1 FILLER_38_2259 ();
 sg13g2_fill_1 FILLER_38_2270 ();
 sg13g2_decap_8 FILLER_38_2291 ();
 sg13g2_decap_8 FILLER_38_2298 ();
 sg13g2_decap_4 FILLER_38_2305 ();
 sg13g2_fill_2 FILLER_38_2309 ();
 sg13g2_fill_1 FILLER_38_2337 ();
 sg13g2_fill_1 FILLER_38_2344 ();
 sg13g2_fill_1 FILLER_38_2349 ();
 sg13g2_decap_8 FILLER_38_2364 ();
 sg13g2_decap_8 FILLER_38_2371 ();
 sg13g2_fill_2 FILLER_38_2378 ();
 sg13g2_fill_1 FILLER_38_2380 ();
 sg13g2_decap_4 FILLER_38_2395 ();
 sg13g2_decap_8 FILLER_38_2429 ();
 sg13g2_decap_8 FILLER_38_2436 ();
 sg13g2_decap_8 FILLER_38_2443 ();
 sg13g2_fill_1 FILLER_38_2450 ();
 sg13g2_decap_4 FILLER_38_2455 ();
 sg13g2_fill_1 FILLER_38_2459 ();
 sg13g2_decap_8 FILLER_38_2464 ();
 sg13g2_fill_2 FILLER_38_2471 ();
 sg13g2_fill_1 FILLER_38_2473 ();
 sg13g2_decap_8 FILLER_38_2491 ();
 sg13g2_fill_1 FILLER_38_2498 ();
 sg13g2_fill_2 FILLER_38_2502 ();
 sg13g2_decap_4 FILLER_38_2509 ();
 sg13g2_fill_1 FILLER_38_2529 ();
 sg13g2_fill_2 FILLER_38_2535 ();
 sg13g2_fill_2 FILLER_38_2544 ();
 sg13g2_fill_2 FILLER_38_2634 ();
 sg13g2_fill_2 FILLER_38_2668 ();
 sg13g2_fill_2 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_62 ();
 sg13g2_fill_1 FILLER_39_103 ();
 sg13g2_fill_2 FILLER_39_124 ();
 sg13g2_fill_1 FILLER_39_126 ();
 sg13g2_fill_2 FILLER_39_131 ();
 sg13g2_decap_8 FILLER_39_138 ();
 sg13g2_decap_8 FILLER_39_145 ();
 sg13g2_fill_1 FILLER_39_152 ();
 sg13g2_decap_8 FILLER_39_157 ();
 sg13g2_decap_8 FILLER_39_164 ();
 sg13g2_fill_2 FILLER_39_240 ();
 sg13g2_fill_1 FILLER_39_242 ();
 sg13g2_decap_8 FILLER_39_248 ();
 sg13g2_decap_8 FILLER_39_255 ();
 sg13g2_decap_8 FILLER_39_262 ();
 sg13g2_fill_2 FILLER_39_284 ();
 sg13g2_fill_2 FILLER_39_296 ();
 sg13g2_fill_2 FILLER_39_303 ();
 sg13g2_fill_1 FILLER_39_305 ();
 sg13g2_fill_2 FILLER_39_313 ();
 sg13g2_decap_4 FILLER_39_322 ();
 sg13g2_fill_2 FILLER_39_326 ();
 sg13g2_fill_1 FILLER_39_402 ();
 sg13g2_fill_2 FILLER_39_456 ();
 sg13g2_fill_2 FILLER_39_462 ();
 sg13g2_fill_1 FILLER_39_464 ();
 sg13g2_decap_8 FILLER_39_469 ();
 sg13g2_fill_2 FILLER_39_476 ();
 sg13g2_decap_4 FILLER_39_482 ();
 sg13g2_fill_1 FILLER_39_486 ();
 sg13g2_fill_1 FILLER_39_500 ();
 sg13g2_fill_1 FILLER_39_514 ();
 sg13g2_decap_8 FILLER_39_520 ();
 sg13g2_decap_4 FILLER_39_527 ();
 sg13g2_fill_1 FILLER_39_531 ();
 sg13g2_fill_1 FILLER_39_536 ();
 sg13g2_fill_2 FILLER_39_547 ();
 sg13g2_fill_1 FILLER_39_616 ();
 sg13g2_fill_1 FILLER_39_622 ();
 sg13g2_fill_1 FILLER_39_627 ();
 sg13g2_fill_1 FILLER_39_633 ();
 sg13g2_fill_2 FILLER_39_639 ();
 sg13g2_fill_1 FILLER_39_682 ();
 sg13g2_fill_1 FILLER_39_689 ();
 sg13g2_fill_1 FILLER_39_721 ();
 sg13g2_fill_2 FILLER_39_740 ();
 sg13g2_fill_1 FILLER_39_755 ();
 sg13g2_fill_1 FILLER_39_782 ();
 sg13g2_fill_2 FILLER_39_804 ();
 sg13g2_fill_1 FILLER_39_806 ();
 sg13g2_fill_2 FILLER_39_812 ();
 sg13g2_fill_1 FILLER_39_814 ();
 sg13g2_fill_2 FILLER_39_825 ();
 sg13g2_fill_2 FILLER_39_837 ();
 sg13g2_decap_8 FILLER_39_904 ();
 sg13g2_decap_8 FILLER_39_911 ();
 sg13g2_decap_8 FILLER_39_918 ();
 sg13g2_decap_8 FILLER_39_925 ();
 sg13g2_fill_2 FILLER_39_932 ();
 sg13g2_fill_2 FILLER_39_943 ();
 sg13g2_fill_2 FILLER_39_1048 ();
 sg13g2_fill_1 FILLER_39_1055 ();
 sg13g2_fill_2 FILLER_39_1078 ();
 sg13g2_fill_1 FILLER_39_1080 ();
 sg13g2_decap_8 FILLER_39_1127 ();
 sg13g2_decap_8 FILLER_39_1134 ();
 sg13g2_fill_2 FILLER_39_1141 ();
 sg13g2_decap_8 FILLER_39_1147 ();
 sg13g2_decap_8 FILLER_39_1154 ();
 sg13g2_decap_8 FILLER_39_1161 ();
 sg13g2_fill_1 FILLER_39_1168 ();
 sg13g2_fill_1 FILLER_39_1174 ();
 sg13g2_fill_2 FILLER_39_1180 ();
 sg13g2_decap_4 FILLER_39_1186 ();
 sg13g2_fill_1 FILLER_39_1190 ();
 sg13g2_fill_1 FILLER_39_1195 ();
 sg13g2_fill_1 FILLER_39_1238 ();
 sg13g2_fill_1 FILLER_39_1247 ();
 sg13g2_decap_8 FILLER_39_1252 ();
 sg13g2_decap_8 FILLER_39_1259 ();
 sg13g2_decap_4 FILLER_39_1266 ();
 sg13g2_fill_1 FILLER_39_1270 ();
 sg13g2_decap_8 FILLER_39_1282 ();
 sg13g2_decap_8 FILLER_39_1289 ();
 sg13g2_fill_2 FILLER_39_1296 ();
 sg13g2_fill_2 FILLER_39_1316 ();
 sg13g2_fill_2 FILLER_39_1331 ();
 sg13g2_decap_4 FILLER_39_1421 ();
 sg13g2_decap_4 FILLER_39_1429 ();
 sg13g2_fill_1 FILLER_39_1433 ();
 sg13g2_decap_4 FILLER_39_1439 ();
 sg13g2_fill_1 FILLER_39_1443 ();
 sg13g2_fill_2 FILLER_39_1450 ();
 sg13g2_fill_1 FILLER_39_1452 ();
 sg13g2_fill_2 FILLER_39_1482 ();
 sg13g2_fill_2 FILLER_39_1497 ();
 sg13g2_fill_1 FILLER_39_1520 ();
 sg13g2_fill_2 FILLER_39_1526 ();
 sg13g2_fill_2 FILLER_39_1572 ();
 sg13g2_decap_4 FILLER_39_1582 ();
 sg13g2_fill_1 FILLER_39_1586 ();
 sg13g2_fill_2 FILLER_39_1597 ();
 sg13g2_fill_1 FILLER_39_1634 ();
 sg13g2_fill_2 FILLER_39_1670 ();
 sg13g2_fill_1 FILLER_39_1672 ();
 sg13g2_fill_1 FILLER_39_1677 ();
 sg13g2_decap_4 FILLER_39_1704 ();
 sg13g2_fill_1 FILLER_39_1734 ();
 sg13g2_fill_1 FILLER_39_1754 ();
 sg13g2_fill_2 FILLER_39_1780 ();
 sg13g2_fill_1 FILLER_39_1782 ();
 sg13g2_decap_4 FILLER_39_1787 ();
 sg13g2_fill_1 FILLER_39_1795 ();
 sg13g2_decap_8 FILLER_39_1808 ();
 sg13g2_decap_4 FILLER_39_1815 ();
 sg13g2_fill_1 FILLER_39_1819 ();
 sg13g2_fill_2 FILLER_39_1884 ();
 sg13g2_decap_8 FILLER_39_1914 ();
 sg13g2_decap_8 FILLER_39_1921 ();
 sg13g2_fill_2 FILLER_39_1937 ();
 sg13g2_fill_1 FILLER_39_1944 ();
 sg13g2_fill_1 FILLER_39_1950 ();
 sg13g2_fill_2 FILLER_39_1955 ();
 sg13g2_fill_1 FILLER_39_2002 ();
 sg13g2_fill_2 FILLER_39_2006 ();
 sg13g2_fill_1 FILLER_39_2008 ();
 sg13g2_fill_1 FILLER_39_2019 ();
 sg13g2_decap_8 FILLER_39_2029 ();
 sg13g2_decap_8 FILLER_39_2036 ();
 sg13g2_decap_4 FILLER_39_2043 ();
 sg13g2_decap_4 FILLER_39_2089 ();
 sg13g2_fill_1 FILLER_39_2103 ();
 sg13g2_fill_2 FILLER_39_2130 ();
 sg13g2_decap_8 FILLER_39_2142 ();
 sg13g2_fill_1 FILLER_39_2207 ();
 sg13g2_fill_1 FILLER_39_2222 ();
 sg13g2_decap_8 FILLER_39_2227 ();
 sg13g2_fill_2 FILLER_39_2234 ();
 sg13g2_decap_4 FILLER_39_2279 ();
 sg13g2_fill_1 FILLER_39_2283 ();
 sg13g2_fill_2 FILLER_39_2314 ();
 sg13g2_decap_8 FILLER_39_2347 ();
 sg13g2_decap_8 FILLER_39_2354 ();
 sg13g2_decap_8 FILLER_39_2361 ();
 sg13g2_decap_8 FILLER_39_2368 ();
 sg13g2_fill_2 FILLER_39_2375 ();
 sg13g2_fill_1 FILLER_39_2403 ();
 sg13g2_fill_2 FILLER_39_2414 ();
 sg13g2_decap_8 FILLER_39_2467 ();
 sg13g2_decap_8 FILLER_39_2474 ();
 sg13g2_decap_4 FILLER_39_2481 ();
 sg13g2_fill_1 FILLER_39_2485 ();
 sg13g2_fill_1 FILLER_39_2490 ();
 sg13g2_fill_2 FILLER_39_2502 ();
 sg13g2_fill_1 FILLER_39_2510 ();
 sg13g2_fill_2 FILLER_39_2545 ();
 sg13g2_fill_1 FILLER_39_2551 ();
 sg13g2_fill_1 FILLER_39_2558 ();
 sg13g2_fill_2 FILLER_39_2565 ();
 sg13g2_fill_2 FILLER_39_2637 ();
 sg13g2_fill_1 FILLER_39_2665 ();
 sg13g2_fill_1 FILLER_39_2669 ();
 sg13g2_fill_2 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_85 ();
 sg13g2_fill_1 FILLER_40_90 ();
 sg13g2_decap_8 FILLER_40_131 ();
 sg13g2_decap_8 FILLER_40_138 ();
 sg13g2_fill_2 FILLER_40_145 ();
 sg13g2_fill_2 FILLER_40_174 ();
 sg13g2_fill_1 FILLER_40_206 ();
 sg13g2_fill_2 FILLER_40_211 ();
 sg13g2_decap_4 FILLER_40_239 ();
 sg13g2_fill_2 FILLER_40_243 ();
 sg13g2_decap_8 FILLER_40_249 ();
 sg13g2_decap_8 FILLER_40_256 ();
 sg13g2_fill_2 FILLER_40_263 ();
 sg13g2_fill_1 FILLER_40_265 ();
 sg13g2_fill_1 FILLER_40_274 ();
 sg13g2_fill_2 FILLER_40_290 ();
 sg13g2_decap_4 FILLER_40_318 ();
 sg13g2_decap_4 FILLER_40_325 ();
 sg13g2_decap_8 FILLER_40_334 ();
 sg13g2_fill_2 FILLER_40_341 ();
 sg13g2_fill_1 FILLER_40_343 ();
 sg13g2_fill_1 FILLER_40_374 ();
 sg13g2_fill_2 FILLER_40_378 ();
 sg13g2_fill_2 FILLER_40_384 ();
 sg13g2_fill_1 FILLER_40_398 ();
 sg13g2_fill_2 FILLER_40_404 ();
 sg13g2_fill_1 FILLER_40_427 ();
 sg13g2_decap_4 FILLER_40_443 ();
 sg13g2_fill_2 FILLER_40_465 ();
 sg13g2_fill_1 FILLER_40_467 ();
 sg13g2_decap_8 FILLER_40_478 ();
 sg13g2_fill_1 FILLER_40_489 ();
 sg13g2_fill_1 FILLER_40_495 ();
 sg13g2_decap_8 FILLER_40_506 ();
 sg13g2_decap_8 FILLER_40_513 ();
 sg13g2_decap_8 FILLER_40_520 ();
 sg13g2_fill_1 FILLER_40_536 ();
 sg13g2_decap_4 FILLER_40_551 ();
 sg13g2_fill_2 FILLER_40_559 ();
 sg13g2_fill_1 FILLER_40_561 ();
 sg13g2_fill_2 FILLER_40_566 ();
 sg13g2_fill_1 FILLER_40_568 ();
 sg13g2_fill_2 FILLER_40_573 ();
 sg13g2_fill_1 FILLER_40_575 ();
 sg13g2_fill_2 FILLER_40_626 ();
 sg13g2_decap_4 FILLER_40_636 ();
 sg13g2_fill_2 FILLER_40_640 ();
 sg13g2_fill_2 FILLER_40_646 ();
 sg13g2_fill_1 FILLER_40_648 ();
 sg13g2_decap_4 FILLER_40_666 ();
 sg13g2_fill_2 FILLER_40_670 ();
 sg13g2_fill_1 FILLER_40_677 ();
 sg13g2_decap_8 FILLER_40_683 ();
 sg13g2_decap_8 FILLER_40_690 ();
 sg13g2_decap_8 FILLER_40_697 ();
 sg13g2_fill_1 FILLER_40_724 ();
 sg13g2_fill_2 FILLER_40_747 ();
 sg13g2_fill_1 FILLER_40_778 ();
 sg13g2_fill_2 FILLER_40_784 ();
 sg13g2_fill_2 FILLER_40_791 ();
 sg13g2_fill_1 FILLER_40_824 ();
 sg13g2_fill_2 FILLER_40_896 ();
 sg13g2_fill_1 FILLER_40_898 ();
 sg13g2_decap_8 FILLER_40_909 ();
 sg13g2_decap_8 FILLER_40_920 ();
 sg13g2_decap_4 FILLER_40_927 ();
 sg13g2_decap_8 FILLER_40_966 ();
 sg13g2_fill_1 FILLER_40_973 ();
 sg13g2_decap_8 FILLER_40_991 ();
 sg13g2_decap_4 FILLER_40_1003 ();
 sg13g2_fill_1 FILLER_40_1007 ();
 sg13g2_fill_1 FILLER_40_1012 ();
 sg13g2_fill_2 FILLER_40_1096 ();
 sg13g2_fill_1 FILLER_40_1098 ();
 sg13g2_fill_2 FILLER_40_1104 ();
 sg13g2_fill_2 FILLER_40_1115 ();
 sg13g2_fill_2 FILLER_40_1169 ();
 sg13g2_decap_8 FILLER_40_1201 ();
 sg13g2_decap_4 FILLER_40_1239 ();
 sg13g2_decap_4 FILLER_40_1247 ();
 sg13g2_fill_2 FILLER_40_1251 ();
 sg13g2_decap_8 FILLER_40_1293 ();
 sg13g2_fill_1 FILLER_40_1300 ();
 sg13g2_fill_2 FILLER_40_1318 ();
 sg13g2_decap_8 FILLER_40_1352 ();
 sg13g2_decap_4 FILLER_40_1359 ();
 sg13g2_decap_4 FILLER_40_1377 ();
 sg13g2_fill_1 FILLER_40_1381 ();
 sg13g2_fill_2 FILLER_40_1387 ();
 sg13g2_fill_1 FILLER_40_1389 ();
 sg13g2_fill_2 FILLER_40_1459 ();
 sg13g2_fill_2 FILLER_40_1474 ();
 sg13g2_fill_1 FILLER_40_1489 ();
 sg13g2_fill_1 FILLER_40_1536 ();
 sg13g2_fill_1 FILLER_40_1552 ();
 sg13g2_fill_2 FILLER_40_1564 ();
 sg13g2_fill_1 FILLER_40_1578 ();
 sg13g2_fill_1 FILLER_40_1588 ();
 sg13g2_fill_1 FILLER_40_1605 ();
 sg13g2_fill_1 FILLER_40_1614 ();
 sg13g2_fill_1 FILLER_40_1636 ();
 sg13g2_fill_1 FILLER_40_1645 ();
 sg13g2_fill_1 FILLER_40_1650 ();
 sg13g2_fill_2 FILLER_40_1656 ();
 sg13g2_fill_2 FILLER_40_1684 ();
 sg13g2_decap_4 FILLER_40_1712 ();
 sg13g2_decap_8 FILLER_40_1720 ();
 sg13g2_fill_2 FILLER_40_1727 ();
 sg13g2_fill_2 FILLER_40_1756 ();
 sg13g2_fill_1 FILLER_40_1767 ();
 sg13g2_decap_4 FILLER_40_1812 ();
 sg13g2_fill_1 FILLER_40_1821 ();
 sg13g2_fill_1 FILLER_40_1838 ();
 sg13g2_fill_2 FILLER_40_1857 ();
 sg13g2_fill_1 FILLER_40_1859 ();
 sg13g2_fill_2 FILLER_40_1872 ();
 sg13g2_decap_8 FILLER_40_1877 ();
 sg13g2_decap_8 FILLER_40_1892 ();
 sg13g2_fill_2 FILLER_40_1903 ();
 sg13g2_fill_1 FILLER_40_1905 ();
 sg13g2_fill_2 FILLER_40_1910 ();
 sg13g2_fill_1 FILLER_40_1912 ();
 sg13g2_fill_2 FILLER_40_1935 ();
 sg13g2_decap_4 FILLER_40_1948 ();
 sg13g2_fill_2 FILLER_40_1972 ();
 sg13g2_fill_2 FILLER_40_1984 ();
 sg13g2_fill_2 FILLER_40_2009 ();
 sg13g2_decap_4 FILLER_40_2020 ();
 sg13g2_fill_2 FILLER_40_2082 ();
 sg13g2_fill_1 FILLER_40_2103 ();
 sg13g2_decap_8 FILLER_40_2217 ();
 sg13g2_decap_8 FILLER_40_2224 ();
 sg13g2_decap_8 FILLER_40_2231 ();
 sg13g2_decap_4 FILLER_40_2238 ();
 sg13g2_fill_2 FILLER_40_2242 ();
 sg13g2_fill_2 FILLER_40_2280 ();
 sg13g2_decap_8 FILLER_40_2296 ();
 sg13g2_decap_8 FILLER_40_2303 ();
 sg13g2_decap_4 FILLER_40_2310 ();
 sg13g2_fill_2 FILLER_40_2314 ();
 sg13g2_fill_1 FILLER_40_2320 ();
 sg13g2_decap_8 FILLER_40_2325 ();
 sg13g2_decap_8 FILLER_40_2332 ();
 sg13g2_decap_8 FILLER_40_2339 ();
 sg13g2_decap_8 FILLER_40_2346 ();
 sg13g2_fill_2 FILLER_40_2363 ();
 sg13g2_fill_1 FILLER_40_2365 ();
 sg13g2_decap_4 FILLER_40_2412 ();
 sg13g2_fill_2 FILLER_40_2416 ();
 sg13g2_decap_4 FILLER_40_2424 ();
 sg13g2_fill_2 FILLER_40_2432 ();
 sg13g2_fill_1 FILLER_40_2522 ();
 sg13g2_fill_1 FILLER_40_2551 ();
 sg13g2_fill_2 FILLER_40_2581 ();
 sg13g2_decap_4 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_4 ();
 sg13g2_fill_1 FILLER_41_44 ();
 sg13g2_fill_1 FILLER_41_49 ();
 sg13g2_fill_1 FILLER_41_53 ();
 sg13g2_fill_2 FILLER_41_58 ();
 sg13g2_fill_1 FILLER_41_60 ();
 sg13g2_fill_1 FILLER_41_83 ();
 sg13g2_fill_2 FILLER_41_89 ();
 sg13g2_fill_2 FILLER_41_101 ();
 sg13g2_fill_1 FILLER_41_103 ();
 sg13g2_fill_2 FILLER_41_108 ();
 sg13g2_fill_2 FILLER_41_115 ();
 sg13g2_fill_1 FILLER_41_117 ();
 sg13g2_fill_2 FILLER_41_144 ();
 sg13g2_fill_1 FILLER_41_146 ();
 sg13g2_fill_2 FILLER_41_156 ();
 sg13g2_fill_1 FILLER_41_158 ();
 sg13g2_fill_2 FILLER_41_164 ();
 sg13g2_decap_8 FILLER_41_171 ();
 sg13g2_decap_8 FILLER_41_178 ();
 sg13g2_fill_1 FILLER_41_185 ();
 sg13g2_fill_1 FILLER_41_212 ();
 sg13g2_fill_2 FILLER_41_230 ();
 sg13g2_decap_8 FILLER_41_258 ();
 sg13g2_fill_2 FILLER_41_265 ();
 sg13g2_fill_1 FILLER_41_267 ();
 sg13g2_fill_1 FILLER_41_288 ();
 sg13g2_fill_2 FILLER_41_328 ();
 sg13g2_fill_2 FILLER_41_356 ();
 sg13g2_fill_1 FILLER_41_362 ();
 sg13g2_fill_2 FILLER_41_371 ();
 sg13g2_fill_2 FILLER_41_378 ();
 sg13g2_fill_2 FILLER_41_384 ();
 sg13g2_fill_1 FILLER_41_386 ();
 sg13g2_fill_1 FILLER_41_406 ();
 sg13g2_fill_2 FILLER_41_463 ();
 sg13g2_fill_1 FILLER_41_465 ();
 sg13g2_decap_4 FILLER_41_479 ();
 sg13g2_fill_2 FILLER_41_496 ();
 sg13g2_decap_4 FILLER_41_502 ();
 sg13g2_fill_1 FILLER_41_506 ();
 sg13g2_decap_8 FILLER_41_511 ();
 sg13g2_fill_1 FILLER_41_518 ();
 sg13g2_fill_1 FILLER_41_536 ();
 sg13g2_decap_8 FILLER_41_541 ();
 sg13g2_decap_8 FILLER_41_548 ();
 sg13g2_decap_8 FILLER_41_555 ();
 sg13g2_decap_4 FILLER_41_562 ();
 sg13g2_fill_2 FILLER_41_566 ();
 sg13g2_decap_4 FILLER_41_572 ();
 sg13g2_fill_2 FILLER_41_576 ();
 sg13g2_fill_1 FILLER_41_582 ();
 sg13g2_fill_2 FILLER_41_592 ();
 sg13g2_fill_2 FILLER_41_599 ();
 sg13g2_fill_2 FILLER_41_605 ();
 sg13g2_fill_1 FILLER_41_611 ();
 sg13g2_decap_4 FILLER_41_616 ();
 sg13g2_fill_2 FILLER_41_638 ();
 sg13g2_fill_1 FILLER_41_640 ();
 sg13g2_fill_2 FILLER_41_646 ();
 sg13g2_fill_2 FILLER_41_657 ();
 sg13g2_fill_2 FILLER_41_664 ();
 sg13g2_fill_1 FILLER_41_666 ();
 sg13g2_decap_8 FILLER_41_675 ();
 sg13g2_fill_2 FILLER_41_682 ();
 sg13g2_fill_1 FILLER_41_684 ();
 sg13g2_decap_8 FILLER_41_689 ();
 sg13g2_decap_8 FILLER_41_696 ();
 sg13g2_fill_1 FILLER_41_749 ();
 sg13g2_fill_1 FILLER_41_766 ();
 sg13g2_fill_2 FILLER_41_786 ();
 sg13g2_fill_2 FILLER_41_800 ();
 sg13g2_fill_2 FILLER_41_832 ();
 sg13g2_fill_2 FILLER_41_883 ();
 sg13g2_fill_1 FILLER_41_885 ();
 sg13g2_fill_1 FILLER_41_890 ();
 sg13g2_decap_4 FILLER_41_904 ();
 sg13g2_fill_1 FILLER_41_908 ();
 sg13g2_decap_8 FILLER_41_961 ();
 sg13g2_decap_8 FILLER_41_968 ();
 sg13g2_fill_2 FILLER_41_975 ();
 sg13g2_fill_2 FILLER_41_982 ();
 sg13g2_decap_4 FILLER_41_1001 ();
 sg13g2_decap_4 FILLER_41_1049 ();
 sg13g2_decap_8 FILLER_41_1057 ();
 sg13g2_decap_8 FILLER_41_1068 ();
 sg13g2_fill_2 FILLER_41_1075 ();
 sg13g2_fill_1 FILLER_41_1077 ();
 sg13g2_decap_8 FILLER_41_1082 ();
 sg13g2_decap_8 FILLER_41_1089 ();
 sg13g2_fill_1 FILLER_41_1096 ();
 sg13g2_fill_2 FILLER_41_1188 ();
 sg13g2_fill_1 FILLER_41_1190 ();
 sg13g2_fill_1 FILLER_41_1217 ();
 sg13g2_fill_2 FILLER_41_1244 ();
 sg13g2_fill_1 FILLER_41_1246 ();
 sg13g2_fill_2 FILLER_41_1263 ();
 sg13g2_fill_1 FILLER_41_1269 ();
 sg13g2_fill_1 FILLER_41_1280 ();
 sg13g2_fill_1 FILLER_41_1307 ();
 sg13g2_fill_1 FILLER_41_1313 ();
 sg13g2_fill_1 FILLER_41_1323 ();
 sg13g2_decap_8 FILLER_41_1344 ();
 sg13g2_decap_8 FILLER_41_1351 ();
 sg13g2_decap_8 FILLER_41_1358 ();
 sg13g2_decap_8 FILLER_41_1365 ();
 sg13g2_decap_8 FILLER_41_1372 ();
 sg13g2_fill_2 FILLER_41_1379 ();
 sg13g2_fill_2 FILLER_41_1399 ();
 sg13g2_decap_4 FILLER_41_1405 ();
 sg13g2_fill_2 FILLER_41_1409 ();
 sg13g2_decap_8 FILLER_41_1421 ();
 sg13g2_decap_4 FILLER_41_1428 ();
 sg13g2_fill_2 FILLER_41_1432 ();
 sg13g2_fill_2 FILLER_41_1444 ();
 sg13g2_fill_1 FILLER_41_1459 ();
 sg13g2_fill_2 FILLER_41_1512 ();
 sg13g2_fill_1 FILLER_41_1572 ();
 sg13g2_fill_1 FILLER_41_1578 ();
 sg13g2_fill_1 FILLER_41_1584 ();
 sg13g2_fill_1 FILLER_41_1610 ();
 sg13g2_fill_1 FILLER_41_1620 ();
 sg13g2_fill_1 FILLER_41_1632 ();
 sg13g2_decap_4 FILLER_41_1648 ();
 sg13g2_decap_4 FILLER_41_1662 ();
 sg13g2_decap_8 FILLER_41_1670 ();
 sg13g2_decap_8 FILLER_41_1677 ();
 sg13g2_decap_8 FILLER_41_1724 ();
 sg13g2_fill_2 FILLER_41_1731 ();
 sg13g2_fill_1 FILLER_41_1743 ();
 sg13g2_fill_1 FILLER_41_1770 ();
 sg13g2_fill_2 FILLER_41_1823 ();
 sg13g2_fill_2 FILLER_41_1844 ();
 sg13g2_fill_2 FILLER_41_1866 ();
 sg13g2_fill_1 FILLER_41_1868 ();
 sg13g2_fill_1 FILLER_41_1874 ();
 sg13g2_fill_2 FILLER_41_1879 ();
 sg13g2_fill_1 FILLER_41_1886 ();
 sg13g2_fill_1 FILLER_41_1892 ();
 sg13g2_fill_1 FILLER_41_1896 ();
 sg13g2_fill_1 FILLER_41_1902 ();
 sg13g2_fill_1 FILLER_41_1908 ();
 sg13g2_fill_1 FILLER_41_1915 ();
 sg13g2_fill_1 FILLER_41_1920 ();
 sg13g2_fill_2 FILLER_41_1932 ();
 sg13g2_fill_1 FILLER_41_1947 ();
 sg13g2_fill_2 FILLER_41_2018 ();
 sg13g2_decap_8 FILLER_41_2027 ();
 sg13g2_decap_8 FILLER_41_2038 ();
 sg13g2_fill_2 FILLER_41_2045 ();
 sg13g2_fill_1 FILLER_41_2047 ();
 sg13g2_fill_1 FILLER_41_2053 ();
 sg13g2_fill_1 FILLER_41_2059 ();
 sg13g2_fill_2 FILLER_41_2118 ();
 sg13g2_fill_1 FILLER_41_2193 ();
 sg13g2_decap_8 FILLER_41_2219 ();
 sg13g2_decap_8 FILLER_41_2226 ();
 sg13g2_fill_2 FILLER_41_2233 ();
 sg13g2_fill_2 FILLER_41_2270 ();
 sg13g2_fill_1 FILLER_41_2272 ();
 sg13g2_decap_4 FILLER_41_2282 ();
 sg13g2_fill_2 FILLER_41_2286 ();
 sg13g2_decap_4 FILLER_41_2301 ();
 sg13g2_decap_8 FILLER_41_2331 ();
 sg13g2_decap_8 FILLER_41_2338 ();
 sg13g2_fill_2 FILLER_41_2345 ();
 sg13g2_fill_1 FILLER_41_2351 ();
 sg13g2_decap_4 FILLER_41_2401 ();
 sg13g2_fill_2 FILLER_41_2415 ();
 sg13g2_fill_1 FILLER_41_2417 ();
 sg13g2_decap_4 FILLER_41_2428 ();
 sg13g2_fill_2 FILLER_41_2432 ();
 sg13g2_fill_2 FILLER_41_2470 ();
 sg13g2_fill_1 FILLER_41_2472 ();
 sg13g2_decap_4 FILLER_41_2503 ();
 sg13g2_fill_2 FILLER_41_2511 ();
 sg13g2_fill_1 FILLER_41_2513 ();
 sg13g2_fill_2 FILLER_41_2518 ();
 sg13g2_fill_1 FILLER_41_2592 ();
 sg13g2_fill_1 FILLER_41_2645 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_4 FILLER_42_29 ();
 sg13g2_fill_1 FILLER_42_43 ();
 sg13g2_fill_2 FILLER_42_48 ();
 sg13g2_fill_1 FILLER_42_58 ();
 sg13g2_decap_4 FILLER_42_97 ();
 sg13g2_fill_1 FILLER_42_101 ();
 sg13g2_decap_4 FILLER_42_106 ();
 sg13g2_fill_1 FILLER_42_115 ();
 sg13g2_fill_2 FILLER_42_125 ();
 sg13g2_fill_1 FILLER_42_136 ();
 sg13g2_fill_2 FILLER_42_173 ();
 sg13g2_fill_1 FILLER_42_175 ();
 sg13g2_fill_1 FILLER_42_179 ();
 sg13g2_fill_1 FILLER_42_192 ();
 sg13g2_fill_2 FILLER_42_206 ();
 sg13g2_fill_2 FILLER_42_239 ();
 sg13g2_fill_2 FILLER_42_248 ();
 sg13g2_decap_8 FILLER_42_257 ();
 sg13g2_decap_4 FILLER_42_264 ();
 sg13g2_fill_2 FILLER_42_277 ();
 sg13g2_fill_1 FILLER_42_279 ();
 sg13g2_decap_8 FILLER_42_292 ();
 sg13g2_fill_2 FILLER_42_299 ();
 sg13g2_fill_1 FILLER_42_301 ();
 sg13g2_fill_2 FILLER_42_316 ();
 sg13g2_fill_1 FILLER_42_318 ();
 sg13g2_decap_4 FILLER_42_324 ();
 sg13g2_fill_2 FILLER_42_336 ();
 sg13g2_decap_8 FILLER_42_345 ();
 sg13g2_fill_1 FILLER_42_352 ();
 sg13g2_fill_2 FILLER_42_381 ();
 sg13g2_fill_1 FILLER_42_383 ();
 sg13g2_fill_2 FILLER_42_401 ();
 sg13g2_fill_1 FILLER_42_421 ();
 sg13g2_fill_2 FILLER_42_427 ();
 sg13g2_decap_8 FILLER_42_449 ();
 sg13g2_fill_2 FILLER_42_460 ();
 sg13g2_fill_1 FILLER_42_462 ();
 sg13g2_fill_1 FILLER_42_541 ();
 sg13g2_decap_8 FILLER_42_551 ();
 sg13g2_fill_1 FILLER_42_558 ();
 sg13g2_fill_2 FILLER_42_568 ();
 sg13g2_decap_4 FILLER_42_579 ();
 sg13g2_fill_1 FILLER_42_583 ();
 sg13g2_decap_4 FILLER_42_589 ();
 sg13g2_fill_2 FILLER_42_593 ();
 sg13g2_decap_4 FILLER_42_599 ();
 sg13g2_fill_1 FILLER_42_607 ();
 sg13g2_fill_1 FILLER_42_612 ();
 sg13g2_fill_1 FILLER_42_639 ();
 sg13g2_fill_2 FILLER_42_644 ();
 sg13g2_fill_2 FILLER_42_656 ();
 sg13g2_decap_4 FILLER_42_662 ();
 sg13g2_fill_2 FILLER_42_670 ();
 sg13g2_decap_8 FILLER_42_676 ();
 sg13g2_fill_2 FILLER_42_683 ();
 sg13g2_fill_2 FILLER_42_695 ();
 sg13g2_fill_2 FILLER_42_707 ();
 sg13g2_fill_2 FILLER_42_753 ();
 sg13g2_decap_4 FILLER_42_769 ();
 sg13g2_fill_1 FILLER_42_773 ();
 sg13g2_fill_1 FILLER_42_779 ();
 sg13g2_fill_1 FILLER_42_795 ();
 sg13g2_fill_1 FILLER_42_808 ();
 sg13g2_fill_2 FILLER_42_838 ();
 sg13g2_fill_1 FILLER_42_873 ();
 sg13g2_decap_8 FILLER_42_915 ();
 sg13g2_decap_8 FILLER_42_922 ();
 sg13g2_decap_8 FILLER_42_929 ();
 sg13g2_decap_4 FILLER_42_936 ();
 sg13g2_fill_2 FILLER_42_940 ();
 sg13g2_decap_8 FILLER_42_950 ();
 sg13g2_fill_2 FILLER_42_957 ();
 sg13g2_decap_8 FILLER_42_1006 ();
 sg13g2_decap_8 FILLER_42_1013 ();
 sg13g2_fill_2 FILLER_42_1020 ();
 sg13g2_fill_1 FILLER_42_1022 ();
 sg13g2_decap_8 FILLER_42_1031 ();
 sg13g2_decap_8 FILLER_42_1038 ();
 sg13g2_decap_8 FILLER_42_1045 ();
 sg13g2_decap_8 FILLER_42_1052 ();
 sg13g2_fill_1 FILLER_42_1063 ();
 sg13g2_fill_1 FILLER_42_1077 ();
 sg13g2_fill_2 FILLER_42_1082 ();
 sg13g2_fill_1 FILLER_42_1084 ();
 sg13g2_fill_1 FILLER_42_1111 ();
 sg13g2_fill_2 FILLER_42_1116 ();
 sg13g2_decap_4 FILLER_42_1149 ();
 sg13g2_fill_2 FILLER_42_1157 ();
 sg13g2_decap_8 FILLER_42_1185 ();
 sg13g2_decap_4 FILLER_42_1192 ();
 sg13g2_fill_2 FILLER_42_1196 ();
 sg13g2_decap_8 FILLER_42_1202 ();
 sg13g2_decap_4 FILLER_42_1219 ();
 sg13g2_fill_1 FILLER_42_1223 ();
 sg13g2_decap_8 FILLER_42_1228 ();
 sg13g2_decap_8 FILLER_42_1235 ();
 sg13g2_decap_4 FILLER_42_1242 ();
 sg13g2_fill_1 FILLER_42_1246 ();
 sg13g2_fill_1 FILLER_42_1258 ();
 sg13g2_decap_4 FILLER_42_1285 ();
 sg13g2_fill_2 FILLER_42_1299 ();
 sg13g2_fill_1 FILLER_42_1301 ();
 sg13g2_decap_4 FILLER_42_1342 ();
 sg13g2_decap_4 FILLER_42_1350 ();
 sg13g2_decap_8 FILLER_42_1357 ();
 sg13g2_decap_4 FILLER_42_1364 ();
 sg13g2_fill_1 FILLER_42_1368 ();
 sg13g2_fill_2 FILLER_42_1388 ();
 sg13g2_fill_1 FILLER_42_1390 ();
 sg13g2_decap_8 FILLER_42_1401 ();
 sg13g2_decap_8 FILLER_42_1408 ();
 sg13g2_decap_8 FILLER_42_1415 ();
 sg13g2_decap_4 FILLER_42_1422 ();
 sg13g2_fill_1 FILLER_42_1426 ();
 sg13g2_fill_2 FILLER_42_1492 ();
 sg13g2_fill_1 FILLER_42_1520 ();
 sg13g2_fill_2 FILLER_42_1541 ();
 sg13g2_fill_1 FILLER_42_1574 ();
 sg13g2_fill_2 FILLER_42_1613 ();
 sg13g2_fill_1 FILLER_42_1628 ();
 sg13g2_fill_2 FILLER_42_1636 ();
 sg13g2_decap_8 FILLER_42_1673 ();
 sg13g2_decap_8 FILLER_42_1680 ();
 sg13g2_decap_8 FILLER_42_1687 ();
 sg13g2_decap_8 FILLER_42_1694 ();
 sg13g2_fill_1 FILLER_42_1701 ();
 sg13g2_decap_4 FILLER_42_1749 ();
 sg13g2_decap_8 FILLER_42_1793 ();
 sg13g2_fill_1 FILLER_42_1807 ();
 sg13g2_decap_8 FILLER_42_1813 ();
 sg13g2_decap_8 FILLER_42_1820 ();
 sg13g2_fill_2 FILLER_42_1827 ();
 sg13g2_fill_2 FILLER_42_1833 ();
 sg13g2_decap_8 FILLER_42_1839 ();
 sg13g2_decap_8 FILLER_42_1846 ();
 sg13g2_decap_8 FILLER_42_1853 ();
 sg13g2_decap_8 FILLER_42_1860 ();
 sg13g2_decap_8 FILLER_42_1867 ();
 sg13g2_decap_4 FILLER_42_1874 ();
 sg13g2_fill_1 FILLER_42_1909 ();
 sg13g2_fill_1 FILLER_42_1938 ();
 sg13g2_fill_1 FILLER_42_1960 ();
 sg13g2_fill_1 FILLER_42_1965 ();
 sg13g2_fill_2 FILLER_42_2001 ();
 sg13g2_decap_4 FILLER_42_2022 ();
 sg13g2_fill_1 FILLER_42_2026 ();
 sg13g2_fill_1 FILLER_42_2057 ();
 sg13g2_decap_4 FILLER_42_2063 ();
 sg13g2_decap_8 FILLER_42_2093 ();
 sg13g2_fill_1 FILLER_42_2100 ();
 sg13g2_fill_2 FILLER_42_2166 ();
 sg13g2_fill_1 FILLER_42_2255 ();
 sg13g2_fill_1 FILLER_42_2266 ();
 sg13g2_decap_4 FILLER_42_2285 ();
 sg13g2_fill_2 FILLER_42_2289 ();
 sg13g2_decap_8 FILLER_42_2311 ();
 sg13g2_fill_2 FILLER_42_2318 ();
 sg13g2_fill_2 FILLER_42_2334 ();
 sg13g2_fill_2 FILLER_42_2341 ();
 sg13g2_fill_1 FILLER_42_2343 ();
 sg13g2_fill_2 FILLER_42_2348 ();
 sg13g2_fill_1 FILLER_42_2392 ();
 sg13g2_fill_2 FILLER_42_2445 ();
 sg13g2_fill_1 FILLER_42_2447 ();
 sg13g2_fill_1 FILLER_42_2474 ();
 sg13g2_fill_1 FILLER_42_2529 ();
 sg13g2_fill_1 FILLER_42_2537 ();
 sg13g2_fill_2 FILLER_42_2550 ();
 sg13g2_fill_1 FILLER_42_2552 ();
 sg13g2_fill_2 FILLER_42_2557 ();
 sg13g2_decap_8 FILLER_42_2573 ();
 sg13g2_decap_8 FILLER_42_2580 ();
 sg13g2_decap_8 FILLER_42_2587 ();
 sg13g2_decap_8 FILLER_42_2604 ();
 sg13g2_decap_4 FILLER_42_2611 ();
 sg13g2_fill_2 FILLER_42_2615 ();
 sg13g2_fill_2 FILLER_42_2630 ();
 sg13g2_fill_2 FILLER_42_2668 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_fill_1 FILLER_43_14 ();
 sg13g2_fill_1 FILLER_43_27 ();
 sg13g2_fill_1 FILLER_43_41 ();
 sg13g2_fill_1 FILLER_43_50 ();
 sg13g2_fill_1 FILLER_43_70 ();
 sg13g2_fill_2 FILLER_43_94 ();
 sg13g2_fill_2 FILLER_43_100 ();
 sg13g2_fill_1 FILLER_43_106 ();
 sg13g2_fill_2 FILLER_43_135 ();
 sg13g2_fill_1 FILLER_43_137 ();
 sg13g2_fill_2 FILLER_43_168 ();
 sg13g2_fill_2 FILLER_43_174 ();
 sg13g2_fill_1 FILLER_43_223 ();
 sg13g2_decap_8 FILLER_43_262 ();
 sg13g2_fill_1 FILLER_43_283 ();
 sg13g2_decap_8 FILLER_43_291 ();
 sg13g2_decap_4 FILLER_43_298 ();
 sg13g2_decap_4 FILLER_43_325 ();
 sg13g2_fill_1 FILLER_43_334 ();
 sg13g2_fill_1 FILLER_43_354 ();
 sg13g2_fill_1 FILLER_43_360 ();
 sg13g2_decap_8 FILLER_43_366 ();
 sg13g2_fill_2 FILLER_43_398 ();
 sg13g2_decap_4 FILLER_43_408 ();
 sg13g2_fill_2 FILLER_43_416 ();
 sg13g2_fill_1 FILLER_43_425 ();
 sg13g2_fill_2 FILLER_43_468 ();
 sg13g2_fill_1 FILLER_43_470 ();
 sg13g2_fill_1 FILLER_43_538 ();
 sg13g2_fill_1 FILLER_43_608 ();
 sg13g2_fill_1 FILLER_43_614 ();
 sg13g2_fill_1 FILLER_43_626 ();
 sg13g2_decap_8 FILLER_43_658 ();
 sg13g2_fill_1 FILLER_43_665 ();
 sg13g2_fill_2 FILLER_43_702 ();
 sg13g2_fill_2 FILLER_43_747 ();
 sg13g2_decap_4 FILLER_43_761 ();
 sg13g2_fill_1 FILLER_43_775 ();
 sg13g2_fill_1 FILLER_43_784 ();
 sg13g2_fill_2 FILLER_43_792 ();
 sg13g2_fill_2 FILLER_43_823 ();
 sg13g2_fill_1 FILLER_43_843 ();
 sg13g2_fill_1 FILLER_43_860 ();
 sg13g2_fill_1 FILLER_43_902 ();
 sg13g2_decap_8 FILLER_43_929 ();
 sg13g2_decap_8 FILLER_43_936 ();
 sg13g2_decap_8 FILLER_43_943 ();
 sg13g2_fill_1 FILLER_43_950 ();
 sg13g2_fill_1 FILLER_43_991 ();
 sg13g2_fill_1 FILLER_43_996 ();
 sg13g2_decap_4 FILLER_43_1023 ();
 sg13g2_fill_1 FILLER_43_1027 ();
 sg13g2_decap_4 FILLER_43_1033 ();
 sg13g2_fill_1 FILLER_43_1037 ();
 sg13g2_decap_4 FILLER_43_1098 ();
 sg13g2_decap_8 FILLER_43_1107 ();
 sg13g2_decap_8 FILLER_43_1114 ();
 sg13g2_fill_1 FILLER_43_1121 ();
 sg13g2_fill_2 FILLER_43_1139 ();
 sg13g2_fill_2 FILLER_43_1145 ();
 sg13g2_fill_1 FILLER_43_1152 ();
 sg13g2_decap_8 FILLER_43_1157 ();
 sg13g2_decap_8 FILLER_43_1164 ();
 sg13g2_fill_1 FILLER_43_1174 ();
 sg13g2_decap_4 FILLER_43_1180 ();
 sg13g2_fill_2 FILLER_43_1184 ();
 sg13g2_fill_2 FILLER_43_1196 ();
 sg13g2_fill_2 FILLER_43_1203 ();
 sg13g2_decap_8 FILLER_43_1210 ();
 sg13g2_decap_8 FILLER_43_1217 ();
 sg13g2_fill_2 FILLER_43_1248 ();
 sg13g2_fill_1 FILLER_43_1259 ();
 sg13g2_fill_1 FILLER_43_1270 ();
 sg13g2_decap_8 FILLER_43_1344 ();
 sg13g2_decap_8 FILLER_43_1351 ();
 sg13g2_decap_8 FILLER_43_1358 ();
 sg13g2_fill_1 FILLER_43_1365 ();
 sg13g2_fill_1 FILLER_43_1409 ();
 sg13g2_fill_2 FILLER_43_1420 ();
 sg13g2_fill_1 FILLER_43_1422 ();
 sg13g2_decap_4 FILLER_43_1432 ();
 sg13g2_fill_1 FILLER_43_1436 ();
 sg13g2_fill_1 FILLER_43_1455 ();
 sg13g2_fill_1 FILLER_43_1459 ();
 sg13g2_fill_2 FILLER_43_1485 ();
 sg13g2_fill_1 FILLER_43_1487 ();
 sg13g2_fill_1 FILLER_43_1497 ();
 sg13g2_fill_1 FILLER_43_1503 ();
 sg13g2_fill_1 FILLER_43_1509 ();
 sg13g2_fill_2 FILLER_43_1521 ();
 sg13g2_fill_1 FILLER_43_1554 ();
 sg13g2_fill_2 FILLER_43_1581 ();
 sg13g2_fill_2 FILLER_43_1601 ();
 sg13g2_decap_4 FILLER_43_1607 ();
 sg13g2_fill_2 FILLER_43_1615 ();
 sg13g2_fill_1 FILLER_43_1652 ();
 sg13g2_decap_8 FILLER_43_1657 ();
 sg13g2_decap_8 FILLER_43_1672 ();
 sg13g2_fill_2 FILLER_43_1679 ();
 sg13g2_fill_1 FILLER_43_1681 ();
 sg13g2_decap_8 FILLER_43_1687 ();
 sg13g2_decap_8 FILLER_43_1694 ();
 sg13g2_decap_8 FILLER_43_1701 ();
 sg13g2_fill_2 FILLER_43_1708 ();
 sg13g2_fill_1 FILLER_43_1710 ();
 sg13g2_decap_8 FILLER_43_1715 ();
 sg13g2_decap_4 FILLER_43_1722 ();
 sg13g2_fill_2 FILLER_43_1726 ();
 sg13g2_fill_2 FILLER_43_1762 ();
 sg13g2_fill_1 FILLER_43_1764 ();
 sg13g2_fill_1 FILLER_43_1791 ();
 sg13g2_decap_4 FILLER_43_1841 ();
 sg13g2_fill_2 FILLER_43_1845 ();
 sg13g2_decap_8 FILLER_43_1856 ();
 sg13g2_decap_4 FILLER_43_1863 ();
 sg13g2_fill_1 FILLER_43_1877 ();
 sg13g2_decap_8 FILLER_43_1885 ();
 sg13g2_decap_8 FILLER_43_1892 ();
 sg13g2_decap_4 FILLER_43_1899 ();
 sg13g2_decap_8 FILLER_43_1907 ();
 sg13g2_decap_4 FILLER_43_1914 ();
 sg13g2_fill_2 FILLER_43_1923 ();
 sg13g2_fill_1 FILLER_43_1925 ();
 sg13g2_decap_8 FILLER_43_1929 ();
 sg13g2_fill_2 FILLER_43_1936 ();
 sg13g2_fill_1 FILLER_43_1938 ();
 sg13g2_fill_1 FILLER_43_1949 ();
 sg13g2_fill_1 FILLER_43_1955 ();
 sg13g2_fill_1 FILLER_43_1982 ();
 sg13g2_decap_8 FILLER_43_1988 ();
 sg13g2_fill_2 FILLER_43_1995 ();
 sg13g2_decap_8 FILLER_43_2002 ();
 sg13g2_fill_2 FILLER_43_2071 ();
 sg13g2_fill_1 FILLER_43_2077 ();
 sg13g2_fill_2 FILLER_43_2113 ();
 sg13g2_fill_1 FILLER_43_2115 ();
 sg13g2_fill_2 FILLER_43_2120 ();
 sg13g2_fill_1 FILLER_43_2122 ();
 sg13g2_fill_2 FILLER_43_2188 ();
 sg13g2_fill_2 FILLER_43_2206 ();
 sg13g2_fill_2 FILLER_43_2234 ();
 sg13g2_fill_1 FILLER_43_2236 ();
 sg13g2_fill_2 FILLER_43_2241 ();
 sg13g2_fill_1 FILLER_43_2243 ();
 sg13g2_decap_4 FILLER_43_2293 ();
 sg13g2_fill_2 FILLER_43_2297 ();
 sg13g2_decap_4 FILLER_43_2343 ();
 sg13g2_fill_2 FILLER_43_2353 ();
 sg13g2_fill_1 FILLER_43_2355 ();
 sg13g2_fill_1 FILLER_43_2376 ();
 sg13g2_decap_8 FILLER_43_2407 ();
 sg13g2_fill_2 FILLER_43_2429 ();
 sg13g2_fill_2 FILLER_43_2436 ();
 sg13g2_fill_1 FILLER_43_2444 ();
 sg13g2_decap_8 FILLER_43_2463 ();
 sg13g2_fill_2 FILLER_43_2474 ();
 sg13g2_fill_1 FILLER_43_2476 ();
 sg13g2_fill_2 FILLER_43_2509 ();
 sg13g2_fill_2 FILLER_43_2525 ();
 sg13g2_fill_1 FILLER_43_2540 ();
 sg13g2_decap_4 FILLER_43_2547 ();
 sg13g2_fill_2 FILLER_43_2551 ();
 sg13g2_decap_8 FILLER_43_2562 ();
 sg13g2_decap_4 FILLER_43_2569 ();
 sg13g2_fill_2 FILLER_43_2573 ();
 sg13g2_decap_8 FILLER_43_2579 ();
 sg13g2_decap_8 FILLER_43_2586 ();
 sg13g2_decap_8 FILLER_43_2593 ();
 sg13g2_decap_4 FILLER_43_2600 ();
 sg13g2_fill_2 FILLER_43_2604 ();
 sg13g2_decap_8 FILLER_43_2653 ();
 sg13g2_decap_8 FILLER_43_2660 ();
 sg13g2_fill_2 FILLER_43_2667 ();
 sg13g2_fill_1 FILLER_43_2669 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_4 FILLER_44_7 ();
 sg13g2_fill_2 FILLER_44_11 ();
 sg13g2_fill_1 FILLER_44_36 ();
 sg13g2_fill_2 FILLER_44_67 ();
 sg13g2_fill_1 FILLER_44_79 ();
 sg13g2_fill_2 FILLER_44_90 ();
 sg13g2_fill_2 FILLER_44_102 ();
 sg13g2_fill_1 FILLER_44_133 ();
 sg13g2_fill_2 FILLER_44_143 ();
 sg13g2_fill_1 FILLER_44_179 ();
 sg13g2_fill_1 FILLER_44_201 ();
 sg13g2_fill_1 FILLER_44_238 ();
 sg13g2_fill_1 FILLER_44_244 ();
 sg13g2_fill_2 FILLER_44_255 ();
 sg13g2_fill_1 FILLER_44_257 ();
 sg13g2_decap_4 FILLER_44_276 ();
 sg13g2_fill_1 FILLER_44_290 ();
 sg13g2_decap_8 FILLER_44_294 ();
 sg13g2_fill_2 FILLER_44_307 ();
 sg13g2_fill_1 FILLER_44_309 ();
 sg13g2_fill_2 FILLER_44_330 ();
 sg13g2_fill_2 FILLER_44_344 ();
 sg13g2_fill_1 FILLER_44_346 ();
 sg13g2_fill_1 FILLER_44_355 ();
 sg13g2_fill_1 FILLER_44_364 ();
 sg13g2_fill_1 FILLER_44_369 ();
 sg13g2_fill_1 FILLER_44_403 ();
 sg13g2_fill_2 FILLER_44_447 ();
 sg13g2_fill_1 FILLER_44_449 ();
 sg13g2_decap_4 FILLER_44_474 ();
 sg13g2_fill_1 FILLER_44_493 ();
 sg13g2_decap_4 FILLER_44_519 ();
 sg13g2_fill_1 FILLER_44_559 ();
 sg13g2_fill_1 FILLER_44_564 ();
 sg13g2_fill_1 FILLER_44_596 ();
 sg13g2_fill_1 FILLER_44_628 ();
 sg13g2_fill_1 FILLER_44_668 ();
 sg13g2_fill_1 FILLER_44_695 ();
 sg13g2_fill_1 FILLER_44_709 ();
 sg13g2_fill_1 FILLER_44_720 ();
 sg13g2_fill_1 FILLER_44_729 ();
 sg13g2_decap_4 FILLER_44_753 ();
 sg13g2_fill_1 FILLER_44_769 ();
 sg13g2_fill_1 FILLER_44_812 ();
 sg13g2_fill_1 FILLER_44_855 ();
 sg13g2_fill_1 FILLER_44_877 ();
 sg13g2_fill_2 FILLER_44_883 ();
 sg13g2_fill_2 FILLER_44_922 ();
 sg13g2_fill_1 FILLER_44_924 ();
 sg13g2_decap_4 FILLER_44_951 ();
 sg13g2_fill_1 FILLER_44_962 ();
 sg13g2_decap_4 FILLER_44_971 ();
 sg13g2_fill_1 FILLER_44_975 ();
 sg13g2_decap_8 FILLER_44_990 ();
 sg13g2_fill_1 FILLER_44_1002 ();
 sg13g2_fill_2 FILLER_44_1038 ();
 sg13g2_fill_2 FILLER_44_1092 ();
 sg13g2_decap_8 FILLER_44_1120 ();
 sg13g2_decap_8 FILLER_44_1127 ();
 sg13g2_decap_8 FILLER_44_1134 ();
 sg13g2_decap_8 FILLER_44_1141 ();
 sg13g2_decap_8 FILLER_44_1148 ();
 sg13g2_fill_2 FILLER_44_1155 ();
 sg13g2_fill_1 FILLER_44_1157 ();
 sg13g2_decap_8 FILLER_44_1210 ();
 sg13g2_decap_8 FILLER_44_1217 ();
 sg13g2_fill_1 FILLER_44_1224 ();
 sg13g2_decap_8 FILLER_44_1229 ();
 sg13g2_decap_4 FILLER_44_1236 ();
 sg13g2_fill_2 FILLER_44_1240 ();
 sg13g2_fill_1 FILLER_44_1255 ();
 sg13g2_fill_1 FILLER_44_1266 ();
 sg13g2_fill_2 FILLER_44_1293 ();
 sg13g2_fill_1 FILLER_44_1310 ();
 sg13g2_fill_1 FILLER_44_1322 ();
 sg13g2_fill_1 FILLER_44_1328 ();
 sg13g2_fill_1 FILLER_44_1355 ();
 sg13g2_fill_1 FILLER_44_1361 ();
 sg13g2_fill_1 FILLER_44_1367 ();
 sg13g2_fill_1 FILLER_44_1374 ();
 sg13g2_fill_1 FILLER_44_1380 ();
 sg13g2_fill_2 FILLER_44_1401 ();
 sg13g2_fill_1 FILLER_44_1418 ();
 sg13g2_fill_1 FILLER_44_1429 ();
 sg13g2_fill_1 FILLER_44_1434 ();
 sg13g2_fill_2 FILLER_44_1439 ();
 sg13g2_fill_2 FILLER_44_1450 ();
 sg13g2_fill_1 FILLER_44_1465 ();
 sg13g2_decap_4 FILLER_44_1492 ();
 sg13g2_fill_2 FILLER_44_1496 ();
 sg13g2_fill_1 FILLER_44_1502 ();
 sg13g2_fill_2 FILLER_44_1545 ();
 sg13g2_fill_1 FILLER_44_1547 ();
 sg13g2_decap_8 FILLER_44_1552 ();
 sg13g2_fill_2 FILLER_44_1559 ();
 sg13g2_fill_1 FILLER_44_1561 ();
 sg13g2_fill_2 FILLER_44_1566 ();
 sg13g2_decap_8 FILLER_44_1581 ();
 sg13g2_fill_1 FILLER_44_1588 ();
 sg13g2_decap_4 FILLER_44_1598 ();
 sg13g2_fill_2 FILLER_44_1607 ();
 sg13g2_fill_1 FILLER_44_1609 ();
 sg13g2_fill_1 FILLER_44_1632 ();
 sg13g2_decap_8 FILLER_44_1711 ();
 sg13g2_decap_4 FILLER_44_1718 ();
 sg13g2_fill_1 FILLER_44_1722 ();
 sg13g2_fill_2 FILLER_44_1753 ();
 sg13g2_fill_1 FILLER_44_1755 ();
 sg13g2_decap_8 FILLER_44_1763 ();
 sg13g2_fill_1 FILLER_44_1770 ();
 sg13g2_decap_4 FILLER_44_1775 ();
 sg13g2_fill_2 FILLER_44_1783 ();
 sg13g2_fill_1 FILLER_44_1785 ();
 sg13g2_fill_1 FILLER_44_1799 ();
 sg13g2_decap_4 FILLER_44_1804 ();
 sg13g2_fill_1 FILLER_44_1808 ();
 sg13g2_fill_2 FILLER_44_1816 ();
 sg13g2_decap_8 FILLER_44_1900 ();
 sg13g2_decap_8 FILLER_44_1907 ();
 sg13g2_decap_8 FILLER_44_1914 ();
 sg13g2_decap_8 FILLER_44_1921 ();
 sg13g2_decap_8 FILLER_44_1928 ();
 sg13g2_decap_8 FILLER_44_1935 ();
 sg13g2_decap_8 FILLER_44_1942 ();
 sg13g2_decap_8 FILLER_44_1949 ();
 sg13g2_decap_8 FILLER_44_1956 ();
 sg13g2_decap_8 FILLER_44_1963 ();
 sg13g2_decap_8 FILLER_44_1970 ();
 sg13g2_decap_4 FILLER_44_1977 ();
 sg13g2_fill_1 FILLER_44_1981 ();
 sg13g2_decap_4 FILLER_44_1986 ();
 sg13g2_decap_8 FILLER_44_1995 ();
 sg13g2_fill_1 FILLER_44_2002 ();
 sg13g2_decap_8 FILLER_44_2007 ();
 sg13g2_decap_4 FILLER_44_2014 ();
 sg13g2_decap_8 FILLER_44_2029 ();
 sg13g2_fill_2 FILLER_44_2036 ();
 sg13g2_decap_4 FILLER_44_2042 ();
 sg13g2_fill_1 FILLER_44_2046 ();
 sg13g2_fill_2 FILLER_44_2051 ();
 sg13g2_fill_1 FILLER_44_2053 ();
 sg13g2_decap_4 FILLER_44_2129 ();
 sg13g2_fill_1 FILLER_44_2150 ();
 sg13g2_decap_4 FILLER_44_2187 ();
 sg13g2_fill_2 FILLER_44_2191 ();
 sg13g2_decap_8 FILLER_44_2196 ();
 sg13g2_decap_8 FILLER_44_2203 ();
 sg13g2_decap_8 FILLER_44_2210 ();
 sg13g2_decap_8 FILLER_44_2221 ();
 sg13g2_decap_8 FILLER_44_2228 ();
 sg13g2_decap_8 FILLER_44_2235 ();
 sg13g2_decap_4 FILLER_44_2242 ();
 sg13g2_fill_1 FILLER_44_2246 ();
 sg13g2_decap_8 FILLER_44_2281 ();
 sg13g2_decap_4 FILLER_44_2292 ();
 sg13g2_fill_2 FILLER_44_2296 ();
 sg13g2_decap_4 FILLER_44_2321 ();
 sg13g2_fill_1 FILLER_44_2370 ();
 sg13g2_fill_2 FILLER_44_2381 ();
 sg13g2_fill_1 FILLER_44_2383 ();
 sg13g2_fill_2 FILLER_44_2388 ();
 sg13g2_decap_8 FILLER_44_2403 ();
 sg13g2_decap_4 FILLER_44_2410 ();
 sg13g2_fill_2 FILLER_44_2414 ();
 sg13g2_fill_2 FILLER_44_2451 ();
 sg13g2_decap_4 FILLER_44_2459 ();
 sg13g2_fill_2 FILLER_44_2463 ();
 sg13g2_fill_1 FILLER_44_2482 ();
 sg13g2_fill_2 FILLER_44_2530 ();
 sg13g2_decap_8 FILLER_44_2537 ();
 sg13g2_decap_8 FILLER_44_2544 ();
 sg13g2_decap_4 FILLER_44_2551 ();
 sg13g2_decap_4 FILLER_44_2591 ();
 sg13g2_fill_2 FILLER_44_2595 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_4 FILLER_45_7 ();
 sg13g2_fill_1 FILLER_45_44 ();
 sg13g2_decap_8 FILLER_45_54 ();
 sg13g2_decap_4 FILLER_45_61 ();
 sg13g2_fill_1 FILLER_45_69 ();
 sg13g2_fill_1 FILLER_45_84 ();
 sg13g2_fill_1 FILLER_45_89 ();
 sg13g2_fill_1 FILLER_45_100 ();
 sg13g2_fill_1 FILLER_45_159 ();
 sg13g2_fill_2 FILLER_45_286 ();
 sg13g2_fill_2 FILLER_45_297 ();
 sg13g2_fill_2 FILLER_45_303 ();
 sg13g2_fill_2 FILLER_45_339 ();
 sg13g2_fill_2 FILLER_45_372 ();
 sg13g2_decap_4 FILLER_45_422 ();
 sg13g2_fill_1 FILLER_45_431 ();
 sg13g2_fill_1 FILLER_45_444 ();
 sg13g2_decap_4 FILLER_45_453 ();
 sg13g2_fill_1 FILLER_45_457 ();
 sg13g2_decap_4 FILLER_45_468 ();
 sg13g2_fill_1 FILLER_45_472 ();
 sg13g2_fill_1 FILLER_45_478 ();
 sg13g2_decap_8 FILLER_45_493 ();
 sg13g2_decap_8 FILLER_45_500 ();
 sg13g2_decap_8 FILLER_45_507 ();
 sg13g2_fill_2 FILLER_45_514 ();
 sg13g2_fill_1 FILLER_45_516 ();
 sg13g2_fill_2 FILLER_45_526 ();
 sg13g2_fill_1 FILLER_45_528 ();
 sg13g2_fill_2 FILLER_45_538 ();
 sg13g2_decap_4 FILLER_45_544 ();
 sg13g2_fill_1 FILLER_45_548 ();
 sg13g2_decap_4 FILLER_45_559 ();
 sg13g2_fill_1 FILLER_45_563 ();
 sg13g2_decap_4 FILLER_45_569 ();
 sg13g2_fill_2 FILLER_45_578 ();
 sg13g2_fill_2 FILLER_45_606 ();
 sg13g2_fill_2 FILLER_45_612 ();
 sg13g2_fill_1 FILLER_45_614 ();
 sg13g2_fill_2 FILLER_45_630 ();
 sg13g2_fill_1 FILLER_45_632 ();
 sg13g2_fill_1 FILLER_45_642 ();
 sg13g2_decap_8 FILLER_45_658 ();
 sg13g2_fill_1 FILLER_45_665 ();
 sg13g2_decap_4 FILLER_45_671 ();
 sg13g2_fill_1 FILLER_45_675 ();
 sg13g2_decap_8 FILLER_45_695 ();
 sg13g2_fill_2 FILLER_45_702 ();
 sg13g2_decap_4 FILLER_45_710 ();
 sg13g2_fill_1 FILLER_45_749 ();
 sg13g2_decap_8 FILLER_45_755 ();
 sg13g2_decap_8 FILLER_45_762 ();
 sg13g2_fill_2 FILLER_45_769 ();
 sg13g2_fill_1 FILLER_45_785 ();
 sg13g2_fill_2 FILLER_45_793 ();
 sg13g2_fill_1 FILLER_45_800 ();
 sg13g2_fill_2 FILLER_45_813 ();
 sg13g2_fill_1 FILLER_45_834 ();
 sg13g2_fill_1 FILLER_45_842 ();
 sg13g2_fill_1 FILLER_45_847 ();
 sg13g2_fill_2 FILLER_45_870 ();
 sg13g2_fill_1 FILLER_45_914 ();
 sg13g2_fill_1 FILLER_45_949 ();
 sg13g2_fill_2 FILLER_45_956 ();
 sg13g2_fill_2 FILLER_45_965 ();
 sg13g2_fill_1 FILLER_45_967 ();
 sg13g2_decap_4 FILLER_45_1001 ();
 sg13g2_fill_2 FILLER_45_1005 ();
 sg13g2_decap_4 FILLER_45_1046 ();
 sg13g2_fill_2 FILLER_45_1063 ();
 sg13g2_fill_2 FILLER_45_1070 ();
 sg13g2_decap_4 FILLER_45_1098 ();
 sg13g2_fill_1 FILLER_45_1110 ();
 sg13g2_fill_1 FILLER_45_1116 ();
 sg13g2_fill_1 FILLER_45_1147 ();
 sg13g2_decap_8 FILLER_45_1155 ();
 sg13g2_fill_2 FILLER_45_1162 ();
 sg13g2_fill_1 FILLER_45_1168 ();
 sg13g2_fill_1 FILLER_45_1195 ();
 sg13g2_decap_8 FILLER_45_1211 ();
 sg13g2_fill_1 FILLER_45_1218 ();
 sg13g2_decap_8 FILLER_45_1248 ();
 sg13g2_decap_8 FILLER_45_1255 ();
 sg13g2_fill_1 FILLER_45_1262 ();
 sg13g2_fill_1 FILLER_45_1344 ();
 sg13g2_fill_1 FILLER_45_1350 ();
 sg13g2_fill_1 FILLER_45_1360 ();
 sg13g2_fill_2 FILLER_45_1389 ();
 sg13g2_fill_2 FILLER_45_1413 ();
 sg13g2_decap_4 FILLER_45_1453 ();
 sg13g2_fill_1 FILLER_45_1457 ();
 sg13g2_fill_2 FILLER_45_1477 ();
 sg13g2_fill_1 FILLER_45_1479 ();
 sg13g2_fill_2 FILLER_45_1485 ();
 sg13g2_fill_1 FILLER_45_1487 ();
 sg13g2_fill_2 FILLER_45_1492 ();
 sg13g2_fill_1 FILLER_45_1502 ();
 sg13g2_fill_1 FILLER_45_1515 ();
 sg13g2_fill_2 FILLER_45_1521 ();
 sg13g2_decap_4 FILLER_45_1549 ();
 sg13g2_fill_2 FILLER_45_1553 ();
 sg13g2_decap_4 FILLER_45_1581 ();
 sg13g2_fill_2 FILLER_45_1637 ();
 sg13g2_fill_2 FILLER_45_1682 ();
 sg13g2_decap_4 FILLER_45_1720 ();
 sg13g2_fill_1 FILLER_45_1732 ();
 sg13g2_fill_1 FILLER_45_1743 ();
 sg13g2_decap_8 FILLER_45_1749 ();
 sg13g2_fill_1 FILLER_45_1770 ();
 sg13g2_fill_2 FILLER_45_1793 ();
 sg13g2_fill_1 FILLER_45_1795 ();
 sg13g2_fill_2 FILLER_45_1813 ();
 sg13g2_fill_1 FILLER_45_1815 ();
 sg13g2_fill_2 FILLER_45_1832 ();
 sg13g2_fill_1 FILLER_45_1834 ();
 sg13g2_decap_4 FILLER_45_1865 ();
 sg13g2_fill_2 FILLER_45_1869 ();
 sg13g2_decap_8 FILLER_45_1908 ();
 sg13g2_decap_8 FILLER_45_1915 ();
 sg13g2_decap_8 FILLER_45_1922 ();
 sg13g2_decap_8 FILLER_45_1929 ();
 sg13g2_decap_8 FILLER_45_1936 ();
 sg13g2_decap_8 FILLER_45_1943 ();
 sg13g2_decap_8 FILLER_45_1950 ();
 sg13g2_fill_2 FILLER_45_1957 ();
 sg13g2_fill_1 FILLER_45_1959 ();
 sg13g2_fill_2 FILLER_45_1970 ();
 sg13g2_fill_1 FILLER_45_1972 ();
 sg13g2_decap_8 FILLER_45_1977 ();
 sg13g2_decap_4 FILLER_45_1984 ();
 sg13g2_fill_1 FILLER_45_1988 ();
 sg13g2_decap_4 FILLER_45_1992 ();
 sg13g2_fill_1 FILLER_45_1996 ();
 sg13g2_decap_8 FILLER_45_2032 ();
 sg13g2_decap_8 FILLER_45_2039 ();
 sg13g2_decap_4 FILLER_45_2046 ();
 sg13g2_decap_8 FILLER_45_2056 ();
 sg13g2_fill_2 FILLER_45_2067 ();
 sg13g2_fill_2 FILLER_45_2072 ();
 sg13g2_fill_1 FILLER_45_2078 ();
 sg13g2_fill_2 FILLER_45_2083 ();
 sg13g2_fill_2 FILLER_45_2094 ();
 sg13g2_decap_8 FILLER_45_2147 ();
 sg13g2_decap_4 FILLER_45_2154 ();
 sg13g2_fill_1 FILLER_45_2158 ();
 sg13g2_decap_8 FILLER_45_2176 ();
 sg13g2_fill_2 FILLER_45_2183 ();
 sg13g2_decap_8 FILLER_45_2221 ();
 sg13g2_decap_8 FILLER_45_2228 ();
 sg13g2_decap_8 FILLER_45_2235 ();
 sg13g2_fill_2 FILLER_45_2242 ();
 sg13g2_fill_1 FILLER_45_2248 ();
 sg13g2_fill_2 FILLER_45_2253 ();
 sg13g2_fill_1 FILLER_45_2255 ();
 sg13g2_fill_2 FILLER_45_2260 ();
 sg13g2_decap_4 FILLER_45_2285 ();
 sg13g2_decap_8 FILLER_45_2293 ();
 sg13g2_decap_8 FILLER_45_2300 ();
 sg13g2_decap_4 FILLER_45_2307 ();
 sg13g2_fill_1 FILLER_45_2311 ();
 sg13g2_decap_8 FILLER_45_2316 ();
 sg13g2_fill_2 FILLER_45_2387 ();
 sg13g2_fill_1 FILLER_45_2420 ();
 sg13g2_fill_1 FILLER_45_2437 ();
 sg13g2_fill_2 FILLER_45_2484 ();
 sg13g2_decap_8 FILLER_45_2537 ();
 sg13g2_fill_1 FILLER_45_2544 ();
 sg13g2_decap_4 FILLER_45_2581 ();
 sg13g2_fill_2 FILLER_45_2585 ();
 sg13g2_fill_1 FILLER_45_2634 ();
 sg13g2_fill_2 FILLER_45_2668 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_fill_2 FILLER_46_7 ();
 sg13g2_decap_4 FILLER_46_13 ();
 sg13g2_fill_1 FILLER_46_17 ();
 sg13g2_fill_2 FILLER_46_22 ();
 sg13g2_decap_8 FILLER_46_33 ();
 sg13g2_decap_8 FILLER_46_45 ();
 sg13g2_decap_8 FILLER_46_52 ();
 sg13g2_decap_8 FILLER_46_59 ();
 sg13g2_fill_1 FILLER_46_66 ();
 sg13g2_fill_2 FILLER_46_72 ();
 sg13g2_decap_8 FILLER_46_78 ();
 sg13g2_decap_4 FILLER_46_85 ();
 sg13g2_fill_1 FILLER_46_145 ();
 sg13g2_fill_2 FILLER_46_194 ();
 sg13g2_fill_1 FILLER_46_201 ();
 sg13g2_fill_2 FILLER_46_243 ();
 sg13g2_fill_2 FILLER_46_344 ();
 sg13g2_fill_2 FILLER_46_376 ();
 sg13g2_decap_4 FILLER_46_417 ();
 sg13g2_fill_1 FILLER_46_421 ();
 sg13g2_fill_2 FILLER_46_439 ();
 sg13g2_fill_1 FILLER_46_467 ();
 sg13g2_fill_2 FILLER_46_473 ();
 sg13g2_fill_2 FILLER_46_480 ();
 sg13g2_decap_8 FILLER_46_506 ();
 sg13g2_fill_1 FILLER_46_513 ();
 sg13g2_decap_8 FILLER_46_518 ();
 sg13g2_fill_2 FILLER_46_525 ();
 sg13g2_fill_1 FILLER_46_536 ();
 sg13g2_decap_4 FILLER_46_541 ();
 sg13g2_decap_8 FILLER_46_549 ();
 sg13g2_fill_2 FILLER_46_556 ();
 sg13g2_fill_1 FILLER_46_558 ();
 sg13g2_decap_4 FILLER_46_568 ();
 sg13g2_decap_4 FILLER_46_581 ();
 sg13g2_fill_1 FILLER_46_585 ();
 sg13g2_fill_1 FILLER_46_604 ();
 sg13g2_decap_4 FILLER_46_609 ();
 sg13g2_decap_8 FILLER_46_631 ();
 sg13g2_decap_4 FILLER_46_638 ();
 sg13g2_decap_8 FILLER_46_659 ();
 sg13g2_decap_8 FILLER_46_666 ();
 sg13g2_fill_2 FILLER_46_673 ();
 sg13g2_fill_2 FILLER_46_679 ();
 sg13g2_fill_1 FILLER_46_681 ();
 sg13g2_decap_8 FILLER_46_696 ();
 sg13g2_fill_1 FILLER_46_718 ();
 sg13g2_fill_1 FILLER_46_723 ();
 sg13g2_fill_1 FILLER_46_734 ();
 sg13g2_fill_2 FILLER_46_763 ();
 sg13g2_fill_1 FILLER_46_765 ();
 sg13g2_fill_1 FILLER_46_770 ();
 sg13g2_fill_2 FILLER_46_796 ();
 sg13g2_fill_2 FILLER_46_806 ();
 sg13g2_fill_1 FILLER_46_843 ();
 sg13g2_fill_1 FILLER_46_886 ();
 sg13g2_fill_1 FILLER_46_897 ();
 sg13g2_fill_2 FILLER_46_924 ();
 sg13g2_fill_1 FILLER_46_967 ();
 sg13g2_decap_4 FILLER_46_973 ();
 sg13g2_fill_2 FILLER_46_981 ();
 sg13g2_fill_2 FILLER_46_1016 ();
 sg13g2_fill_1 FILLER_46_1023 ();
 sg13g2_fill_2 FILLER_46_1032 ();
 sg13g2_decap_4 FILLER_46_1065 ();
 sg13g2_fill_2 FILLER_46_1069 ();
 sg13g2_fill_1 FILLER_46_1080 ();
 sg13g2_decap_8 FILLER_46_1090 ();
 sg13g2_decap_8 FILLER_46_1097 ();
 sg13g2_decap_8 FILLER_46_1104 ();
 sg13g2_decap_8 FILLER_46_1111 ();
 sg13g2_fill_2 FILLER_46_1157 ();
 sg13g2_fill_2 FILLER_46_1164 ();
 sg13g2_fill_1 FILLER_46_1196 ();
 sg13g2_fill_1 FILLER_46_1223 ();
 sg13g2_decap_4 FILLER_46_1276 ();
 sg13g2_fill_2 FILLER_46_1280 ();
 sg13g2_decap_4 FILLER_46_1286 ();
 sg13g2_decap_4 FILLER_46_1303 ();
 sg13g2_fill_1 FILLER_46_1333 ();
 sg13g2_fill_2 FILLER_46_1339 ();
 sg13g2_decap_4 FILLER_46_1345 ();
 sg13g2_fill_2 FILLER_46_1349 ();
 sg13g2_decap_8 FILLER_46_1356 ();
 sg13g2_fill_1 FILLER_46_1376 ();
 sg13g2_fill_1 FILLER_46_1388 ();
 sg13g2_fill_1 FILLER_46_1396 ();
 sg13g2_fill_1 FILLER_46_1403 ();
 sg13g2_decap_8 FILLER_46_1423 ();
 sg13g2_decap_4 FILLER_46_1448 ();
 sg13g2_decap_4 FILLER_46_1467 ();
 sg13g2_fill_1 FILLER_46_1471 ();
 sg13g2_decap_4 FILLER_46_1476 ();
 sg13g2_fill_2 FILLER_46_1480 ();
 sg13g2_fill_1 FILLER_46_1490 ();
 sg13g2_fill_1 FILLER_46_1499 ();
 sg13g2_decap_4 FILLER_46_1517 ();
 sg13g2_fill_2 FILLER_46_1521 ();
 sg13g2_decap_8 FILLER_46_1542 ();
 sg13g2_decap_4 FILLER_46_1549 ();
 sg13g2_fill_1 FILLER_46_1553 ();
 sg13g2_fill_1 FILLER_46_1561 ();
 sg13g2_decap_8 FILLER_46_1566 ();
 sg13g2_fill_2 FILLER_46_1573 ();
 sg13g2_fill_1 FILLER_46_1575 ();
 sg13g2_fill_2 FILLER_46_1580 ();
 sg13g2_fill_2 FILLER_46_1620 ();
 sg13g2_fill_2 FILLER_46_1637 ();
 sg13g2_fill_1 FILLER_46_1650 ();
 sg13g2_fill_2 FILLER_46_1683 ();
 sg13g2_fill_2 FILLER_46_1692 ();
 sg13g2_decap_8 FILLER_46_1720 ();
 sg13g2_decap_4 FILLER_46_1727 ();
 sg13g2_fill_1 FILLER_46_1731 ();
 sg13g2_fill_2 FILLER_46_1742 ();
 sg13g2_fill_1 FILLER_46_1744 ();
 sg13g2_fill_1 FILLER_46_1755 ();
 sg13g2_decap_8 FILLER_46_1761 ();
 sg13g2_decap_4 FILLER_46_1768 ();
 sg13g2_decap_4 FILLER_46_1780 ();
 sg13g2_fill_1 FILLER_46_1784 ();
 sg13g2_fill_2 FILLER_46_1801 ();
 sg13g2_fill_1 FILLER_46_1803 ();
 sg13g2_fill_1 FILLER_46_1808 ();
 sg13g2_fill_1 FILLER_46_1825 ();
 sg13g2_fill_2 FILLER_46_1840 ();
 sg13g2_decap_4 FILLER_46_1846 ();
 sg13g2_fill_2 FILLER_46_1850 ();
 sg13g2_decap_4 FILLER_46_1878 ();
 sg13g2_fill_1 FILLER_46_1886 ();
 sg13g2_fill_2 FILLER_46_1891 ();
 sg13g2_fill_1 FILLER_46_1893 ();
 sg13g2_decap_8 FILLER_46_1898 ();
 sg13g2_fill_2 FILLER_46_1905 ();
 sg13g2_fill_1 FILLER_46_1907 ();
 sg13g2_decap_8 FILLER_46_1960 ();
 sg13g2_decap_8 FILLER_46_1997 ();
 sg13g2_decap_8 FILLER_46_2008 ();
 sg13g2_fill_2 FILLER_46_2015 ();
 sg13g2_decap_4 FILLER_46_2022 ();
 sg13g2_fill_1 FILLER_46_2035 ();
 sg13g2_decap_4 FILLER_46_2040 ();
 sg13g2_fill_1 FILLER_46_2044 ();
 sg13g2_decap_8 FILLER_46_2064 ();
 sg13g2_fill_2 FILLER_46_2071 ();
 sg13g2_decap_4 FILLER_46_2078 ();
 sg13g2_fill_1 FILLER_46_2082 ();
 sg13g2_decap_8 FILLER_46_2086 ();
 sg13g2_decap_8 FILLER_46_2093 ();
 sg13g2_fill_2 FILLER_46_2100 ();
 sg13g2_fill_1 FILLER_46_2102 ();
 sg13g2_decap_8 FILLER_46_2139 ();
 sg13g2_decap_4 FILLER_46_2146 ();
 sg13g2_decap_8 FILLER_46_2160 ();
 sg13g2_decap_8 FILLER_46_2177 ();
 sg13g2_decap_8 FILLER_46_2184 ();
 sg13g2_fill_1 FILLER_46_2191 ();
 sg13g2_fill_1 FILLER_46_2202 ();
 sg13g2_decap_8 FILLER_46_2228 ();
 sg13g2_decap_4 FILLER_46_2235 ();
 sg13g2_fill_2 FILLER_46_2239 ();
 sg13g2_fill_2 FILLER_46_2321 ();
 sg13g2_fill_1 FILLER_46_2323 ();
 sg13g2_fill_2 FILLER_46_2347 ();
 sg13g2_fill_1 FILLER_46_2349 ();
 sg13g2_fill_2 FILLER_46_2360 ();
 sg13g2_fill_2 FILLER_46_2402 ();
 sg13g2_fill_1 FILLER_46_2445 ();
 sg13g2_fill_1 FILLER_46_2456 ();
 sg13g2_fill_1 FILLER_46_2473 ();
 sg13g2_decap_4 FILLER_46_2480 ();
 sg13g2_fill_2 FILLER_46_2500 ();
 sg13g2_fill_1 FILLER_46_2502 ();
 sg13g2_fill_1 FILLER_46_2523 ();
 sg13g2_fill_1 FILLER_46_2528 ();
 sg13g2_fill_1 FILLER_46_2535 ();
 sg13g2_fill_2 FILLER_46_2546 ();
 sg13g2_fill_1 FILLER_46_2552 ();
 sg13g2_fill_1 FILLER_46_2557 ();
 sg13g2_fill_1 FILLER_46_2562 ();
 sg13g2_fill_2 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_38 ();
 sg13g2_decap_4 FILLER_47_45 ();
 sg13g2_fill_1 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_54 ();
 sg13g2_decap_4 FILLER_47_61 ();
 sg13g2_fill_2 FILLER_47_81 ();
 sg13g2_fill_1 FILLER_47_83 ();
 sg13g2_decap_8 FILLER_47_94 ();
 sg13g2_decap_8 FILLER_47_101 ();
 sg13g2_decap_8 FILLER_47_108 ();
 sg13g2_fill_2 FILLER_47_115 ();
 sg13g2_fill_2 FILLER_47_124 ();
 sg13g2_fill_1 FILLER_47_146 ();
 sg13g2_fill_1 FILLER_47_159 ();
 sg13g2_fill_2 FILLER_47_206 ();
 sg13g2_decap_8 FILLER_47_216 ();
 sg13g2_decap_8 FILLER_47_257 ();
 sg13g2_fill_1 FILLER_47_268 ();
 sg13g2_fill_2 FILLER_47_289 ();
 sg13g2_fill_1 FILLER_47_353 ();
 sg13g2_fill_2 FILLER_47_358 ();
 sg13g2_fill_2 FILLER_47_364 ();
 sg13g2_fill_1 FILLER_47_393 ();
 sg13g2_fill_2 FILLER_47_408 ();
 sg13g2_fill_2 FILLER_47_426 ();
 sg13g2_fill_1 FILLER_47_428 ();
 sg13g2_fill_1 FILLER_47_433 ();
 sg13g2_fill_1 FILLER_47_505 ();
 sg13g2_fill_1 FILLER_47_515 ();
 sg13g2_fill_2 FILLER_47_522 ();
 sg13g2_fill_1 FILLER_47_524 ();
 sg13g2_fill_1 FILLER_47_540 ();
 sg13g2_fill_1 FILLER_47_582 ();
 sg13g2_fill_1 FILLER_47_588 ();
 sg13g2_fill_2 FILLER_47_594 ();
 sg13g2_fill_1 FILLER_47_596 ();
 sg13g2_fill_2 FILLER_47_614 ();
 sg13g2_fill_1 FILLER_47_616 ();
 sg13g2_fill_2 FILLER_47_650 ();
 sg13g2_fill_2 FILLER_47_667 ();
 sg13g2_fill_1 FILLER_47_669 ();
 sg13g2_fill_1 FILLER_47_706 ();
 sg13g2_fill_1 FILLER_47_740 ();
 sg13g2_fill_2 FILLER_47_746 ();
 sg13g2_fill_1 FILLER_47_748 ();
 sg13g2_fill_2 FILLER_47_805 ();
 sg13g2_fill_2 FILLER_47_812 ();
 sg13g2_fill_1 FILLER_47_818 ();
 sg13g2_fill_2 FILLER_47_823 ();
 sg13g2_fill_2 FILLER_47_898 ();
 sg13g2_fill_2 FILLER_47_916 ();
 sg13g2_fill_1 FILLER_47_946 ();
 sg13g2_fill_1 FILLER_47_960 ();
 sg13g2_fill_1 FILLER_47_999 ();
 sg13g2_decap_8 FILLER_47_1030 ();
 sg13g2_fill_1 FILLER_47_1037 ();
 sg13g2_fill_2 FILLER_47_1041 ();
 sg13g2_fill_1 FILLER_47_1043 ();
 sg13g2_decap_8 FILLER_47_1071 ();
 sg13g2_fill_2 FILLER_47_1078 ();
 sg13g2_fill_1 FILLER_47_1080 ();
 sg13g2_fill_2 FILLER_47_1112 ();
 sg13g2_fill_1 FILLER_47_1114 ();
 sg13g2_fill_1 FILLER_47_1177 ();
 sg13g2_fill_1 FILLER_47_1199 ();
 sg13g2_fill_2 FILLER_47_1203 ();
 sg13g2_decap_4 FILLER_47_1271 ();
 sg13g2_fill_2 FILLER_47_1295 ();
 sg13g2_fill_1 FILLER_47_1297 ();
 sg13g2_fill_1 FILLER_47_1312 ();
 sg13g2_fill_2 FILLER_47_1323 ();
 sg13g2_fill_1 FILLER_47_1325 ();
 sg13g2_decap_8 FILLER_47_1333 ();
 sg13g2_fill_2 FILLER_47_1340 ();
 sg13g2_fill_2 FILLER_47_1347 ();
 sg13g2_fill_2 FILLER_47_1354 ();
 sg13g2_fill_1 FILLER_47_1356 ();
 sg13g2_fill_1 FILLER_47_1362 ();
 sg13g2_fill_2 FILLER_47_1368 ();
 sg13g2_fill_1 FILLER_47_1375 ();
 sg13g2_decap_8 FILLER_47_1386 ();
 sg13g2_fill_1 FILLER_47_1398 ();
 sg13g2_fill_2 FILLER_47_1424 ();
 sg13g2_decap_8 FILLER_47_1442 ();
 sg13g2_decap_4 FILLER_47_1449 ();
 sg13g2_fill_1 FILLER_47_1453 ();
 sg13g2_decap_8 FILLER_47_1485 ();
 sg13g2_decap_4 FILLER_47_1492 ();
 sg13g2_fill_1 FILLER_47_1496 ();
 sg13g2_decap_8 FILLER_47_1505 ();
 sg13g2_decap_4 FILLER_47_1512 ();
 sg13g2_fill_2 FILLER_47_1543 ();
 sg13g2_decap_8 FILLER_47_1563 ();
 sg13g2_fill_1 FILLER_47_1570 ();
 sg13g2_decap_8 FILLER_47_1576 ();
 sg13g2_decap_8 FILLER_47_1583 ();
 sg13g2_decap_8 FILLER_47_1597 ();
 sg13g2_decap_8 FILLER_47_1604 ();
 sg13g2_decap_4 FILLER_47_1611 ();
 sg13g2_decap_8 FILLER_47_1620 ();
 sg13g2_fill_2 FILLER_47_1627 ();
 sg13g2_fill_1 FILLER_47_1638 ();
 sg13g2_fill_1 FILLER_47_1642 ();
 sg13g2_fill_2 FILLER_47_1648 ();
 sg13g2_fill_1 FILLER_47_1709 ();
 sg13g2_decap_8 FILLER_47_1714 ();
 sg13g2_decap_8 FILLER_47_1721 ();
 sg13g2_fill_2 FILLER_47_1728 ();
 sg13g2_fill_1 FILLER_47_1730 ();
 sg13g2_fill_2 FILLER_47_1736 ();
 sg13g2_fill_1 FILLER_47_1738 ();
 sg13g2_fill_2 FILLER_47_1744 ();
 sg13g2_fill_1 FILLER_47_1746 ();
 sg13g2_fill_2 FILLER_47_1752 ();
 sg13g2_fill_1 FILLER_47_1754 ();
 sg13g2_decap_4 FILLER_47_1765 ();
 sg13g2_fill_2 FILLER_47_1769 ();
 sg13g2_fill_2 FILLER_47_1781 ();
 sg13g2_fill_2 FILLER_47_1787 ();
 sg13g2_fill_2 FILLER_47_1799 ();
 sg13g2_fill_1 FILLER_47_1801 ();
 sg13g2_decap_4 FILLER_47_1845 ();
 sg13g2_fill_2 FILLER_47_1849 ();
 sg13g2_fill_2 FILLER_47_1855 ();
 sg13g2_fill_1 FILLER_47_1857 ();
 sg13g2_fill_2 FILLER_47_1862 ();
 sg13g2_fill_1 FILLER_47_1864 ();
 sg13g2_decap_8 FILLER_47_1882 ();
 sg13g2_decap_8 FILLER_47_1889 ();
 sg13g2_decap_8 FILLER_47_1896 ();
 sg13g2_decap_4 FILLER_47_1903 ();
 sg13g2_fill_2 FILLER_47_1907 ();
 sg13g2_fill_2 FILLER_47_1920 ();
 sg13g2_fill_1 FILLER_47_1927 ();
 sg13g2_fill_2 FILLER_47_1932 ();
 sg13g2_fill_1 FILLER_47_1938 ();
 sg13g2_decap_8 FILLER_47_1969 ();
 sg13g2_decap_8 FILLER_47_1976 ();
 sg13g2_fill_2 FILLER_47_1983 ();
 sg13g2_fill_1 FILLER_47_1985 ();
 sg13g2_decap_4 FILLER_47_2017 ();
 sg13g2_fill_2 FILLER_47_2025 ();
 sg13g2_decap_8 FILLER_47_2031 ();
 sg13g2_decap_4 FILLER_47_2038 ();
 sg13g2_fill_2 FILLER_47_2042 ();
 sg13g2_fill_1 FILLER_47_2069 ();
 sg13g2_decap_8 FILLER_47_2074 ();
 sg13g2_decap_8 FILLER_47_2081 ();
 sg13g2_decap_8 FILLER_47_2088 ();
 sg13g2_decap_4 FILLER_47_2095 ();
 sg13g2_fill_2 FILLER_47_2099 ();
 sg13g2_fill_2 FILLER_47_2141 ();
 sg13g2_fill_1 FILLER_47_2147 ();
 sg13g2_fill_2 FILLER_47_2224 ();
 sg13g2_decap_4 FILLER_47_2266 ();
 sg13g2_fill_2 FILLER_47_2274 ();
 sg13g2_fill_2 FILLER_47_2285 ();
 sg13g2_fill_1 FILLER_47_2302 ();
 sg13g2_fill_2 FILLER_47_2318 ();
 sg13g2_fill_1 FILLER_47_2359 ();
 sg13g2_decap_4 FILLER_47_2366 ();
 sg13g2_fill_2 FILLER_47_2370 ();
 sg13g2_fill_2 FILLER_47_2376 ();
 sg13g2_fill_2 FILLER_47_2387 ();
 sg13g2_fill_2 FILLER_47_2399 ();
 sg13g2_decap_8 FILLER_47_2405 ();
 sg13g2_fill_1 FILLER_47_2438 ();
 sg13g2_fill_2 FILLER_47_2465 ();
 sg13g2_fill_1 FILLER_47_2493 ();
 sg13g2_fill_2 FILLER_47_2499 ();
 sg13g2_decap_8 FILLER_47_2506 ();
 sg13g2_fill_2 FILLER_47_2513 ();
 sg13g2_fill_1 FILLER_47_2515 ();
 sg13g2_fill_2 FILLER_47_2521 ();
 sg13g2_fill_1 FILLER_47_2523 ();
 sg13g2_fill_2 FILLER_47_2529 ();
 sg13g2_fill_1 FILLER_47_2567 ();
 sg13g2_decap_4 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_4 ();
 sg13g2_decap_4 FILLER_48_55 ();
 sg13g2_decap_4 FILLER_48_63 ();
 sg13g2_fill_1 FILLER_48_67 ();
 sg13g2_decap_4 FILLER_48_102 ();
 sg13g2_fill_2 FILLER_48_106 ();
 sg13g2_fill_2 FILLER_48_112 ();
 sg13g2_fill_2 FILLER_48_118 ();
 sg13g2_fill_1 FILLER_48_145 ();
 sg13g2_fill_1 FILLER_48_153 ();
 sg13g2_fill_1 FILLER_48_163 ();
 sg13g2_fill_2 FILLER_48_171 ();
 sg13g2_fill_2 FILLER_48_182 ();
 sg13g2_decap_8 FILLER_48_216 ();
 sg13g2_fill_1 FILLER_48_223 ();
 sg13g2_decap_8 FILLER_48_229 ();
 sg13g2_fill_2 FILLER_48_236 ();
 sg13g2_fill_1 FILLER_48_238 ();
 sg13g2_decap_8 FILLER_48_243 ();
 sg13g2_fill_2 FILLER_48_250 ();
 sg13g2_fill_2 FILLER_48_261 ();
 sg13g2_fill_2 FILLER_48_270 ();
 sg13g2_fill_1 FILLER_48_281 ();
 sg13g2_fill_1 FILLER_48_306 ();
 sg13g2_fill_2 FILLER_48_310 ();
 sg13g2_fill_2 FILLER_48_377 ();
 sg13g2_fill_2 FILLER_48_392 ();
 sg13g2_fill_1 FILLER_48_439 ();
 sg13g2_fill_2 FILLER_48_449 ();
 sg13g2_fill_1 FILLER_48_455 ();
 sg13g2_fill_1 FILLER_48_508 ();
 sg13g2_fill_2 FILLER_48_602 ();
 sg13g2_fill_1 FILLER_48_604 ();
 sg13g2_decap_8 FILLER_48_635 ();
 sg13g2_fill_2 FILLER_48_707 ();
 sg13g2_decap_8 FILLER_48_720 ();
 sg13g2_fill_2 FILLER_48_749 ();
 sg13g2_fill_1 FILLER_48_751 ();
 sg13g2_decap_4 FILLER_48_778 ();
 sg13g2_fill_1 FILLER_48_782 ();
 sg13g2_fill_2 FILLER_48_787 ();
 sg13g2_fill_2 FILLER_48_801 ();
 sg13g2_fill_2 FILLER_48_811 ();
 sg13g2_fill_1 FILLER_48_825 ();
 sg13g2_fill_1 FILLER_48_854 ();
 sg13g2_fill_2 FILLER_48_920 ();
 sg13g2_fill_1 FILLER_48_966 ();
 sg13g2_fill_2 FILLER_48_1001 ();
 sg13g2_decap_8 FILLER_48_1033 ();
 sg13g2_decap_8 FILLER_48_1040 ();
 sg13g2_fill_2 FILLER_48_1047 ();
 sg13g2_decap_4 FILLER_48_1056 ();
 sg13g2_fill_2 FILLER_48_1122 ();
 sg13g2_fill_1 FILLER_48_1124 ();
 sg13g2_fill_2 FILLER_48_1151 ();
 sg13g2_decap_8 FILLER_48_1293 ();
 sg13g2_decap_4 FILLER_48_1300 ();
 sg13g2_fill_1 FILLER_48_1304 ();
 sg13g2_fill_2 FILLER_48_1357 ();
 sg13g2_fill_1 FILLER_48_1359 ();
 sg13g2_fill_2 FILLER_48_1380 ();
 sg13g2_fill_2 FILLER_48_1403 ();
 sg13g2_decap_8 FILLER_48_1409 ();
 sg13g2_fill_1 FILLER_48_1416 ();
 sg13g2_fill_2 FILLER_48_1439 ();
 sg13g2_fill_2 FILLER_48_1451 ();
 sg13g2_decap_8 FILLER_48_1457 ();
 sg13g2_decap_8 FILLER_48_1468 ();
 sg13g2_decap_8 FILLER_48_1475 ();
 sg13g2_decap_4 FILLER_48_1482 ();
 sg13g2_decap_8 FILLER_48_1495 ();
 sg13g2_decap_8 FILLER_48_1502 ();
 sg13g2_fill_1 FILLER_48_1509 ();
 sg13g2_fill_1 FILLER_48_1547 ();
 sg13g2_fill_1 FILLER_48_1555 ();
 sg13g2_fill_1 FILLER_48_1582 ();
 sg13g2_fill_2 FILLER_48_1616 ();
 sg13g2_fill_1 FILLER_48_1618 ();
 sg13g2_fill_1 FILLER_48_1624 ();
 sg13g2_fill_1 FILLER_48_1636 ();
 sg13g2_decap_4 FILLER_48_1645 ();
 sg13g2_fill_2 FILLER_48_1649 ();
 sg13g2_fill_1 FILLER_48_1689 ();
 sg13g2_decap_8 FILLER_48_1703 ();
 sg13g2_decap_8 FILLER_48_1710 ();
 sg13g2_decap_8 FILLER_48_1717 ();
 sg13g2_decap_4 FILLER_48_1724 ();
 sg13g2_decap_4 FILLER_48_1737 ();
 sg13g2_decap_8 FILLER_48_1752 ();
 sg13g2_decap_8 FILLER_48_1759 ();
 sg13g2_decap_4 FILLER_48_1766 ();
 sg13g2_fill_2 FILLER_48_1770 ();
 sg13g2_fill_2 FILLER_48_1776 ();
 sg13g2_fill_1 FILLER_48_1778 ();
 sg13g2_decap_4 FILLER_48_1789 ();
 sg13g2_fill_1 FILLER_48_1793 ();
 sg13g2_fill_2 FILLER_48_1801 ();
 sg13g2_decap_8 FILLER_48_1838 ();
 sg13g2_decap_8 FILLER_48_1845 ();
 sg13g2_fill_1 FILLER_48_1852 ();
 sg13g2_decap_4 FILLER_48_1857 ();
 sg13g2_fill_2 FILLER_48_1861 ();
 sg13g2_fill_2 FILLER_48_1882 ();
 sg13g2_decap_8 FILLER_48_1895 ();
 sg13g2_fill_2 FILLER_48_1902 ();
 sg13g2_fill_1 FILLER_48_1904 ();
 sg13g2_fill_1 FILLER_48_1934 ();
 sg13g2_fill_2 FILLER_48_1945 ();
 sg13g2_fill_1 FILLER_48_1956 ();
 sg13g2_decap_8 FILLER_48_1962 ();
 sg13g2_decap_8 FILLER_48_1969 ();
 sg13g2_fill_2 FILLER_48_1976 ();
 sg13g2_fill_1 FILLER_48_1978 ();
 sg13g2_fill_1 FILLER_48_1984 ();
 sg13g2_fill_1 FILLER_48_2081 ();
 sg13g2_decap_8 FILLER_48_2089 ();
 sg13g2_fill_1 FILLER_48_2096 ();
 sg13g2_decap_8 FILLER_48_2101 ();
 sg13g2_fill_2 FILLER_48_2108 ();
 sg13g2_fill_1 FILLER_48_2110 ();
 sg13g2_fill_2 FILLER_48_2115 ();
 sg13g2_fill_1 FILLER_48_2117 ();
 sg13g2_fill_2 FILLER_48_2122 ();
 sg13g2_fill_1 FILLER_48_2124 ();
 sg13g2_fill_2 FILLER_48_2174 ();
 sg13g2_fill_1 FILLER_48_2197 ();
 sg13g2_decap_8 FILLER_48_2227 ();
 sg13g2_fill_2 FILLER_48_2234 ();
 sg13g2_fill_1 FILLER_48_2236 ();
 sg13g2_decap_4 FILLER_48_2246 ();
 sg13g2_fill_1 FILLER_48_2269 ();
 sg13g2_fill_1 FILLER_48_2290 ();
 sg13g2_fill_1 FILLER_48_2306 ();
 sg13g2_fill_1 FILLER_48_2320 ();
 sg13g2_fill_1 FILLER_48_2327 ();
 sg13g2_fill_1 FILLER_48_2374 ();
 sg13g2_decap_8 FILLER_48_2424 ();
 sg13g2_fill_2 FILLER_48_2431 ();
 sg13g2_fill_2 FILLER_48_2443 ();
 sg13g2_fill_1 FILLER_48_2445 ();
 sg13g2_decap_4 FILLER_48_2464 ();
 sg13g2_fill_2 FILLER_48_2512 ();
 sg13g2_fill_1 FILLER_48_2514 ();
 sg13g2_fill_1 FILLER_48_2523 ();
 sg13g2_decap_4 FILLER_48_2540 ();
 sg13g2_fill_2 FILLER_48_2544 ();
 sg13g2_decap_8 FILLER_48_2550 ();
 sg13g2_decap_8 FILLER_48_2557 ();
 sg13g2_decap_8 FILLER_48_2564 ();
 sg13g2_fill_2 FILLER_48_2668 ();
 sg13g2_fill_1 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_27 ();
 sg13g2_fill_2 FILLER_49_32 ();
 sg13g2_fill_1 FILLER_49_38 ();
 sg13g2_decap_8 FILLER_49_43 ();
 sg13g2_fill_2 FILLER_49_50 ();
 sg13g2_fill_1 FILLER_49_52 ();
 sg13g2_fill_2 FILLER_49_66 ();
 sg13g2_decap_8 FILLER_49_85 ();
 sg13g2_fill_2 FILLER_49_97 ();
 sg13g2_fill_2 FILLER_49_116 ();
 sg13g2_fill_1 FILLER_49_148 ();
 sg13g2_fill_2 FILLER_49_182 ();
 sg13g2_fill_2 FILLER_49_194 ();
 sg13g2_decap_8 FILLER_49_229 ();
 sg13g2_fill_2 FILLER_49_254 ();
 sg13g2_fill_1 FILLER_49_256 ();
 sg13g2_fill_1 FILLER_49_349 ();
 sg13g2_fill_2 FILLER_49_470 ();
 sg13g2_fill_2 FILLER_49_481 ();
 sg13g2_fill_1 FILLER_49_487 ();
 sg13g2_fill_2 FILLER_49_510 ();
 sg13g2_fill_2 FILLER_49_538 ();
 sg13g2_fill_1 FILLER_49_646 ();
 sg13g2_fill_1 FILLER_49_652 ();
 sg13g2_fill_1 FILLER_49_689 ();
 sg13g2_fill_2 FILLER_49_699 ();
 sg13g2_fill_1 FILLER_49_701 ();
 sg13g2_decap_8 FILLER_49_720 ();
 sg13g2_decap_4 FILLER_49_727 ();
 sg13g2_fill_2 FILLER_49_731 ();
 sg13g2_decap_8 FILLER_49_737 ();
 sg13g2_decap_8 FILLER_49_749 ();
 sg13g2_decap_8 FILLER_49_764 ();
 sg13g2_decap_4 FILLER_49_771 ();
 sg13g2_fill_2 FILLER_49_775 ();
 sg13g2_decap_4 FILLER_49_782 ();
 sg13g2_fill_2 FILLER_49_786 ();
 sg13g2_fill_1 FILLER_49_848 ();
 sg13g2_fill_1 FILLER_49_858 ();
 sg13g2_fill_1 FILLER_49_888 ();
 sg13g2_fill_2 FILLER_49_892 ();
 sg13g2_fill_1 FILLER_49_909 ();
 sg13g2_decap_4 FILLER_49_913 ();
 sg13g2_fill_1 FILLER_49_917 ();
 sg13g2_decap_4 FILLER_49_979 ();
 sg13g2_fill_1 FILLER_49_983 ();
 sg13g2_fill_2 FILLER_49_989 ();
 sg13g2_fill_1 FILLER_49_991 ();
 sg13g2_fill_2 FILLER_49_1065 ();
 sg13g2_fill_1 FILLER_49_1067 ();
 sg13g2_fill_2 FILLER_49_1072 ();
 sg13g2_fill_2 FILLER_49_1148 ();
 sg13g2_fill_2 FILLER_49_1165 ();
 sg13g2_fill_1 FILLER_49_1175 ();
 sg13g2_fill_1 FILLER_49_1180 ();
 sg13g2_fill_2 FILLER_49_1194 ();
 sg13g2_fill_2 FILLER_49_1208 ();
 sg13g2_fill_2 FILLER_49_1244 ();
 sg13g2_fill_2 FILLER_49_1263 ();
 sg13g2_fill_2 FILLER_49_1291 ();
 sg13g2_fill_1 FILLER_49_1293 ();
 sg13g2_fill_2 FILLER_49_1312 ();
 sg13g2_decap_4 FILLER_49_1319 ();
 sg13g2_fill_1 FILLER_49_1323 ();
 sg13g2_decap_8 FILLER_49_1341 ();
 sg13g2_decap_4 FILLER_49_1348 ();
 sg13g2_fill_1 FILLER_49_1352 ();
 sg13g2_fill_2 FILLER_49_1369 ();
 sg13g2_fill_1 FILLER_49_1371 ();
 sg13g2_fill_1 FILLER_49_1377 ();
 sg13g2_fill_1 FILLER_49_1385 ();
 sg13g2_fill_1 FILLER_49_1393 ();
 sg13g2_fill_2 FILLER_49_1400 ();
 sg13g2_fill_1 FILLER_49_1402 ();
 sg13g2_decap_8 FILLER_49_1409 ();
 sg13g2_decap_4 FILLER_49_1434 ();
 sg13g2_fill_2 FILLER_49_1438 ();
 sg13g2_decap_8 FILLER_49_1448 ();
 sg13g2_fill_1 FILLER_49_1455 ();
 sg13g2_fill_2 FILLER_49_1461 ();
 sg13g2_fill_1 FILLER_49_1463 ();
 sg13g2_decap_4 FILLER_49_1474 ();
 sg13g2_fill_1 FILLER_49_1493 ();
 sg13g2_fill_2 FILLER_49_1530 ();
 sg13g2_decap_4 FILLER_49_1601 ();
 sg13g2_fill_1 FILLER_49_1605 ();
 sg13g2_fill_2 FILLER_49_1632 ();
 sg13g2_fill_1 FILLER_49_1634 ();
 sg13g2_decap_8 FILLER_49_1640 ();
 sg13g2_fill_2 FILLER_49_1656 ();
 sg13g2_fill_2 FILLER_49_1690 ();
 sg13g2_decap_8 FILLER_49_1722 ();
 sg13g2_fill_1 FILLER_49_1729 ();
 sg13g2_fill_1 FILLER_49_1736 ();
 sg13g2_fill_1 FILLER_49_1740 ();
 sg13g2_fill_2 FILLER_49_1753 ();
 sg13g2_fill_1 FILLER_49_1755 ();
 sg13g2_decap_4 FILLER_49_1788 ();
 sg13g2_decap_8 FILLER_49_1796 ();
 sg13g2_fill_1 FILLER_49_1803 ();
 sg13g2_fill_1 FILLER_49_1809 ();
 sg13g2_decap_8 FILLER_49_1823 ();
 sg13g2_decap_8 FILLER_49_1830 ();
 sg13g2_decap_4 FILLER_49_1837 ();
 sg13g2_decap_8 FILLER_49_1846 ();
 sg13g2_decap_4 FILLER_49_1853 ();
 sg13g2_fill_2 FILLER_49_1857 ();
 sg13g2_fill_1 FILLER_49_1882 ();
 sg13g2_decap_4 FILLER_49_1930 ();
 sg13g2_fill_1 FILLER_49_1942 ();
 sg13g2_fill_2 FILLER_49_1955 ();
 sg13g2_decap_8 FILLER_49_1961 ();
 sg13g2_decap_8 FILLER_49_1968 ();
 sg13g2_decap_4 FILLER_49_1975 ();
 sg13g2_fill_2 FILLER_49_1979 ();
 sg13g2_fill_2 FILLER_49_1993 ();
 sg13g2_fill_2 FILLER_49_1999 ();
 sg13g2_fill_1 FILLER_49_2001 ();
 sg13g2_fill_2 FILLER_49_2037 ();
 sg13g2_fill_1 FILLER_49_2056 ();
 sg13g2_fill_1 FILLER_49_2062 ();
 sg13g2_decap_8 FILLER_49_2091 ();
 sg13g2_decap_8 FILLER_49_2098 ();
 sg13g2_decap_8 FILLER_49_2105 ();
 sg13g2_fill_2 FILLER_49_2152 ();
 sg13g2_fill_1 FILLER_49_2154 ();
 sg13g2_decap_8 FILLER_49_2159 ();
 sg13g2_decap_8 FILLER_49_2166 ();
 sg13g2_decap_8 FILLER_49_2173 ();
 sg13g2_fill_2 FILLER_49_2180 ();
 sg13g2_decap_8 FILLER_49_2196 ();
 sg13g2_fill_2 FILLER_49_2203 ();
 sg13g2_decap_8 FILLER_49_2209 ();
 sg13g2_fill_1 FILLER_49_2216 ();
 sg13g2_decap_4 FILLER_49_2222 ();
 sg13g2_decap_4 FILLER_49_2268 ();
 sg13g2_decap_4 FILLER_49_2302 ();
 sg13g2_fill_1 FILLER_49_2306 ();
 sg13g2_fill_2 FILLER_49_2350 ();
 sg13g2_fill_1 FILLER_49_2357 ();
 sg13g2_decap_4 FILLER_49_2368 ();
 sg13g2_fill_1 FILLER_49_2382 ();
 sg13g2_fill_1 FILLER_49_2409 ();
 sg13g2_fill_2 FILLER_49_2414 ();
 sg13g2_fill_2 FILLER_49_2421 ();
 sg13g2_fill_2 FILLER_49_2427 ();
 sg13g2_fill_1 FILLER_49_2429 ();
 sg13g2_decap_8 FILLER_49_2450 ();
 sg13g2_decap_8 FILLER_49_2457 ();
 sg13g2_decap_4 FILLER_49_2464 ();
 sg13g2_fill_2 FILLER_49_2468 ();
 sg13g2_fill_2 FILLER_49_2528 ();
 sg13g2_fill_1 FILLER_49_2530 ();
 sg13g2_fill_2 FILLER_49_2561 ();
 sg13g2_fill_1 FILLER_49_2563 ();
 sg13g2_fill_1 FILLER_49_2646 ();
 sg13g2_fill_2 FILLER_49_2651 ();
 sg13g2_decap_4 FILLER_49_2657 ();
 sg13g2_fill_1 FILLER_49_2661 ();
 sg13g2_fill_2 FILLER_49_2665 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_4 FILLER_50_7 ();
 sg13g2_fill_2 FILLER_50_34 ();
 sg13g2_fill_1 FILLER_50_36 ();
 sg13g2_fill_2 FILLER_50_42 ();
 sg13g2_fill_1 FILLER_50_60 ();
 sg13g2_fill_2 FILLER_50_66 ();
 sg13g2_fill_2 FILLER_50_81 ();
 sg13g2_fill_2 FILLER_50_160 ();
 sg13g2_fill_2 FILLER_50_166 ();
 sg13g2_fill_2 FILLER_50_171 ();
 sg13g2_decap_4 FILLER_50_177 ();
 sg13g2_fill_1 FILLER_50_181 ();
 sg13g2_fill_1 FILLER_50_195 ();
 sg13g2_fill_1 FILLER_50_245 ();
 sg13g2_fill_2 FILLER_50_302 ();
 sg13g2_fill_2 FILLER_50_310 ();
 sg13g2_fill_2 FILLER_50_315 ();
 sg13g2_fill_1 FILLER_50_324 ();
 sg13g2_fill_1 FILLER_50_353 ();
 sg13g2_fill_1 FILLER_50_364 ();
 sg13g2_fill_1 FILLER_50_372 ();
 sg13g2_fill_2 FILLER_50_377 ();
 sg13g2_fill_1 FILLER_50_434 ();
 sg13g2_decap_8 FILLER_50_479 ();
 sg13g2_decap_8 FILLER_50_490 ();
 sg13g2_decap_4 FILLER_50_497 ();
 sg13g2_fill_1 FILLER_50_501 ();
 sg13g2_decap_4 FILLER_50_524 ();
 sg13g2_fill_2 FILLER_50_528 ();
 sg13g2_decap_8 FILLER_50_535 ();
 sg13g2_decap_8 FILLER_50_542 ();
 sg13g2_fill_1 FILLER_50_549 ();
 sg13g2_fill_2 FILLER_50_563 ();
 sg13g2_fill_1 FILLER_50_565 ();
 sg13g2_fill_1 FILLER_50_571 ();
 sg13g2_fill_2 FILLER_50_581 ();
 sg13g2_decap_8 FILLER_50_593 ();
 sg13g2_decap_4 FILLER_50_600 ();
 sg13g2_fill_2 FILLER_50_625 ();
 sg13g2_decap_8 FILLER_50_631 ();
 sg13g2_fill_2 FILLER_50_638 ();
 sg13g2_fill_2 FILLER_50_644 ();
 sg13g2_fill_1 FILLER_50_646 ();
 sg13g2_decap_8 FILLER_50_651 ();
 sg13g2_fill_2 FILLER_50_658 ();
 sg13g2_fill_2 FILLER_50_664 ();
 sg13g2_fill_1 FILLER_50_666 ();
 sg13g2_decap_4 FILLER_50_672 ();
 sg13g2_fill_1 FILLER_50_676 ();
 sg13g2_fill_1 FILLER_50_686 ();
 sg13g2_decap_4 FILLER_50_691 ();
 sg13g2_fill_1 FILLER_50_695 ();
 sg13g2_fill_2 FILLER_50_700 ();
 sg13g2_fill_1 FILLER_50_702 ();
 sg13g2_decap_8 FILLER_50_716 ();
 sg13g2_decap_8 FILLER_50_723 ();
 sg13g2_fill_1 FILLER_50_730 ();
 sg13g2_fill_1 FILLER_50_738 ();
 sg13g2_decap_4 FILLER_50_749 ();
 sg13g2_fill_1 FILLER_50_753 ();
 sg13g2_decap_8 FILLER_50_771 ();
 sg13g2_fill_2 FILLER_50_778 ();
 sg13g2_fill_1 FILLER_50_876 ();
 sg13g2_fill_1 FILLER_50_884 ();
 sg13g2_fill_1 FILLER_50_929 ();
 sg13g2_fill_2 FILLER_50_945 ();
 sg13g2_decap_4 FILLER_50_972 ();
 sg13g2_fill_2 FILLER_50_1002 ();
 sg13g2_fill_2 FILLER_50_1008 ();
 sg13g2_fill_1 FILLER_50_1014 ();
 sg13g2_fill_2 FILLER_50_1023 ();
 sg13g2_decap_4 FILLER_50_1037 ();
 sg13g2_fill_2 FILLER_50_1041 ();
 sg13g2_fill_2 FILLER_50_1058 ();
 sg13g2_fill_2 FILLER_50_1065 ();
 sg13g2_fill_1 FILLER_50_1087 ();
 sg13g2_fill_2 FILLER_50_1158 ();
 sg13g2_fill_1 FILLER_50_1228 ();
 sg13g2_fill_1 FILLER_50_1258 ();
 sg13g2_fill_2 FILLER_50_1272 ();
 sg13g2_fill_1 FILLER_50_1278 ();
 sg13g2_fill_2 FILLER_50_1282 ();
 sg13g2_decap_8 FILLER_50_1313 ();
 sg13g2_decap_4 FILLER_50_1320 ();
 sg13g2_fill_1 FILLER_50_1345 ();
 sg13g2_decap_8 FILLER_50_1361 ();
 sg13g2_fill_1 FILLER_50_1373 ();
 sg13g2_fill_1 FILLER_50_1402 ();
 sg13g2_fill_1 FILLER_50_1424 ();
 sg13g2_decap_8 FILLER_50_1430 ();
 sg13g2_fill_2 FILLER_50_1450 ();
 sg13g2_fill_1 FILLER_50_1452 ();
 sg13g2_fill_2 FILLER_50_1458 ();
 sg13g2_fill_1 FILLER_50_1460 ();
 sg13g2_fill_2 FILLER_50_1465 ();
 sg13g2_fill_1 FILLER_50_1477 ();
 sg13g2_fill_2 FILLER_50_1490 ();
 sg13g2_fill_1 FILLER_50_1505 ();
 sg13g2_fill_1 FILLER_50_1531 ();
 sg13g2_fill_1 FILLER_50_1537 ();
 sg13g2_fill_1 FILLER_50_1542 ();
 sg13g2_fill_1 FILLER_50_1589 ();
 sg13g2_fill_2 FILLER_50_1603 ();
 sg13g2_fill_1 FILLER_50_1605 ();
 sg13g2_fill_1 FILLER_50_1611 ();
 sg13g2_fill_1 FILLER_50_1676 ();
 sg13g2_fill_2 FILLER_50_1683 ();
 sg13g2_fill_2 FILLER_50_1715 ();
 sg13g2_fill_2 FILLER_50_1721 ();
 sg13g2_fill_1 FILLER_50_1727 ();
 sg13g2_fill_1 FILLER_50_1751 ();
 sg13g2_decap_8 FILLER_50_1765 ();
 sg13g2_decap_8 FILLER_50_1772 ();
 sg13g2_fill_2 FILLER_50_1779 ();
 sg13g2_decap_8 FILLER_50_1791 ();
 sg13g2_decap_4 FILLER_50_1798 ();
 sg13g2_decap_4 FILLER_50_1815 ();
 sg13g2_fill_1 FILLER_50_1819 ();
 sg13g2_decap_4 FILLER_50_1837 ();
 sg13g2_fill_2 FILLER_50_1841 ();
 sg13g2_decap_8 FILLER_50_1848 ();
 sg13g2_fill_2 FILLER_50_1855 ();
 sg13g2_fill_1 FILLER_50_1869 ();
 sg13g2_fill_1 FILLER_50_1936 ();
 sg13g2_fill_1 FILLER_50_1961 ();
 sg13g2_decap_8 FILLER_50_1977 ();
 sg13g2_fill_1 FILLER_50_1984 ();
 sg13g2_decap_4 FILLER_50_1990 ();
 sg13g2_fill_1 FILLER_50_1999 ();
 sg13g2_fill_1 FILLER_50_2019 ();
 sg13g2_decap_4 FILLER_50_2029 ();
 sg13g2_fill_2 FILLER_50_2037 ();
 sg13g2_fill_1 FILLER_50_2039 ();
 sg13g2_fill_1 FILLER_50_2046 ();
 sg13g2_fill_2 FILLER_50_2053 ();
 sg13g2_fill_1 FILLER_50_2055 ();
 sg13g2_fill_2 FILLER_50_2074 ();
 sg13g2_fill_2 FILLER_50_2087 ();
 sg13g2_fill_1 FILLER_50_2099 ();
 sg13g2_fill_1 FILLER_50_2105 ();
 sg13g2_decap_8 FILLER_50_2112 ();
 sg13g2_decap_8 FILLER_50_2119 ();
 sg13g2_decap_8 FILLER_50_2126 ();
 sg13g2_decap_8 FILLER_50_2133 ();
 sg13g2_decap_8 FILLER_50_2181 ();
 sg13g2_fill_1 FILLER_50_2188 ();
 sg13g2_fill_1 FILLER_50_2223 ();
 sg13g2_decap_8 FILLER_50_2264 ();
 sg13g2_decap_8 FILLER_50_2271 ();
 sg13g2_fill_2 FILLER_50_2278 ();
 sg13g2_fill_1 FILLER_50_2280 ();
 sg13g2_fill_2 FILLER_50_2288 ();
 sg13g2_fill_1 FILLER_50_2290 ();
 sg13g2_decap_8 FILLER_50_2301 ();
 sg13g2_fill_1 FILLER_50_2308 ();
 sg13g2_decap_4 FILLER_50_2328 ();
 sg13g2_fill_2 FILLER_50_2340 ();
 sg13g2_fill_2 FILLER_50_2352 ();
 sg13g2_decap_8 FILLER_50_2359 ();
 sg13g2_fill_2 FILLER_50_2366 ();
 sg13g2_fill_1 FILLER_50_2368 ();
 sg13g2_fill_1 FILLER_50_2378 ();
 sg13g2_fill_2 FILLER_50_2392 ();
 sg13g2_fill_1 FILLER_50_2402 ();
 sg13g2_fill_1 FILLER_50_2413 ();
 sg13g2_fill_1 FILLER_50_2419 ();
 sg13g2_fill_2 FILLER_50_2424 ();
 sg13g2_fill_2 FILLER_50_2430 ();
 sg13g2_fill_2 FILLER_50_2436 ();
 sg13g2_fill_1 FILLER_50_2438 ();
 sg13g2_fill_1 FILLER_50_2465 ();
 sg13g2_fill_2 FILLER_50_2487 ();
 sg13g2_fill_1 FILLER_50_2489 ();
 sg13g2_fill_1 FILLER_50_2495 ();
 sg13g2_fill_2 FILLER_50_2501 ();
 sg13g2_fill_1 FILLER_50_2503 ();
 sg13g2_decap_4 FILLER_50_2530 ();
 sg13g2_fill_1 FILLER_50_2534 ();
 sg13g2_decap_8 FILLER_50_2561 ();
 sg13g2_fill_2 FILLER_50_2568 ();
 sg13g2_fill_1 FILLER_50_2570 ();
 sg13g2_decap_4 FILLER_50_2576 ();
 sg13g2_fill_1 FILLER_50_2604 ();
 sg13g2_fill_2 FILLER_50_2617 ();
 sg13g2_fill_1 FILLER_50_2625 ();
 sg13g2_fill_1 FILLER_50_2641 ();
 sg13g2_fill_2 FILLER_50_2668 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_fill_1 FILLER_51_14 ();
 sg13g2_fill_1 FILLER_51_45 ();
 sg13g2_fill_1 FILLER_51_50 ();
 sg13g2_fill_2 FILLER_51_68 ();
 sg13g2_fill_1 FILLER_51_88 ();
 sg13g2_decap_4 FILLER_51_105 ();
 sg13g2_fill_1 FILLER_51_128 ();
 sg13g2_fill_2 FILLER_51_154 ();
 sg13g2_decap_8 FILLER_51_162 ();
 sg13g2_fill_2 FILLER_51_169 ();
 sg13g2_fill_1 FILLER_51_187 ();
 sg13g2_fill_2 FILLER_51_196 ();
 sg13g2_fill_1 FILLER_51_205 ();
 sg13g2_fill_2 FILLER_51_226 ();
 sg13g2_fill_1 FILLER_51_232 ();
 sg13g2_fill_2 FILLER_51_274 ();
 sg13g2_fill_1 FILLER_51_282 ();
 sg13g2_fill_1 FILLER_51_293 ();
 sg13g2_fill_2 FILLER_51_304 ();
 sg13g2_fill_1 FILLER_51_351 ();
 sg13g2_fill_2 FILLER_51_403 ();
 sg13g2_fill_1 FILLER_51_443 ();
 sg13g2_fill_1 FILLER_51_481 ();
 sg13g2_fill_2 FILLER_51_486 ();
 sg13g2_decap_4 FILLER_51_492 ();
 sg13g2_decap_8 FILLER_51_500 ();
 sg13g2_fill_2 FILLER_51_507 ();
 sg13g2_decap_8 FILLER_51_523 ();
 sg13g2_decap_8 FILLER_51_542 ();
 sg13g2_fill_2 FILLER_51_558 ();
 sg13g2_fill_1 FILLER_51_560 ();
 sg13g2_fill_2 FILLER_51_566 ();
 sg13g2_fill_1 FILLER_51_578 ();
 sg13g2_decap_4 FILLER_51_583 ();
 sg13g2_decap_8 FILLER_51_590 ();
 sg13g2_decap_8 FILLER_51_597 ();
 sg13g2_decap_8 FILLER_51_604 ();
 sg13g2_decap_8 FILLER_51_615 ();
 sg13g2_decap_8 FILLER_51_622 ();
 sg13g2_fill_2 FILLER_51_629 ();
 sg13g2_fill_1 FILLER_51_631 ();
 sg13g2_decap_4 FILLER_51_637 ();
 sg13g2_fill_1 FILLER_51_641 ();
 sg13g2_fill_2 FILLER_51_660 ();
 sg13g2_fill_2 FILLER_51_697 ();
 sg13g2_fill_2 FILLER_51_719 ();
 sg13g2_fill_1 FILLER_51_773 ();
 sg13g2_decap_4 FILLER_51_779 ();
 sg13g2_fill_1 FILLER_51_783 ();
 sg13g2_fill_1 FILLER_51_847 ();
 sg13g2_fill_1 FILLER_51_935 ();
 sg13g2_decap_8 FILLER_51_970 ();
 sg13g2_decap_4 FILLER_51_977 ();
 sg13g2_decap_8 FILLER_51_989 ();
 sg13g2_decap_4 FILLER_51_996 ();
 sg13g2_fill_2 FILLER_51_1000 ();
 sg13g2_decap_8 FILLER_51_1026 ();
 sg13g2_decap_8 FILLER_51_1033 ();
 sg13g2_decap_8 FILLER_51_1040 ();
 sg13g2_fill_2 FILLER_51_1073 ();
 sg13g2_fill_1 FILLER_51_1075 ();
 sg13g2_decap_4 FILLER_51_1110 ();
 sg13g2_fill_2 FILLER_51_1114 ();
 sg13g2_fill_2 FILLER_51_1192 ();
 sg13g2_fill_1 FILLER_51_1318 ();
 sg13g2_decap_8 FILLER_51_1355 ();
 sg13g2_decap_8 FILLER_51_1362 ();
 sg13g2_decap_8 FILLER_51_1369 ();
 sg13g2_fill_1 FILLER_51_1376 ();
 sg13g2_fill_1 FILLER_51_1381 ();
 sg13g2_fill_2 FILLER_51_1387 ();
 sg13g2_decap_4 FILLER_51_1394 ();
 sg13g2_fill_1 FILLER_51_1408 ();
 sg13g2_fill_1 FILLER_51_1413 ();
 sg13g2_fill_2 FILLER_51_1423 ();
 sg13g2_decap_4 FILLER_51_1431 ();
 sg13g2_fill_1 FILLER_51_1435 ();
 sg13g2_fill_2 FILLER_51_1450 ();
 sg13g2_fill_1 FILLER_51_1452 ();
 sg13g2_decap_8 FILLER_51_1458 ();
 sg13g2_fill_2 FILLER_51_1465 ();
 sg13g2_fill_2 FILLER_51_1471 ();
 sg13g2_fill_2 FILLER_51_1478 ();
 sg13g2_decap_8 FILLER_51_1523 ();
 sg13g2_decap_4 FILLER_51_1534 ();
 sg13g2_fill_2 FILLER_51_1543 ();
 sg13g2_fill_1 FILLER_51_1545 ();
 sg13g2_fill_1 FILLER_51_1551 ();
 sg13g2_decap_8 FILLER_51_1570 ();
 sg13g2_decap_8 FILLER_51_1577 ();
 sg13g2_decap_8 FILLER_51_1584 ();
 sg13g2_decap_4 FILLER_51_1591 ();
 sg13g2_fill_1 FILLER_51_1595 ();
 sg13g2_decap_8 FILLER_51_1608 ();
 sg13g2_decap_8 FILLER_51_1615 ();
 sg13g2_decap_8 FILLER_51_1622 ();
 sg13g2_fill_1 FILLER_51_1629 ();
 sg13g2_fill_1 FILLER_51_1658 ();
 sg13g2_fill_1 FILLER_51_1667 ();
 sg13g2_fill_2 FILLER_51_1716 ();
 sg13g2_fill_1 FILLER_51_1718 ();
 sg13g2_fill_2 FILLER_51_1755 ();
 sg13g2_decap_8 FILLER_51_1808 ();
 sg13g2_fill_1 FILLER_51_1815 ();
 sg13g2_decap_4 FILLER_51_1824 ();
 sg13g2_fill_2 FILLER_51_1846 ();
 sg13g2_fill_1 FILLER_51_1848 ();
 sg13g2_fill_2 FILLER_51_1854 ();
 sg13g2_fill_1 FILLER_51_1856 ();
 sg13g2_fill_2 FILLER_51_1862 ();
 sg13g2_fill_2 FILLER_51_1872 ();
 sg13g2_fill_2 FILLER_51_1880 ();
 sg13g2_fill_2 FILLER_51_1887 ();
 sg13g2_fill_1 FILLER_51_1889 ();
 sg13g2_decap_4 FILLER_51_1896 ();
 sg13g2_fill_2 FILLER_51_1979 ();
 sg13g2_decap_4 FILLER_51_1990 ();
 sg13g2_fill_2 FILLER_51_1994 ();
 sg13g2_fill_1 FILLER_51_2001 ();
 sg13g2_fill_1 FILLER_51_2016 ();
 sg13g2_fill_1 FILLER_51_2021 ();
 sg13g2_fill_2 FILLER_51_2026 ();
 sg13g2_fill_2 FILLER_51_2048 ();
 sg13g2_fill_1 FILLER_51_2055 ();
 sg13g2_fill_1 FILLER_51_2078 ();
 sg13g2_fill_1 FILLER_51_2106 ();
 sg13g2_decap_8 FILLER_51_2111 ();
 sg13g2_decap_8 FILLER_51_2118 ();
 sg13g2_decap_8 FILLER_51_2125 ();
 sg13g2_decap_8 FILLER_51_2132 ();
 sg13g2_decap_8 FILLER_51_2139 ();
 sg13g2_fill_2 FILLER_51_2146 ();
 sg13g2_decap_4 FILLER_51_2152 ();
 sg13g2_fill_2 FILLER_51_2156 ();
 sg13g2_decap_4 FILLER_51_2162 ();
 sg13g2_fill_2 FILLER_51_2206 ();
 sg13g2_decap_8 FILLER_51_2269 ();
 sg13g2_fill_1 FILLER_51_2307 ();
 sg13g2_fill_2 FILLER_51_2312 ();
 sg13g2_fill_1 FILLER_51_2314 ();
 sg13g2_fill_2 FILLER_51_2319 ();
 sg13g2_decap_8 FILLER_51_2351 ();
 sg13g2_fill_2 FILLER_51_2358 ();
 sg13g2_fill_2 FILLER_51_2376 ();
 sg13g2_fill_1 FILLER_51_2388 ();
 sg13g2_fill_2 FILLER_51_2399 ();
 sg13g2_fill_2 FILLER_51_2411 ();
 sg13g2_fill_1 FILLER_51_2413 ();
 sg13g2_fill_1 FILLER_51_2418 ();
 sg13g2_fill_1 FILLER_51_2427 ();
 sg13g2_fill_2 FILLER_51_2468 ();
 sg13g2_fill_2 FILLER_51_2480 ();
 sg13g2_fill_1 FILLER_51_2482 ();
 sg13g2_decap_8 FILLER_51_2560 ();
 sg13g2_decap_8 FILLER_51_2567 ();
 sg13g2_decap_8 FILLER_51_2574 ();
 sg13g2_decap_4 FILLER_51_2581 ();
 sg13g2_fill_1 FILLER_51_2585 ();
 sg13g2_decap_4 FILLER_51_2591 ();
 sg13g2_fill_2 FILLER_51_2609 ();
 sg13g2_decap_8 FILLER_51_2657 ();
 sg13g2_decap_4 FILLER_51_2664 ();
 sg13g2_fill_2 FILLER_51_2668 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_fill_2 FILLER_52_7 ();
 sg13g2_fill_2 FILLER_52_40 ();
 sg13g2_fill_2 FILLER_52_55 ();
 sg13g2_fill_1 FILLER_52_57 ();
 sg13g2_fill_2 FILLER_52_102 ();
 sg13g2_fill_1 FILLER_52_108 ();
 sg13g2_fill_2 FILLER_52_113 ();
 sg13g2_fill_1 FILLER_52_155 ();
 sg13g2_fill_1 FILLER_52_174 ();
 sg13g2_fill_1 FILLER_52_180 ();
 sg13g2_fill_2 FILLER_52_185 ();
 sg13g2_fill_1 FILLER_52_191 ();
 sg13g2_fill_1 FILLER_52_196 ();
 sg13g2_decap_4 FILLER_52_201 ();
 sg13g2_decap_4 FILLER_52_225 ();
 sg13g2_fill_1 FILLER_52_229 ();
 sg13g2_fill_2 FILLER_52_236 ();
 sg13g2_fill_2 FILLER_52_258 ();
 sg13g2_fill_1 FILLER_52_260 ();
 sg13g2_fill_1 FILLER_52_296 ();
 sg13g2_fill_2 FILLER_52_310 ();
 sg13g2_fill_1 FILLER_52_315 ();
 sg13g2_fill_2 FILLER_52_366 ();
 sg13g2_fill_1 FILLER_52_392 ();
 sg13g2_fill_2 FILLER_52_400 ();
 sg13g2_fill_1 FILLER_52_459 ();
 sg13g2_fill_2 FILLER_52_472 ();
 sg13g2_fill_1 FILLER_52_514 ();
 sg13g2_fill_1 FILLER_52_540 ();
 sg13g2_decap_8 FILLER_52_546 ();
 sg13g2_fill_1 FILLER_52_553 ();
 sg13g2_decap_8 FILLER_52_598 ();
 sg13g2_decap_8 FILLER_52_605 ();
 sg13g2_decap_8 FILLER_52_612 ();
 sg13g2_decap_8 FILLER_52_685 ();
 sg13g2_decap_4 FILLER_52_692 ();
 sg13g2_fill_2 FILLER_52_696 ();
 sg13g2_fill_2 FILLER_52_770 ();
 sg13g2_fill_1 FILLER_52_772 ();
 sg13g2_fill_1 FILLER_52_830 ();
 sg13g2_fill_1 FILLER_52_924 ();
 sg13g2_fill_2 FILLER_52_936 ();
 sg13g2_fill_1 FILLER_52_941 ();
 sg13g2_fill_1 FILLER_52_956 ();
 sg13g2_decap_8 FILLER_52_987 ();
 sg13g2_decap_8 FILLER_52_994 ();
 sg13g2_decap_8 FILLER_52_1001 ();
 sg13g2_decap_8 FILLER_52_1008 ();
 sg13g2_fill_1 FILLER_52_1015 ();
 sg13g2_decap_8 FILLER_52_1047 ();
 sg13g2_fill_1 FILLER_52_1054 ();
 sg13g2_decap_8 FILLER_52_1059 ();
 sg13g2_decap_8 FILLER_52_1066 ();
 sg13g2_decap_8 FILLER_52_1073 ();
 sg13g2_decap_4 FILLER_52_1080 ();
 sg13g2_decap_8 FILLER_52_1088 ();
 sg13g2_decap_8 FILLER_52_1095 ();
 sg13g2_fill_2 FILLER_52_1102 ();
 sg13g2_decap_4 FILLER_52_1111 ();
 sg13g2_fill_1 FILLER_52_1115 ();
 sg13g2_fill_1 FILLER_52_1172 ();
 sg13g2_decap_8 FILLER_52_1205 ();
 sg13g2_decap_8 FILLER_52_1212 ();
 sg13g2_decap_8 FILLER_52_1219 ();
 sg13g2_fill_1 FILLER_52_1226 ();
 sg13g2_decap_8 FILLER_52_1232 ();
 sg13g2_fill_1 FILLER_52_1275 ();
 sg13g2_fill_2 FILLER_52_1282 ();
 sg13g2_fill_2 FILLER_52_1296 ();
 sg13g2_decap_4 FILLER_52_1317 ();
 sg13g2_fill_1 FILLER_52_1321 ();
 sg13g2_fill_2 FILLER_52_1348 ();
 sg13g2_decap_8 FILLER_52_1354 ();
 sg13g2_fill_2 FILLER_52_1361 ();
 sg13g2_fill_2 FILLER_52_1367 ();
 sg13g2_fill_2 FILLER_52_1373 ();
 sg13g2_fill_2 FILLER_52_1402 ();
 sg13g2_fill_1 FILLER_52_1404 ();
 sg13g2_fill_2 FILLER_52_1409 ();
 sg13g2_decap_4 FILLER_52_1421 ();
 sg13g2_fill_2 FILLER_52_1425 ();
 sg13g2_fill_2 FILLER_52_1431 ();
 sg13g2_fill_1 FILLER_52_1450 ();
 sg13g2_fill_1 FILLER_52_1461 ();
 sg13g2_fill_1 FILLER_52_1467 ();
 sg13g2_fill_1 FILLER_52_1498 ();
 sg13g2_fill_1 FILLER_52_1503 ();
 sg13g2_fill_1 FILLER_52_1513 ();
 sg13g2_fill_1 FILLER_52_1530 ();
 sg13g2_fill_1 FILLER_52_1540 ();
 sg13g2_fill_2 FILLER_52_1545 ();
 sg13g2_fill_1 FILLER_52_1547 ();
 sg13g2_fill_2 FILLER_52_1552 ();
 sg13g2_decap_8 FILLER_52_1558 ();
 sg13g2_decap_8 FILLER_52_1565 ();
 sg13g2_decap_4 FILLER_52_1572 ();
 sg13g2_fill_2 FILLER_52_1576 ();
 sg13g2_decap_8 FILLER_52_1604 ();
 sg13g2_decap_8 FILLER_52_1611 ();
 sg13g2_fill_2 FILLER_52_1618 ();
 sg13g2_fill_1 FILLER_52_1635 ();
 sg13g2_fill_2 FILLER_52_1641 ();
 sg13g2_fill_2 FILLER_52_1657 ();
 sg13g2_fill_1 FILLER_52_1692 ();
 sg13g2_fill_2 FILLER_52_1701 ();
 sg13g2_fill_1 FILLER_52_1740 ();
 sg13g2_fill_1 FILLER_52_1757 ();
 sg13g2_fill_1 FILLER_52_1787 ();
 sg13g2_fill_1 FILLER_52_1798 ();
 sg13g2_fill_1 FILLER_52_1804 ();
 sg13g2_decap_4 FILLER_52_1812 ();
 sg13g2_fill_1 FILLER_52_1816 ();
 sg13g2_fill_2 FILLER_52_1821 ();
 sg13g2_decap_4 FILLER_52_1838 ();
 sg13g2_fill_2 FILLER_52_1842 ();
 sg13g2_decap_8 FILLER_52_1848 ();
 sg13g2_decap_4 FILLER_52_1868 ();
 sg13g2_fill_2 FILLER_52_1872 ();
 sg13g2_decap_8 FILLER_52_1894 ();
 sg13g2_fill_2 FILLER_52_1901 ();
 sg13g2_fill_1 FILLER_52_1915 ();
 sg13g2_decap_4 FILLER_52_1921 ();
 sg13g2_fill_1 FILLER_52_1934 ();
 sg13g2_fill_1 FILLER_52_1940 ();
 sg13g2_decap_4 FILLER_52_1973 ();
 sg13g2_fill_2 FILLER_52_1977 ();
 sg13g2_fill_2 FILLER_52_1983 ();
 sg13g2_fill_2 FILLER_52_1990 ();
 sg13g2_fill_1 FILLER_52_1992 ();
 sg13g2_decap_8 FILLER_52_2001 ();
 sg13g2_decap_8 FILLER_52_2012 ();
 sg13g2_fill_1 FILLER_52_2019 ();
 sg13g2_fill_1 FILLER_52_2024 ();
 sg13g2_decap_8 FILLER_52_2030 ();
 sg13g2_fill_1 FILLER_52_2037 ();
 sg13g2_fill_2 FILLER_52_2051 ();
 sg13g2_fill_1 FILLER_52_2053 ();
 sg13g2_fill_2 FILLER_52_2072 ();
 sg13g2_fill_1 FILLER_52_2074 ();
 sg13g2_decap_8 FILLER_52_2105 ();
 sg13g2_decap_8 FILLER_52_2112 ();
 sg13g2_decap_8 FILLER_52_2119 ();
 sg13g2_decap_8 FILLER_52_2126 ();
 sg13g2_fill_1 FILLER_52_2133 ();
 sg13g2_fill_1 FILLER_52_2138 ();
 sg13g2_fill_2 FILLER_52_2226 ();
 sg13g2_fill_1 FILLER_52_2254 ();
 sg13g2_decap_8 FILLER_52_2265 ();
 sg13g2_fill_2 FILLER_52_2272 ();
 sg13g2_fill_1 FILLER_52_2274 ();
 sg13g2_decap_8 FILLER_52_2279 ();
 sg13g2_fill_1 FILLER_52_2286 ();
 sg13g2_decap_8 FILLER_52_2291 ();
 sg13g2_fill_2 FILLER_52_2298 ();
 sg13g2_decap_4 FILLER_52_2304 ();
 sg13g2_decap_8 FILLER_52_2422 ();
 sg13g2_fill_1 FILLER_52_2429 ();
 sg13g2_fill_2 FILLER_52_2440 ();
 sg13g2_decap_8 FILLER_52_2450 ();
 sg13g2_decap_8 FILLER_52_2457 ();
 sg13g2_decap_4 FILLER_52_2468 ();
 sg13g2_fill_2 FILLER_52_2490 ();
 sg13g2_fill_1 FILLER_52_2492 ();
 sg13g2_fill_1 FILLER_52_2535 ();
 sg13g2_decap_8 FILLER_52_2545 ();
 sg13g2_fill_2 FILLER_52_2552 ();
 sg13g2_decap_4 FILLER_52_2560 ();
 sg13g2_fill_2 FILLER_52_2604 ();
 sg13g2_fill_1 FILLER_52_2609 ();
 sg13g2_fill_2 FILLER_52_2667 ();
 sg13g2_fill_1 FILLER_52_2669 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_4 FILLER_53_7 ();
 sg13g2_fill_1 FILLER_53_41 ();
 sg13g2_decap_4 FILLER_53_47 ();
 sg13g2_decap_8 FILLER_53_60 ();
 sg13g2_decap_4 FILLER_53_67 ();
 sg13g2_fill_2 FILLER_53_71 ();
 sg13g2_fill_1 FILLER_53_78 ();
 sg13g2_fill_1 FILLER_53_84 ();
 sg13g2_fill_2 FILLER_53_89 ();
 sg13g2_fill_2 FILLER_53_101 ();
 sg13g2_fill_1 FILLER_53_103 ();
 sg13g2_fill_2 FILLER_53_108 ();
 sg13g2_fill_1 FILLER_53_110 ();
 sg13g2_fill_1 FILLER_53_116 ();
 sg13g2_fill_2 FILLER_53_121 ();
 sg13g2_fill_1 FILLER_53_161 ();
 sg13g2_fill_1 FILLER_53_167 ();
 sg13g2_fill_1 FILLER_53_187 ();
 sg13g2_fill_1 FILLER_53_197 ();
 sg13g2_fill_1 FILLER_53_203 ();
 sg13g2_decap_8 FILLER_53_218 ();
 sg13g2_decap_8 FILLER_53_225 ();
 sg13g2_decap_8 FILLER_53_232 ();
 sg13g2_decap_8 FILLER_53_239 ();
 sg13g2_decap_8 FILLER_53_246 ();
 sg13g2_decap_8 FILLER_53_253 ();
 sg13g2_fill_1 FILLER_53_260 ();
 sg13g2_fill_1 FILLER_53_272 ();
 sg13g2_fill_2 FILLER_53_341 ();
 sg13g2_fill_2 FILLER_53_354 ();
 sg13g2_fill_1 FILLER_53_361 ();
 sg13g2_fill_2 FILLER_53_391 ();
 sg13g2_fill_2 FILLER_53_397 ();
 sg13g2_fill_1 FILLER_53_477 ();
 sg13g2_fill_1 FILLER_53_590 ();
 sg13g2_fill_2 FILLER_53_598 ();
 sg13g2_fill_1 FILLER_53_609 ();
 sg13g2_fill_1 FILLER_53_621 ();
 sg13g2_decap_8 FILLER_53_630 ();
 sg13g2_decap_4 FILLER_53_645 ();
 sg13g2_fill_2 FILLER_53_649 ();
 sg13g2_fill_1 FILLER_53_655 ();
 sg13g2_fill_1 FILLER_53_659 ();
 sg13g2_fill_2 FILLER_53_668 ();
 sg13g2_fill_2 FILLER_53_709 ();
 sg13g2_fill_1 FILLER_53_730 ();
 sg13g2_fill_1 FILLER_53_782 ();
 sg13g2_decap_8 FILLER_53_788 ();
 sg13g2_decap_8 FILLER_53_799 ();
 sg13g2_fill_1 FILLER_53_819 ();
 sg13g2_fill_1 FILLER_53_862 ();
 sg13g2_fill_2 FILLER_53_973 ();
 sg13g2_fill_2 FILLER_53_984 ();
 sg13g2_decap_4 FILLER_53_998 ();
 sg13g2_fill_2 FILLER_53_1002 ();
 sg13g2_fill_2 FILLER_53_1035 ();
 sg13g2_decap_8 FILLER_53_1073 ();
 sg13g2_decap_4 FILLER_53_1080 ();
 sg13g2_decap_4 FILLER_53_1090 ();
 sg13g2_fill_2 FILLER_53_1102 ();
 sg13g2_decap_4 FILLER_53_1124 ();
 sg13g2_fill_1 FILLER_53_1183 ();
 sg13g2_decap_8 FILLER_53_1214 ();
 sg13g2_decap_8 FILLER_53_1221 ();
 sg13g2_decap_8 FILLER_53_1228 ();
 sg13g2_fill_2 FILLER_53_1235 ();
 sg13g2_fill_1 FILLER_53_1237 ();
 sg13g2_decap_4 FILLER_53_1246 ();
 sg13g2_fill_1 FILLER_53_1260 ();
 sg13g2_fill_2 FILLER_53_1313 ();
 sg13g2_fill_1 FILLER_53_1326 ();
 sg13g2_decap_4 FILLER_53_1349 ();
 sg13g2_fill_1 FILLER_53_1353 ();
 sg13g2_fill_2 FILLER_53_1358 ();
 sg13g2_fill_1 FILLER_53_1373 ();
 sg13g2_fill_2 FILLER_53_1405 ();
 sg13g2_decap_8 FILLER_53_1411 ();
 sg13g2_fill_2 FILLER_53_1418 ();
 sg13g2_fill_1 FILLER_53_1420 ();
 sg13g2_fill_2 FILLER_53_1435 ();
 sg13g2_decap_4 FILLER_53_1442 ();
 sg13g2_fill_2 FILLER_53_1446 ();
 sg13g2_decap_8 FILLER_53_1453 ();
 sg13g2_decap_8 FILLER_53_1460 ();
 sg13g2_decap_4 FILLER_53_1467 ();
 sg13g2_fill_2 FILLER_53_1476 ();
 sg13g2_fill_1 FILLER_53_1483 ();
 sg13g2_fill_2 FILLER_53_1490 ();
 sg13g2_fill_1 FILLER_53_1499 ();
 sg13g2_decap_8 FILLER_53_1509 ();
 sg13g2_fill_2 FILLER_53_1582 ();
 sg13g2_fill_2 FILLER_53_1596 ();
 sg13g2_decap_8 FILLER_53_1602 ();
 sg13g2_decap_8 FILLER_53_1622 ();
 sg13g2_decap_4 FILLER_53_1634 ();
 sg13g2_decap_4 FILLER_53_1655 ();
 sg13g2_fill_1 FILLER_53_1676 ();
 sg13g2_decap_8 FILLER_53_1697 ();
 sg13g2_decap_8 FILLER_53_1704 ();
 sg13g2_decap_8 FILLER_53_1711 ();
 sg13g2_fill_1 FILLER_53_1718 ();
 sg13g2_fill_1 FILLER_53_1736 ();
 sg13g2_fill_1 FILLER_53_1742 ();
 sg13g2_fill_2 FILLER_53_1760 ();
 sg13g2_fill_1 FILLER_53_1785 ();
 sg13g2_fill_1 FILLER_53_1806 ();
 sg13g2_decap_8 FILLER_53_1842 ();
 sg13g2_decap_8 FILLER_53_1849 ();
 sg13g2_decap_8 FILLER_53_1856 ();
 sg13g2_decap_8 FILLER_53_1863 ();
 sg13g2_decap_8 FILLER_53_1870 ();
 sg13g2_decap_8 FILLER_53_1877 ();
 sg13g2_fill_2 FILLER_53_1884 ();
 sg13g2_fill_2 FILLER_53_1911 ();
 sg13g2_decap_4 FILLER_53_1939 ();
 sg13g2_fill_2 FILLER_53_1947 ();
 sg13g2_decap_4 FILLER_53_1966 ();
 sg13g2_fill_2 FILLER_53_1970 ();
 sg13g2_fill_2 FILLER_53_1981 ();
 sg13g2_decap_4 FILLER_53_1990 ();
 sg13g2_fill_2 FILLER_53_1994 ();
 sg13g2_decap_8 FILLER_53_2001 ();
 sg13g2_decap_8 FILLER_53_2008 ();
 sg13g2_decap_4 FILLER_53_2019 ();
 sg13g2_fill_1 FILLER_53_2039 ();
 sg13g2_fill_1 FILLER_53_2056 ();
 sg13g2_fill_2 FILLER_53_2087 ();
 sg13g2_fill_1 FILLER_53_2089 ();
 sg13g2_fill_2 FILLER_53_2094 ();
 sg13g2_fill_1 FILLER_53_2096 ();
 sg13g2_fill_2 FILLER_53_2106 ();
 sg13g2_decap_8 FILLER_53_2113 ();
 sg13g2_decap_8 FILLER_53_2120 ();
 sg13g2_fill_1 FILLER_53_2127 ();
 sg13g2_decap_8 FILLER_53_2174 ();
 sg13g2_fill_2 FILLER_53_2181 ();
 sg13g2_decap_8 FILLER_53_2187 ();
 sg13g2_fill_1 FILLER_53_2194 ();
 sg13g2_decap_8 FILLER_53_2200 ();
 sg13g2_fill_2 FILLER_53_2207 ();
 sg13g2_fill_2 FILLER_53_2213 ();
 sg13g2_fill_1 FILLER_53_2215 ();
 sg13g2_decap_4 FILLER_53_2238 ();
 sg13g2_fill_1 FILLER_53_2242 ();
 sg13g2_fill_1 FILLER_53_2294 ();
 sg13g2_decap_8 FILLER_53_2312 ();
 sg13g2_decap_4 FILLER_53_2319 ();
 sg13g2_decap_4 FILLER_53_2337 ();
 sg13g2_fill_2 FILLER_53_2372 ();
 sg13g2_fill_2 FILLER_53_2404 ();
 sg13g2_fill_1 FILLER_53_2406 ();
 sg13g2_fill_2 FILLER_53_2439 ();
 sg13g2_fill_2 FILLER_53_2451 ();
 sg13g2_fill_1 FILLER_53_2453 ();
 sg13g2_fill_2 FILLER_53_2458 ();
 sg13g2_fill_1 FILLER_53_2460 ();
 sg13g2_fill_2 FILLER_53_2466 ();
 sg13g2_fill_1 FILLER_53_2468 ();
 sg13g2_fill_2 FILLER_53_2532 ();
 sg13g2_fill_2 FILLER_53_2540 ();
 sg13g2_decap_4 FILLER_53_2546 ();
 sg13g2_fill_1 FILLER_53_2550 ();
 sg13g2_fill_2 FILLER_53_2587 ();
 sg13g2_decap_8 FILLER_53_2640 ();
 sg13g2_fill_1 FILLER_53_2647 ();
 sg13g2_decap_8 FILLER_53_2652 ();
 sg13g2_decap_8 FILLER_53_2659 ();
 sg13g2_decap_4 FILLER_53_2666 ();
 sg13g2_fill_2 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_77 ();
 sg13g2_fill_1 FILLER_54_79 ();
 sg13g2_fill_2 FILLER_54_90 ();
 sg13g2_fill_1 FILLER_54_92 ();
 sg13g2_fill_1 FILLER_54_139 ();
 sg13g2_fill_2 FILLER_54_144 ();
 sg13g2_fill_2 FILLER_54_173 ();
 sg13g2_decap_4 FILLER_54_198 ();
 sg13g2_fill_2 FILLER_54_206 ();
 sg13g2_fill_1 FILLER_54_208 ();
 sg13g2_fill_2 FILLER_54_230 ();
 sg13g2_decap_4 FILLER_54_242 ();
 sg13g2_fill_2 FILLER_54_246 ();
 sg13g2_fill_2 FILLER_54_258 ();
 sg13g2_fill_1 FILLER_54_260 ();
 sg13g2_fill_1 FILLER_54_271 ();
 sg13g2_fill_2 FILLER_54_354 ();
 sg13g2_fill_1 FILLER_54_378 ();
 sg13g2_fill_1 FILLER_54_412 ();
 sg13g2_fill_1 FILLER_54_434 ();
 sg13g2_fill_1 FILLER_54_439 ();
 sg13g2_fill_1 FILLER_54_497 ();
 sg13g2_fill_2 FILLER_54_522 ();
 sg13g2_fill_1 FILLER_54_533 ();
 sg13g2_decap_4 FILLER_54_542 ();
 sg13g2_fill_1 FILLER_54_565 ();
 sg13g2_fill_1 FILLER_54_575 ();
 sg13g2_fill_2 FILLER_54_613 ();
 sg13g2_fill_1 FILLER_54_615 ();
 sg13g2_fill_2 FILLER_54_628 ();
 sg13g2_fill_1 FILLER_54_630 ();
 sg13g2_fill_2 FILLER_54_635 ();
 sg13g2_fill_1 FILLER_54_641 ();
 sg13g2_decap_4 FILLER_54_647 ();
 sg13g2_fill_1 FILLER_54_651 ();
 sg13g2_fill_1 FILLER_54_668 ();
 sg13g2_decap_4 FILLER_54_678 ();
 sg13g2_fill_1 FILLER_54_694 ();
 sg13g2_fill_2 FILLER_54_740 ();
 sg13g2_decap_8 FILLER_54_759 ();
 sg13g2_decap_4 FILLER_54_766 ();
 sg13g2_decap_8 FILLER_54_775 ();
 sg13g2_fill_1 FILLER_54_782 ();
 sg13g2_fill_2 FILLER_54_788 ();
 sg13g2_fill_1 FILLER_54_790 ();
 sg13g2_decap_8 FILLER_54_800 ();
 sg13g2_decap_4 FILLER_54_807 ();
 sg13g2_fill_1 FILLER_54_811 ();
 sg13g2_fill_1 FILLER_54_820 ();
 sg13g2_fill_2 FILLER_54_918 ();
 sg13g2_fill_1 FILLER_54_964 ();
 sg13g2_decap_4 FILLER_54_1000 ();
 sg13g2_fill_2 FILLER_54_1004 ();
 sg13g2_fill_2 FILLER_54_1015 ();
 sg13g2_fill_1 FILLER_54_1017 ();
 sg13g2_decap_8 FILLER_54_1076 ();
 sg13g2_fill_1 FILLER_54_1083 ();
 sg13g2_decap_8 FILLER_54_1088 ();
 sg13g2_fill_1 FILLER_54_1095 ();
 sg13g2_decap_8 FILLER_54_1112 ();
 sg13g2_decap_4 FILLER_54_1119 ();
 sg13g2_fill_1 FILLER_54_1123 ();
 sg13g2_decap_4 FILLER_54_1136 ();
 sg13g2_fill_1 FILLER_54_1140 ();
 sg13g2_fill_2 FILLER_54_1162 ();
 sg13g2_fill_2 FILLER_54_1179 ();
 sg13g2_decap_4 FILLER_54_1188 ();
 sg13g2_fill_2 FILLER_54_1192 ();
 sg13g2_decap_8 FILLER_54_1218 ();
 sg13g2_fill_2 FILLER_54_1248 ();
 sg13g2_fill_1 FILLER_54_1257 ();
 sg13g2_fill_2 FILLER_54_1291 ();
 sg13g2_fill_2 FILLER_54_1315 ();
 sg13g2_fill_1 FILLER_54_1317 ();
 sg13g2_fill_2 FILLER_54_1323 ();
 sg13g2_decap_8 FILLER_54_1329 ();
 sg13g2_fill_1 FILLER_54_1341 ();
 sg13g2_decap_8 FILLER_54_1352 ();
 sg13g2_decap_4 FILLER_54_1359 ();
 sg13g2_fill_1 FILLER_54_1374 ();
 sg13g2_fill_1 FILLER_54_1386 ();
 sg13g2_fill_1 FILLER_54_1397 ();
 sg13g2_fill_2 FILLER_54_1404 ();
 sg13g2_fill_1 FILLER_54_1416 ();
 sg13g2_fill_1 FILLER_54_1442 ();
 sg13g2_fill_2 FILLER_54_1453 ();
 sg13g2_fill_1 FILLER_54_1455 ();
 sg13g2_decap_8 FILLER_54_1461 ();
 sg13g2_fill_1 FILLER_54_1483 ();
 sg13g2_fill_1 FILLER_54_1492 ();
 sg13g2_decap_8 FILLER_54_1497 ();
 sg13g2_decap_4 FILLER_54_1601 ();
 sg13g2_fill_2 FILLER_54_1605 ();
 sg13g2_decap_4 FILLER_54_1633 ();
 sg13g2_fill_2 FILLER_54_1637 ();
 sg13g2_decap_4 FILLER_54_1653 ();
 sg13g2_fill_1 FILLER_54_1657 ();
 sg13g2_fill_2 FILLER_54_1664 ();
 sg13g2_decap_8 FILLER_54_1710 ();
 sg13g2_decap_8 FILLER_54_1717 ();
 sg13g2_decap_4 FILLER_54_1724 ();
 sg13g2_fill_1 FILLER_54_1728 ();
 sg13g2_fill_1 FILLER_54_1772 ();
 sg13g2_decap_4 FILLER_54_1779 ();
 sg13g2_fill_1 FILLER_54_1783 ();
 sg13g2_fill_1 FILLER_54_1793 ();
 sg13g2_fill_1 FILLER_54_1823 ();
 sg13g2_fill_1 FILLER_54_1829 ();
 sg13g2_fill_2 FILLER_54_1839 ();
 sg13g2_fill_1 FILLER_54_1841 ();
 sg13g2_fill_1 FILLER_54_1846 ();
 sg13g2_fill_2 FILLER_54_1855 ();
 sg13g2_fill_1 FILLER_54_1862 ();
 sg13g2_fill_2 FILLER_54_1868 ();
 sg13g2_fill_2 FILLER_54_1875 ();
 sg13g2_fill_2 FILLER_54_1885 ();
 sg13g2_fill_1 FILLER_54_1887 ();
 sg13g2_decap_8 FILLER_54_1898 ();
 sg13g2_fill_1 FILLER_54_1905 ();
 sg13g2_decap_4 FILLER_54_1911 ();
 sg13g2_fill_1 FILLER_54_1915 ();
 sg13g2_decap_8 FILLER_54_1921 ();
 sg13g2_fill_1 FILLER_54_1928 ();
 sg13g2_decap_8 FILLER_54_1935 ();
 sg13g2_fill_2 FILLER_54_1951 ();
 sg13g2_fill_1 FILLER_54_1953 ();
 sg13g2_fill_1 FILLER_54_1967 ();
 sg13g2_decap_4 FILLER_54_1973 ();
 sg13g2_fill_2 FILLER_54_1977 ();
 sg13g2_decap_8 FILLER_54_1988 ();
 sg13g2_fill_2 FILLER_54_1995 ();
 sg13g2_decap_4 FILLER_54_2014 ();
 sg13g2_fill_1 FILLER_54_2022 ();
 sg13g2_fill_2 FILLER_54_2028 ();
 sg13g2_fill_2 FILLER_54_2086 ();
 sg13g2_decap_8 FILLER_54_2105 ();
 sg13g2_fill_2 FILLER_54_2112 ();
 sg13g2_decap_4 FILLER_54_2118 ();
 sg13g2_decap_4 FILLER_54_2126 ();
 sg13g2_fill_2 FILLER_54_2130 ();
 sg13g2_decap_8 FILLER_54_2202 ();
 sg13g2_decap_4 FILLER_54_2209 ();
 sg13g2_fill_2 FILLER_54_2213 ();
 sg13g2_fill_2 FILLER_54_2227 ();
 sg13g2_fill_1 FILLER_54_2229 ();
 sg13g2_decap_4 FILLER_54_2291 ();
 sg13g2_decap_8 FILLER_54_2325 ();
 sg13g2_decap_8 FILLER_54_2332 ();
 sg13g2_decap_8 FILLER_54_2339 ();
 sg13g2_fill_1 FILLER_54_2346 ();
 sg13g2_fill_1 FILLER_54_2359 ();
 sg13g2_decap_8 FILLER_54_2368 ();
 sg13g2_fill_2 FILLER_54_2375 ();
 sg13g2_fill_1 FILLER_54_2377 ();
 sg13g2_decap_4 FILLER_54_2403 ();
 sg13g2_fill_2 FILLER_54_2407 ();
 sg13g2_fill_1 FILLER_54_2444 ();
 sg13g2_fill_1 FILLER_54_2471 ();
 sg13g2_fill_1 FILLER_54_2537 ();
 sg13g2_fill_1 FILLER_54_2543 ();
 sg13g2_fill_2 FILLER_54_2549 ();
 sg13g2_fill_2 FILLER_54_2557 ();
 sg13g2_fill_1 FILLER_54_2615 ();
 sg13g2_fill_2 FILLER_54_2667 ();
 sg13g2_fill_1 FILLER_54_2669 ();
 sg13g2_decap_4 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_4 ();
 sg13g2_decap_4 FILLER_55_31 ();
 sg13g2_fill_2 FILLER_55_35 ();
 sg13g2_fill_1 FILLER_55_47 ();
 sg13g2_fill_1 FILLER_55_52 ();
 sg13g2_fill_2 FILLER_55_101 ();
 sg13g2_fill_1 FILLER_55_103 ();
 sg13g2_fill_2 FILLER_55_122 ();
 sg13g2_fill_2 FILLER_55_129 ();
 sg13g2_fill_2 FILLER_55_135 ();
 sg13g2_decap_4 FILLER_55_146 ();
 sg13g2_fill_1 FILLER_55_233 ();
 sg13g2_decap_4 FILLER_55_260 ();
 sg13g2_fill_2 FILLER_55_286 ();
 sg13g2_fill_1 FILLER_55_299 ();
 sg13g2_fill_1 FILLER_55_338 ();
 sg13g2_fill_1 FILLER_55_374 ();
 sg13g2_fill_2 FILLER_55_399 ();
 sg13g2_fill_1 FILLER_55_422 ();
 sg13g2_fill_1 FILLER_55_434 ();
 sg13g2_fill_1 FILLER_55_445 ();
 sg13g2_decap_4 FILLER_55_479 ();
 sg13g2_decap_4 FILLER_55_502 ();
 sg13g2_fill_2 FILLER_55_506 ();
 sg13g2_decap_8 FILLER_55_513 ();
 sg13g2_fill_2 FILLER_55_520 ();
 sg13g2_fill_2 FILLER_55_528 ();
 sg13g2_decap_8 FILLER_55_554 ();
 sg13g2_fill_1 FILLER_55_575 ();
 sg13g2_decap_4 FILLER_55_602 ();
 sg13g2_fill_1 FILLER_55_634 ();
 sg13g2_fill_1 FILLER_55_641 ();
 sg13g2_fill_1 FILLER_55_655 ();
 sg13g2_fill_2 FILLER_55_673 ();
 sg13g2_fill_2 FILLER_55_684 ();
 sg13g2_fill_2 FILLER_55_711 ();
 sg13g2_fill_2 FILLER_55_718 ();
 sg13g2_fill_1 FILLER_55_724 ();
 sg13g2_decap_4 FILLER_55_734 ();
 sg13g2_fill_2 FILLER_55_738 ();
 sg13g2_decap_8 FILLER_55_748 ();
 sg13g2_decap_4 FILLER_55_755 ();
 sg13g2_fill_2 FILLER_55_759 ();
 sg13g2_fill_2 FILLER_55_766 ();
 sg13g2_fill_1 FILLER_55_768 ();
 sg13g2_decap_8 FILLER_55_777 ();
 sg13g2_decap_4 FILLER_55_784 ();
 sg13g2_fill_2 FILLER_55_793 ();
 sg13g2_decap_8 FILLER_55_807 ();
 sg13g2_decap_4 FILLER_55_814 ();
 sg13g2_fill_1 FILLER_55_826 ();
 sg13g2_fill_1 FILLER_55_832 ();
 sg13g2_fill_2 FILLER_55_838 ();
 sg13g2_fill_2 FILLER_55_877 ();
 sg13g2_fill_2 FILLER_55_892 ();
 sg13g2_decap_8 FILLER_55_899 ();
 sg13g2_decap_4 FILLER_55_906 ();
 sg13g2_fill_1 FILLER_55_910 ();
 sg13g2_fill_1 FILLER_55_928 ();
 sg13g2_fill_1 FILLER_55_934 ();
 sg13g2_fill_1 FILLER_55_940 ();
 sg13g2_fill_1 FILLER_55_969 ();
 sg13g2_fill_1 FILLER_55_984 ();
 sg13g2_fill_1 FILLER_55_1010 ();
 sg13g2_fill_2 FILLER_55_1019 ();
 sg13g2_fill_1 FILLER_55_1021 ();
 sg13g2_decap_4 FILLER_55_1026 ();
 sg13g2_fill_1 FILLER_55_1034 ();
 sg13g2_decap_4 FILLER_55_1052 ();
 sg13g2_fill_2 FILLER_55_1117 ();
 sg13g2_fill_1 FILLER_55_1137 ();
 sg13g2_fill_1 FILLER_55_1142 ();
 sg13g2_decap_8 FILLER_55_1175 ();
 sg13g2_fill_2 FILLER_55_1182 ();
 sg13g2_decap_4 FILLER_55_1214 ();
 sg13g2_fill_1 FILLER_55_1228 ();
 sg13g2_fill_1 FILLER_55_1258 ();
 sg13g2_fill_2 FILLER_55_1263 ();
 sg13g2_fill_2 FILLER_55_1280 ();
 sg13g2_fill_1 FILLER_55_1291 ();
 sg13g2_fill_2 FILLER_55_1299 ();
 sg13g2_fill_2 FILLER_55_1311 ();
 sg13g2_fill_2 FILLER_55_1323 ();
 sg13g2_decap_8 FILLER_55_1350 ();
 sg13g2_decap_8 FILLER_55_1357 ();
 sg13g2_decap_4 FILLER_55_1364 ();
 sg13g2_fill_2 FILLER_55_1368 ();
 sg13g2_fill_2 FILLER_55_1395 ();
 sg13g2_decap_8 FILLER_55_1403 ();
 sg13g2_fill_1 FILLER_55_1410 ();
 sg13g2_decap_4 FILLER_55_1415 ();
 sg13g2_fill_2 FILLER_55_1434 ();
 sg13g2_fill_1 FILLER_55_1436 ();
 sg13g2_fill_2 FILLER_55_1504 ();
 sg13g2_fill_1 FILLER_55_1506 ();
 sg13g2_fill_2 FILLER_55_1517 ();
 sg13g2_fill_1 FILLER_55_1519 ();
 sg13g2_fill_1 FILLER_55_1556 ();
 sg13g2_fill_2 FILLER_55_1583 ();
 sg13g2_fill_1 FILLER_55_1611 ();
 sg13g2_decap_8 FILLER_55_1646 ();
 sg13g2_decap_4 FILLER_55_1653 ();
 sg13g2_fill_2 FILLER_55_1657 ();
 sg13g2_decap_4 FILLER_55_1664 ();
 sg13g2_decap_4 FILLER_55_1678 ();
 sg13g2_fill_2 FILLER_55_1690 ();
 sg13g2_decap_8 FILLER_55_1696 ();
 sg13g2_fill_2 FILLER_55_1703 ();
 sg13g2_fill_2 FILLER_55_1708 ();
 sg13g2_fill_1 FILLER_55_1715 ();
 sg13g2_fill_1 FILLER_55_1720 ();
 sg13g2_fill_1 FILLER_55_1726 ();
 sg13g2_fill_2 FILLER_55_1731 ();
 sg13g2_fill_2 FILLER_55_1743 ();
 sg13g2_fill_1 FILLER_55_1773 ();
 sg13g2_fill_2 FILLER_55_1814 ();
 sg13g2_fill_1 FILLER_55_1826 ();
 sg13g2_decap_8 FILLER_55_1837 ();
 sg13g2_fill_2 FILLER_55_1844 ();
 sg13g2_fill_1 FILLER_55_1846 ();
 sg13g2_fill_2 FILLER_55_1870 ();
 sg13g2_fill_1 FILLER_55_1872 ();
 sg13g2_fill_2 FILLER_55_1908 ();
 sg13g2_fill_1 FILLER_55_1910 ();
 sg13g2_decap_4 FILLER_55_1915 ();
 sg13g2_fill_1 FILLER_55_1924 ();
 sg13g2_fill_1 FILLER_55_1931 ();
 sg13g2_fill_2 FILLER_55_1940 ();
 sg13g2_decap_8 FILLER_55_1973 ();
 sg13g2_decap_8 FILLER_55_1980 ();
 sg13g2_decap_4 FILLER_55_1987 ();
 sg13g2_fill_1 FILLER_55_2036 ();
 sg13g2_fill_1 FILLER_55_2051 ();
 sg13g2_fill_2 FILLER_55_2069 ();
 sg13g2_fill_1 FILLER_55_2071 ();
 sg13g2_fill_1 FILLER_55_2081 ();
 sg13g2_fill_1 FILLER_55_2095 ();
 sg13g2_fill_2 FILLER_55_2105 ();
 sg13g2_fill_1 FILLER_55_2107 ();
 sg13g2_fill_1 FILLER_55_2117 ();
 sg13g2_decap_8 FILLER_55_2127 ();
 sg13g2_fill_2 FILLER_55_2134 ();
 sg13g2_fill_1 FILLER_55_2136 ();
 sg13g2_decap_4 FILLER_55_2142 ();
 sg13g2_fill_1 FILLER_55_2154 ();
 sg13g2_fill_1 FILLER_55_2160 ();
 sg13g2_fill_2 FILLER_55_2171 ();
 sg13g2_decap_8 FILLER_55_2204 ();
 sg13g2_fill_1 FILLER_55_2211 ();
 sg13g2_fill_2 FILLER_55_2238 ();
 sg13g2_fill_1 FILLER_55_2253 ();
 sg13g2_fill_1 FILLER_55_2268 ();
 sg13g2_fill_1 FILLER_55_2274 ();
 sg13g2_fill_1 FILLER_55_2284 ();
 sg13g2_fill_2 FILLER_55_2295 ();
 sg13g2_fill_1 FILLER_55_2297 ();
 sg13g2_decap_8 FILLER_55_2324 ();
 sg13g2_decap_8 FILLER_55_2331 ();
 sg13g2_decap_8 FILLER_55_2338 ();
 sg13g2_fill_2 FILLER_55_2345 ();
 sg13g2_fill_1 FILLER_55_2347 ();
 sg13g2_decap_8 FILLER_55_2378 ();
 sg13g2_decap_8 FILLER_55_2385 ();
 sg13g2_decap_8 FILLER_55_2392 ();
 sg13g2_decap_4 FILLER_55_2399 ();
 sg13g2_fill_1 FILLER_55_2403 ();
 sg13g2_fill_2 FILLER_55_2408 ();
 sg13g2_fill_1 FILLER_55_2410 ();
 sg13g2_decap_4 FILLER_55_2416 ();
 sg13g2_fill_2 FILLER_55_2420 ();
 sg13g2_fill_1 FILLER_55_2426 ();
 sg13g2_fill_2 FILLER_55_2446 ();
 sg13g2_decap_8 FILLER_55_2452 ();
 sg13g2_decap_8 FILLER_55_2459 ();
 sg13g2_fill_1 FILLER_55_2466 ();
 sg13g2_fill_2 FILLER_55_2485 ();
 sg13g2_decap_4 FILLER_55_2493 ();
 sg13g2_fill_2 FILLER_55_2567 ();
 sg13g2_fill_1 FILLER_55_2569 ();
 sg13g2_fill_2 FILLER_55_2574 ();
 sg13g2_fill_2 FILLER_55_2580 ();
 sg13g2_fill_1 FILLER_55_2582 ();
 sg13g2_fill_1 FILLER_55_2587 ();
 sg13g2_fill_2 FILLER_55_2627 ();
 sg13g2_decap_4 FILLER_56_0 ();
 sg13g2_decap_4 FILLER_56_30 ();
 sg13g2_fill_2 FILLER_56_34 ();
 sg13g2_decap_4 FILLER_56_62 ();
 sg13g2_decap_8 FILLER_56_74 ();
 sg13g2_decap_4 FILLER_56_81 ();
 sg13g2_fill_1 FILLER_56_85 ();
 sg13g2_decap_8 FILLER_56_95 ();
 sg13g2_decap_8 FILLER_56_102 ();
 sg13g2_fill_2 FILLER_56_118 ();
 sg13g2_fill_1 FILLER_56_120 ();
 sg13g2_fill_1 FILLER_56_141 ();
 sg13g2_fill_2 FILLER_56_153 ();
 sg13g2_fill_1 FILLER_56_170 ();
 sg13g2_fill_2 FILLER_56_190 ();
 sg13g2_fill_2 FILLER_56_206 ();
 sg13g2_fill_1 FILLER_56_212 ();
 sg13g2_decap_4 FILLER_56_217 ();
 sg13g2_fill_2 FILLER_56_221 ();
 sg13g2_fill_2 FILLER_56_267 ();
 sg13g2_fill_2 FILLER_56_297 ();
 sg13g2_fill_2 FILLER_56_338 ();
 sg13g2_fill_2 FILLER_56_349 ();
 sg13g2_fill_2 FILLER_56_381 ();
 sg13g2_fill_1 FILLER_56_400 ();
 sg13g2_fill_2 FILLER_56_414 ();
 sg13g2_fill_1 FILLER_56_442 ();
 sg13g2_fill_1 FILLER_56_448 ();
 sg13g2_decap_4 FILLER_56_460 ();
 sg13g2_decap_8 FILLER_56_478 ();
 sg13g2_decap_8 FILLER_56_485 ();
 sg13g2_decap_8 FILLER_56_492 ();
 sg13g2_decap_4 FILLER_56_499 ();
 sg13g2_fill_1 FILLER_56_503 ();
 sg13g2_fill_2 FILLER_56_517 ();
 sg13g2_fill_1 FILLER_56_519 ();
 sg13g2_fill_1 FILLER_56_530 ();
 sg13g2_fill_1 FILLER_56_535 ();
 sg13g2_decap_8 FILLER_56_541 ();
 sg13g2_decap_8 FILLER_56_548 ();
 sg13g2_decap_8 FILLER_56_555 ();
 sg13g2_decap_4 FILLER_56_562 ();
 sg13g2_fill_1 FILLER_56_566 ();
 sg13g2_decap_4 FILLER_56_577 ();
 sg13g2_fill_2 FILLER_56_581 ();
 sg13g2_fill_2 FILLER_56_591 ();
 sg13g2_decap_4 FILLER_56_625 ();
 sg13g2_fill_1 FILLER_56_629 ();
 sg13g2_fill_1 FILLER_56_644 ();
 sg13g2_fill_2 FILLER_56_650 ();
 sg13g2_fill_2 FILLER_56_657 ();
 sg13g2_fill_2 FILLER_56_663 ();
 sg13g2_fill_2 FILLER_56_674 ();
 sg13g2_fill_1 FILLER_56_676 ();
 sg13g2_decap_8 FILLER_56_713 ();
 sg13g2_fill_2 FILLER_56_720 ();
 sg13g2_fill_1 FILLER_56_722 ();
 sg13g2_fill_2 FILLER_56_753 ();
 sg13g2_fill_1 FILLER_56_755 ();
 sg13g2_fill_1 FILLER_56_830 ();
 sg13g2_fill_1 FILLER_56_841 ();
 sg13g2_fill_2 FILLER_56_858 ();
 sg13g2_fill_1 FILLER_56_877 ();
 sg13g2_decap_4 FILLER_56_903 ();
 sg13g2_fill_2 FILLER_56_911 ();
 sg13g2_fill_1 FILLER_56_913 ();
 sg13g2_decap_8 FILLER_56_918 ();
 sg13g2_decap_4 FILLER_56_925 ();
 sg13g2_decap_8 FILLER_56_934 ();
 sg13g2_fill_1 FILLER_56_948 ();
 sg13g2_fill_2 FILLER_56_969 ();
 sg13g2_fill_1 FILLER_56_975 ();
 sg13g2_decap_8 FILLER_56_994 ();
 sg13g2_fill_1 FILLER_56_1010 ();
 sg13g2_decap_8 FILLER_56_1015 ();
 sg13g2_decap_4 FILLER_56_1022 ();
 sg13g2_decap_8 FILLER_56_1031 ();
 sg13g2_decap_4 FILLER_56_1038 ();
 sg13g2_decap_8 FILLER_56_1045 ();
 sg13g2_decap_4 FILLER_56_1052 ();
 sg13g2_fill_1 FILLER_56_1056 ();
 sg13g2_fill_1 FILLER_56_1064 ();
 sg13g2_decap_4 FILLER_56_1085 ();
 sg13g2_fill_1 FILLER_56_1119 ();
 sg13g2_decap_4 FILLER_56_1156 ();
 sg13g2_fill_1 FILLER_56_1190 ();
 sg13g2_decap_8 FILLER_56_1199 ();
 sg13g2_decap_4 FILLER_56_1206 ();
 sg13g2_fill_1 FILLER_56_1210 ();
 sg13g2_fill_1 FILLER_56_1215 ();
 sg13g2_fill_1 FILLER_56_1252 ();
 sg13g2_decap_4 FILLER_56_1263 ();
 sg13g2_fill_2 FILLER_56_1296 ();
 sg13g2_fill_1 FILLER_56_1308 ();
 sg13g2_fill_2 FILLER_56_1315 ();
 sg13g2_fill_1 FILLER_56_1317 ();
 sg13g2_fill_1 FILLER_56_1332 ();
 sg13g2_fill_2 FILLER_56_1338 ();
 sg13g2_decap_8 FILLER_56_1346 ();
 sg13g2_fill_2 FILLER_56_1353 ();
 sg13g2_decap_8 FILLER_56_1361 ();
 sg13g2_decap_4 FILLER_56_1391 ();
 sg13g2_fill_1 FILLER_56_1395 ();
 sg13g2_fill_1 FILLER_56_1405 ();
 sg13g2_decap_4 FILLER_56_1418 ();
 sg13g2_fill_2 FILLER_56_1422 ();
 sg13g2_fill_2 FILLER_56_1446 ();
 sg13g2_fill_2 FILLER_56_1452 ();
 sg13g2_decap_8 FILLER_56_1465 ();
 sg13g2_decap_4 FILLER_56_1472 ();
 sg13g2_fill_1 FILLER_56_1476 ();
 sg13g2_decap_8 FILLER_56_1487 ();
 sg13g2_decap_4 FILLER_56_1494 ();
 sg13g2_fill_1 FILLER_56_1498 ();
 sg13g2_fill_2 FILLER_56_1544 ();
 sg13g2_fill_2 FILLER_56_1574 ();
 sg13g2_fill_1 FILLER_56_1576 ();
 sg13g2_fill_2 FILLER_56_1608 ();
 sg13g2_fill_2 FILLER_56_1659 ();
 sg13g2_fill_1 FILLER_56_1661 ();
 sg13g2_fill_2 FILLER_56_1744 ();
 sg13g2_fill_1 FILLER_56_1746 ();
 sg13g2_fill_2 FILLER_56_1752 ();
 sg13g2_fill_1 FILLER_56_1754 ();
 sg13g2_fill_1 FILLER_56_1763 ();
 sg13g2_decap_4 FILLER_56_1775 ();
 sg13g2_fill_2 FILLER_56_1779 ();
 sg13g2_decap_4 FILLER_56_1826 ();
 sg13g2_fill_1 FILLER_56_1838 ();
 sg13g2_fill_1 FILLER_56_1843 ();
 sg13g2_decap_4 FILLER_56_1857 ();
 sg13g2_fill_1 FILLER_56_1870 ();
 sg13g2_decap_4 FILLER_56_1907 ();
 sg13g2_fill_2 FILLER_56_1915 ();
 sg13g2_decap_4 FILLER_56_1945 ();
 sg13g2_fill_1 FILLER_56_1949 ();
 sg13g2_decap_8 FILLER_56_1958 ();
 sg13g2_decap_8 FILLER_56_1965 ();
 sg13g2_decap_8 FILLER_56_1972 ();
 sg13g2_decap_8 FILLER_56_1979 ();
 sg13g2_fill_2 FILLER_56_1991 ();
 sg13g2_fill_1 FILLER_56_1993 ();
 sg13g2_fill_1 FILLER_56_2026 ();
 sg13g2_fill_1 FILLER_56_2031 ();
 sg13g2_fill_1 FILLER_56_2045 ();
 sg13g2_fill_2 FILLER_56_2052 ();
 sg13g2_fill_1 FILLER_56_2054 ();
 sg13g2_fill_1 FILLER_56_2060 ();
 sg13g2_fill_1 FILLER_56_2075 ();
 sg13g2_fill_1 FILLER_56_2084 ();
 sg13g2_fill_1 FILLER_56_2090 ();
 sg13g2_fill_2 FILLER_56_2110 ();
 sg13g2_fill_1 FILLER_56_2112 ();
 sg13g2_decap_8 FILLER_56_2123 ();
 sg13g2_decap_8 FILLER_56_2130 ();
 sg13g2_decap_8 FILLER_56_2137 ();
 sg13g2_decap_8 FILLER_56_2144 ();
 sg13g2_decap_4 FILLER_56_2151 ();
 sg13g2_fill_1 FILLER_56_2155 ();
 sg13g2_fill_2 FILLER_56_2166 ();
 sg13g2_fill_1 FILLER_56_2168 ();
 sg13g2_decap_8 FILLER_56_2208 ();
 sg13g2_decap_8 FILLER_56_2215 ();
 sg13g2_fill_2 FILLER_56_2222 ();
 sg13g2_fill_1 FILLER_56_2232 ();
 sg13g2_fill_1 FILLER_56_2237 ();
 sg13g2_fill_1 FILLER_56_2242 ();
 sg13g2_fill_2 FILLER_56_2247 ();
 sg13g2_fill_2 FILLER_56_2262 ();
 sg13g2_decap_4 FILLER_56_2334 ();
 sg13g2_decap_8 FILLER_56_2369 ();
 sg13g2_decap_8 FILLER_56_2376 ();
 sg13g2_decap_8 FILLER_56_2383 ();
 sg13g2_decap_8 FILLER_56_2390 ();
 sg13g2_decap_4 FILLER_56_2397 ();
 sg13g2_fill_1 FILLER_56_2431 ();
 sg13g2_fill_2 FILLER_56_2440 ();
 sg13g2_decap_4 FILLER_56_2446 ();
 sg13g2_decap_8 FILLER_56_2459 ();
 sg13g2_decap_8 FILLER_56_2466 ();
 sg13g2_decap_8 FILLER_56_2473 ();
 sg13g2_decap_8 FILLER_56_2480 ();
 sg13g2_decap_4 FILLER_56_2487 ();
 sg13g2_fill_2 FILLER_56_2491 ();
 sg13g2_decap_4 FILLER_56_2503 ();
 sg13g2_fill_2 FILLER_56_2511 ();
 sg13g2_fill_1 FILLER_56_2549 ();
 sg13g2_fill_2 FILLER_56_2586 ();
 sg13g2_fill_1 FILLER_56_2588 ();
 sg13g2_fill_1 FILLER_56_2607 ();
 sg13g2_fill_2 FILLER_56_2629 ();
 sg13g2_fill_1 FILLER_56_2644 ();
 sg13g2_decap_8 FILLER_56_2663 ();
 sg13g2_fill_2 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_2 ();
 sg13g2_fill_2 FILLER_57_33 ();
 sg13g2_decap_4 FILLER_57_39 ();
 sg13g2_fill_2 FILLER_57_43 ();
 sg13g2_fill_2 FILLER_57_49 ();
 sg13g2_fill_2 FILLER_57_55 ();
 sg13g2_fill_1 FILLER_57_57 ();
 sg13g2_decap_8 FILLER_57_62 ();
 sg13g2_decap_4 FILLER_57_69 ();
 sg13g2_fill_1 FILLER_57_73 ();
 sg13g2_decap_4 FILLER_57_88 ();
 sg13g2_decap_4 FILLER_57_126 ();
 sg13g2_fill_1 FILLER_57_130 ();
 sg13g2_fill_1 FILLER_57_180 ();
 sg13g2_fill_2 FILLER_57_213 ();
 sg13g2_fill_2 FILLER_57_241 ();
 sg13g2_fill_1 FILLER_57_243 ();
 sg13g2_decap_8 FILLER_57_248 ();
 sg13g2_fill_2 FILLER_57_255 ();
 sg13g2_fill_1 FILLER_57_257 ();
 sg13g2_fill_1 FILLER_57_277 ();
 sg13g2_fill_1 FILLER_57_292 ();
 sg13g2_fill_2 FILLER_57_302 ();
 sg13g2_fill_2 FILLER_57_317 ();
 sg13g2_fill_2 FILLER_57_322 ();
 sg13g2_fill_1 FILLER_57_400 ();
 sg13g2_fill_2 FILLER_57_442 ();
 sg13g2_fill_1 FILLER_57_475 ();
 sg13g2_fill_1 FILLER_57_481 ();
 sg13g2_fill_2 FILLER_57_492 ();
 sg13g2_fill_1 FILLER_57_494 ();
 sg13g2_fill_1 FILLER_57_549 ();
 sg13g2_decap_4 FILLER_57_566 ();
 sg13g2_fill_2 FILLER_57_570 ();
 sg13g2_decap_8 FILLER_57_578 ();
 sg13g2_fill_1 FILLER_57_585 ();
 sg13g2_fill_1 FILLER_57_590 ();
 sg13g2_fill_2 FILLER_57_596 ();
 sg13g2_fill_2 FILLER_57_602 ();
 sg13g2_fill_2 FILLER_57_614 ();
 sg13g2_fill_2 FILLER_57_642 ();
 sg13g2_fill_1 FILLER_57_644 ();
 sg13g2_decap_8 FILLER_57_648 ();
 sg13g2_decap_8 FILLER_57_655 ();
 sg13g2_fill_1 FILLER_57_673 ();
 sg13g2_fill_1 FILLER_57_682 ();
 sg13g2_fill_1 FILLER_57_711 ();
 sg13g2_fill_1 FILLER_57_717 ();
 sg13g2_fill_2 FILLER_57_722 ();
 sg13g2_fill_1 FILLER_57_728 ();
 sg13g2_decap_4 FILLER_57_755 ();
 sg13g2_fill_1 FILLER_57_766 ();
 sg13g2_fill_2 FILLER_57_806 ();
 sg13g2_decap_8 FILLER_57_812 ();
 sg13g2_fill_2 FILLER_57_819 ();
 sg13g2_decap_8 FILLER_57_829 ();
 sg13g2_fill_2 FILLER_57_836 ();
 sg13g2_fill_1 FILLER_57_851 ();
 sg13g2_fill_1 FILLER_57_863 ();
 sg13g2_fill_1 FILLER_57_872 ();
 sg13g2_fill_2 FILLER_57_882 ();
 sg13g2_decap_4 FILLER_57_931 ();
 sg13g2_fill_1 FILLER_57_935 ();
 sg13g2_fill_2 FILLER_57_962 ();
 sg13g2_fill_1 FILLER_57_977 ();
 sg13g2_fill_1 FILLER_57_1042 ();
 sg13g2_fill_2 FILLER_57_1048 ();
 sg13g2_fill_1 FILLER_57_1074 ();
 sg13g2_decap_8 FILLER_57_1111 ();
 sg13g2_fill_2 FILLER_57_1118 ();
 sg13g2_fill_1 FILLER_57_1123 ();
 sg13g2_fill_2 FILLER_57_1155 ();
 sg13g2_fill_1 FILLER_57_1157 ();
 sg13g2_decap_8 FILLER_57_1184 ();
 sg13g2_decap_8 FILLER_57_1191 ();
 sg13g2_decap_4 FILLER_57_1198 ();
 sg13g2_fill_2 FILLER_57_1202 ();
 sg13g2_fill_2 FILLER_57_1240 ();
 sg13g2_fill_1 FILLER_57_1246 ();
 sg13g2_fill_1 FILLER_57_1273 ();
 sg13g2_fill_1 FILLER_57_1324 ();
 sg13g2_decap_8 FILLER_57_1343 ();
 sg13g2_decap_8 FILLER_57_1350 ();
 sg13g2_decap_8 FILLER_57_1357 ();
 sg13g2_fill_1 FILLER_57_1364 ();
 sg13g2_decap_8 FILLER_57_1371 ();
 sg13g2_decap_8 FILLER_57_1378 ();
 sg13g2_decap_4 FILLER_57_1385 ();
 sg13g2_fill_2 FILLER_57_1389 ();
 sg13g2_decap_8 FILLER_57_1395 ();
 sg13g2_decap_8 FILLER_57_1402 ();
 sg13g2_decap_4 FILLER_57_1409 ();
 sg13g2_fill_1 FILLER_57_1413 ();
 sg13g2_fill_2 FILLER_57_1418 ();
 sg13g2_fill_1 FILLER_57_1420 ();
 sg13g2_fill_2 FILLER_57_1434 ();
 sg13g2_decap_8 FILLER_57_1459 ();
 sg13g2_fill_1 FILLER_57_1466 ();
 sg13g2_fill_1 FILLER_57_1473 ();
 sg13g2_fill_1 FILLER_57_1484 ();
 sg13g2_decap_8 FILLER_57_1511 ();
 sg13g2_fill_2 FILLER_57_1518 ();
 sg13g2_fill_1 FILLER_57_1520 ();
 sg13g2_decap_4 FILLER_57_1525 ();
 sg13g2_fill_1 FILLER_57_1529 ();
 sg13g2_decap_8 FILLER_57_1570 ();
 sg13g2_decap_8 FILLER_57_1577 ();
 sg13g2_fill_2 FILLER_57_1584 ();
 sg13g2_decap_8 FILLER_57_1590 ();
 sg13g2_decap_4 FILLER_57_1597 ();
 sg13g2_fill_1 FILLER_57_1621 ();
 sg13g2_fill_1 FILLER_57_1627 ();
 sg13g2_fill_1 FILLER_57_1633 ();
 sg13g2_fill_1 FILLER_57_1638 ();
 sg13g2_fill_2 FILLER_57_1647 ();
 sg13g2_fill_2 FILLER_57_1657 ();
 sg13g2_fill_2 FILLER_57_1663 ();
 sg13g2_fill_1 FILLER_57_1665 ();
 sg13g2_fill_1 FILLER_57_1677 ();
 sg13g2_fill_1 FILLER_57_1683 ();
 sg13g2_fill_2 FILLER_57_1693 ();
 sg13g2_fill_1 FILLER_57_1695 ();
 sg13g2_decap_4 FILLER_57_1700 ();
 sg13g2_fill_1 FILLER_57_1704 ();
 sg13g2_decap_4 FILLER_57_1710 ();
 sg13g2_fill_1 FILLER_57_1714 ();
 sg13g2_decap_8 FILLER_57_1718 ();
 sg13g2_decap_4 FILLER_57_1725 ();
 sg13g2_fill_1 FILLER_57_1729 ();
 sg13g2_decap_4 FILLER_57_1734 ();
 sg13g2_fill_2 FILLER_57_1738 ();
 sg13g2_fill_2 FILLER_57_1744 ();
 sg13g2_fill_1 FILLER_57_1746 ();
 sg13g2_decap_8 FILLER_57_1751 ();
 sg13g2_decap_8 FILLER_57_1758 ();
 sg13g2_fill_2 FILLER_57_1765 ();
 sg13g2_decap_4 FILLER_57_1771 ();
 sg13g2_fill_2 FILLER_57_1794 ();
 sg13g2_fill_1 FILLER_57_1796 ();
 sg13g2_fill_2 FILLER_57_1817 ();
 sg13g2_fill_1 FILLER_57_1824 ();
 sg13g2_decap_4 FILLER_57_1835 ();
 sg13g2_fill_1 FILLER_57_1839 ();
 sg13g2_decap_4 FILLER_57_1845 ();
 sg13g2_decap_4 FILLER_57_1861 ();
 sg13g2_decap_4 FILLER_57_1869 ();
 sg13g2_fill_1 FILLER_57_1916 ();
 sg13g2_fill_1 FILLER_57_1944 ();
 sg13g2_decap_8 FILLER_57_1950 ();
 sg13g2_decap_4 FILLER_57_1957 ();
 sg13g2_fill_1 FILLER_57_1961 ();
 sg13g2_decap_8 FILLER_57_1967 ();
 sg13g2_fill_1 FILLER_57_1974 ();
 sg13g2_decap_8 FILLER_57_1984 ();
 sg13g2_decap_8 FILLER_57_1991 ();
 sg13g2_decap_4 FILLER_57_1998 ();
 sg13g2_fill_1 FILLER_57_2002 ();
 sg13g2_decap_4 FILLER_57_2007 ();
 sg13g2_fill_1 FILLER_57_2032 ();
 sg13g2_fill_1 FILLER_57_2060 ();
 sg13g2_fill_1 FILLER_57_2065 ();
 sg13g2_fill_1 FILLER_57_2076 ();
 sg13g2_fill_1 FILLER_57_2083 ();
 sg13g2_fill_1 FILLER_57_2090 ();
 sg13g2_fill_1 FILLER_57_2096 ();
 sg13g2_fill_2 FILLER_57_2111 ();
 sg13g2_decap_8 FILLER_57_2126 ();
 sg13g2_decap_8 FILLER_57_2133 ();
 sg13g2_fill_2 FILLER_57_2140 ();
 sg13g2_decap_8 FILLER_57_2146 ();
 sg13g2_decap_8 FILLER_57_2153 ();
 sg13g2_decap_4 FILLER_57_2160 ();
 sg13g2_fill_1 FILLER_57_2164 ();
 sg13g2_decap_8 FILLER_57_2201 ();
 sg13g2_decap_4 FILLER_57_2208 ();
 sg13g2_fill_1 FILLER_57_2212 ();
 sg13g2_fill_1 FILLER_57_2226 ();
 sg13g2_decap_8 FILLER_57_2277 ();
 sg13g2_decap_8 FILLER_57_2284 ();
 sg13g2_decap_8 FILLER_57_2291 ();
 sg13g2_fill_2 FILLER_57_2298 ();
 sg13g2_fill_1 FILLER_57_2326 ();
 sg13g2_fill_1 FILLER_57_2374 ();
 sg13g2_fill_1 FILLER_57_2406 ();
 sg13g2_decap_4 FILLER_57_2420 ();
 sg13g2_fill_2 FILLER_57_2424 ();
 sg13g2_fill_1 FILLER_57_2434 ();
 sg13g2_fill_2 FILLER_57_2439 ();
 sg13g2_fill_2 FILLER_57_2467 ();
 sg13g2_decap_4 FILLER_57_2478 ();
 sg13g2_decap_8 FILLER_57_2486 ();
 sg13g2_decap_8 FILLER_57_2493 ();
 sg13g2_decap_8 FILLER_57_2500 ();
 sg13g2_decap_8 FILLER_57_2507 ();
 sg13g2_decap_8 FILLER_57_2514 ();
 sg13g2_fill_2 FILLER_57_2525 ();
 sg13g2_fill_1 FILLER_57_2527 ();
 sg13g2_fill_2 FILLER_57_2532 ();
 sg13g2_fill_1 FILLER_57_2534 ();
 sg13g2_fill_2 FILLER_57_2539 ();
 sg13g2_decap_8 FILLER_57_2545 ();
 sg13g2_decap_4 FILLER_57_2552 ();
 sg13g2_fill_1 FILLER_57_2556 ();
 sg13g2_fill_2 FILLER_57_2593 ();
 sg13g2_fill_1 FILLER_57_2595 ();
 sg13g2_fill_1 FILLER_57_2630 ();
 sg13g2_fill_1 FILLER_57_2634 ();
 sg13g2_fill_2 FILLER_57_2668 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_fill_2 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_17 ();
 sg13g2_decap_8 FILLER_58_24 ();
 sg13g2_decap_8 FILLER_58_31 ();
 sg13g2_decap_8 FILLER_58_38 ();
 sg13g2_decap_4 FILLER_58_45 ();
 sg13g2_fill_2 FILLER_58_49 ();
 sg13g2_fill_2 FILLER_58_66 ();
 sg13g2_fill_1 FILLER_58_68 ();
 sg13g2_decap_4 FILLER_58_74 ();
 sg13g2_fill_1 FILLER_58_78 ();
 sg13g2_fill_2 FILLER_58_105 ();
 sg13g2_decap_4 FILLER_58_116 ();
 sg13g2_fill_2 FILLER_58_130 ();
 sg13g2_fill_1 FILLER_58_132 ();
 sg13g2_fill_1 FILLER_58_171 ();
 sg13g2_fill_2 FILLER_58_176 ();
 sg13g2_fill_2 FILLER_58_185 ();
 sg13g2_fill_1 FILLER_58_201 ();
 sg13g2_fill_2 FILLER_58_213 ();
 sg13g2_decap_8 FILLER_58_245 ();
 sg13g2_fill_2 FILLER_58_252 ();
 sg13g2_fill_1 FILLER_58_292 ();
 sg13g2_fill_1 FILLER_58_381 ();
 sg13g2_fill_2 FILLER_58_430 ();
 sg13g2_fill_1 FILLER_58_440 ();
 sg13g2_fill_1 FILLER_58_448 ();
 sg13g2_fill_2 FILLER_58_464 ();
 sg13g2_fill_1 FILLER_58_496 ();
 sg13g2_decap_4 FILLER_58_615 ();
 sg13g2_fill_2 FILLER_58_619 ();
 sg13g2_decap_4 FILLER_58_625 ();
 sg13g2_fill_2 FILLER_58_629 ();
 sg13g2_fill_1 FILLER_58_635 ();
 sg13g2_fill_2 FILLER_58_646 ();
 sg13g2_decap_4 FILLER_58_704 ();
 sg13g2_fill_1 FILLER_58_789 ();
 sg13g2_fill_2 FILLER_58_794 ();
 sg13g2_fill_1 FILLER_58_804 ();
 sg13g2_fill_2 FILLER_58_815 ();
 sg13g2_decap_8 FILLER_58_821 ();
 sg13g2_decap_4 FILLER_58_828 ();
 sg13g2_fill_2 FILLER_58_832 ();
 sg13g2_fill_1 FILLER_58_842 ();
 sg13g2_fill_1 FILLER_58_852 ();
 sg13g2_fill_1 FILLER_58_861 ();
 sg13g2_fill_2 FILLER_58_915 ();
 sg13g2_fill_2 FILLER_58_947 ();
 sg13g2_fill_1 FILLER_58_1000 ();
 sg13g2_fill_2 FILLER_58_1006 ();
 sg13g2_fill_1 FILLER_58_1008 ();
 sg13g2_fill_2 FILLER_58_1013 ();
 sg13g2_fill_1 FILLER_58_1015 ();
 sg13g2_fill_1 FILLER_58_1121 ();
 sg13g2_fill_1 FILLER_58_1132 ();
 sg13g2_fill_1 FILLER_58_1159 ();
 sg13g2_fill_2 FILLER_58_1165 ();
 sg13g2_fill_1 FILLER_58_1171 ();
 sg13g2_fill_2 FILLER_58_1211 ();
 sg13g2_fill_1 FILLER_58_1213 ();
 sg13g2_fill_2 FILLER_58_1231 ();
 sg13g2_fill_1 FILLER_58_1233 ();
 sg13g2_decap_8 FILLER_58_1244 ();
 sg13g2_fill_2 FILLER_58_1251 ();
 sg13g2_decap_4 FILLER_58_1279 ();
 sg13g2_fill_1 FILLER_58_1294 ();
 sg13g2_fill_2 FILLER_58_1302 ();
 sg13g2_fill_2 FILLER_58_1312 ();
 sg13g2_fill_1 FILLER_58_1328 ();
 sg13g2_fill_1 FILLER_58_1342 ();
 sg13g2_decap_4 FILLER_58_1348 ();
 sg13g2_fill_1 FILLER_58_1352 ();
 sg13g2_fill_1 FILLER_58_1374 ();
 sg13g2_decap_4 FILLER_58_1399 ();
 sg13g2_fill_1 FILLER_58_1403 ();
 sg13g2_decap_8 FILLER_58_1419 ();
 sg13g2_fill_2 FILLER_58_1426 ();
 sg13g2_decap_8 FILLER_58_1436 ();
 sg13g2_decap_8 FILLER_58_1443 ();
 sg13g2_fill_2 FILLER_58_1470 ();
 sg13g2_fill_1 FILLER_58_1477 ();
 sg13g2_fill_1 FILLER_58_1483 ();
 sg13g2_fill_2 FILLER_58_1492 ();
 sg13g2_decap_8 FILLER_58_1524 ();
 sg13g2_decap_8 FILLER_58_1531 ();
 sg13g2_decap_8 FILLER_58_1538 ();
 sg13g2_decap_4 FILLER_58_1545 ();
 sg13g2_fill_1 FILLER_58_1554 ();
 sg13g2_decap_8 FILLER_58_1559 ();
 sg13g2_decap_8 FILLER_58_1566 ();
 sg13g2_decap_8 FILLER_58_1573 ();
 sg13g2_decap_8 FILLER_58_1580 ();
 sg13g2_decap_8 FILLER_58_1587 ();
 sg13g2_decap_8 FILLER_58_1594 ();
 sg13g2_decap_4 FILLER_58_1606 ();
 sg13g2_fill_1 FILLER_58_1623 ();
 sg13g2_decap_8 FILLER_58_1629 ();
 sg13g2_decap_4 FILLER_58_1636 ();
 sg13g2_fill_2 FILLER_58_1640 ();
 sg13g2_decap_4 FILLER_58_1645 ();
 sg13g2_decap_8 FILLER_58_1652 ();
 sg13g2_fill_2 FILLER_58_1659 ();
 sg13g2_fill_1 FILLER_58_1661 ();
 sg13g2_fill_2 FILLER_58_1665 ();
 sg13g2_fill_2 FILLER_58_1673 ();
 sg13g2_fill_2 FILLER_58_1699 ();
 sg13g2_fill_1 FILLER_58_1701 ();
 sg13g2_decap_8 FILLER_58_1706 ();
 sg13g2_decap_8 FILLER_58_1713 ();
 sg13g2_decap_8 FILLER_58_1725 ();
 sg13g2_fill_1 FILLER_58_1737 ();
 sg13g2_fill_2 FILLER_58_1743 ();
 sg13g2_fill_2 FILLER_58_1750 ();
 sg13g2_fill_2 FILLER_58_1773 ();
 sg13g2_decap_8 FILLER_58_1779 ();
 sg13g2_decap_8 FILLER_58_1786 ();
 sg13g2_decap_8 FILLER_58_1793 ();
 sg13g2_decap_4 FILLER_58_1800 ();
 sg13g2_fill_1 FILLER_58_1812 ();
 sg13g2_fill_1 FILLER_58_1824 ();
 sg13g2_decap_4 FILLER_58_1833 ();
 sg13g2_fill_1 FILLER_58_1837 ();
 sg13g2_fill_1 FILLER_58_1842 ();
 sg13g2_fill_1 FILLER_58_1853 ();
 sg13g2_decap_8 FILLER_58_1862 ();
 sg13g2_decap_4 FILLER_58_1869 ();
 sg13g2_fill_2 FILLER_58_1873 ();
 sg13g2_fill_1 FILLER_58_1885 ();
 sg13g2_fill_1 FILLER_58_1891 ();
 sg13g2_fill_1 FILLER_58_1896 ();
 sg13g2_fill_1 FILLER_58_1902 ();
 sg13g2_fill_2 FILLER_58_1935 ();
 sg13g2_fill_1 FILLER_58_1937 ();
 sg13g2_decap_8 FILLER_58_1954 ();
 sg13g2_fill_2 FILLER_58_1961 ();
 sg13g2_fill_1 FILLER_58_1963 ();
 sg13g2_decap_8 FILLER_58_1983 ();
 sg13g2_fill_2 FILLER_58_1990 ();
 sg13g2_fill_2 FILLER_58_2000 ();
 sg13g2_fill_2 FILLER_58_2007 ();
 sg13g2_fill_1 FILLER_58_2026 ();
 sg13g2_fill_2 FILLER_58_2031 ();
 sg13g2_fill_1 FILLER_58_2033 ();
 sg13g2_fill_2 FILLER_58_2038 ();
 sg13g2_fill_2 FILLER_58_2044 ();
 sg13g2_fill_1 FILLER_58_2046 ();
 sg13g2_decap_8 FILLER_58_2076 ();
 sg13g2_decap_4 FILLER_58_2102 ();
 sg13g2_fill_1 FILLER_58_2106 ();
 sg13g2_fill_1 FILLER_58_2146 ();
 sg13g2_fill_1 FILLER_58_2152 ();
 sg13g2_fill_2 FILLER_58_2163 ();
 sg13g2_fill_1 FILLER_58_2165 ();
 sg13g2_decap_4 FILLER_58_2187 ();
 sg13g2_fill_1 FILLER_58_2191 ();
 sg13g2_decap_4 FILLER_58_2222 ();
 sg13g2_decap_4 FILLER_58_2231 ();
 sg13g2_fill_1 FILLER_58_2235 ();
 sg13g2_fill_1 FILLER_58_2262 ();
 sg13g2_fill_1 FILLER_58_2267 ();
 sg13g2_fill_2 FILLER_58_2272 ();
 sg13g2_fill_2 FILLER_58_2279 ();
 sg13g2_fill_1 FILLER_58_2281 ();
 sg13g2_decap_4 FILLER_58_2304 ();
 sg13g2_fill_2 FILLER_58_2313 ();
 sg13g2_fill_2 FILLER_58_2345 ();
 sg13g2_fill_1 FILLER_58_2347 ();
 sg13g2_fill_2 FILLER_58_2379 ();
 sg13g2_fill_1 FILLER_58_2386 ();
 sg13g2_fill_2 FILLER_58_2391 ();
 sg13g2_fill_2 FILLER_58_2397 ();
 sg13g2_fill_2 FILLER_58_2403 ();
 sg13g2_fill_1 FILLER_58_2411 ();
 sg13g2_fill_1 FILLER_58_2425 ();
 sg13g2_fill_2 FILLER_58_2430 ();
 sg13g2_fill_1 FILLER_58_2432 ();
 sg13g2_decap_4 FILLER_58_2467 ();
 sg13g2_fill_1 FILLER_58_2506 ();
 sg13g2_decap_8 FILLER_58_2516 ();
 sg13g2_decap_8 FILLER_58_2523 ();
 sg13g2_decap_8 FILLER_58_2530 ();
 sg13g2_fill_1 FILLER_58_2537 ();
 sg13g2_decap_8 FILLER_58_2546 ();
 sg13g2_decap_8 FILLER_58_2553 ();
 sg13g2_decap_8 FILLER_58_2560 ();
 sg13g2_fill_2 FILLER_58_2571 ();
 sg13g2_decap_8 FILLER_58_2581 ();
 sg13g2_fill_2 FILLER_58_2588 ();
 sg13g2_fill_1 FILLER_58_2590 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_4 FILLER_59_14 ();
 sg13g2_fill_2 FILLER_59_18 ();
 sg13g2_fill_1 FILLER_59_30 ();
 sg13g2_fill_1 FILLER_59_61 ();
 sg13g2_decap_8 FILLER_59_66 ();
 sg13g2_fill_1 FILLER_59_73 ();
 sg13g2_decap_4 FILLER_59_126 ();
 sg13g2_decap_4 FILLER_59_134 ();
 sg13g2_fill_1 FILLER_59_138 ();
 sg13g2_fill_2 FILLER_59_155 ();
 sg13g2_fill_2 FILLER_59_168 ();
 sg13g2_fill_2 FILLER_59_174 ();
 sg13g2_fill_1 FILLER_59_176 ();
 sg13g2_fill_1 FILLER_59_198 ();
 sg13g2_fill_2 FILLER_59_222 ();
 sg13g2_decap_8 FILLER_59_228 ();
 sg13g2_decap_8 FILLER_59_235 ();
 sg13g2_decap_8 FILLER_59_242 ();
 sg13g2_fill_1 FILLER_59_280 ();
 sg13g2_fill_1 FILLER_59_311 ();
 sg13g2_fill_2 FILLER_59_321 ();
 sg13g2_fill_1 FILLER_59_327 ();
 sg13g2_fill_2 FILLER_59_333 ();
 sg13g2_fill_1 FILLER_59_366 ();
 sg13g2_fill_2 FILLER_59_372 ();
 sg13g2_fill_2 FILLER_59_382 ();
 sg13g2_fill_1 FILLER_59_395 ();
 sg13g2_fill_2 FILLER_59_405 ();
 sg13g2_fill_2 FILLER_59_410 ();
 sg13g2_fill_1 FILLER_59_441 ();
 sg13g2_fill_1 FILLER_59_484 ();
 sg13g2_decap_8 FILLER_59_552 ();
 sg13g2_decap_4 FILLER_59_569 ();
 sg13g2_fill_1 FILLER_59_573 ();
 sg13g2_fill_2 FILLER_59_584 ();
 sg13g2_fill_1 FILLER_59_591 ();
 sg13g2_decap_8 FILLER_59_598 ();
 sg13g2_decap_8 FILLER_59_605 ();
 sg13g2_decap_4 FILLER_59_612 ();
 sg13g2_fill_1 FILLER_59_616 ();
 sg13g2_decap_8 FILLER_59_623 ();
 sg13g2_decap_4 FILLER_59_630 ();
 sg13g2_fill_1 FILLER_59_640 ();
 sg13g2_fill_2 FILLER_59_689 ();
 sg13g2_fill_1 FILLER_59_691 ();
 sg13g2_fill_1 FILLER_59_828 ();
 sg13g2_fill_1 FILLER_59_837 ();
 sg13g2_fill_1 FILLER_59_842 ();
 sg13g2_fill_2 FILLER_59_886 ();
 sg13g2_fill_1 FILLER_59_971 ();
 sg13g2_fill_1 FILLER_59_994 ();
 sg13g2_fill_2 FILLER_59_1000 ();
 sg13g2_decap_4 FILLER_59_1009 ();
 sg13g2_fill_1 FILLER_59_1013 ();
 sg13g2_fill_1 FILLER_59_1029 ();
 sg13g2_fill_2 FILLER_59_1068 ();
 sg13g2_fill_1 FILLER_59_1070 ();
 sg13g2_decap_4 FILLER_59_1081 ();
 sg13g2_fill_2 FILLER_59_1085 ();
 sg13g2_fill_2 FILLER_59_1091 ();
 sg13g2_fill_1 FILLER_59_1104 ();
 sg13g2_decap_8 FILLER_59_1144 ();
 sg13g2_fill_2 FILLER_59_1151 ();
 sg13g2_fill_1 FILLER_59_1153 ();
 sg13g2_decap_8 FILLER_59_1163 ();
 sg13g2_decap_8 FILLER_59_1170 ();
 sg13g2_decap_8 FILLER_59_1177 ();
 sg13g2_fill_1 FILLER_59_1184 ();
 sg13g2_fill_2 FILLER_59_1195 ();
 sg13g2_fill_1 FILLER_59_1197 ();
 sg13g2_fill_1 FILLER_59_1224 ();
 sg13g2_decap_8 FILLER_59_1251 ();
 sg13g2_decap_4 FILLER_59_1258 ();
 sg13g2_decap_8 FILLER_59_1266 ();
 sg13g2_decap_8 FILLER_59_1283 ();
 sg13g2_decap_4 FILLER_59_1306 ();
 sg13g2_fill_2 FILLER_59_1310 ();
 sg13g2_fill_1 FILLER_59_1321 ();
 sg13g2_fill_1 FILLER_59_1337 ();
 sg13g2_fill_1 FILLER_59_1358 ();
 sg13g2_fill_2 FILLER_59_1365 ();
 sg13g2_fill_1 FILLER_59_1388 ();
 sg13g2_decap_4 FILLER_59_1415 ();
 sg13g2_fill_1 FILLER_59_1419 ();
 sg13g2_fill_1 FILLER_59_1452 ();
 sg13g2_fill_1 FILLER_59_1461 ();
 sg13g2_fill_2 FILLER_59_1487 ();
 sg13g2_decap_8 FILLER_59_1499 ();
 sg13g2_decap_4 FILLER_59_1506 ();
 sg13g2_decap_8 FILLER_59_1556 ();
 sg13g2_fill_1 FILLER_59_1563 ();
 sg13g2_fill_1 FILLER_59_1622 ();
 sg13g2_fill_2 FILLER_59_1631 ();
 sg13g2_decap_4 FILLER_59_1642 ();
 sg13g2_fill_2 FILLER_59_1646 ();
 sg13g2_fill_2 FILLER_59_1663 ();
 sg13g2_fill_2 FILLER_59_1670 ();
 sg13g2_fill_1 FILLER_59_1709 ();
 sg13g2_fill_2 FILLER_59_1718 ();
 sg13g2_fill_2 FILLER_59_1746 ();
 sg13g2_fill_2 FILLER_59_1790 ();
 sg13g2_fill_1 FILLER_59_1792 ();
 sg13g2_decap_4 FILLER_59_1797 ();
 sg13g2_fill_2 FILLER_59_1801 ();
 sg13g2_decap_4 FILLER_59_1815 ();
 sg13g2_fill_2 FILLER_59_1819 ();
 sg13g2_fill_2 FILLER_59_1825 ();
 sg13g2_fill_1 FILLER_59_1827 ();
 sg13g2_fill_2 FILLER_59_1832 ();
 sg13g2_decap_8 FILLER_59_1860 ();
 sg13g2_decap_8 FILLER_59_1867 ();
 sg13g2_fill_2 FILLER_59_1874 ();
 sg13g2_fill_1 FILLER_59_1885 ();
 sg13g2_fill_1 FILLER_59_1891 ();
 sg13g2_fill_2 FILLER_59_1920 ();
 sg13g2_fill_1 FILLER_59_1922 ();
 sg13g2_fill_1 FILLER_59_1932 ();
 sg13g2_decap_4 FILLER_59_1959 ();
 sg13g2_fill_2 FILLER_59_1963 ();
 sg13g2_decap_4 FILLER_59_1971 ();
 sg13g2_fill_2 FILLER_59_1975 ();
 sg13g2_fill_1 FILLER_59_1987 ();
 sg13g2_fill_1 FILLER_59_1992 ();
 sg13g2_fill_2 FILLER_59_2025 ();
 sg13g2_fill_2 FILLER_59_2031 ();
 sg13g2_decap_8 FILLER_59_2037 ();
 sg13g2_decap_8 FILLER_59_2044 ();
 sg13g2_fill_1 FILLER_59_2051 ();
 sg13g2_decap_8 FILLER_59_2066 ();
 sg13g2_fill_2 FILLER_59_2073 ();
 sg13g2_fill_2 FILLER_59_2080 ();
 sg13g2_fill_1 FILLER_59_2082 ();
 sg13g2_fill_1 FILLER_59_2135 ();
 sg13g2_decap_4 FILLER_59_2155 ();
 sg13g2_fill_2 FILLER_59_2185 ();
 sg13g2_fill_2 FILLER_59_2213 ();
 sg13g2_fill_2 FILLER_59_2224 ();
 sg13g2_fill_1 FILLER_59_2231 ();
 sg13g2_fill_1 FILLER_59_2236 ();
 sg13g2_fill_2 FILLER_59_2242 ();
 sg13g2_fill_1 FILLER_59_2244 ();
 sg13g2_fill_1 FILLER_59_2271 ();
 sg13g2_decap_8 FILLER_59_2303 ();
 sg13g2_decap_4 FILLER_59_2310 ();
 sg13g2_fill_2 FILLER_59_2314 ();
 sg13g2_decap_4 FILLER_59_2348 ();
 sg13g2_fill_2 FILLER_59_2361 ();
 sg13g2_fill_1 FILLER_59_2363 ();
 sg13g2_fill_1 FILLER_59_2374 ();
 sg13g2_fill_1 FILLER_59_2379 ();
 sg13g2_fill_2 FILLER_59_2392 ();
 sg13g2_fill_1 FILLER_59_2394 ();
 sg13g2_fill_2 FILLER_59_2400 ();
 sg13g2_fill_1 FILLER_59_2402 ();
 sg13g2_fill_2 FILLER_59_2429 ();
 sg13g2_fill_1 FILLER_59_2431 ();
 sg13g2_decap_4 FILLER_59_2465 ();
 sg13g2_fill_1 FILLER_59_2473 ();
 sg13g2_fill_1 FILLER_59_2480 ();
 sg13g2_fill_2 FILLER_59_2496 ();
 sg13g2_fill_2 FILLER_59_2528 ();
 sg13g2_fill_2 FILLER_59_2562 ();
 sg13g2_fill_2 FILLER_59_2568 ();
 sg13g2_fill_1 FILLER_59_2570 ();
 sg13g2_decap_8 FILLER_59_2594 ();
 sg13g2_fill_2 FILLER_59_2601 ();
 sg13g2_decap_8 FILLER_59_2607 ();
 sg13g2_fill_2 FILLER_59_2622 ();
 sg13g2_decap_4 FILLER_59_2664 ();
 sg13g2_fill_2 FILLER_59_2668 ();
 sg13g2_fill_1 FILLER_60_0 ();
 sg13g2_fill_1 FILLER_60_27 ();
 sg13g2_fill_1 FILLER_60_38 ();
 sg13g2_fill_1 FILLER_60_44 ();
 sg13g2_fill_1 FILLER_60_49 ();
 sg13g2_fill_1 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_93 ();
 sg13g2_decap_4 FILLER_60_100 ();
 sg13g2_fill_2 FILLER_60_104 ();
 sg13g2_decap_8 FILLER_60_128 ();
 sg13g2_decap_8 FILLER_60_135 ();
 sg13g2_fill_1 FILLER_60_142 ();
 sg13g2_decap_4 FILLER_60_168 ();
 sg13g2_fill_1 FILLER_60_172 ();
 sg13g2_fill_2 FILLER_60_213 ();
 sg13g2_decap_8 FILLER_60_221 ();
 sg13g2_decap_8 FILLER_60_228 ();
 sg13g2_decap_4 FILLER_60_235 ();
 sg13g2_fill_1 FILLER_60_239 ();
 sg13g2_fill_2 FILLER_60_250 ();
 sg13g2_fill_1 FILLER_60_295 ();
 sg13g2_fill_1 FILLER_60_397 ();
 sg13g2_fill_1 FILLER_60_406 ();
 sg13g2_fill_1 FILLER_60_429 ();
 sg13g2_fill_1 FILLER_60_435 ();
 sg13g2_fill_2 FILLER_60_444 ();
 sg13g2_fill_2 FILLER_60_460 ();
 sg13g2_decap_8 FILLER_60_469 ();
 sg13g2_decap_8 FILLER_60_476 ();
 sg13g2_fill_2 FILLER_60_483 ();
 sg13g2_fill_1 FILLER_60_485 ();
 sg13g2_fill_1 FILLER_60_505 ();
 sg13g2_fill_1 FILLER_60_511 ();
 sg13g2_decap_4 FILLER_60_553 ();
 sg13g2_decap_4 FILLER_60_607 ();
 sg13g2_decap_8 FILLER_60_628 ();
 sg13g2_fill_1 FILLER_60_635 ();
 sg13g2_fill_1 FILLER_60_641 ();
 sg13g2_decap_8 FILLER_60_685 ();
 sg13g2_decap_4 FILLER_60_692 ();
 sg13g2_fill_2 FILLER_60_696 ();
 sg13g2_decap_4 FILLER_60_709 ();
 sg13g2_fill_2 FILLER_60_767 ();
 sg13g2_fill_1 FILLER_60_837 ();
 sg13g2_fill_1 FILLER_60_843 ();
 sg13g2_fill_1 FILLER_60_860 ();
 sg13g2_fill_1 FILLER_60_866 ();
 sg13g2_fill_2 FILLER_60_875 ();
 sg13g2_fill_2 FILLER_60_907 ();
 sg13g2_fill_1 FILLER_60_913 ();
 sg13g2_fill_1 FILLER_60_940 ();
 sg13g2_fill_1 FILLER_60_951 ();
 sg13g2_fill_1 FILLER_60_956 ();
 sg13g2_fill_1 FILLER_60_961 ();
 sg13g2_fill_1 FILLER_60_967 ();
 sg13g2_fill_1 FILLER_60_1011 ();
 sg13g2_fill_1 FILLER_60_1025 ();
 sg13g2_fill_2 FILLER_60_1031 ();
 sg13g2_decap_8 FILLER_60_1057 ();
 sg13g2_fill_2 FILLER_60_1112 ();
 sg13g2_fill_1 FILLER_60_1191 ();
 sg13g2_fill_2 FILLER_60_1232 ();
 sg13g2_decap_8 FILLER_60_1238 ();
 sg13g2_fill_2 FILLER_60_1245 ();
 sg13g2_fill_1 FILLER_60_1247 ();
 sg13g2_decap_8 FILLER_60_1258 ();
 sg13g2_decap_8 FILLER_60_1265 ();
 sg13g2_fill_2 FILLER_60_1272 ();
 sg13g2_fill_1 FILLER_60_1274 ();
 sg13g2_fill_1 FILLER_60_1283 ();
 sg13g2_decap_8 FILLER_60_1308 ();
 sg13g2_fill_2 FILLER_60_1315 ();
 sg13g2_fill_1 FILLER_60_1317 ();
 sg13g2_fill_1 FILLER_60_1337 ();
 sg13g2_decap_4 FILLER_60_1352 ();
 sg13g2_fill_2 FILLER_60_1356 ();
 sg13g2_fill_2 FILLER_60_1363 ();
 sg13g2_fill_1 FILLER_60_1365 ();
 sg13g2_fill_1 FILLER_60_1392 ();
 sg13g2_fill_1 FILLER_60_1398 ();
 sg13g2_decap_4 FILLER_60_1402 ();
 sg13g2_fill_1 FILLER_60_1414 ();
 sg13g2_decap_4 FILLER_60_1420 ();
 sg13g2_fill_2 FILLER_60_1424 ();
 sg13g2_decap_4 FILLER_60_1439 ();
 sg13g2_fill_1 FILLER_60_1443 ();
 sg13g2_fill_2 FILLER_60_1453 ();
 sg13g2_fill_1 FILLER_60_1455 ();
 sg13g2_fill_1 FILLER_60_1468 ();
 sg13g2_fill_2 FILLER_60_1479 ();
 sg13g2_fill_1 FILLER_60_1481 ();
 sg13g2_fill_2 FILLER_60_1486 ();
 sg13g2_fill_2 FILLER_60_1507 ();
 sg13g2_decap_8 FILLER_60_1514 ();
 sg13g2_decap_8 FILLER_60_1561 ();
 sg13g2_decap_4 FILLER_60_1568 ();
 sg13g2_fill_2 FILLER_60_1572 ();
 sg13g2_decap_4 FILLER_60_1578 ();
 sg13g2_fill_1 FILLER_60_1582 ();
 sg13g2_fill_1 FILLER_60_1588 ();
 sg13g2_fill_2 FILLER_60_1607 ();
 sg13g2_fill_2 FILLER_60_1617 ();
 sg13g2_fill_1 FILLER_60_1623 ();
 sg13g2_fill_2 FILLER_60_1642 ();
 sg13g2_fill_2 FILLER_60_1655 ();
 sg13g2_fill_1 FILLER_60_1663 ();
 sg13g2_fill_1 FILLER_60_1696 ();
 sg13g2_fill_2 FILLER_60_1701 ();
 sg13g2_fill_1 FILLER_60_1703 ();
 sg13g2_fill_1 FILLER_60_1730 ();
 sg13g2_fill_1 FILLER_60_1735 ();
 sg13g2_decap_4 FILLER_60_1740 ();
 sg13g2_fill_1 FILLER_60_1744 ();
 sg13g2_fill_2 FILLER_60_1769 ();
 sg13g2_fill_1 FILLER_60_1788 ();
 sg13g2_fill_1 FILLER_60_1797 ();
 sg13g2_fill_2 FILLER_60_1802 ();
 sg13g2_fill_1 FILLER_60_1804 ();
 sg13g2_fill_2 FILLER_60_1809 ();
 sg13g2_fill_1 FILLER_60_1811 ();
 sg13g2_decap_4 FILLER_60_1829 ();
 sg13g2_fill_2 FILLER_60_1833 ();
 sg13g2_fill_2 FILLER_60_1843 ();
 sg13g2_fill_1 FILLER_60_1845 ();
 sg13g2_decap_8 FILLER_60_1850 ();
 sg13g2_decap_8 FILLER_60_1857 ();
 sg13g2_decap_8 FILLER_60_1864 ();
 sg13g2_decap_8 FILLER_60_1871 ();
 sg13g2_fill_1 FILLER_60_1878 ();
 sg13g2_fill_1 FILLER_60_1883 ();
 sg13g2_fill_1 FILLER_60_1897 ();
 sg13g2_fill_2 FILLER_60_1903 ();
 sg13g2_fill_1 FILLER_60_1905 ();
 sg13g2_fill_2 FILLER_60_1915 ();
 sg13g2_fill_1 FILLER_60_1922 ();
 sg13g2_fill_2 FILLER_60_1936 ();
 sg13g2_fill_2 FILLER_60_1945 ();
 sg13g2_fill_1 FILLER_60_1947 ();
 sg13g2_decap_8 FILLER_60_1952 ();
 sg13g2_decap_4 FILLER_60_1959 ();
 sg13g2_fill_2 FILLER_60_1963 ();
 sg13g2_decap_4 FILLER_60_1986 ();
 sg13g2_fill_1 FILLER_60_1990 ();
 sg13g2_fill_2 FILLER_60_1996 ();
 sg13g2_fill_2 FILLER_60_2025 ();
 sg13g2_fill_1 FILLER_60_2027 ();
 sg13g2_decap_8 FILLER_60_2045 ();
 sg13g2_decap_8 FILLER_60_2057 ();
 sg13g2_fill_1 FILLER_60_2064 ();
 sg13g2_decap_4 FILLER_60_2070 ();
 sg13g2_decap_8 FILLER_60_2079 ();
 sg13g2_fill_1 FILLER_60_2086 ();
 sg13g2_fill_1 FILLER_60_2092 ();
 sg13g2_fill_1 FILLER_60_2143 ();
 sg13g2_decap_4 FILLER_60_2164 ();
 sg13g2_fill_1 FILLER_60_2172 ();
 sg13g2_decap_8 FILLER_60_2177 ();
 sg13g2_decap_8 FILLER_60_2184 ();
 sg13g2_decap_8 FILLER_60_2191 ();
 sg13g2_fill_2 FILLER_60_2198 ();
 sg13g2_fill_2 FILLER_60_2204 ();
 sg13g2_fill_1 FILLER_60_2256 ();
 sg13g2_decap_8 FILLER_60_2261 ();
 sg13g2_fill_2 FILLER_60_2268 ();
 sg13g2_fill_1 FILLER_60_2270 ();
 sg13g2_fill_2 FILLER_60_2302 ();
 sg13g2_fill_1 FILLER_60_2304 ();
 sg13g2_decap_4 FILLER_60_2311 ();
 sg13g2_fill_2 FILLER_60_2324 ();
 sg13g2_decap_8 FILLER_60_2330 ();
 sg13g2_fill_2 FILLER_60_2337 ();
 sg13g2_decap_8 FILLER_60_2348 ();
 sg13g2_fill_2 FILLER_60_2355 ();
 sg13g2_fill_1 FILLER_60_2357 ();
 sg13g2_fill_2 FILLER_60_2362 ();
 sg13g2_decap_8 FILLER_60_2439 ();
 sg13g2_decap_4 FILLER_60_2459 ();
 sg13g2_fill_1 FILLER_60_2463 ();
 sg13g2_decap_4 FILLER_60_2469 ();
 sg13g2_fill_1 FILLER_60_2473 ();
 sg13g2_fill_2 FILLER_60_2479 ();
 sg13g2_fill_1 FILLER_60_2486 ();
 sg13g2_decap_4 FILLER_60_2499 ();
 sg13g2_fill_2 FILLER_60_2503 ();
 sg13g2_fill_2 FILLER_60_2511 ();
 sg13g2_fill_1 FILLER_60_2549 ();
 sg13g2_fill_2 FILLER_60_2555 ();
 sg13g2_decap_8 FILLER_60_2583 ();
 sg13g2_fill_2 FILLER_60_2590 ();
 sg13g2_decap_8 FILLER_60_2601 ();
 sg13g2_fill_2 FILLER_60_2608 ();
 sg13g2_fill_1 FILLER_60_2610 ();
 sg13g2_fill_1 FILLER_60_2637 ();
 sg13g2_decap_8 FILLER_60_2645 ();
 sg13g2_decap_8 FILLER_60_2652 ();
 sg13g2_decap_8 FILLER_60_2659 ();
 sg13g2_decap_4 FILLER_60_2666 ();
 sg13g2_fill_2 FILLER_61_0 ();
 sg13g2_fill_2 FILLER_61_28 ();
 sg13g2_fill_2 FILLER_61_56 ();
 sg13g2_fill_1 FILLER_61_58 ();
 sg13g2_decap_4 FILLER_61_69 ();
 sg13g2_fill_1 FILLER_61_73 ();
 sg13g2_decap_8 FILLER_61_78 ();
 sg13g2_decap_8 FILLER_61_85 ();
 sg13g2_decap_8 FILLER_61_92 ();
 sg13g2_decap_8 FILLER_61_99 ();
 sg13g2_fill_2 FILLER_61_106 ();
 sg13g2_fill_2 FILLER_61_111 ();
 sg13g2_fill_2 FILLER_61_142 ();
 sg13g2_decap_8 FILLER_61_184 ();
 sg13g2_decap_8 FILLER_61_191 ();
 sg13g2_decap_8 FILLER_61_198 ();
 sg13g2_fill_2 FILLER_61_205 ();
 sg13g2_decap_8 FILLER_61_213 ();
 sg13g2_decap_8 FILLER_61_220 ();
 sg13g2_decap_4 FILLER_61_227 ();
 sg13g2_decap_4 FILLER_61_245 ();
 sg13g2_fill_2 FILLER_61_249 ();
 sg13g2_fill_1 FILLER_61_299 ();
 sg13g2_fill_1 FILLER_61_317 ();
 sg13g2_fill_1 FILLER_61_332 ();
 sg13g2_fill_2 FILLER_61_337 ();
 sg13g2_fill_2 FILLER_61_350 ();
 sg13g2_fill_1 FILLER_61_375 ();
 sg13g2_fill_2 FILLER_61_428 ();
 sg13g2_fill_2 FILLER_61_438 ();
 sg13g2_fill_2 FILLER_61_444 ();
 sg13g2_fill_2 FILLER_61_460 ();
 sg13g2_decap_8 FILLER_61_466 ();
 sg13g2_fill_2 FILLER_61_473 ();
 sg13g2_fill_1 FILLER_61_475 ();
 sg13g2_fill_2 FILLER_61_486 ();
 sg13g2_fill_1 FILLER_61_498 ();
 sg13g2_fill_2 FILLER_61_516 ();
 sg13g2_fill_2 FILLER_61_523 ();
 sg13g2_fill_2 FILLER_61_530 ();
 sg13g2_fill_1 FILLER_61_532 ();
 sg13g2_decap_8 FILLER_61_548 ();
 sg13g2_decap_8 FILLER_61_555 ();
 sg13g2_decap_8 FILLER_61_562 ();
 sg13g2_fill_2 FILLER_61_569 ();
 sg13g2_decap_8 FILLER_61_629 ();
 sg13g2_fill_1 FILLER_61_636 ();
 sg13g2_fill_2 FILLER_61_641 ();
 sg13g2_fill_1 FILLER_61_643 ();
 sg13g2_fill_1 FILLER_61_649 ();
 sg13g2_fill_2 FILLER_61_655 ();
 sg13g2_fill_2 FILLER_61_702 ();
 sg13g2_fill_2 FILLER_61_716 ();
 sg13g2_decap_4 FILLER_61_739 ();
 sg13g2_fill_1 FILLER_61_743 ();
 sg13g2_fill_1 FILLER_61_795 ();
 sg13g2_fill_1 FILLER_61_810 ();
 sg13g2_fill_2 FILLER_61_823 ();
 sg13g2_fill_1 FILLER_61_886 ();
 sg13g2_fill_2 FILLER_61_916 ();
 sg13g2_fill_1 FILLER_61_931 ();
 sg13g2_fill_1 FILLER_61_996 ();
 sg13g2_fill_1 FILLER_61_1021 ();
 sg13g2_fill_1 FILLER_61_1030 ();
 sg13g2_fill_1 FILLER_61_1035 ();
 sg13g2_fill_2 FILLER_61_1044 ();
 sg13g2_fill_1 FILLER_61_1055 ();
 sg13g2_decap_4 FILLER_61_1065 ();
 sg13g2_fill_1 FILLER_61_1069 ();
 sg13g2_decap_4 FILLER_61_1117 ();
 sg13g2_fill_1 FILLER_61_1121 ();
 sg13g2_fill_1 FILLER_61_1132 ();
 sg13g2_fill_1 FILLER_61_1159 ();
 sg13g2_fill_2 FILLER_61_1169 ();
 sg13g2_fill_2 FILLER_61_1175 ();
 sg13g2_fill_1 FILLER_61_1177 ();
 sg13g2_fill_2 FILLER_61_1204 ();
 sg13g2_decap_4 FILLER_61_1220 ();
 sg13g2_decap_8 FILLER_61_1276 ();
 sg13g2_fill_2 FILLER_61_1316 ();
 sg13g2_fill_2 FILLER_61_1324 ();
 sg13g2_fill_1 FILLER_61_1326 ();
 sg13g2_fill_2 FILLER_61_1332 ();
 sg13g2_fill_1 FILLER_61_1334 ();
 sg13g2_fill_1 FILLER_61_1340 ();
 sg13g2_decap_8 FILLER_61_1345 ();
 sg13g2_fill_2 FILLER_61_1352 ();
 sg13g2_fill_1 FILLER_61_1360 ();
 sg13g2_fill_1 FILLER_61_1367 ();
 sg13g2_fill_1 FILLER_61_1373 ();
 sg13g2_fill_2 FILLER_61_1389 ();
 sg13g2_decap_8 FILLER_61_1397 ();
 sg13g2_fill_2 FILLER_61_1404 ();
 sg13g2_fill_2 FILLER_61_1412 ();
 sg13g2_fill_2 FILLER_61_1428 ();
 sg13g2_fill_2 FILLER_61_1440 ();
 sg13g2_decap_8 FILLER_61_1447 ();
 sg13g2_decap_8 FILLER_61_1458 ();
 sg13g2_fill_2 FILLER_61_1465 ();
 sg13g2_fill_2 FILLER_61_1494 ();
 sg13g2_fill_1 FILLER_61_1511 ();
 sg13g2_fill_2 FILLER_61_1516 ();
 sg13g2_fill_1 FILLER_61_1518 ();
 sg13g2_decap_4 FILLER_61_1536 ();
 sg13g2_fill_2 FILLER_61_1570 ();
 sg13g2_decap_4 FILLER_61_1589 ();
 sg13g2_fill_2 FILLER_61_1593 ();
 sg13g2_fill_1 FILLER_61_1606 ();
 sg13g2_decap_4 FILLER_61_1642 ();
 sg13g2_fill_2 FILLER_61_1646 ();
 sg13g2_fill_1 FILLER_61_1679 ();
 sg13g2_fill_1 FILLER_61_1703 ();
 sg13g2_fill_2 FILLER_61_1707 ();
 sg13g2_fill_1 FILLER_61_1709 ();
 sg13g2_decap_4 FILLER_61_1717 ();
 sg13g2_fill_1 FILLER_61_1721 ();
 sg13g2_fill_2 FILLER_61_1739 ();
 sg13g2_fill_1 FILLER_61_1741 ();
 sg13g2_decap_8 FILLER_61_1753 ();
 sg13g2_decap_8 FILLER_61_1760 ();
 sg13g2_fill_2 FILLER_61_1767 ();
 sg13g2_fill_1 FILLER_61_1790 ();
 sg13g2_fill_2 FILLER_61_1820 ();
 sg13g2_decap_4 FILLER_61_1856 ();
 sg13g2_fill_2 FILLER_61_1860 ();
 sg13g2_decap_8 FILLER_61_1867 ();
 sg13g2_fill_2 FILLER_61_1874 ();
 sg13g2_fill_2 FILLER_61_1881 ();
 sg13g2_fill_1 FILLER_61_1883 ();
 sg13g2_fill_1 FILLER_61_1897 ();
 sg13g2_fill_1 FILLER_61_1902 ();
 sg13g2_fill_1 FILLER_61_1915 ();
 sg13g2_fill_1 FILLER_61_1947 ();
 sg13g2_fill_1 FILLER_61_1980 ();
 sg13g2_fill_2 FILLER_61_1989 ();
 sg13g2_fill_1 FILLER_61_2000 ();
 sg13g2_fill_1 FILLER_61_2006 ();
 sg13g2_fill_2 FILLER_61_2011 ();
 sg13g2_fill_1 FILLER_61_2021 ();
 sg13g2_decap_8 FILLER_61_2031 ();
 sg13g2_decap_4 FILLER_61_2038 ();
 sg13g2_fill_2 FILLER_61_2046 ();
 sg13g2_fill_1 FILLER_61_2048 ();
 sg13g2_decap_8 FILLER_61_2057 ();
 sg13g2_decap_8 FILLER_61_2064 ();
 sg13g2_decap_8 FILLER_61_2071 ();
 sg13g2_decap_8 FILLER_61_2078 ();
 sg13g2_fill_2 FILLER_61_2085 ();
 sg13g2_fill_2 FILLER_61_2103 ();
 sg13g2_fill_1 FILLER_61_2105 ();
 sg13g2_decap_4 FILLER_61_2111 ();
 sg13g2_fill_1 FILLER_61_2115 ();
 sg13g2_decap_4 FILLER_61_2151 ();
 sg13g2_fill_2 FILLER_61_2155 ();
 sg13g2_decap_8 FILLER_61_2187 ();
 sg13g2_decap_4 FILLER_61_2194 ();
 sg13g2_fill_2 FILLER_61_2232 ();
 sg13g2_fill_1 FILLER_61_2234 ();
 sg13g2_fill_2 FILLER_61_2245 ();
 sg13g2_decap_8 FILLER_61_2251 ();
 sg13g2_decap_8 FILLER_61_2258 ();
 sg13g2_decap_4 FILLER_61_2265 ();
 sg13g2_fill_1 FILLER_61_2269 ();
 sg13g2_fill_1 FILLER_61_2275 ();
 sg13g2_fill_1 FILLER_61_2280 ();
 sg13g2_decap_4 FILLER_61_2326 ();
 sg13g2_decap_8 FILLER_61_2336 ();
 sg13g2_decap_8 FILLER_61_2343 ();
 sg13g2_decap_4 FILLER_61_2385 ();
 sg13g2_fill_2 FILLER_61_2389 ();
 sg13g2_decap_8 FILLER_61_2396 ();
 sg13g2_decap_4 FILLER_61_2471 ();
 sg13g2_fill_1 FILLER_61_2501 ();
 sg13g2_fill_1 FILLER_61_2508 ();
 sg13g2_fill_2 FILLER_61_2513 ();
 sg13g2_fill_1 FILLER_61_2519 ();
 sg13g2_fill_1 FILLER_61_2530 ();
 sg13g2_fill_1 FILLER_61_2535 ();
 sg13g2_fill_2 FILLER_61_2540 ();
 sg13g2_fill_2 FILLER_61_2582 ();
 sg13g2_fill_2 FILLER_61_2588 ();
 sg13g2_decap_8 FILLER_61_2616 ();
 sg13g2_decap_4 FILLER_61_2623 ();
 sg13g2_fill_1 FILLER_61_2627 ();
 sg13g2_decap_8 FILLER_61_2634 ();
 sg13g2_decap_8 FILLER_61_2641 ();
 sg13g2_decap_8 FILLER_61_2648 ();
 sg13g2_decap_8 FILLER_61_2655 ();
 sg13g2_decap_8 FILLER_61_2662 ();
 sg13g2_fill_1 FILLER_61_2669 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_15 ();
 sg13g2_fill_1 FILLER_62_26 ();
 sg13g2_fill_1 FILLER_62_37 ();
 sg13g2_fill_1 FILLER_62_42 ();
 sg13g2_fill_2 FILLER_62_92 ();
 sg13g2_fill_1 FILLER_62_94 ();
 sg13g2_fill_1 FILLER_62_108 ();
 sg13g2_fill_1 FILLER_62_113 ();
 sg13g2_fill_2 FILLER_62_148 ();
 sg13g2_fill_1 FILLER_62_150 ();
 sg13g2_decap_4 FILLER_62_249 ();
 sg13g2_fill_2 FILLER_62_253 ();
 sg13g2_fill_1 FILLER_62_290 ();
 sg13g2_fill_1 FILLER_62_342 ();
 sg13g2_fill_2 FILLER_62_376 ();
 sg13g2_fill_1 FILLER_62_401 ();
 sg13g2_fill_1 FILLER_62_428 ();
 sg13g2_fill_1 FILLER_62_455 ();
 sg13g2_fill_2 FILLER_62_495 ();
 sg13g2_decap_4 FILLER_62_564 ();
 sg13g2_fill_1 FILLER_62_568 ();
 sg13g2_decap_4 FILLER_62_577 ();
 sg13g2_fill_2 FILLER_62_581 ();
 sg13g2_fill_2 FILLER_62_619 ();
 sg13g2_fill_1 FILLER_62_621 ();
 sg13g2_fill_2 FILLER_62_694 ();
 sg13g2_decap_8 FILLER_62_709 ();
 sg13g2_fill_2 FILLER_62_716 ();
 sg13g2_decap_8 FILLER_62_723 ();
 sg13g2_fill_2 FILLER_62_744 ();
 sg13g2_fill_1 FILLER_62_746 ();
 sg13g2_fill_1 FILLER_62_763 ();
 sg13g2_fill_1 FILLER_62_770 ();
 sg13g2_fill_1 FILLER_62_775 ();
 sg13g2_fill_2 FILLER_62_806 ();
 sg13g2_fill_2 FILLER_62_916 ();
 sg13g2_fill_2 FILLER_62_949 ();
 sg13g2_fill_2 FILLER_62_976 ();
 sg13g2_fill_1 FILLER_62_1052 ();
 sg13g2_decap_4 FILLER_62_1068 ();
 sg13g2_fill_2 FILLER_62_1072 ();
 sg13g2_decap_8 FILLER_62_1114 ();
 sg13g2_fill_2 FILLER_62_1121 ();
 sg13g2_fill_1 FILLER_62_1153 ();
 sg13g2_fill_1 FILLER_62_1185 ();
 sg13g2_decap_4 FILLER_62_1213 ();
 sg13g2_decap_4 FILLER_62_1253 ();
 sg13g2_fill_1 FILLER_62_1257 ();
 sg13g2_decap_8 FILLER_62_1262 ();
 sg13g2_decap_8 FILLER_62_1269 ();
 sg13g2_fill_2 FILLER_62_1276 ();
 sg13g2_decap_4 FILLER_62_1293 ();
 sg13g2_fill_2 FILLER_62_1309 ();
 sg13g2_fill_1 FILLER_62_1315 ();
 sg13g2_fill_1 FILLER_62_1321 ();
 sg13g2_fill_1 FILLER_62_1329 ();
 sg13g2_decap_4 FILLER_62_1345 ();
 sg13g2_fill_2 FILLER_62_1354 ();
 sg13g2_fill_1 FILLER_62_1356 ();
 sg13g2_decap_8 FILLER_62_1362 ();
 sg13g2_decap_4 FILLER_62_1369 ();
 sg13g2_decap_4 FILLER_62_1378 ();
 sg13g2_fill_2 FILLER_62_1382 ();
 sg13g2_decap_4 FILLER_62_1387 ();
 sg13g2_fill_1 FILLER_62_1391 ();
 sg13g2_decap_4 FILLER_62_1402 ();
 sg13g2_fill_2 FILLER_62_1406 ();
 sg13g2_fill_2 FILLER_62_1417 ();
 sg13g2_decap_8 FILLER_62_1422 ();
 sg13g2_decap_4 FILLER_62_1429 ();
 sg13g2_fill_1 FILLER_62_1433 ();
 sg13g2_fill_1 FILLER_62_1446 ();
 sg13g2_fill_2 FILLER_62_1452 ();
 sg13g2_fill_1 FILLER_62_1454 ();
 sg13g2_fill_2 FILLER_62_1460 ();
 sg13g2_fill_2 FILLER_62_1467 ();
 sg13g2_fill_1 FILLER_62_1483 ();
 sg13g2_fill_1 FILLER_62_1510 ();
 sg13g2_fill_1 FILLER_62_1516 ();
 sg13g2_fill_2 FILLER_62_1522 ();
 sg13g2_fill_2 FILLER_62_1528 ();
 sg13g2_fill_2 FILLER_62_1540 ();
 sg13g2_fill_1 FILLER_62_1542 ();
 sg13g2_decap_4 FILLER_62_1551 ();
 sg13g2_decap_8 FILLER_62_1559 ();
 sg13g2_decap_4 FILLER_62_1566 ();
 sg13g2_fill_2 FILLER_62_1570 ();
 sg13g2_fill_1 FILLER_62_1585 ();
 sg13g2_decap_8 FILLER_62_1593 ();
 sg13g2_fill_2 FILLER_62_1600 ();
 sg13g2_decap_4 FILLER_62_1607 ();
 sg13g2_fill_2 FILLER_62_1611 ();
 sg13g2_fill_1 FILLER_62_1616 ();
 sg13g2_fill_1 FILLER_62_1622 ();
 sg13g2_decap_8 FILLER_62_1663 ();
 sg13g2_decap_4 FILLER_62_1670 ();
 sg13g2_fill_2 FILLER_62_1674 ();
 sg13g2_fill_1 FILLER_62_1705 ();
 sg13g2_decap_8 FILLER_62_1710 ();
 sg13g2_decap_8 FILLER_62_1717 ();
 sg13g2_decap_8 FILLER_62_1724 ();
 sg13g2_decap_4 FILLER_62_1731 ();
 sg13g2_fill_1 FILLER_62_1747 ();
 sg13g2_decap_4 FILLER_62_1765 ();
 sg13g2_fill_2 FILLER_62_1806 ();
 sg13g2_fill_1 FILLER_62_1808 ();
 sg13g2_fill_2 FILLER_62_1830 ();
 sg13g2_fill_1 FILLER_62_1843 ();
 sg13g2_fill_1 FILLER_62_1852 ();
 sg13g2_decap_8 FILLER_62_1858 ();
 sg13g2_decap_8 FILLER_62_1865 ();
 sg13g2_fill_2 FILLER_62_1872 ();
 sg13g2_fill_1 FILLER_62_1874 ();
 sg13g2_fill_1 FILLER_62_1887 ();
 sg13g2_fill_2 FILLER_62_1893 ();
 sg13g2_fill_1 FILLER_62_1899 ();
 sg13g2_fill_2 FILLER_62_1905 ();
 sg13g2_fill_2 FILLER_62_1928 ();
 sg13g2_fill_1 FILLER_62_1930 ();
 sg13g2_decap_4 FILLER_62_1935 ();
 sg13g2_fill_1 FILLER_62_1939 ();
 sg13g2_decap_8 FILLER_62_1944 ();
 sg13g2_decap_8 FILLER_62_1951 ();
 sg13g2_fill_2 FILLER_62_1958 ();
 sg13g2_decap_8 FILLER_62_1973 ();
 sg13g2_decap_8 FILLER_62_1980 ();
 sg13g2_decap_8 FILLER_62_1987 ();
 sg13g2_decap_4 FILLER_62_1994 ();
 sg13g2_fill_2 FILLER_62_1998 ();
 sg13g2_decap_8 FILLER_62_2015 ();
 sg13g2_fill_2 FILLER_62_2037 ();
 sg13g2_decap_4 FILLER_62_2073 ();
 sg13g2_fill_2 FILLER_62_2077 ();
 sg13g2_fill_2 FILLER_62_2088 ();
 sg13g2_fill_2 FILLER_62_2118 ();
 sg13g2_fill_1 FILLER_62_2130 ();
 sg13g2_fill_2 FILLER_62_2136 ();
 sg13g2_fill_1 FILLER_62_2143 ();
 sg13g2_fill_2 FILLER_62_2148 ();
 sg13g2_decap_8 FILLER_62_2154 ();
 sg13g2_decap_8 FILLER_62_2161 ();
 sg13g2_decap_8 FILLER_62_2168 ();
 sg13g2_decap_8 FILLER_62_2175 ();
 sg13g2_decap_8 FILLER_62_2182 ();
 sg13g2_fill_2 FILLER_62_2189 ();
 sg13g2_decap_4 FILLER_62_2217 ();
 sg13g2_fill_1 FILLER_62_2221 ();
 sg13g2_fill_2 FILLER_62_2238 ();
 sg13g2_fill_1 FILLER_62_2240 ();
 sg13g2_fill_1 FILLER_62_2249 ();
 sg13g2_fill_2 FILLER_62_2263 ();
 sg13g2_fill_2 FILLER_62_2268 ();
 sg13g2_fill_1 FILLER_62_2270 ();
 sg13g2_decap_4 FILLER_62_2276 ();
 sg13g2_fill_1 FILLER_62_2280 ();
 sg13g2_fill_2 FILLER_62_2291 ();
 sg13g2_fill_1 FILLER_62_2293 ();
 sg13g2_fill_2 FILLER_62_2298 ();
 sg13g2_fill_1 FILLER_62_2300 ();
 sg13g2_fill_2 FILLER_62_2305 ();
 sg13g2_fill_1 FILLER_62_2307 ();
 sg13g2_decap_4 FILLER_62_2334 ();
 sg13g2_fill_2 FILLER_62_2338 ();
 sg13g2_decap_4 FILLER_62_2377 ();
 sg13g2_fill_2 FILLER_62_2381 ();
 sg13g2_decap_4 FILLER_62_2408 ();
 sg13g2_fill_1 FILLER_62_2421 ();
 sg13g2_fill_1 FILLER_62_2479 ();
 sg13g2_decap_4 FILLER_62_2515 ();
 sg13g2_fill_1 FILLER_62_2523 ();
 sg13g2_fill_2 FILLER_62_2554 ();
 sg13g2_fill_1 FILLER_62_2561 ();
 sg13g2_fill_1 FILLER_62_2566 ();
 sg13g2_fill_1 FILLER_62_2593 ();
 sg13g2_fill_1 FILLER_62_2604 ();
 sg13g2_decap_4 FILLER_62_2615 ();
 sg13g2_decap_8 FILLER_62_2627 ();
 sg13g2_decap_8 FILLER_62_2634 ();
 sg13g2_decap_8 FILLER_62_2641 ();
 sg13g2_decap_8 FILLER_62_2648 ();
 sg13g2_decap_8 FILLER_62_2655 ();
 sg13g2_decap_8 FILLER_62_2662 ();
 sg13g2_fill_1 FILLER_62_2669 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_fill_1 FILLER_63_14 ();
 sg13g2_fill_1 FILLER_63_62 ();
 sg13g2_fill_2 FILLER_63_67 ();
 sg13g2_fill_1 FILLER_63_100 ();
 sg13g2_fill_1 FILLER_63_106 ();
 sg13g2_fill_2 FILLER_63_145 ();
 sg13g2_fill_1 FILLER_63_152 ();
 sg13g2_fill_2 FILLER_63_157 ();
 sg13g2_fill_1 FILLER_63_159 ();
 sg13g2_decap_8 FILLER_63_164 ();
 sg13g2_decap_4 FILLER_63_171 ();
 sg13g2_fill_2 FILLER_63_179 ();
 sg13g2_fill_1 FILLER_63_181 ();
 sg13g2_fill_2 FILLER_63_244 ();
 sg13g2_fill_1 FILLER_63_246 ();
 sg13g2_fill_2 FILLER_63_315 ();
 sg13g2_fill_2 FILLER_63_336 ();
 sg13g2_fill_2 FILLER_63_371 ();
 sg13g2_fill_2 FILLER_63_423 ();
 sg13g2_fill_1 FILLER_63_431 ();
 sg13g2_fill_1 FILLER_63_436 ();
 sg13g2_fill_1 FILLER_63_442 ();
 sg13g2_fill_1 FILLER_63_479 ();
 sg13g2_fill_1 FILLER_63_494 ();
 sg13g2_fill_1 FILLER_63_500 ();
 sg13g2_fill_1 FILLER_63_520 ();
 sg13g2_fill_1 FILLER_63_525 ();
 sg13g2_fill_1 FILLER_63_531 ();
 sg13g2_fill_1 FILLER_63_558 ();
 sg13g2_fill_1 FILLER_63_568 ();
 sg13g2_fill_2 FILLER_63_574 ();
 sg13g2_fill_1 FILLER_63_576 ();
 sg13g2_decap_8 FILLER_63_581 ();
 sg13g2_fill_2 FILLER_63_588 ();
 sg13g2_fill_1 FILLER_63_590 ();
 sg13g2_decap_4 FILLER_63_605 ();
 sg13g2_fill_2 FILLER_63_615 ();
 sg13g2_fill_1 FILLER_63_622 ();
 sg13g2_fill_1 FILLER_63_652 ();
 sg13g2_fill_1 FILLER_63_707 ();
 sg13g2_decap_4 FILLER_63_721 ();
 sg13g2_fill_2 FILLER_63_725 ();
 sg13g2_fill_1 FILLER_63_735 ();
 sg13g2_fill_2 FILLER_63_742 ();
 sg13g2_fill_2 FILLER_63_750 ();
 sg13g2_fill_2 FILLER_63_757 ();
 sg13g2_fill_1 FILLER_63_766 ();
 sg13g2_decap_4 FILLER_63_780 ();
 sg13g2_fill_2 FILLER_63_794 ();
 sg13g2_fill_1 FILLER_63_796 ();
 sg13g2_fill_1 FILLER_63_826 ();
 sg13g2_fill_1 FILLER_63_872 ();
 sg13g2_fill_1 FILLER_63_883 ();
 sg13g2_fill_1 FILLER_63_894 ();
 sg13g2_fill_1 FILLER_63_940 ();
 sg13g2_fill_2 FILLER_63_1006 ();
 sg13g2_decap_8 FILLER_63_1039 ();
 sg13g2_decap_4 FILLER_63_1046 ();
 sg13g2_fill_1 FILLER_63_1050 ();
 sg13g2_fill_2 FILLER_63_1055 ();
 sg13g2_fill_1 FILLER_63_1057 ();
 sg13g2_decap_8 FILLER_63_1115 ();
 sg13g2_decap_8 FILLER_63_1122 ();
 sg13g2_fill_2 FILLER_63_1133 ();
 sg13g2_decap_8 FILLER_63_1165 ();
 sg13g2_decap_8 FILLER_63_1172 ();
 sg13g2_decap_8 FILLER_63_1179 ();
 sg13g2_fill_2 FILLER_63_1186 ();
 sg13g2_decap_8 FILLER_63_1221 ();
 sg13g2_fill_1 FILLER_63_1228 ();
 sg13g2_decap_8 FILLER_63_1247 ();
 sg13g2_decap_8 FILLER_63_1254 ();
 sg13g2_decap_8 FILLER_63_1261 ();
 sg13g2_decap_4 FILLER_63_1268 ();
 sg13g2_fill_1 FILLER_63_1272 ();
 sg13g2_fill_1 FILLER_63_1288 ();
 sg13g2_fill_2 FILLER_63_1300 ();
 sg13g2_fill_2 FILLER_63_1329 ();
 sg13g2_fill_1 FILLER_63_1331 ();
 sg13g2_fill_1 FILLER_63_1346 ();
 sg13g2_decap_8 FILLER_63_1353 ();
 sg13g2_decap_8 FILLER_63_1360 ();
 sg13g2_decap_8 FILLER_63_1367 ();
 sg13g2_fill_1 FILLER_63_1396 ();
 sg13g2_fill_2 FILLER_63_1404 ();
 sg13g2_fill_1 FILLER_63_1422 ();
 sg13g2_fill_2 FILLER_63_1432 ();
 sg13g2_fill_2 FILLER_63_1444 ();
 sg13g2_fill_1 FILLER_63_1526 ();
 sg13g2_fill_2 FILLER_63_1532 ();
 sg13g2_fill_1 FILLER_63_1547 ();
 sg13g2_fill_2 FILLER_63_1574 ();
 sg13g2_fill_2 FILLER_63_1580 ();
 sg13g2_fill_1 FILLER_63_1585 ();
 sg13g2_fill_2 FILLER_63_1609 ();
 sg13g2_fill_2 FILLER_63_1653 ();
 sg13g2_fill_1 FILLER_63_1655 ();
 sg13g2_fill_2 FILLER_63_1682 ();
 sg13g2_decap_8 FILLER_63_1697 ();
 sg13g2_decap_4 FILLER_63_1704 ();
 sg13g2_fill_2 FILLER_63_1708 ();
 sg13g2_decap_4 FILLER_63_1714 ();
 sg13g2_fill_1 FILLER_63_1722 ();
 sg13g2_fill_1 FILLER_63_1735 ();
 sg13g2_fill_2 FILLER_63_1760 ();
 sg13g2_fill_1 FILLER_63_1768 ();
 sg13g2_decap_4 FILLER_63_1782 ();
 sg13g2_fill_1 FILLER_63_1806 ();
 sg13g2_fill_1 FILLER_63_1815 ();
 sg13g2_fill_1 FILLER_63_1829 ();
 sg13g2_fill_2 FILLER_63_1840 ();
 sg13g2_decap_8 FILLER_63_1851 ();
 sg13g2_decap_8 FILLER_63_1858 ();
 sg13g2_decap_8 FILLER_63_1865 ();
 sg13g2_fill_2 FILLER_63_1872 ();
 sg13g2_decap_8 FILLER_63_1932 ();
 sg13g2_decap_8 FILLER_63_1939 ();
 sg13g2_decap_8 FILLER_63_1946 ();
 sg13g2_fill_2 FILLER_63_1953 ();
 sg13g2_fill_1 FILLER_63_1955 ();
 sg13g2_decap_8 FILLER_63_1960 ();
 sg13g2_decap_4 FILLER_63_1971 ();
 sg13g2_fill_2 FILLER_63_1975 ();
 sg13g2_fill_2 FILLER_63_2012 ();
 sg13g2_fill_1 FILLER_63_2014 ();
 sg13g2_fill_2 FILLER_63_2028 ();
 sg13g2_fill_1 FILLER_63_2030 ();
 sg13g2_fill_2 FILLER_63_2036 ();
 sg13g2_fill_2 FILLER_63_2049 ();
 sg13g2_fill_1 FILLER_63_2051 ();
 sg13g2_fill_1 FILLER_63_2070 ();
 sg13g2_decap_4 FILLER_63_2076 ();
 sg13g2_fill_2 FILLER_63_2080 ();
 sg13g2_fill_1 FILLER_63_2100 ();
 sg13g2_fill_2 FILLER_63_2111 ();
 sg13g2_fill_1 FILLER_63_2113 ();
 sg13g2_fill_1 FILLER_63_2127 ();
 sg13g2_decap_8 FILLER_63_2150 ();
 sg13g2_decap_8 FILLER_63_2157 ();
 sg13g2_decap_8 FILLER_63_2164 ();
 sg13g2_decap_8 FILLER_63_2171 ();
 sg13g2_decap_8 FILLER_63_2178 ();
 sg13g2_decap_4 FILLER_63_2185 ();
 sg13g2_decap_4 FILLER_63_2229 ();
 sg13g2_fill_2 FILLER_63_2233 ();
 sg13g2_decap_4 FILLER_63_2240 ();
 sg13g2_decap_4 FILLER_63_2276 ();
 sg13g2_fill_2 FILLER_63_2280 ();
 sg13g2_fill_1 FILLER_63_2291 ();
 sg13g2_fill_1 FILLER_63_2300 ();
 sg13g2_fill_2 FILLER_63_2333 ();
 sg13g2_decap_4 FILLER_63_2344 ();
 sg13g2_fill_1 FILLER_63_2348 ();
 sg13g2_fill_1 FILLER_63_2353 ();
 sg13g2_fill_1 FILLER_63_2358 ();
 sg13g2_fill_2 FILLER_63_2368 ();
 sg13g2_decap_8 FILLER_63_2374 ();
 sg13g2_fill_1 FILLER_63_2381 ();
 sg13g2_decap_4 FILLER_63_2412 ();
 sg13g2_fill_2 FILLER_63_2424 ();
 sg13g2_fill_1 FILLER_63_2426 ();
 sg13g2_fill_2 FILLER_63_2431 ();
 sg13g2_fill_2 FILLER_63_2437 ();
 sg13g2_fill_2 FILLER_63_2444 ();
 sg13g2_fill_1 FILLER_63_2446 ();
 sg13g2_fill_1 FILLER_63_2451 ();
 sg13g2_fill_2 FILLER_63_2457 ();
 sg13g2_fill_1 FILLER_63_2459 ();
 sg13g2_fill_1 FILLER_63_2468 ();
 sg13g2_decap_4 FILLER_63_2473 ();
 sg13g2_fill_2 FILLER_63_2477 ();
 sg13g2_fill_1 FILLER_63_2484 ();
 sg13g2_decap_4 FILLER_63_2494 ();
 sg13g2_fill_1 FILLER_63_2498 ();
 sg13g2_fill_1 FILLER_63_2508 ();
 sg13g2_fill_2 FILLER_63_2518 ();
 sg13g2_fill_1 FILLER_63_2520 ();
 sg13g2_fill_2 FILLER_63_2525 ();
 sg13g2_fill_1 FILLER_63_2531 ();
 sg13g2_fill_1 FILLER_63_2536 ();
 sg13g2_decap_8 FILLER_63_2546 ();
 sg13g2_decap_8 FILLER_63_2553 ();
 sg13g2_decap_8 FILLER_63_2560 ();
 sg13g2_fill_2 FILLER_63_2567 ();
 sg13g2_fill_1 FILLER_63_2569 ();
 sg13g2_decap_4 FILLER_63_2579 ();
 sg13g2_fill_1 FILLER_63_2583 ();
 sg13g2_decap_8 FILLER_63_2630 ();
 sg13g2_decap_8 FILLER_63_2637 ();
 sg13g2_decap_8 FILLER_63_2644 ();
 sg13g2_decap_8 FILLER_63_2651 ();
 sg13g2_decap_8 FILLER_63_2658 ();
 sg13g2_decap_4 FILLER_63_2665 ();
 sg13g2_fill_1 FILLER_63_2669 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_4 FILLER_64_7 ();
 sg13g2_decap_4 FILLER_64_15 ();
 sg13g2_fill_1 FILLER_64_24 ();
 sg13g2_fill_1 FILLER_64_35 ();
 sg13g2_fill_1 FILLER_64_41 ();
 sg13g2_decap_4 FILLER_64_50 ();
 sg13g2_fill_1 FILLER_64_54 ();
 sg13g2_decap_4 FILLER_64_59 ();
 sg13g2_fill_2 FILLER_64_63 ();
 sg13g2_decap_4 FILLER_64_87 ();
 sg13g2_decap_8 FILLER_64_126 ();
 sg13g2_decap_8 FILLER_64_133 ();
 sg13g2_decap_8 FILLER_64_140 ();
 sg13g2_decap_8 FILLER_64_147 ();
 sg13g2_decap_8 FILLER_64_154 ();
 sg13g2_decap_8 FILLER_64_161 ();
 sg13g2_decap_8 FILLER_64_168 ();
 sg13g2_fill_2 FILLER_64_175 ();
 sg13g2_fill_2 FILLER_64_192 ();
 sg13g2_fill_1 FILLER_64_194 ();
 sg13g2_fill_1 FILLER_64_244 ();
 sg13g2_decap_8 FILLER_64_250 ();
 sg13g2_decap_4 FILLER_64_257 ();
 sg13g2_fill_1 FILLER_64_261 ();
 sg13g2_fill_1 FILLER_64_301 ();
 sg13g2_fill_1 FILLER_64_310 ();
 sg13g2_fill_1 FILLER_64_347 ();
 sg13g2_fill_2 FILLER_64_401 ();
 sg13g2_fill_1 FILLER_64_410 ();
 sg13g2_fill_1 FILLER_64_419 ();
 sg13g2_decap_8 FILLER_64_428 ();
 sg13g2_fill_1 FILLER_64_435 ();
 sg13g2_fill_2 FILLER_64_452 ();
 sg13g2_fill_1 FILLER_64_454 ();
 sg13g2_fill_1 FILLER_64_464 ();
 sg13g2_fill_2 FILLER_64_478 ();
 sg13g2_fill_1 FILLER_64_480 ();
 sg13g2_decap_4 FILLER_64_545 ();
 sg13g2_decap_8 FILLER_64_575 ();
 sg13g2_decap_8 FILLER_64_582 ();
 sg13g2_fill_2 FILLER_64_589 ();
 sg13g2_fill_1 FILLER_64_600 ();
 sg13g2_decap_4 FILLER_64_606 ();
 sg13g2_fill_1 FILLER_64_676 ();
 sg13g2_fill_1 FILLER_64_681 ();
 sg13g2_fill_2 FILLER_64_708 ();
 sg13g2_fill_2 FILLER_64_714 ();
 sg13g2_decap_8 FILLER_64_751 ();
 sg13g2_decap_8 FILLER_64_758 ();
 sg13g2_fill_2 FILLER_64_777 ();
 sg13g2_fill_1 FILLER_64_835 ();
 sg13g2_fill_2 FILLER_64_878 ();
 sg13g2_fill_1 FILLER_64_893 ();
 sg13g2_fill_1 FILLER_64_953 ();
 sg13g2_fill_2 FILLER_64_997 ();
 sg13g2_fill_2 FILLER_64_1008 ();
 sg13g2_fill_2 FILLER_64_1050 ();
 sg13g2_fill_1 FILLER_64_1082 ();
 sg13g2_decap_4 FILLER_64_1088 ();
 sg13g2_fill_2 FILLER_64_1122 ();
 sg13g2_fill_1 FILLER_64_1124 ();
 sg13g2_fill_2 FILLER_64_1130 ();
 sg13g2_fill_1 FILLER_64_1132 ();
 sg13g2_decap_8 FILLER_64_1143 ();
 sg13g2_fill_1 FILLER_64_1150 ();
 sg13g2_decap_4 FILLER_64_1157 ();
 sg13g2_decap_8 FILLER_64_1165 ();
 sg13g2_decap_8 FILLER_64_1172 ();
 sg13g2_decap_8 FILLER_64_1179 ();
 sg13g2_decap_8 FILLER_64_1186 ();
 sg13g2_decap_8 FILLER_64_1193 ();
 sg13g2_fill_1 FILLER_64_1200 ();
 sg13g2_decap_8 FILLER_64_1205 ();
 sg13g2_decap_4 FILLER_64_1212 ();
 sg13g2_decap_8 FILLER_64_1256 ();
 sg13g2_decap_4 FILLER_64_1263 ();
 sg13g2_fill_1 FILLER_64_1267 ();
 sg13g2_fill_1 FILLER_64_1326 ();
 sg13g2_decap_8 FILLER_64_1355 ();
 sg13g2_fill_2 FILLER_64_1362 ();
 sg13g2_fill_1 FILLER_64_1364 ();
 sg13g2_fill_2 FILLER_64_1378 ();
 sg13g2_fill_1 FILLER_64_1389 ();
 sg13g2_fill_1 FILLER_64_1400 ();
 sg13g2_fill_1 FILLER_64_1410 ();
 sg13g2_decap_8 FILLER_64_1423 ();
 sg13g2_fill_1 FILLER_64_1456 ();
 sg13g2_fill_2 FILLER_64_1465 ();
 sg13g2_fill_1 FILLER_64_1477 ();
 sg13g2_fill_1 FILLER_64_1482 ();
 sg13g2_decap_8 FILLER_64_1554 ();
 sg13g2_decap_8 FILLER_64_1561 ();
 sg13g2_decap_4 FILLER_64_1568 ();
 sg13g2_fill_2 FILLER_64_1576 ();
 sg13g2_fill_1 FILLER_64_1578 ();
 sg13g2_fill_1 FILLER_64_1589 ();
 sg13g2_fill_1 FILLER_64_1593 ();
 sg13g2_decap_8 FILLER_64_1613 ();
 sg13g2_fill_2 FILLER_64_1620 ();
 sg13g2_fill_1 FILLER_64_1622 ();
 sg13g2_fill_2 FILLER_64_1632 ();
 sg13g2_fill_1 FILLER_64_1634 ();
 sg13g2_fill_2 FILLER_64_1638 ();
 sg13g2_decap_8 FILLER_64_1650 ();
 sg13g2_decap_8 FILLER_64_1657 ();
 sg13g2_decap_4 FILLER_64_1664 ();
 sg13g2_decap_8 FILLER_64_1671 ();
 sg13g2_decap_8 FILLER_64_1678 ();
 sg13g2_decap_4 FILLER_64_1685 ();
 sg13g2_fill_2 FILLER_64_1689 ();
 sg13g2_decap_4 FILLER_64_1765 ();
 sg13g2_fill_2 FILLER_64_1769 ();
 sg13g2_fill_1 FILLER_64_1775 ();
 sg13g2_fill_1 FILLER_64_1782 ();
 sg13g2_fill_1 FILLER_64_1788 ();
 sg13g2_fill_1 FILLER_64_1797 ();
 sg13g2_fill_1 FILLER_64_1803 ();
 sg13g2_fill_2 FILLER_64_1809 ();
 sg13g2_fill_1 FILLER_64_1820 ();
 sg13g2_fill_2 FILLER_64_1826 ();
 sg13g2_fill_1 FILLER_64_1843 ();
 sg13g2_decap_4 FILLER_64_1849 ();
 sg13g2_fill_2 FILLER_64_1853 ();
 sg13g2_decap_8 FILLER_64_1860 ();
 sg13g2_decap_4 FILLER_64_1867 ();
 sg13g2_fill_1 FILLER_64_1871 ();
 sg13g2_fill_1 FILLER_64_1877 ();
 sg13g2_fill_2 FILLER_64_1882 ();
 sg13g2_fill_1 FILLER_64_1901 ();
 sg13g2_fill_1 FILLER_64_1907 ();
 sg13g2_fill_1 FILLER_64_1913 ();
 sg13g2_fill_1 FILLER_64_1919 ();
 sg13g2_decap_8 FILLER_64_1925 ();
 sg13g2_decap_4 FILLER_64_1932 ();
 sg13g2_decap_8 FILLER_64_1945 ();
 sg13g2_decap_8 FILLER_64_1961 ();
 sg13g2_fill_2 FILLER_64_1972 ();
 sg13g2_decap_4 FILLER_64_1979 ();
 sg13g2_fill_1 FILLER_64_1983 ();
 sg13g2_decap_8 FILLER_64_1988 ();
 sg13g2_fill_2 FILLER_64_1999 ();
 sg13g2_fill_1 FILLER_64_2001 ();
 sg13g2_decap_8 FILLER_64_2014 ();
 sg13g2_fill_2 FILLER_64_2021 ();
 sg13g2_fill_1 FILLER_64_2037 ();
 sg13g2_fill_2 FILLER_64_2042 ();
 sg13g2_fill_1 FILLER_64_2048 ();
 sg13g2_fill_2 FILLER_64_2053 ();
 sg13g2_fill_2 FILLER_64_2060 ();
 sg13g2_fill_2 FILLER_64_2066 ();
 sg13g2_fill_1 FILLER_64_2072 ();
 sg13g2_fill_1 FILLER_64_2077 ();
 sg13g2_fill_1 FILLER_64_2088 ();
 sg13g2_fill_2 FILLER_64_2097 ();
 sg13g2_fill_2 FILLER_64_2137 ();
 sg13g2_fill_1 FILLER_64_2159 ();
 sg13g2_decap_8 FILLER_64_2170 ();
 sg13g2_decap_8 FILLER_64_2177 ();
 sg13g2_fill_1 FILLER_64_2228 ();
 sg13g2_fill_2 FILLER_64_2300 ();
 sg13g2_fill_1 FILLER_64_2306 ();
 sg13g2_decap_8 FILLER_64_2321 ();
 sg13g2_decap_8 FILLER_64_2363 ();
 sg13g2_decap_4 FILLER_64_2370 ();
 sg13g2_fill_1 FILLER_64_2405 ();
 sg13g2_decap_8 FILLER_64_2414 ();
 sg13g2_decap_8 FILLER_64_2421 ();
 sg13g2_decap_4 FILLER_64_2428 ();
 sg13g2_fill_2 FILLER_64_2432 ();
 sg13g2_fill_1 FILLER_64_2444 ();
 sg13g2_fill_2 FILLER_64_2479 ();
 sg13g2_fill_2 FILLER_64_2485 ();
 sg13g2_fill_1 FILLER_64_2487 ();
 sg13g2_fill_1 FILLER_64_2493 ();
 sg13g2_fill_1 FILLER_64_2498 ();
 sg13g2_fill_1 FILLER_64_2537 ();
 sg13g2_decap_4 FILLER_64_2568 ();
 sg13g2_decap_8 FILLER_64_2633 ();
 sg13g2_decap_8 FILLER_64_2640 ();
 sg13g2_decap_8 FILLER_64_2647 ();
 sg13g2_decap_8 FILLER_64_2654 ();
 sg13g2_decap_8 FILLER_64_2661 ();
 sg13g2_fill_2 FILLER_64_2668 ();
 sg13g2_fill_2 FILLER_65_0 ();
 sg13g2_fill_2 FILLER_65_32 ();
 sg13g2_decap_8 FILLER_65_41 ();
 sg13g2_fill_1 FILLER_65_48 ();
 sg13g2_fill_2 FILLER_65_60 ();
 sg13g2_fill_1 FILLER_65_70 ();
 sg13g2_fill_1 FILLER_65_107 ();
 sg13g2_decap_8 FILLER_65_137 ();
 sg13g2_decap_8 FILLER_65_157 ();
 sg13g2_decap_8 FILLER_65_164 ();
 sg13g2_fill_1 FILLER_65_171 ();
 sg13g2_fill_2 FILLER_65_190 ();
 sg13g2_fill_2 FILLER_65_200 ();
 sg13g2_fill_1 FILLER_65_202 ();
 sg13g2_fill_2 FILLER_65_212 ();
 sg13g2_decap_8 FILLER_65_218 ();
 sg13g2_decap_4 FILLER_65_225 ();
 sg13g2_fill_1 FILLER_65_229 ();
 sg13g2_decap_8 FILLER_65_240 ();
 sg13g2_decap_8 FILLER_65_247 ();
 sg13g2_decap_8 FILLER_65_254 ();
 sg13g2_fill_2 FILLER_65_266 ();
 sg13g2_fill_1 FILLER_65_287 ();
 sg13g2_fill_2 FILLER_65_309 ();
 sg13g2_fill_1 FILLER_65_330 ();
 sg13g2_fill_2 FILLER_65_336 ();
 sg13g2_fill_1 FILLER_65_351 ();
 sg13g2_fill_2 FILLER_65_355 ();
 sg13g2_fill_1 FILLER_65_391 ();
 sg13g2_fill_1 FILLER_65_410 ();
 sg13g2_decap_8 FILLER_65_419 ();
 sg13g2_fill_2 FILLER_65_431 ();
 sg13g2_decap_8 FILLER_65_445 ();
 sg13g2_decap_8 FILLER_65_452 ();
 sg13g2_decap_8 FILLER_65_459 ();
 sg13g2_fill_1 FILLER_65_466 ();
 sg13g2_decap_4 FILLER_65_472 ();
 sg13g2_decap_8 FILLER_65_532 ();
 sg13g2_decap_8 FILLER_65_539 ();
 sg13g2_decap_4 FILLER_65_546 ();
 sg13g2_fill_2 FILLER_65_577 ();
 sg13g2_fill_1 FILLER_65_610 ();
 sg13g2_decap_8 FILLER_65_615 ();
 sg13g2_decap_4 FILLER_65_622 ();
 sg13g2_fill_1 FILLER_65_634 ();
 sg13g2_fill_1 FILLER_65_640 ();
 sg13g2_fill_2 FILLER_65_646 ();
 sg13g2_fill_1 FILLER_65_648 ();
 sg13g2_fill_1 FILLER_65_669 ();
 sg13g2_fill_1 FILLER_65_678 ();
 sg13g2_decap_8 FILLER_65_683 ();
 sg13g2_fill_1 FILLER_65_690 ();
 sg13g2_fill_1 FILLER_65_695 ();
 sg13g2_decap_8 FILLER_65_699 ();
 sg13g2_decap_4 FILLER_65_706 ();
 sg13g2_fill_2 FILLER_65_714 ();
 sg13g2_fill_1 FILLER_65_716 ();
 sg13g2_decap_8 FILLER_65_721 ();
 sg13g2_decap_4 FILLER_65_728 ();
 sg13g2_fill_2 FILLER_65_732 ();
 sg13g2_decap_4 FILLER_65_740 ();
 sg13g2_fill_1 FILLER_65_744 ();
 sg13g2_decap_8 FILLER_65_759 ();
 sg13g2_decap_4 FILLER_65_766 ();
 sg13g2_fill_2 FILLER_65_770 ();
 sg13g2_fill_1 FILLER_65_796 ();
 sg13g2_decap_4 FILLER_65_805 ();
 sg13g2_decap_8 FILLER_65_812 ();
 sg13g2_fill_1 FILLER_65_819 ();
 sg13g2_fill_1 FILLER_65_862 ();
 sg13g2_fill_1 FILLER_65_898 ();
 sg13g2_fill_2 FILLER_65_912 ();
 sg13g2_fill_2 FILLER_65_955 ();
 sg13g2_fill_2 FILLER_65_961 ();
 sg13g2_fill_2 FILLER_65_972 ();
 sg13g2_fill_2 FILLER_65_978 ();
 sg13g2_fill_2 FILLER_65_984 ();
 sg13g2_fill_2 FILLER_65_990 ();
 sg13g2_fill_2 FILLER_65_1000 ();
 sg13g2_fill_1 FILLER_65_1002 ();
 sg13g2_decap_4 FILLER_65_1007 ();
 sg13g2_fill_2 FILLER_65_1011 ();
 sg13g2_decap_4 FILLER_65_1017 ();
 sg13g2_decap_8 FILLER_65_1030 ();
 sg13g2_decap_8 FILLER_65_1037 ();
 sg13g2_decap_4 FILLER_65_1044 ();
 sg13g2_fill_2 FILLER_65_1058 ();
 sg13g2_decap_4 FILLER_65_1074 ();
 sg13g2_fill_1 FILLER_65_1078 ();
 sg13g2_fill_1 FILLER_65_1084 ();
 sg13g2_decap_4 FILLER_65_1095 ();
 sg13g2_fill_1 FILLER_65_1099 ();
 sg13g2_fill_2 FILLER_65_1105 ();
 sg13g2_fill_1 FILLER_65_1107 ();
 sg13g2_fill_1 FILLER_65_1113 ();
 sg13g2_decap_8 FILLER_65_1124 ();
 sg13g2_fill_1 FILLER_65_1135 ();
 sg13g2_fill_1 FILLER_65_1146 ();
 sg13g2_fill_1 FILLER_65_1156 ();
 sg13g2_decap_4 FILLER_65_1161 ();
 sg13g2_fill_2 FILLER_65_1165 ();
 sg13g2_fill_2 FILLER_65_1172 ();
 sg13g2_fill_1 FILLER_65_1174 ();
 sg13g2_decap_8 FILLER_65_1206 ();
 sg13g2_decap_8 FILLER_65_1213 ();
 sg13g2_fill_1 FILLER_65_1220 ();
 sg13g2_fill_1 FILLER_65_1231 ();
 sg13g2_decap_4 FILLER_65_1262 ();
 sg13g2_fill_1 FILLER_65_1266 ();
 sg13g2_fill_1 FILLER_65_1291 ();
 sg13g2_fill_1 FILLER_65_1311 ();
 sg13g2_fill_1 FILLER_65_1318 ();
 sg13g2_fill_1 FILLER_65_1330 ();
 sg13g2_fill_2 FILLER_65_1355 ();
 sg13g2_fill_2 FILLER_65_1366 ();
 sg13g2_fill_2 FILLER_65_1396 ();
 sg13g2_decap_4 FILLER_65_1420 ();
 sg13g2_fill_1 FILLER_65_1424 ();
 sg13g2_fill_2 FILLER_65_1447 ();
 sg13g2_fill_1 FILLER_65_1471 ();
 sg13g2_fill_1 FILLER_65_1494 ();
 sg13g2_fill_2 FILLER_65_1505 ();
 sg13g2_fill_1 FILLER_65_1507 ();
 sg13g2_decap_4 FILLER_65_1519 ();
 sg13g2_fill_1 FILLER_65_1523 ();
 sg13g2_decap_8 FILLER_65_1529 ();
 sg13g2_fill_1 FILLER_65_1536 ();
 sg13g2_decap_8 FILLER_65_1571 ();
 sg13g2_fill_2 FILLER_65_1578 ();
 sg13g2_fill_1 FILLER_65_1580 ();
 sg13g2_fill_1 FILLER_65_1585 ();
 sg13g2_fill_2 FILLER_65_1599 ();
 sg13g2_fill_2 FILLER_65_1627 ();
 sg13g2_fill_1 FILLER_65_1629 ();
 sg13g2_fill_2 FILLER_65_1643 ();
 sg13g2_decap_4 FILLER_65_1662 ();
 sg13g2_fill_2 FILLER_65_1666 ();
 sg13g2_decap_8 FILLER_65_1678 ();
 sg13g2_decap_4 FILLER_65_1685 ();
 sg13g2_decap_8 FILLER_65_1699 ();
 sg13g2_decap_8 FILLER_65_1706 ();
 sg13g2_fill_1 FILLER_65_1713 ();
 sg13g2_fill_1 FILLER_65_1719 ();
 sg13g2_fill_1 FILLER_65_1729 ();
 sg13g2_fill_1 FILLER_65_1735 ();
 sg13g2_fill_2 FILLER_65_1749 ();
 sg13g2_fill_1 FILLER_65_1756 ();
 sg13g2_fill_1 FILLER_65_1762 ();
 sg13g2_fill_2 FILLER_65_1771 ();
 sg13g2_fill_1 FILLER_65_1773 ();
 sg13g2_fill_2 FILLER_65_1777 ();
 sg13g2_fill_1 FILLER_65_1779 ();
 sg13g2_fill_1 FILLER_65_1799 ();
 sg13g2_decap_8 FILLER_65_1808 ();
 sg13g2_decap_4 FILLER_65_1815 ();
 sg13g2_decap_8 FILLER_65_1844 ();
 sg13g2_fill_2 FILLER_65_1851 ();
 sg13g2_decap_8 FILLER_65_1866 ();
 sg13g2_fill_2 FILLER_65_1873 ();
 sg13g2_decap_8 FILLER_65_1879 ();
 sg13g2_decap_8 FILLER_65_1886 ();
 sg13g2_fill_1 FILLER_65_1893 ();
 sg13g2_fill_2 FILLER_65_1916 ();
 sg13g2_fill_1 FILLER_65_1918 ();
 sg13g2_decap_8 FILLER_65_1963 ();
 sg13g2_fill_1 FILLER_65_1970 ();
 sg13g2_decap_8 FILLER_65_1975 ();
 sg13g2_fill_1 FILLER_65_1982 ();
 sg13g2_fill_1 FILLER_65_1991 ();
 sg13g2_fill_1 FILLER_65_1997 ();
 sg13g2_fill_1 FILLER_65_2002 ();
 sg13g2_fill_2 FILLER_65_2007 ();
 sg13g2_fill_1 FILLER_65_2025 ();
 sg13g2_decap_8 FILLER_65_2036 ();
 sg13g2_fill_2 FILLER_65_2043 ();
 sg13g2_decap_4 FILLER_65_2055 ();
 sg13g2_fill_1 FILLER_65_2063 ();
 sg13g2_fill_1 FILLER_65_2073 ();
 sg13g2_fill_2 FILLER_65_2085 ();
 sg13g2_fill_1 FILLER_65_2126 ();
 sg13g2_fill_1 FILLER_65_2133 ();
 sg13g2_fill_1 FILLER_65_2167 ();
 sg13g2_fill_1 FILLER_65_2194 ();
 sg13g2_fill_2 FILLER_65_2199 ();
 sg13g2_fill_1 FILLER_65_2217 ();
 sg13g2_fill_1 FILLER_65_2223 ();
 sg13g2_fill_2 FILLER_65_2229 ();
 sg13g2_fill_1 FILLER_65_2239 ();
 sg13g2_fill_1 FILLER_65_2251 ();
 sg13g2_fill_2 FILLER_65_2270 ();
 sg13g2_fill_1 FILLER_65_2276 ();
 sg13g2_fill_1 FILLER_65_2281 ();
 sg13g2_decap_4 FILLER_65_2314 ();
 sg13g2_decap_8 FILLER_65_2321 ();
 sg13g2_fill_1 FILLER_65_2394 ();
 sg13g2_fill_1 FILLER_65_2524 ();
 sg13g2_decap_8 FILLER_65_2529 ();
 sg13g2_fill_2 FILLER_65_2536 ();
 sg13g2_decap_4 FILLER_65_2542 ();
 sg13g2_fill_2 FILLER_65_2546 ();
 sg13g2_fill_2 FILLER_65_2583 ();
 sg13g2_fill_2 FILLER_65_2589 ();
 sg13g2_fill_1 FILLER_65_2591 ();
 sg13g2_decap_4 FILLER_65_2608 ();
 sg13g2_fill_2 FILLER_65_2616 ();
 sg13g2_fill_1 FILLER_65_2618 ();
 sg13g2_decap_8 FILLER_65_2623 ();
 sg13g2_decap_8 FILLER_65_2630 ();
 sg13g2_decap_8 FILLER_65_2637 ();
 sg13g2_decap_8 FILLER_65_2644 ();
 sg13g2_decap_8 FILLER_65_2651 ();
 sg13g2_decap_8 FILLER_65_2658 ();
 sg13g2_decap_4 FILLER_65_2665 ();
 sg13g2_fill_1 FILLER_65_2669 ();
 sg13g2_fill_2 FILLER_66_0 ();
 sg13g2_fill_1 FILLER_66_28 ();
 sg13g2_decap_4 FILLER_66_33 ();
 sg13g2_fill_1 FILLER_66_37 ();
 sg13g2_decap_8 FILLER_66_65 ();
 sg13g2_fill_2 FILLER_66_72 ();
 sg13g2_fill_1 FILLER_66_104 ();
 sg13g2_decap_4 FILLER_66_114 ();
 sg13g2_decap_8 FILLER_66_122 ();
 sg13g2_decap_4 FILLER_66_129 ();
 sg13g2_fill_1 FILLER_66_133 ();
 sg13g2_decap_4 FILLER_66_138 ();
 sg13g2_decap_4 FILLER_66_217 ();
 sg13g2_fill_1 FILLER_66_221 ();
 sg13g2_decap_4 FILLER_66_226 ();
 sg13g2_decap_8 FILLER_66_260 ();
 sg13g2_fill_2 FILLER_66_267 ();
 sg13g2_fill_2 FILLER_66_275 ();
 sg13g2_fill_1 FILLER_66_283 ();
 sg13g2_fill_1 FILLER_66_297 ();
 sg13g2_fill_1 FILLER_66_328 ();
 sg13g2_fill_2 FILLER_66_360 ();
 sg13g2_fill_1 FILLER_66_365 ();
 sg13g2_fill_1 FILLER_66_370 ();
 sg13g2_fill_2 FILLER_66_451 ();
 sg13g2_decap_8 FILLER_66_457 ();
 sg13g2_decap_8 FILLER_66_464 ();
 sg13g2_decap_8 FILLER_66_471 ();
 sg13g2_decap_4 FILLER_66_478 ();
 sg13g2_decap_8 FILLER_66_486 ();
 sg13g2_fill_2 FILLER_66_493 ();
 sg13g2_decap_8 FILLER_66_515 ();
 sg13g2_decap_8 FILLER_66_522 ();
 sg13g2_decap_8 FILLER_66_529 ();
 sg13g2_decap_8 FILLER_66_536 ();
 sg13g2_decap_4 FILLER_66_543 ();
 sg13g2_fill_1 FILLER_66_547 ();
 sg13g2_fill_1 FILLER_66_578 ();
 sg13g2_fill_1 FILLER_66_583 ();
 sg13g2_fill_1 FILLER_66_589 ();
 sg13g2_fill_1 FILLER_66_595 ();
 sg13g2_fill_2 FILLER_66_622 ();
 sg13g2_fill_1 FILLER_66_624 ();
 sg13g2_fill_1 FILLER_66_639 ();
 sg13g2_decap_4 FILLER_66_653 ();
 sg13g2_fill_1 FILLER_66_657 ();
 sg13g2_fill_2 FILLER_66_663 ();
 sg13g2_fill_1 FILLER_66_668 ();
 sg13g2_decap_8 FILLER_66_674 ();
 sg13g2_decap_8 FILLER_66_681 ();
 sg13g2_decap_8 FILLER_66_688 ();
 sg13g2_decap_8 FILLER_66_695 ();
 sg13g2_fill_1 FILLER_66_702 ();
 sg13g2_decap_4 FILLER_66_737 ();
 sg13g2_fill_1 FILLER_66_741 ();
 sg13g2_decap_4 FILLER_66_813 ();
 sg13g2_fill_1 FILLER_66_899 ();
 sg13g2_fill_2 FILLER_66_960 ();
 sg13g2_fill_1 FILLER_66_962 ();
 sg13g2_decap_4 FILLER_66_997 ();
 sg13g2_decap_8 FILLER_66_1007 ();
 sg13g2_fill_1 FILLER_66_1014 ();
 sg13g2_fill_2 FILLER_66_1021 ();
 sg13g2_fill_1 FILLER_66_1033 ();
 sg13g2_fill_2 FILLER_66_1038 ();
 sg13g2_fill_1 FILLER_66_1040 ();
 sg13g2_fill_2 FILLER_66_1056 ();
 sg13g2_fill_1 FILLER_66_1058 ();
 sg13g2_decap_8 FILLER_66_1063 ();
 sg13g2_fill_1 FILLER_66_1080 ();
 sg13g2_decap_8 FILLER_66_1091 ();
 sg13g2_decap_8 FILLER_66_1098 ();
 sg13g2_fill_1 FILLER_66_1110 ();
 sg13g2_fill_1 FILLER_66_1137 ();
 sg13g2_decap_4 FILLER_66_1170 ();
 sg13g2_fill_1 FILLER_66_1174 ();
 sg13g2_decap_8 FILLER_66_1214 ();
 sg13g2_decap_8 FILLER_66_1221 ();
 sg13g2_decap_8 FILLER_66_1228 ();
 sg13g2_decap_8 FILLER_66_1235 ();
 sg13g2_decap_8 FILLER_66_1242 ();
 sg13g2_fill_1 FILLER_66_1249 ();
 sg13g2_decap_8 FILLER_66_1260 ();
 sg13g2_fill_2 FILLER_66_1267 ();
 sg13g2_fill_1 FILLER_66_1295 ();
 sg13g2_fill_1 FILLER_66_1302 ();
 sg13g2_fill_2 FILLER_66_1338 ();
 sg13g2_fill_1 FILLER_66_1345 ();
 sg13g2_fill_1 FILLER_66_1353 ();
 sg13g2_fill_2 FILLER_66_1358 ();
 sg13g2_fill_1 FILLER_66_1374 ();
 sg13g2_fill_2 FILLER_66_1383 ();
 sg13g2_decap_4 FILLER_66_1415 ();
 sg13g2_fill_1 FILLER_66_1419 ();
 sg13g2_fill_1 FILLER_66_1426 ();
 sg13g2_fill_1 FILLER_66_1471 ();
 sg13g2_fill_1 FILLER_66_1485 ();
 sg13g2_fill_2 FILLER_66_1506 ();
 sg13g2_decap_4 FILLER_66_1543 ();
 sg13g2_decap_4 FILLER_66_1587 ();
 sg13g2_fill_2 FILLER_66_1591 ();
 sg13g2_decap_4 FILLER_66_1598 ();
 sg13g2_fill_1 FILLER_66_1602 ();
 sg13g2_fill_2 FILLER_66_1613 ();
 sg13g2_fill_1 FILLER_66_1615 ();
 sg13g2_decap_8 FILLER_66_1623 ();
 sg13g2_decap_8 FILLER_66_1657 ();
 sg13g2_fill_2 FILLER_66_1664 ();
 sg13g2_decap_4 FILLER_66_1698 ();
 sg13g2_fill_1 FILLER_66_1702 ();
 sg13g2_decap_8 FILLER_66_1708 ();
 sg13g2_decap_8 FILLER_66_1715 ();
 sg13g2_fill_1 FILLER_66_1722 ();
 sg13g2_fill_1 FILLER_66_1731 ();
 sg13g2_fill_1 FILLER_66_1736 ();
 sg13g2_fill_2 FILLER_66_1777 ();
 sg13g2_fill_2 FILLER_66_1789 ();
 sg13g2_fill_1 FILLER_66_1791 ();
 sg13g2_fill_1 FILLER_66_1796 ();
 sg13g2_fill_2 FILLER_66_1806 ();
 sg13g2_decap_8 FILLER_66_1813 ();
 sg13g2_fill_1 FILLER_66_1820 ();
 sg13g2_fill_2 FILLER_66_1859 ();
 sg13g2_fill_2 FILLER_66_1875 ();
 sg13g2_decap_4 FILLER_66_1895 ();
 sg13g2_fill_1 FILLER_66_1899 ();
 sg13g2_decap_4 FILLER_66_1933 ();
 sg13g2_decap_8 FILLER_66_1941 ();
 sg13g2_decap_8 FILLER_66_1948 ();
 sg13g2_decap_4 FILLER_66_1955 ();
 sg13g2_decap_8 FILLER_66_1963 ();
 sg13g2_fill_1 FILLER_66_1970 ();
 sg13g2_fill_2 FILLER_66_1987 ();
 sg13g2_fill_2 FILLER_66_1997 ();
 sg13g2_fill_1 FILLER_66_2004 ();
 sg13g2_decap_4 FILLER_66_2018 ();
 sg13g2_fill_1 FILLER_66_2038 ();
 sg13g2_fill_1 FILLER_66_2058 ();
 sg13g2_fill_1 FILLER_66_2071 ();
 sg13g2_fill_2 FILLER_66_2159 ();
 sg13g2_decap_4 FILLER_66_2171 ();
 sg13g2_fill_2 FILLER_66_2175 ();
 sg13g2_decap_8 FILLER_66_2181 ();
 sg13g2_fill_1 FILLER_66_2224 ();
 sg13g2_decap_8 FILLER_66_2262 ();
 sg13g2_decap_8 FILLER_66_2269 ();
 sg13g2_fill_1 FILLER_66_2276 ();
 sg13g2_fill_1 FILLER_66_2312 ();
 sg13g2_fill_1 FILLER_66_2317 ();
 sg13g2_fill_1 FILLER_66_2376 ();
 sg13g2_fill_1 FILLER_66_2382 ();
 sg13g2_fill_1 FILLER_66_2401 ();
 sg13g2_fill_2 FILLER_66_2463 ();
 sg13g2_decap_4 FILLER_66_2469 ();
 sg13g2_fill_1 FILLER_66_2473 ();
 sg13g2_decap_8 FILLER_66_2478 ();
 sg13g2_fill_2 FILLER_66_2485 ();
 sg13g2_fill_2 FILLER_66_2496 ();
 sg13g2_fill_2 FILLER_66_2503 ();
 sg13g2_fill_1 FILLER_66_2505 ();
 sg13g2_fill_1 FILLER_66_2512 ();
 sg13g2_fill_1 FILLER_66_2523 ();
 sg13g2_fill_2 FILLER_66_2529 ();
 sg13g2_fill_2 FILLER_66_2541 ();
 sg13g2_fill_2 FILLER_66_2603 ();
 sg13g2_fill_1 FILLER_66_2605 ();
 sg13g2_decap_8 FILLER_66_2625 ();
 sg13g2_decap_8 FILLER_66_2632 ();
 sg13g2_decap_8 FILLER_66_2639 ();
 sg13g2_decap_8 FILLER_66_2646 ();
 sg13g2_decap_8 FILLER_66_2653 ();
 sg13g2_decap_8 FILLER_66_2660 ();
 sg13g2_fill_2 FILLER_66_2667 ();
 sg13g2_fill_1 FILLER_66_2669 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_fill_2 FILLER_67_7 ();
 sg13g2_decap_4 FILLER_67_13 ();
 sg13g2_fill_1 FILLER_67_38 ();
 sg13g2_decap_8 FILLER_67_69 ();
 sg13g2_decap_8 FILLER_67_76 ();
 sg13g2_fill_1 FILLER_67_83 ();
 sg13g2_decap_8 FILLER_67_97 ();
 sg13g2_decap_8 FILLER_67_104 ();
 sg13g2_decap_8 FILLER_67_111 ();
 sg13g2_fill_1 FILLER_67_169 ();
 sg13g2_fill_2 FILLER_67_190 ();
 sg13g2_fill_1 FILLER_67_192 ();
 sg13g2_fill_2 FILLER_67_198 ();
 sg13g2_fill_1 FILLER_67_200 ();
 sg13g2_decap_4 FILLER_67_206 ();
 sg13g2_fill_1 FILLER_67_210 ();
 sg13g2_fill_1 FILLER_67_275 ();
 sg13g2_fill_1 FILLER_67_293 ();
 sg13g2_fill_1 FILLER_67_313 ();
 sg13g2_fill_1 FILLER_67_355 ();
 sg13g2_fill_1 FILLER_67_377 ();
 sg13g2_fill_2 FILLER_67_381 ();
 sg13g2_fill_2 FILLER_67_428 ();
 sg13g2_fill_1 FILLER_67_430 ();
 sg13g2_decap_4 FILLER_67_466 ();
 sg13g2_fill_2 FILLER_67_470 ();
 sg13g2_decap_8 FILLER_67_475 ();
 sg13g2_decap_8 FILLER_67_485 ();
 sg13g2_decap_8 FILLER_67_492 ();
 sg13g2_decap_4 FILLER_67_499 ();
 sg13g2_fill_2 FILLER_67_503 ();
 sg13g2_fill_2 FILLER_67_543 ();
 sg13g2_fill_2 FILLER_67_576 ();
 sg13g2_fill_1 FILLER_67_578 ();
 sg13g2_fill_2 FILLER_67_625 ();
 sg13g2_decap_8 FILLER_67_632 ();
 sg13g2_fill_1 FILLER_67_639 ();
 sg13g2_decap_4 FILLER_67_645 ();
 sg13g2_fill_1 FILLER_67_649 ();
 sg13g2_fill_2 FILLER_67_665 ();
 sg13g2_decap_8 FILLER_67_679 ();
 sg13g2_decap_8 FILLER_67_686 ();
 sg13g2_fill_2 FILLER_67_693 ();
 sg13g2_fill_1 FILLER_67_695 ();
 sg13g2_decap_4 FILLER_67_701 ();
 sg13g2_decap_8 FILLER_67_709 ();
 sg13g2_decap_8 FILLER_67_716 ();
 sg13g2_fill_2 FILLER_67_723 ();
 sg13g2_fill_1 FILLER_67_725 ();
 sg13g2_fill_2 FILLER_67_770 ();
 sg13g2_fill_1 FILLER_67_772 ();
 sg13g2_decap_4 FILLER_67_783 ();
 sg13g2_fill_2 FILLER_67_787 ();
 sg13g2_fill_1 FILLER_67_793 ();
 sg13g2_decap_4 FILLER_67_804 ();
 sg13g2_fill_1 FILLER_67_808 ();
 sg13g2_decap_4 FILLER_67_814 ();
 sg13g2_fill_1 FILLER_67_818 ();
 sg13g2_fill_1 FILLER_67_868 ();
 sg13g2_fill_1 FILLER_67_879 ();
 sg13g2_fill_1 FILLER_67_932 ();
 sg13g2_decap_8 FILLER_67_947 ();
 sg13g2_decap_4 FILLER_67_954 ();
 sg13g2_decap_8 FILLER_67_962 ();
 sg13g2_fill_2 FILLER_67_969 ();
 sg13g2_fill_1 FILLER_67_971 ();
 sg13g2_decap_8 FILLER_67_976 ();
 sg13g2_fill_2 FILLER_67_983 ();
 sg13g2_fill_1 FILLER_67_985 ();
 sg13g2_fill_2 FILLER_67_990 ();
 sg13g2_fill_1 FILLER_67_992 ();
 sg13g2_decap_8 FILLER_67_1093 ();
 sg13g2_decap_4 FILLER_67_1104 ();
 sg13g2_fill_1 FILLER_67_1118 ();
 sg13g2_fill_1 FILLER_67_1133 ();
 sg13g2_fill_1 FILLER_67_1198 ();
 sg13g2_fill_2 FILLER_67_1229 ();
 sg13g2_fill_1 FILLER_67_1231 ();
 sg13g2_fill_2 FILLER_67_1236 ();
 sg13g2_fill_1 FILLER_67_1238 ();
 sg13g2_decap_8 FILLER_67_1269 ();
 sg13g2_decap_4 FILLER_67_1276 ();
 sg13g2_fill_1 FILLER_67_1285 ();
 sg13g2_fill_1 FILLER_67_1312 ();
 sg13g2_fill_2 FILLER_67_1319 ();
 sg13g2_fill_1 FILLER_67_1329 ();
 sg13g2_decap_4 FILLER_67_1341 ();
 sg13g2_fill_1 FILLER_67_1345 ();
 sg13g2_decap_8 FILLER_67_1353 ();
 sg13g2_decap_8 FILLER_67_1360 ();
 sg13g2_decap_4 FILLER_67_1367 ();
 sg13g2_fill_1 FILLER_67_1371 ();
 sg13g2_fill_1 FILLER_67_1386 ();
 sg13g2_fill_2 FILLER_67_1417 ();
 sg13g2_fill_2 FILLER_67_1437 ();
 sg13g2_fill_1 FILLER_67_1452 ();
 sg13g2_fill_2 FILLER_67_1476 ();
 sg13g2_fill_1 FILLER_67_1478 ();
 sg13g2_decap_4 FILLER_67_1506 ();
 sg13g2_fill_2 FILLER_67_1510 ();
 sg13g2_decap_8 FILLER_67_1519 ();
 sg13g2_decap_8 FILLER_67_1526 ();
 sg13g2_fill_1 FILLER_67_1533 ();
 sg13g2_decap_4 FILLER_67_1539 ();
 sg13g2_fill_2 FILLER_67_1543 ();
 sg13g2_decap_8 FILLER_67_1581 ();
 sg13g2_decap_4 FILLER_67_1608 ();
 sg13g2_decap_8 FILLER_67_1636 ();
 sg13g2_decap_4 FILLER_67_1643 ();
 sg13g2_fill_2 FILLER_67_1647 ();
 sg13g2_decap_8 FILLER_67_1665 ();
 sg13g2_decap_8 FILLER_67_1672 ();
 sg13g2_decap_4 FILLER_67_1684 ();
 sg13g2_fill_2 FILLER_67_1688 ();
 sg13g2_decap_4 FILLER_67_1695 ();
 sg13g2_fill_1 FILLER_67_1699 ();
 sg13g2_fill_1 FILLER_67_1704 ();
 sg13g2_decap_8 FILLER_67_1711 ();
 sg13g2_decap_4 FILLER_67_1718 ();
 sg13g2_fill_2 FILLER_67_1722 ();
 sg13g2_fill_2 FILLER_67_1744 ();
 sg13g2_fill_1 FILLER_67_1749 ();
 sg13g2_fill_1 FILLER_67_1760 ();
 sg13g2_fill_2 FILLER_67_1788 ();
 sg13g2_fill_1 FILLER_67_1795 ();
 sg13g2_fill_1 FILLER_67_1807 ();
 sg13g2_fill_2 FILLER_67_1820 ();
 sg13g2_decap_4 FILLER_67_1856 ();
 sg13g2_fill_2 FILLER_67_1860 ();
 sg13g2_decap_4 FILLER_67_1867 ();
 sg13g2_fill_1 FILLER_67_1885 ();
 sg13g2_fill_2 FILLER_67_1896 ();
 sg13g2_fill_1 FILLER_67_1898 ();
 sg13g2_decap_8 FILLER_67_1925 ();
 sg13g2_decap_8 FILLER_67_1932 ();
 sg13g2_decap_8 FILLER_67_1939 ();
 sg13g2_decap_4 FILLER_67_1982 ();
 sg13g2_fill_1 FILLER_67_1986 ();
 sg13g2_decap_8 FILLER_67_2011 ();
 sg13g2_decap_8 FILLER_67_2018 ();
 sg13g2_decap_4 FILLER_67_2025 ();
 sg13g2_fill_1 FILLER_67_2029 ();
 sg13g2_fill_1 FILLER_67_2034 ();
 sg13g2_fill_2 FILLER_67_2044 ();
 sg13g2_decap_8 FILLER_67_2050 ();
 sg13g2_decap_8 FILLER_67_2057 ();
 sg13g2_decap_4 FILLER_67_2064 ();
 sg13g2_fill_1 FILLER_67_2068 ();
 sg13g2_fill_1 FILLER_67_2081 ();
 sg13g2_fill_1 FILLER_67_2139 ();
 sg13g2_fill_2 FILLER_67_2156 ();
 sg13g2_fill_1 FILLER_67_2162 ();
 sg13g2_fill_2 FILLER_67_2167 ();
 sg13g2_fill_1 FILLER_67_2195 ();
 sg13g2_fill_1 FILLER_67_2203 ();
 sg13g2_decap_8 FILLER_67_2281 ();
 sg13g2_fill_2 FILLER_67_2293 ();
 sg13g2_fill_1 FILLER_67_2295 ();
 sg13g2_fill_1 FILLER_67_2305 ();
 sg13g2_fill_2 FILLER_67_2316 ();
 sg13g2_fill_2 FILLER_67_2321 ();
 sg13g2_fill_2 FILLER_67_2344 ();
 sg13g2_fill_1 FILLER_67_2346 ();
 sg13g2_decap_4 FILLER_67_2384 ();
 sg13g2_fill_2 FILLER_67_2414 ();
 sg13g2_fill_2 FILLER_67_2457 ();
 sg13g2_fill_1 FILLER_67_2459 ();
 sg13g2_fill_2 FILLER_67_2464 ();
 sg13g2_fill_1 FILLER_67_2502 ();
 sg13g2_fill_1 FILLER_67_2512 ();
 sg13g2_fill_2 FILLER_67_2539 ();
 sg13g2_fill_1 FILLER_67_2541 ();
 sg13g2_fill_2 FILLER_67_2548 ();
 sg13g2_fill_1 FILLER_67_2550 ();
 sg13g2_fill_2 FILLER_67_2555 ();
 sg13g2_fill_1 FILLER_67_2557 ();
 sg13g2_fill_1 FILLER_67_2594 ();
 sg13g2_decap_8 FILLER_67_2621 ();
 sg13g2_decap_8 FILLER_67_2628 ();
 sg13g2_decap_8 FILLER_67_2635 ();
 sg13g2_decap_8 FILLER_67_2642 ();
 sg13g2_decap_8 FILLER_67_2649 ();
 sg13g2_decap_8 FILLER_67_2656 ();
 sg13g2_decap_8 FILLER_67_2663 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_4 FILLER_68_7 ();
 sg13g2_fill_1 FILLER_68_25 ();
 sg13g2_fill_2 FILLER_68_31 ();
 sg13g2_fill_1 FILLER_68_33 ();
 sg13g2_fill_1 FILLER_68_38 ();
 sg13g2_decap_4 FILLER_68_64 ();
 sg13g2_decap_8 FILLER_68_72 ();
 sg13g2_fill_1 FILLER_68_79 ();
 sg13g2_fill_2 FILLER_68_106 ();
 sg13g2_fill_1 FILLER_68_108 ();
 sg13g2_fill_2 FILLER_68_143 ();
 sg13g2_fill_1 FILLER_68_145 ();
 sg13g2_fill_2 FILLER_68_151 ();
 sg13g2_fill_1 FILLER_68_153 ();
 sg13g2_fill_2 FILLER_68_159 ();
 sg13g2_fill_1 FILLER_68_161 ();
 sg13g2_fill_2 FILLER_68_230 ();
 sg13g2_fill_2 FILLER_68_237 ();
 sg13g2_fill_2 FILLER_68_243 ();
 sg13g2_fill_1 FILLER_68_245 ();
 sg13g2_fill_1 FILLER_68_251 ();
 sg13g2_fill_2 FILLER_68_256 ();
 sg13g2_fill_1 FILLER_68_258 ();
 sg13g2_decap_8 FILLER_68_265 ();
 sg13g2_fill_1 FILLER_68_286 ();
 sg13g2_fill_1 FILLER_68_302 ();
 sg13g2_fill_1 FILLER_68_326 ();
 sg13g2_fill_2 FILLER_68_333 ();
 sg13g2_fill_2 FILLER_68_372 ();
 sg13g2_fill_1 FILLER_68_383 ();
 sg13g2_fill_1 FILLER_68_410 ();
 sg13g2_fill_1 FILLER_68_415 ();
 sg13g2_fill_2 FILLER_68_420 ();
 sg13g2_decap_4 FILLER_68_426 ();
 sg13g2_fill_2 FILLER_68_430 ();
 sg13g2_decap_4 FILLER_68_513 ();
 sg13g2_fill_2 FILLER_68_555 ();
 sg13g2_fill_1 FILLER_68_557 ();
 sg13g2_fill_2 FILLER_68_577 ();
 sg13g2_fill_2 FILLER_68_584 ();
 sg13g2_fill_1 FILLER_68_586 ();
 sg13g2_fill_1 FILLER_68_613 ();
 sg13g2_fill_2 FILLER_68_640 ();
 sg13g2_fill_1 FILLER_68_642 ();
 sg13g2_fill_2 FILLER_68_695 ();
 sg13g2_fill_1 FILLER_68_697 ();
 sg13g2_decap_8 FILLER_68_755 ();
 sg13g2_fill_2 FILLER_68_762 ();
 sg13g2_fill_1 FILLER_68_764 ();
 sg13g2_decap_8 FILLER_68_769 ();
 sg13g2_decap_4 FILLER_68_776 ();
 sg13g2_fill_1 FILLER_68_780 ();
 sg13g2_fill_1 FILLER_68_793 ();
 sg13g2_fill_1 FILLER_68_815 ();
 sg13g2_fill_1 FILLER_68_873 ();
 sg13g2_fill_2 FILLER_68_901 ();
 sg13g2_decap_8 FILLER_68_939 ();
 sg13g2_fill_1 FILLER_68_976 ();
 sg13g2_fill_2 FILLER_68_1013 ();
 sg13g2_fill_1 FILLER_68_1015 ();
 sg13g2_fill_1 FILLER_68_1026 ();
 sg13g2_fill_1 FILLER_68_1033 ();
 sg13g2_fill_2 FILLER_68_1060 ();
 sg13g2_fill_1 FILLER_68_1192 ();
 sg13g2_fill_2 FILLER_68_1203 ();
 sg13g2_fill_1 FILLER_68_1205 ();
 sg13g2_fill_2 FILLER_68_1210 ();
 sg13g2_fill_1 FILLER_68_1212 ();
 sg13g2_decap_8 FILLER_68_1249 ();
 sg13g2_fill_2 FILLER_68_1256 ();
 sg13g2_fill_1 FILLER_68_1290 ();
 sg13g2_fill_1 FILLER_68_1318 ();
 sg13g2_fill_1 FILLER_68_1335 ();
 sg13g2_decap_4 FILLER_68_1341 ();
 sg13g2_fill_1 FILLER_68_1345 ();
 sg13g2_decap_8 FILLER_68_1355 ();
 sg13g2_fill_2 FILLER_68_1362 ();
 sg13g2_fill_1 FILLER_68_1364 ();
 sg13g2_decap_8 FILLER_68_1374 ();
 sg13g2_fill_2 FILLER_68_1414 ();
 sg13g2_fill_2 FILLER_68_1445 ();
 sg13g2_fill_1 FILLER_68_1447 ();
 sg13g2_fill_1 FILLER_68_1476 ();
 sg13g2_fill_1 FILLER_68_1491 ();
 sg13g2_decap_8 FILLER_68_1537 ();
 sg13g2_decap_8 FILLER_68_1544 ();
 sg13g2_fill_2 FILLER_68_1551 ();
 sg13g2_fill_1 FILLER_68_1553 ();
 sg13g2_decap_8 FILLER_68_1590 ();
 sg13g2_decap_8 FILLER_68_1597 ();
 sg13g2_decap_8 FILLER_68_1604 ();
 sg13g2_decap_8 FILLER_68_1611 ();
 sg13g2_fill_2 FILLER_68_1641 ();
 sg13g2_fill_1 FILLER_68_1643 ();
 sg13g2_decap_8 FILLER_68_1649 ();
 sg13g2_decap_4 FILLER_68_1656 ();
 sg13g2_fill_2 FILLER_68_1660 ();
 sg13g2_decap_8 FILLER_68_1667 ();
 sg13g2_fill_2 FILLER_68_1684 ();
 sg13g2_fill_1 FILLER_68_1686 ();
 sg13g2_decap_4 FILLER_68_1691 ();
 sg13g2_fill_2 FILLER_68_1695 ();
 sg13g2_decap_4 FILLER_68_1701 ();
 sg13g2_fill_1 FILLER_68_1705 ();
 sg13g2_fill_1 FILLER_68_1739 ();
 sg13g2_fill_1 FILLER_68_1764 ();
 sg13g2_fill_1 FILLER_68_1769 ();
 sg13g2_fill_1 FILLER_68_1783 ();
 sg13g2_fill_1 FILLER_68_1795 ();
 sg13g2_fill_1 FILLER_68_1815 ();
 sg13g2_fill_1 FILLER_68_1835 ();
 sg13g2_decap_8 FILLER_68_1854 ();
 sg13g2_decap_8 FILLER_68_1861 ();
 sg13g2_fill_2 FILLER_68_1868 ();
 sg13g2_decap_4 FILLER_68_1881 ();
 sg13g2_fill_1 FILLER_68_1885 ();
 sg13g2_fill_2 FILLER_68_1909 ();
 sg13g2_decap_4 FILLER_68_1938 ();
 sg13g2_fill_2 FILLER_68_1942 ();
 sg13g2_fill_2 FILLER_68_1949 ();
 sg13g2_fill_2 FILLER_68_1956 ();
 sg13g2_fill_1 FILLER_68_1958 ();
 sg13g2_fill_1 FILLER_68_1972 ();
 sg13g2_fill_1 FILLER_68_2007 ();
 sg13g2_fill_2 FILLER_68_2013 ();
 sg13g2_fill_1 FILLER_68_2019 ();
 sg13g2_fill_2 FILLER_68_2025 ();
 sg13g2_fill_1 FILLER_68_2027 ();
 sg13g2_decap_8 FILLER_68_2049 ();
 sg13g2_decap_4 FILLER_68_2056 ();
 sg13g2_fill_2 FILLER_68_2064 ();
 sg13g2_fill_1 FILLER_68_2085 ();
 sg13g2_fill_1 FILLER_68_2091 ();
 sg13g2_fill_2 FILLER_68_2118 ();
 sg13g2_decap_8 FILLER_68_2164 ();
 sg13g2_decap_4 FILLER_68_2171 ();
 sg13g2_fill_2 FILLER_68_2175 ();
 sg13g2_decap_8 FILLER_68_2181 ();
 sg13g2_fill_1 FILLER_68_2224 ();
 sg13g2_fill_1 FILLER_68_2247 ();
 sg13g2_fill_2 FILLER_68_2270 ();
 sg13g2_fill_1 FILLER_68_2334 ();
 sg13g2_decap_4 FILLER_68_2339 ();
 sg13g2_decap_8 FILLER_68_2348 ();
 sg13g2_decap_4 FILLER_68_2355 ();
 sg13g2_fill_1 FILLER_68_2363 ();
 sg13g2_decap_4 FILLER_68_2369 ();
 sg13g2_fill_1 FILLER_68_2373 ();
 sg13g2_decap_8 FILLER_68_2379 ();
 sg13g2_decap_4 FILLER_68_2386 ();
 sg13g2_fill_1 FILLER_68_2399 ();
 sg13g2_fill_2 FILLER_68_2404 ();
 sg13g2_decap_8 FILLER_68_2457 ();
 sg13g2_decap_8 FILLER_68_2499 ();
 sg13g2_fill_2 FILLER_68_2506 ();
 sg13g2_fill_1 FILLER_68_2508 ();
 sg13g2_decap_8 FILLER_68_2515 ();
 sg13g2_fill_2 FILLER_68_2549 ();
 sg13g2_fill_1 FILLER_68_2551 ();
 sg13g2_fill_1 FILLER_68_2556 ();
 sg13g2_fill_2 FILLER_68_2562 ();
 sg13g2_fill_2 FILLER_68_2568 ();
 sg13g2_fill_2 FILLER_68_2574 ();
 sg13g2_decap_8 FILLER_68_2628 ();
 sg13g2_decap_8 FILLER_68_2635 ();
 sg13g2_decap_8 FILLER_68_2642 ();
 sg13g2_decap_8 FILLER_68_2649 ();
 sg13g2_decap_8 FILLER_68_2656 ();
 sg13g2_decap_8 FILLER_68_2663 ();
 sg13g2_fill_2 FILLER_69_0 ();
 sg13g2_fill_2 FILLER_69_28 ();
 sg13g2_fill_1 FILLER_69_30 ();
 sg13g2_fill_2 FILLER_69_36 ();
 sg13g2_fill_2 FILLER_69_64 ();
 sg13g2_fill_2 FILLER_69_102 ();
 sg13g2_fill_1 FILLER_69_104 ();
 sg13g2_decap_4 FILLER_69_124 ();
 sg13g2_fill_1 FILLER_69_154 ();
 sg13g2_fill_2 FILLER_69_160 ();
 sg13g2_fill_2 FILLER_69_188 ();
 sg13g2_fill_1 FILLER_69_190 ();
 sg13g2_fill_2 FILLER_69_217 ();
 sg13g2_fill_1 FILLER_69_260 ();
 sg13g2_fill_1 FILLER_69_284 ();
 sg13g2_fill_1 FILLER_69_296 ();
 sg13g2_fill_2 FILLER_69_300 ();
 sg13g2_fill_1 FILLER_69_312 ();
 sg13g2_fill_1 FILLER_69_343 ();
 sg13g2_fill_1 FILLER_69_354 ();
 sg13g2_fill_2 FILLER_69_392 ();
 sg13g2_fill_1 FILLER_69_398 ();
 sg13g2_fill_2 FILLER_69_407 ();
 sg13g2_decap_4 FILLER_69_418 ();
 sg13g2_decap_4 FILLER_69_427 ();
 sg13g2_fill_1 FILLER_69_448 ();
 sg13g2_fill_1 FILLER_69_457 ();
 sg13g2_fill_2 FILLER_69_462 ();
 sg13g2_fill_1 FILLER_69_464 ();
 sg13g2_decap_8 FILLER_69_517 ();
 sg13g2_fill_1 FILLER_69_532 ();
 sg13g2_decap_8 FILLER_69_537 ();
 sg13g2_decap_8 FILLER_69_553 ();
 sg13g2_fill_2 FILLER_69_560 ();
 sg13g2_fill_2 FILLER_69_592 ();
 sg13g2_fill_1 FILLER_69_598 ();
 sg13g2_decap_8 FILLER_69_605 ();
 sg13g2_fill_1 FILLER_69_616 ();
 sg13g2_fill_1 FILLER_69_621 ();
 sg13g2_fill_1 FILLER_69_648 ();
 sg13g2_fill_1 FILLER_69_677 ();
 sg13g2_fill_2 FILLER_69_683 ();
 sg13g2_decap_8 FILLER_69_690 ();
 sg13g2_decap_8 FILLER_69_697 ();
 sg13g2_fill_2 FILLER_69_704 ();
 sg13g2_fill_1 FILLER_69_710 ();
 sg13g2_fill_1 FILLER_69_737 ();
 sg13g2_decap_8 FILLER_69_758 ();
 sg13g2_fill_2 FILLER_69_765 ();
 sg13g2_fill_1 FILLER_69_777 ();
 sg13g2_fill_2 FILLER_69_784 ();
 sg13g2_fill_1 FILLER_69_790 ();
 sg13g2_fill_2 FILLER_69_817 ();
 sg13g2_fill_2 FILLER_69_827 ();
 sg13g2_fill_1 FILLER_69_881 ();
 sg13g2_decap_4 FILLER_69_888 ();
 sg13g2_fill_1 FILLER_69_892 ();
 sg13g2_fill_2 FILLER_69_903 ();
 sg13g2_fill_1 FILLER_69_908 ();
 sg13g2_fill_2 FILLER_69_915 ();
 sg13g2_fill_1 FILLER_69_917 ();
 sg13g2_fill_1 FILLER_69_921 ();
 sg13g2_decap_8 FILLER_69_936 ();
 sg13g2_fill_1 FILLER_69_943 ();
 sg13g2_fill_2 FILLER_69_954 ();
 sg13g2_fill_2 FILLER_69_1006 ();
 sg13g2_fill_1 FILLER_69_1008 ();
 sg13g2_fill_2 FILLER_69_1014 ();
 sg13g2_fill_1 FILLER_69_1087 ();
 sg13g2_decap_4 FILLER_69_1092 ();
 sg13g2_fill_2 FILLER_69_1096 ();
 sg13g2_fill_2 FILLER_69_1105 ();
 sg13g2_decap_8 FILLER_69_1187 ();
 sg13g2_decap_8 FILLER_69_1194 ();
 sg13g2_decap_4 FILLER_69_1201 ();
 sg13g2_fill_2 FILLER_69_1215 ();
 sg13g2_fill_2 FILLER_69_1227 ();
 sg13g2_fill_2 FILLER_69_1242 ();
 sg13g2_fill_2 FILLER_69_1270 ();
 sg13g2_fill_1 FILLER_69_1285 ();
 sg13g2_fill_1 FILLER_69_1337 ();
 sg13g2_fill_2 FILLER_69_1355 ();
 sg13g2_fill_1 FILLER_69_1357 ();
 sg13g2_decap_4 FILLER_69_1363 ();
 sg13g2_fill_1 FILLER_69_1388 ();
 sg13g2_fill_2 FILLER_69_1399 ();
 sg13g2_fill_1 FILLER_69_1418 ();
 sg13g2_decap_4 FILLER_69_1425 ();
 sg13g2_fill_2 FILLER_69_1434 ();
 sg13g2_fill_1 FILLER_69_1436 ();
 sg13g2_decap_4 FILLER_69_1444 ();
 sg13g2_fill_1 FILLER_69_1459 ();
 sg13g2_fill_2 FILLER_69_1468 ();
 sg13g2_decap_4 FILLER_69_1475 ();
 sg13g2_fill_2 FILLER_69_1489 ();
 sg13g2_fill_1 FILLER_69_1491 ();
 sg13g2_fill_1 FILLER_69_1497 ();
 sg13g2_fill_1 FILLER_69_1516 ();
 sg13g2_fill_2 FILLER_69_1521 ();
 sg13g2_fill_1 FILLER_69_1523 ();
 sg13g2_fill_2 FILLER_69_1564 ();
 sg13g2_fill_1 FILLER_69_1570 ();
 sg13g2_decap_8 FILLER_69_1579 ();
 sg13g2_decap_8 FILLER_69_1586 ();
 sg13g2_decap_8 FILLER_69_1593 ();
 sg13g2_decap_8 FILLER_69_1600 ();
 sg13g2_decap_8 FILLER_69_1607 ();
 sg13g2_decap_8 FILLER_69_1614 ();
 sg13g2_decap_4 FILLER_69_1621 ();
 sg13g2_decap_8 FILLER_69_1658 ();
 sg13g2_fill_2 FILLER_69_1665 ();
 sg13g2_fill_1 FILLER_69_1667 ();
 sg13g2_fill_1 FILLER_69_1683 ();
 sg13g2_fill_2 FILLER_69_1691 ();
 sg13g2_fill_1 FILLER_69_1693 ();
 sg13g2_fill_1 FILLER_69_1705 ();
 sg13g2_fill_2 FILLER_69_1716 ();
 sg13g2_fill_2 FILLER_69_1744 ();
 sg13g2_fill_1 FILLER_69_1785 ();
 sg13g2_decap_4 FILLER_69_1790 ();
 sg13g2_fill_2 FILLER_69_1794 ();
 sg13g2_fill_2 FILLER_69_1842 ();
 sg13g2_fill_1 FILLER_69_1849 ();
 sg13g2_decap_8 FILLER_69_1855 ();
 sg13g2_decap_4 FILLER_69_1862 ();
 sg13g2_fill_2 FILLER_69_1866 ();
 sg13g2_decap_8 FILLER_69_1877 ();
 sg13g2_decap_4 FILLER_69_1884 ();
 sg13g2_fill_2 FILLER_69_1888 ();
 sg13g2_fill_1 FILLER_69_1894 ();
 sg13g2_fill_1 FILLER_69_1926 ();
 sg13g2_decap_8 FILLER_69_1933 ();
 sg13g2_fill_1 FILLER_69_1950 ();
 sg13g2_fill_2 FILLER_69_1987 ();
 sg13g2_fill_1 FILLER_69_2018 ();
 sg13g2_fill_1 FILLER_69_2024 ();
 sg13g2_decap_8 FILLER_69_2033 ();
 sg13g2_decap_8 FILLER_69_2040 ();
 sg13g2_decap_8 FILLER_69_2047 ();
 sg13g2_decap_8 FILLER_69_2054 ();
 sg13g2_decap_8 FILLER_69_2157 ();
 sg13g2_decap_8 FILLER_69_2164 ();
 sg13g2_fill_1 FILLER_69_2171 ();
 sg13g2_fill_2 FILLER_69_2217 ();
 sg13g2_fill_2 FILLER_69_2257 ();
 sg13g2_fill_2 FILLER_69_2271 ();
 sg13g2_fill_2 FILLER_69_2276 ();
 sg13g2_fill_2 FILLER_69_2282 ();
 sg13g2_fill_1 FILLER_69_2292 ();
 sg13g2_fill_1 FILLER_69_2297 ();
 sg13g2_fill_1 FILLER_69_2304 ();
 sg13g2_fill_1 FILLER_69_2311 ();
 sg13g2_fill_2 FILLER_69_2317 ();
 sg13g2_fill_2 FILLER_69_2323 ();
 sg13g2_fill_1 FILLER_69_2325 ();
 sg13g2_fill_2 FILLER_69_2332 ();
 sg13g2_fill_1 FILLER_69_2334 ();
 sg13g2_decap_4 FILLER_69_2369 ();
 sg13g2_fill_1 FILLER_69_2373 ();
 sg13g2_fill_1 FILLER_69_2379 ();
 sg13g2_fill_2 FILLER_69_2410 ();
 sg13g2_fill_2 FILLER_69_2435 ();
 sg13g2_fill_2 FILLER_69_2467 ();
 sg13g2_fill_2 FILLER_69_2474 ();
 sg13g2_decap_8 FILLER_69_2480 ();
 sg13g2_fill_1 FILLER_69_2487 ();
 sg13g2_fill_2 FILLER_69_2498 ();
 sg13g2_fill_2 FILLER_69_2505 ();
 sg13g2_fill_2 FILLER_69_2606 ();
 sg13g2_decap_8 FILLER_69_2612 ();
 sg13g2_decap_8 FILLER_69_2619 ();
 sg13g2_decap_8 FILLER_69_2626 ();
 sg13g2_decap_8 FILLER_69_2633 ();
 sg13g2_decap_8 FILLER_69_2640 ();
 sg13g2_decap_8 FILLER_69_2647 ();
 sg13g2_decap_8 FILLER_69_2654 ();
 sg13g2_decap_8 FILLER_69_2661 ();
 sg13g2_fill_2 FILLER_69_2668 ();
 sg13g2_fill_2 FILLER_70_0 ();
 sg13g2_fill_2 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_48 ();
 sg13g2_decap_8 FILLER_70_55 ();
 sg13g2_decap_8 FILLER_70_62 ();
 sg13g2_decap_8 FILLER_70_69 ();
 sg13g2_decap_8 FILLER_70_76 ();
 sg13g2_fill_2 FILLER_70_83 ();
 sg13g2_decap_8 FILLER_70_93 ();
 sg13g2_decap_4 FILLER_70_100 ();
 sg13g2_fill_2 FILLER_70_104 ();
 sg13g2_fill_1 FILLER_70_111 ();
 sg13g2_decap_4 FILLER_70_138 ();
 sg13g2_fill_1 FILLER_70_142 ();
 sg13g2_decap_4 FILLER_70_155 ();
 sg13g2_fill_2 FILLER_70_159 ();
 sg13g2_fill_1 FILLER_70_170 ();
 sg13g2_decap_4 FILLER_70_175 ();
 sg13g2_fill_1 FILLER_70_179 ();
 sg13g2_fill_2 FILLER_70_185 ();
 sg13g2_fill_1 FILLER_70_187 ();
 sg13g2_fill_1 FILLER_70_192 ();
 sg13g2_fill_2 FILLER_70_219 ();
 sg13g2_fill_1 FILLER_70_221 ();
 sg13g2_decap_4 FILLER_70_230 ();
 sg13g2_fill_2 FILLER_70_234 ();
 sg13g2_decap_8 FILLER_70_240 ();
 sg13g2_decap_8 FILLER_70_247 ();
 sg13g2_fill_1 FILLER_70_254 ();
 sg13g2_fill_2 FILLER_70_261 ();
 sg13g2_fill_1 FILLER_70_263 ();
 sg13g2_fill_1 FILLER_70_269 ();
 sg13g2_fill_1 FILLER_70_276 ();
 sg13g2_fill_1 FILLER_70_282 ();
 sg13g2_fill_2 FILLER_70_288 ();
 sg13g2_fill_2 FILLER_70_295 ();
 sg13g2_fill_2 FILLER_70_322 ();
 sg13g2_fill_2 FILLER_70_350 ();
 sg13g2_decap_8 FILLER_70_394 ();
 sg13g2_fill_1 FILLER_70_401 ();
 sg13g2_decap_4 FILLER_70_438 ();
 sg13g2_fill_2 FILLER_70_442 ();
 sg13g2_fill_1 FILLER_70_474 ();
 sg13g2_fill_2 FILLER_70_478 ();
 sg13g2_decap_8 FILLER_70_550 ();
 sg13g2_decap_8 FILLER_70_557 ();
 sg13g2_fill_2 FILLER_70_564 ();
 sg13g2_fill_1 FILLER_70_566 ();
 sg13g2_fill_1 FILLER_70_577 ();
 sg13g2_fill_2 FILLER_70_582 ();
 sg13g2_decap_4 FILLER_70_611 ();
 sg13g2_fill_1 FILLER_70_615 ();
 sg13g2_fill_1 FILLER_70_635 ();
 sg13g2_fill_2 FILLER_70_641 ();
 sg13g2_fill_1 FILLER_70_643 ();
 sg13g2_fill_2 FILLER_70_648 ();
 sg13g2_fill_2 FILLER_70_659 ();
 sg13g2_fill_1 FILLER_70_661 ();
 sg13g2_fill_1 FILLER_70_667 ();
 sg13g2_fill_1 FILLER_70_673 ();
 sg13g2_fill_1 FILLER_70_700 ();
 sg13g2_fill_1 FILLER_70_705 ();
 sg13g2_fill_2 FILLER_70_751 ();
 sg13g2_fill_1 FILLER_70_753 ();
 sg13g2_fill_2 FILLER_70_816 ();
 sg13g2_fill_1 FILLER_70_844 ();
 sg13g2_fill_2 FILLER_70_871 ();
 sg13g2_decap_4 FILLER_70_919 ();
 sg13g2_fill_2 FILLER_70_923 ();
 sg13g2_decap_4 FILLER_70_965 ();
 sg13g2_fill_2 FILLER_70_969 ();
 sg13g2_decap_8 FILLER_70_980 ();
 sg13g2_decap_8 FILLER_70_993 ();
 sg13g2_decap_4 FILLER_70_1000 ();
 sg13g2_fill_2 FILLER_70_1004 ();
 sg13g2_decap_4 FILLER_70_1010 ();
 sg13g2_fill_1 FILLER_70_1017 ();
 sg13g2_decap_8 FILLER_70_1028 ();
 sg13g2_fill_1 FILLER_70_1035 ();
 sg13g2_decap_8 FILLER_70_1053 ();
 sg13g2_fill_1 FILLER_70_1060 ();
 sg13g2_fill_2 FILLER_70_1072 ();
 sg13g2_fill_2 FILLER_70_1081 ();
 sg13g2_fill_1 FILLER_70_1093 ();
 sg13g2_fill_1 FILLER_70_1120 ();
 sg13g2_fill_2 FILLER_70_1131 ();
 sg13g2_decap_8 FILLER_70_1185 ();
 sg13g2_decap_8 FILLER_70_1192 ();
 sg13g2_decap_8 FILLER_70_1199 ();
 sg13g2_decap_8 FILLER_70_1206 ();
 sg13g2_decap_4 FILLER_70_1213 ();
 sg13g2_fill_2 FILLER_70_1217 ();
 sg13g2_fill_2 FILLER_70_1249 ();
 sg13g2_decap_4 FILLER_70_1262 ();
 sg13g2_fill_2 FILLER_70_1266 ();
 sg13g2_fill_2 FILLER_70_1301 ();
 sg13g2_fill_1 FILLER_70_1319 ();
 sg13g2_fill_2 FILLER_70_1326 ();
 sg13g2_decap_8 FILLER_70_1362 ();
 sg13g2_decap_8 FILLER_70_1369 ();
 sg13g2_decap_8 FILLER_70_1376 ();
 sg13g2_decap_4 FILLER_70_1383 ();
 sg13g2_fill_2 FILLER_70_1387 ();
 sg13g2_fill_2 FILLER_70_1404 ();
 sg13g2_fill_2 FILLER_70_1417 ();
 sg13g2_decap_4 FILLER_70_1424 ();
 sg13g2_fill_2 FILLER_70_1428 ();
 sg13g2_decap_8 FILLER_70_1440 ();
 sg13g2_fill_2 FILLER_70_1447 ();
 sg13g2_fill_2 FILLER_70_1463 ();
 sg13g2_fill_1 FILLER_70_1465 ();
 sg13g2_fill_1 FILLER_70_1471 ();
 sg13g2_decap_8 FILLER_70_1477 ();
 sg13g2_decap_4 FILLER_70_1484 ();
 sg13g2_fill_2 FILLER_70_1488 ();
 sg13g2_fill_1 FILLER_70_1499 ();
 sg13g2_fill_2 FILLER_70_1503 ();
 sg13g2_fill_1 FILLER_70_1510 ();
 sg13g2_decap_8 FILLER_70_1524 ();
 sg13g2_decap_4 FILLER_70_1531 ();
 sg13g2_decap_8 FILLER_70_1552 ();
 sg13g2_decap_8 FILLER_70_1559 ();
 sg13g2_fill_2 FILLER_70_1566 ();
 sg13g2_fill_1 FILLER_70_1568 ();
 sg13g2_decap_4 FILLER_70_1579 ();
 sg13g2_fill_2 FILLER_70_1583 ();
 sg13g2_decap_8 FILLER_70_1603 ();
 sg13g2_decap_8 FILLER_70_1610 ();
 sg13g2_fill_2 FILLER_70_1617 ();
 sg13g2_fill_1 FILLER_70_1619 ();
 sg13g2_decap_8 FILLER_70_1653 ();
 sg13g2_fill_2 FILLER_70_1660 ();
 sg13g2_decap_8 FILLER_70_1666 ();
 sg13g2_fill_1 FILLER_70_1678 ();
 sg13g2_fill_1 FILLER_70_1683 ();
 sg13g2_fill_1 FILLER_70_1704 ();
 sg13g2_decap_4 FILLER_70_1711 ();
 sg13g2_fill_2 FILLER_70_1719 ();
 sg13g2_fill_2 FILLER_70_1733 ();
 sg13g2_fill_1 FILLER_70_1743 ();
 sg13g2_fill_1 FILLER_70_1783 ();
 sg13g2_decap_8 FILLER_70_1806 ();
 sg13g2_fill_2 FILLER_70_1838 ();
 sg13g2_fill_1 FILLER_70_1840 ();
 sg13g2_fill_2 FILLER_70_1858 ();
 sg13g2_decap_8 FILLER_70_1864 ();
 sg13g2_decap_8 FILLER_70_1871 ();
 sg13g2_decap_4 FILLER_70_1878 ();
 sg13g2_fill_2 FILLER_70_1882 ();
 sg13g2_fill_2 FILLER_70_1916 ();
 sg13g2_fill_2 FILLER_70_1925 ();
 sg13g2_fill_2 FILLER_70_1932 ();
 sg13g2_fill_1 FILLER_70_1934 ();
 sg13g2_fill_2 FILLER_70_1946 ();
 sg13g2_fill_1 FILLER_70_1976 ();
 sg13g2_fill_2 FILLER_70_2015 ();
 sg13g2_fill_1 FILLER_70_2017 ();
 sg13g2_decap_8 FILLER_70_2022 ();
 sg13g2_decap_4 FILLER_70_2029 ();
 sg13g2_fill_1 FILLER_70_2033 ();
 sg13g2_decap_8 FILLER_70_2038 ();
 sg13g2_fill_2 FILLER_70_2045 ();
 sg13g2_fill_1 FILLER_70_2052 ();
 sg13g2_fill_1 FILLER_70_2057 ();
 sg13g2_fill_2 FILLER_70_2067 ();
 sg13g2_fill_1 FILLER_70_2087 ();
 sg13g2_fill_1 FILLER_70_2107 ();
 sg13g2_fill_1 FILLER_70_2113 ();
 sg13g2_fill_1 FILLER_70_2122 ();
 sg13g2_fill_1 FILLER_70_2143 ();
 sg13g2_fill_1 FILLER_70_2149 ();
 sg13g2_decap_8 FILLER_70_2159 ();
 sg13g2_decap_8 FILLER_70_2166 ();
 sg13g2_decap_8 FILLER_70_2173 ();
 sg13g2_decap_4 FILLER_70_2180 ();
 sg13g2_fill_1 FILLER_70_2184 ();
 sg13g2_fill_2 FILLER_70_2189 ();
 sg13g2_fill_2 FILLER_70_2227 ();
 sg13g2_fill_1 FILLER_70_2254 ();
 sg13g2_fill_2 FILLER_70_2333 ();
 sg13g2_fill_1 FILLER_70_2335 ();
 sg13g2_decap_8 FILLER_70_2340 ();
 sg13g2_decap_8 FILLER_70_2347 ();
 sg13g2_fill_1 FILLER_70_2354 ();
 sg13g2_decap_4 FILLER_70_2360 ();
 sg13g2_fill_1 FILLER_70_2364 ();
 sg13g2_fill_1 FILLER_70_2379 ();
 sg13g2_decap_4 FILLER_70_2398 ();
 sg13g2_decap_4 FILLER_70_2416 ();
 sg13g2_fill_2 FILLER_70_2420 ();
 sg13g2_fill_2 FILLER_70_2426 ();
 sg13g2_fill_1 FILLER_70_2466 ();
 sg13g2_fill_1 FILLER_70_2497 ();
 sg13g2_fill_2 FILLER_70_2528 ();
 sg13g2_decap_8 FILLER_70_2543 ();
 sg13g2_decap_8 FILLER_70_2550 ();
 sg13g2_decap_4 FILLER_70_2557 ();
 sg13g2_fill_2 FILLER_70_2587 ();
 sg13g2_fill_1 FILLER_70_2589 ();
 sg13g2_decap_8 FILLER_70_2598 ();
 sg13g2_decap_8 FILLER_70_2605 ();
 sg13g2_decap_8 FILLER_70_2612 ();
 sg13g2_decap_8 FILLER_70_2619 ();
 sg13g2_decap_8 FILLER_70_2626 ();
 sg13g2_decap_8 FILLER_70_2633 ();
 sg13g2_decap_8 FILLER_70_2640 ();
 sg13g2_decap_8 FILLER_70_2647 ();
 sg13g2_decap_8 FILLER_70_2654 ();
 sg13g2_decap_8 FILLER_70_2661 ();
 sg13g2_fill_2 FILLER_70_2668 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_12 ();
 sg13g2_decap_8 FILLER_71_19 ();
 sg13g2_decap_4 FILLER_71_26 ();
 sg13g2_fill_2 FILLER_71_30 ();
 sg13g2_decap_8 FILLER_71_36 ();
 sg13g2_decap_4 FILLER_71_43 ();
 sg13g2_fill_1 FILLER_71_47 ();
 sg13g2_decap_4 FILLER_71_68 ();
 sg13g2_fill_2 FILLER_71_72 ();
 sg13g2_decap_4 FILLER_71_78 ();
 sg13g2_fill_1 FILLER_71_82 ();
 sg13g2_decap_8 FILLER_71_130 ();
 sg13g2_fill_2 FILLER_71_151 ();
 sg13g2_fill_1 FILLER_71_153 ();
 sg13g2_fill_2 FILLER_71_168 ();
 sg13g2_fill_2 FILLER_71_175 ();
 sg13g2_fill_2 FILLER_71_182 ();
 sg13g2_fill_1 FILLER_71_184 ();
 sg13g2_fill_1 FILLER_71_191 ();
 sg13g2_decap_4 FILLER_71_217 ();
 sg13g2_decap_4 FILLER_71_257 ();
 sg13g2_fill_2 FILLER_71_272 ();
 sg13g2_fill_1 FILLER_71_274 ();
 sg13g2_fill_1 FILLER_71_280 ();
 sg13g2_decap_4 FILLER_71_319 ();
 sg13g2_fill_2 FILLER_71_323 ();
 sg13g2_fill_2 FILLER_71_331 ();
 sg13g2_fill_1 FILLER_71_343 ();
 sg13g2_fill_2 FILLER_71_355 ();
 sg13g2_fill_2 FILLER_71_363 ();
 sg13g2_decap_8 FILLER_71_399 ();
 sg13g2_fill_2 FILLER_71_406 ();
 sg13g2_fill_2 FILLER_71_451 ();
 sg13g2_fill_1 FILLER_71_453 ();
 sg13g2_fill_2 FILLER_71_463 ();
 sg13g2_fill_1 FILLER_71_524 ();
 sg13g2_fill_2 FILLER_71_529 ();
 sg13g2_fill_2 FILLER_71_537 ();
 sg13g2_fill_2 FILLER_71_545 ();
 sg13g2_fill_1 FILLER_71_547 ();
 sg13g2_fill_1 FILLER_71_551 ();
 sg13g2_fill_2 FILLER_71_557 ();
 sg13g2_decap_8 FILLER_71_567 ();
 sg13g2_decap_4 FILLER_71_574 ();
 sg13g2_fill_1 FILLER_71_578 ();
 sg13g2_decap_8 FILLER_71_602 ();
 sg13g2_decap_8 FILLER_71_609 ();
 sg13g2_fill_1 FILLER_71_625 ();
 sg13g2_fill_1 FILLER_71_652 ();
 sg13g2_decap_8 FILLER_71_658 ();
 sg13g2_decap_4 FILLER_71_665 ();
 sg13g2_decap_8 FILLER_71_700 ();
 sg13g2_fill_2 FILLER_71_707 ();
 sg13g2_fill_1 FILLER_71_709 ();
 sg13g2_decap_8 FILLER_71_719 ();
 sg13g2_fill_1 FILLER_71_726 ();
 sg13g2_fill_2 FILLER_71_737 ();
 sg13g2_fill_1 FILLER_71_739 ();
 sg13g2_decap_4 FILLER_71_780 ();
 sg13g2_fill_2 FILLER_71_797 ();
 sg13g2_fill_1 FILLER_71_799 ();
 sg13g2_fill_1 FILLER_71_804 ();
 sg13g2_fill_1 FILLER_71_839 ();
 sg13g2_decap_4 FILLER_71_854 ();
 sg13g2_fill_1 FILLER_71_858 ();
 sg13g2_fill_1 FILLER_71_885 ();
 sg13g2_fill_2 FILLER_71_926 ();
 sg13g2_fill_1 FILLER_71_928 ();
 sg13g2_fill_2 FILLER_71_955 ();
 sg13g2_fill_2 FILLER_71_967 ();
 sg13g2_decap_4 FILLER_71_974 ();
 sg13g2_fill_2 FILLER_71_978 ();
 sg13g2_decap_4 FILLER_71_990 ();
 sg13g2_fill_1 FILLER_71_994 ();
 sg13g2_decap_8 FILLER_71_1016 ();
 sg13g2_decap_8 FILLER_71_1023 ();
 sg13g2_fill_1 FILLER_71_1035 ();
 sg13g2_fill_2 FILLER_71_1062 ();
 sg13g2_decap_4 FILLER_71_1070 ();
 sg13g2_decap_4 FILLER_71_1080 ();
 sg13g2_fill_2 FILLER_71_1157 ();
 sg13g2_fill_1 FILLER_71_1189 ();
 sg13g2_fill_2 FILLER_71_1200 ();
 sg13g2_decap_8 FILLER_71_1242 ();
 sg13g2_decap_4 FILLER_71_1249 ();
 sg13g2_fill_2 FILLER_71_1253 ();
 sg13g2_decap_4 FILLER_71_1263 ();
 sg13g2_fill_1 FILLER_71_1267 ();
 sg13g2_fill_1 FILLER_71_1318 ();
 sg13g2_fill_2 FILLER_71_1345 ();
 sg13g2_fill_2 FILLER_71_1350 ();
 sg13g2_decap_4 FILLER_71_1369 ();
 sg13g2_fill_1 FILLER_71_1373 ();
 sg13g2_fill_2 FILLER_71_1384 ();
 sg13g2_fill_1 FILLER_71_1393 ();
 sg13g2_fill_2 FILLER_71_1414 ();
 sg13g2_fill_2 FILLER_71_1421 ();
 sg13g2_fill_1 FILLER_71_1431 ();
 sg13g2_fill_1 FILLER_71_1453 ();
 sg13g2_decap_4 FILLER_71_1511 ();
 sg13g2_fill_2 FILLER_71_1515 ();
 sg13g2_fill_2 FILLER_71_1527 ();
 sg13g2_decap_8 FILLER_71_1555 ();
 sg13g2_decap_8 FILLER_71_1562 ();
 sg13g2_fill_2 FILLER_71_1579 ();
 sg13g2_fill_1 FILLER_71_1581 ();
 sg13g2_decap_8 FILLER_71_1608 ();
 sg13g2_fill_2 FILLER_71_1619 ();
 sg13g2_decap_4 FILLER_71_1634 ();
 sg13g2_fill_2 FILLER_71_1638 ();
 sg13g2_decap_4 FILLER_71_1708 ();
 sg13g2_fill_1 FILLER_71_1712 ();
 sg13g2_fill_1 FILLER_71_1757 ();
 sg13g2_fill_1 FILLER_71_1772 ();
 sg13g2_fill_1 FILLER_71_1777 ();
 sg13g2_decap_8 FILLER_71_1787 ();
 sg13g2_fill_1 FILLER_71_1794 ();
 sg13g2_decap_4 FILLER_71_1800 ();
 sg13g2_fill_1 FILLER_71_1804 ();
 sg13g2_decap_8 FILLER_71_1815 ();
 sg13g2_decap_4 FILLER_71_1822 ();
 sg13g2_fill_1 FILLER_71_1826 ();
 sg13g2_decap_4 FILLER_71_1834 ();
 sg13g2_fill_1 FILLER_71_1838 ();
 sg13g2_decap_8 FILLER_71_1843 ();
 sg13g2_decap_8 FILLER_71_1850 ();
 sg13g2_fill_1 FILLER_71_1891 ();
 sg13g2_fill_2 FILLER_71_1906 ();
 sg13g2_decap_8 FILLER_71_1915 ();
 sg13g2_decap_8 FILLER_71_1922 ();
 sg13g2_fill_2 FILLER_71_1929 ();
 sg13g2_fill_2 FILLER_71_1983 ();
 sg13g2_fill_1 FILLER_71_1998 ();
 sg13g2_decap_8 FILLER_71_2005 ();
 sg13g2_decap_4 FILLER_71_2012 ();
 sg13g2_fill_1 FILLER_71_2016 ();
 sg13g2_fill_1 FILLER_71_2037 ();
 sg13g2_fill_2 FILLER_71_2054 ();
 sg13g2_fill_1 FILLER_71_2056 ();
 sg13g2_fill_2 FILLER_71_2062 ();
 sg13g2_fill_1 FILLER_71_2064 ();
 sg13g2_fill_1 FILLER_71_2072 ();
 sg13g2_fill_2 FILLER_71_2088 ();
 sg13g2_fill_1 FILLER_71_2090 ();
 sg13g2_fill_1 FILLER_71_2115 ();
 sg13g2_fill_1 FILLER_71_2120 ();
 sg13g2_fill_2 FILLER_71_2125 ();
 sg13g2_fill_2 FILLER_71_2131 ();
 sg13g2_fill_1 FILLER_71_2133 ();
 sg13g2_decap_8 FILLER_71_2156 ();
 sg13g2_fill_2 FILLER_71_2163 ();
 sg13g2_fill_2 FILLER_71_2201 ();
 sg13g2_fill_1 FILLER_71_2308 ();
 sg13g2_decap_4 FILLER_71_2335 ();
 sg13g2_fill_1 FILLER_71_2339 ();
 sg13g2_decap_4 FILLER_71_2345 ();
 sg13g2_fill_1 FILLER_71_2349 ();
 sg13g2_fill_2 FILLER_71_2376 ();
 sg13g2_fill_1 FILLER_71_2378 ();
 sg13g2_decap_8 FILLER_71_2414 ();
 sg13g2_decap_4 FILLER_71_2421 ();
 sg13g2_fill_2 FILLER_71_2432 ();
 sg13g2_fill_1 FILLER_71_2460 ();
 sg13g2_fill_2 FILLER_71_2493 ();
 sg13g2_decap_4 FILLER_71_2501 ();
 sg13g2_decap_4 FILLER_71_2509 ();
 sg13g2_decap_4 FILLER_71_2518 ();
 sg13g2_fill_2 FILLER_71_2522 ();
 sg13g2_fill_1 FILLER_71_2540 ();
 sg13g2_fill_1 FILLER_71_2567 ();
 sg13g2_decap_8 FILLER_71_2576 ();
 sg13g2_decap_8 FILLER_71_2583 ();
 sg13g2_decap_8 FILLER_71_2590 ();
 sg13g2_decap_8 FILLER_71_2597 ();
 sg13g2_decap_8 FILLER_71_2604 ();
 sg13g2_decap_8 FILLER_71_2611 ();
 sg13g2_decap_8 FILLER_71_2618 ();
 sg13g2_decap_8 FILLER_71_2625 ();
 sg13g2_decap_8 FILLER_71_2632 ();
 sg13g2_decap_8 FILLER_71_2639 ();
 sg13g2_decap_8 FILLER_71_2646 ();
 sg13g2_decap_8 FILLER_71_2653 ();
 sg13g2_decap_8 FILLER_71_2660 ();
 sg13g2_fill_2 FILLER_71_2667 ();
 sg13g2_fill_1 FILLER_71_2669 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_fill_2 FILLER_72_14 ();
 sg13g2_fill_1 FILLER_72_16 ();
 sg13g2_fill_1 FILLER_72_43 ();
 sg13g2_fill_2 FILLER_72_75 ();
 sg13g2_fill_1 FILLER_72_77 ();
 sg13g2_fill_2 FILLER_72_129 ();
 sg13g2_fill_1 FILLER_72_131 ();
 sg13g2_fill_2 FILLER_72_225 ();
 sg13g2_decap_4 FILLER_72_263 ();
 sg13g2_fill_1 FILLER_72_272 ();
 sg13g2_decap_8 FILLER_72_311 ();
 sg13g2_decap_4 FILLER_72_323 ();
 sg13g2_fill_1 FILLER_72_327 ();
 sg13g2_fill_2 FILLER_72_346 ();
 sg13g2_fill_1 FILLER_72_366 ();
 sg13g2_fill_2 FILLER_72_373 ();
 sg13g2_decap_8 FILLER_72_386 ();
 sg13g2_decap_8 FILLER_72_393 ();
 sg13g2_decap_8 FILLER_72_400 ();
 sg13g2_decap_4 FILLER_72_407 ();
 sg13g2_fill_1 FILLER_72_411 ();
 sg13g2_fill_2 FILLER_72_417 ();
 sg13g2_decap_4 FILLER_72_424 ();
 sg13g2_decap_8 FILLER_72_437 ();
 sg13g2_decap_4 FILLER_72_449 ();
 sg13g2_fill_1 FILLER_72_453 ();
 sg13g2_fill_1 FILLER_72_459 ();
 sg13g2_fill_1 FILLER_72_493 ();
 sg13g2_fill_1 FILLER_72_507 ();
 sg13g2_fill_1 FILLER_72_522 ();
 sg13g2_fill_2 FILLER_72_528 ();
 sg13g2_fill_1 FILLER_72_530 ();
 sg13g2_fill_2 FILLER_72_539 ();
 sg13g2_fill_1 FILLER_72_546 ();
 sg13g2_fill_2 FILLER_72_551 ();
 sg13g2_fill_1 FILLER_72_553 ();
 sg13g2_fill_2 FILLER_72_580 ();
 sg13g2_fill_1 FILLER_72_582 ();
 sg13g2_fill_2 FILLER_72_587 ();
 sg13g2_decap_8 FILLER_72_630 ();
 sg13g2_fill_2 FILLER_72_637 ();
 sg13g2_decap_4 FILLER_72_649 ();
 sg13g2_fill_2 FILLER_72_683 ();
 sg13g2_decap_8 FILLER_72_689 ();
 sg13g2_decap_8 FILLER_72_696 ();
 sg13g2_decap_4 FILLER_72_703 ();
 sg13g2_fill_2 FILLER_72_743 ();
 sg13g2_fill_2 FILLER_72_760 ();
 sg13g2_fill_1 FILLER_72_762 ();
 sg13g2_fill_2 FILLER_72_793 ();
 sg13g2_fill_1 FILLER_72_795 ();
 sg13g2_decap_8 FILLER_72_801 ();
 sg13g2_decap_8 FILLER_72_808 ();
 sg13g2_fill_2 FILLER_72_815 ();
 sg13g2_fill_2 FILLER_72_821 ();
 sg13g2_fill_1 FILLER_72_823 ();
 sg13g2_fill_2 FILLER_72_834 ();
 sg13g2_fill_1 FILLER_72_836 ();
 sg13g2_fill_2 FILLER_72_852 ();
 sg13g2_fill_1 FILLER_72_868 ();
 sg13g2_decap_8 FILLER_72_877 ();
 sg13g2_decap_8 FILLER_72_884 ();
 sg13g2_fill_2 FILLER_72_891 ();
 sg13g2_fill_1 FILLER_72_893 ();
 sg13g2_decap_8 FILLER_72_903 ();
 sg13g2_fill_1 FILLER_72_910 ();
 sg13g2_decap_8 FILLER_72_934 ();
 sg13g2_decap_8 FILLER_72_941 ();
 sg13g2_decap_8 FILLER_72_948 ();
 sg13g2_fill_2 FILLER_72_955 ();
 sg13g2_fill_1 FILLER_72_967 ();
 sg13g2_fill_2 FILLER_72_994 ();
 sg13g2_decap_4 FILLER_72_1006 ();
 sg13g2_fill_1 FILLER_72_1010 ();
 sg13g2_fill_1 FILLER_72_1047 ();
 sg13g2_fill_2 FILLER_72_1084 ();
 sg13g2_fill_1 FILLER_72_1086 ();
 sg13g2_fill_2 FILLER_72_1113 ();
 sg13g2_fill_2 FILLER_72_1186 ();
 sg13g2_fill_1 FILLER_72_1214 ();
 sg13g2_fill_2 FILLER_72_1241 ();
 sg13g2_fill_1 FILLER_72_1269 ();
 sg13g2_decap_4 FILLER_72_1278 ();
 sg13g2_fill_1 FILLER_72_1286 ();
 sg13g2_fill_1 FILLER_72_1296 ();
 sg13g2_fill_1 FILLER_72_1307 ();
 sg13g2_fill_1 FILLER_72_1315 ();
 sg13g2_fill_1 FILLER_72_1324 ();
 sg13g2_fill_2 FILLER_72_1334 ();
 sg13g2_decap_4 FILLER_72_1377 ();
 sg13g2_fill_2 FILLER_72_1395 ();
 sg13g2_decap_4 FILLER_72_1412 ();
 sg13g2_fill_1 FILLER_72_1416 ();
 sg13g2_decap_4 FILLER_72_1430 ();
 sg13g2_fill_1 FILLER_72_1444 ();
 sg13g2_fill_1 FILLER_72_1478 ();
 sg13g2_fill_2 FILLER_72_1485 ();
 sg13g2_decap_4 FILLER_72_1500 ();
 sg13g2_fill_1 FILLER_72_1504 ();
 sg13g2_decap_8 FILLER_72_1518 ();
 sg13g2_decap_8 FILLER_72_1525 ();
 sg13g2_decap_4 FILLER_72_1532 ();
 sg13g2_fill_1 FILLER_72_1536 ();
 sg13g2_decap_8 FILLER_72_1541 ();
 sg13g2_decap_4 FILLER_72_1548 ();
 sg13g2_decap_4 FILLER_72_1556 ();
 sg13g2_fill_2 FILLER_72_1596 ();
 sg13g2_fill_2 FILLER_72_1624 ();
 sg13g2_fill_1 FILLER_72_1626 ();
 sg13g2_fill_2 FILLER_72_1649 ();
 sg13g2_fill_1 FILLER_72_1663 ();
 sg13g2_fill_1 FILLER_72_1700 ();
 sg13g2_decap_4 FILLER_72_1717 ();
 sg13g2_fill_1 FILLER_72_1721 ();
 sg13g2_fill_2 FILLER_72_1733 ();
 sg13g2_decap_4 FILLER_72_1783 ();
 sg13g2_fill_1 FILLER_72_1787 ();
 sg13g2_decap_8 FILLER_72_1796 ();
 sg13g2_decap_4 FILLER_72_1803 ();
 sg13g2_fill_1 FILLER_72_1807 ();
 sg13g2_fill_1 FILLER_72_1817 ();
 sg13g2_decap_8 FILLER_72_1822 ();
 sg13g2_decap_8 FILLER_72_1829 ();
 sg13g2_decap_8 FILLER_72_1836 ();
 sg13g2_decap_8 FILLER_72_1843 ();
 sg13g2_decap_8 FILLER_72_1850 ();
 sg13g2_fill_2 FILLER_72_1857 ();
 sg13g2_fill_2 FILLER_72_1863 ();
 sg13g2_fill_1 FILLER_72_1875 ();
 sg13g2_decap_8 FILLER_72_1888 ();
 sg13g2_decap_8 FILLER_72_1930 ();
 sg13g2_fill_2 FILLER_72_1963 ();
 sg13g2_fill_1 FILLER_72_1969 ();
 sg13g2_fill_1 FILLER_72_1980 ();
 sg13g2_decap_4 FILLER_72_1990 ();
 sg13g2_fill_2 FILLER_72_1998 ();
 sg13g2_fill_2 FILLER_72_2010 ();
 sg13g2_decap_4 FILLER_72_2021 ();
 sg13g2_fill_1 FILLER_72_2038 ();
 sg13g2_fill_1 FILLER_72_2044 ();
 sg13g2_fill_1 FILLER_72_2052 ();
 sg13g2_fill_1 FILLER_72_2061 ();
 sg13g2_fill_2 FILLER_72_2070 ();
 sg13g2_fill_2 FILLER_72_2081 ();
 sg13g2_fill_1 FILLER_72_2093 ();
 sg13g2_decap_8 FILLER_72_2151 ();
 sg13g2_fill_2 FILLER_72_2158 ();
 sg13g2_fill_1 FILLER_72_2160 ();
 sg13g2_fill_1 FILLER_72_2174 ();
 sg13g2_decap_4 FILLER_72_2194 ();
 sg13g2_fill_1 FILLER_72_2198 ();
 sg13g2_fill_1 FILLER_72_2216 ();
 sg13g2_fill_1 FILLER_72_2222 ();
 sg13g2_fill_2 FILLER_72_2228 ();
 sg13g2_fill_1 FILLER_72_2240 ();
 sg13g2_fill_1 FILLER_72_2275 ();
 sg13g2_fill_1 FILLER_72_2299 ();
 sg13g2_fill_2 FILLER_72_2320 ();
 sg13g2_fill_2 FILLER_72_2328 ();
 sg13g2_fill_1 FILLER_72_2330 ();
 sg13g2_decap_4 FILLER_72_2371 ();
 sg13g2_decap_4 FILLER_72_2414 ();
 sg13g2_fill_2 FILLER_72_2418 ();
 sg13g2_decap_4 FILLER_72_2425 ();
 sg13g2_decap_8 FILLER_72_2438 ();
 sg13g2_fill_2 FILLER_72_2445 ();
 sg13g2_fill_2 FILLER_72_2458 ();
 sg13g2_fill_1 FILLER_72_2460 ();
 sg13g2_fill_2 FILLER_72_2466 ();
 sg13g2_fill_1 FILLER_72_2472 ();
 sg13g2_fill_1 FILLER_72_2481 ();
 sg13g2_fill_1 FILLER_72_2491 ();
 sg13g2_fill_1 FILLER_72_2498 ();
 sg13g2_fill_2 FILLER_72_2508 ();
 sg13g2_fill_1 FILLER_72_2524 ();
 sg13g2_decap_8 FILLER_72_2574 ();
 sg13g2_decap_8 FILLER_72_2581 ();
 sg13g2_decap_8 FILLER_72_2588 ();
 sg13g2_decap_8 FILLER_72_2595 ();
 sg13g2_decap_8 FILLER_72_2602 ();
 sg13g2_decap_8 FILLER_72_2609 ();
 sg13g2_decap_8 FILLER_72_2616 ();
 sg13g2_decap_8 FILLER_72_2623 ();
 sg13g2_decap_8 FILLER_72_2630 ();
 sg13g2_decap_8 FILLER_72_2637 ();
 sg13g2_decap_8 FILLER_72_2644 ();
 sg13g2_decap_8 FILLER_72_2651 ();
 sg13g2_decap_8 FILLER_72_2658 ();
 sg13g2_decap_4 FILLER_72_2665 ();
 sg13g2_fill_1 FILLER_72_2669 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_7 ();
 sg13g2_fill_1 FILLER_73_9 ();
 sg13g2_decap_4 FILLER_73_14 ();
 sg13g2_fill_2 FILLER_73_22 ();
 sg13g2_fill_2 FILLER_73_34 ();
 sg13g2_decap_4 FILLER_73_50 ();
 sg13g2_fill_1 FILLER_73_94 ();
 sg13g2_decap_8 FILLER_73_99 ();
 sg13g2_decap_4 FILLER_73_116 ();
 sg13g2_fill_2 FILLER_73_120 ();
 sg13g2_decap_4 FILLER_73_132 ();
 sg13g2_fill_1 FILLER_73_136 ();
 sg13g2_fill_2 FILLER_73_145 ();
 sg13g2_fill_2 FILLER_73_151 ();
 sg13g2_fill_1 FILLER_73_153 ();
 sg13g2_fill_2 FILLER_73_159 ();
 sg13g2_fill_1 FILLER_73_161 ();
 sg13g2_fill_1 FILLER_73_177 ();
 sg13g2_fill_1 FILLER_73_183 ();
 sg13g2_fill_2 FILLER_73_192 ();
 sg13g2_fill_1 FILLER_73_194 ();
 sg13g2_decap_4 FILLER_73_232 ();
 sg13g2_fill_2 FILLER_73_240 ();
 sg13g2_fill_1 FILLER_73_242 ();
 sg13g2_decap_8 FILLER_73_247 ();
 sg13g2_decap_4 FILLER_73_254 ();
 sg13g2_decap_4 FILLER_73_272 ();
 sg13g2_fill_1 FILLER_73_298 ();
 sg13g2_decap_4 FILLER_73_303 ();
 sg13g2_decap_8 FILLER_73_317 ();
 sg13g2_decap_8 FILLER_73_324 ();
 sg13g2_decap_8 FILLER_73_375 ();
 sg13g2_decap_8 FILLER_73_382 ();
 sg13g2_decap_8 FILLER_73_389 ();
 sg13g2_fill_1 FILLER_73_426 ();
 sg13g2_decap_8 FILLER_73_432 ();
 sg13g2_decap_8 FILLER_73_439 ();
 sg13g2_decap_8 FILLER_73_446 ();
 sg13g2_fill_1 FILLER_73_453 ();
 sg13g2_fill_1 FILLER_73_463 ();
 sg13g2_fill_2 FILLER_73_472 ();
 sg13g2_fill_1 FILLER_73_474 ();
 sg13g2_fill_2 FILLER_73_481 ();
 sg13g2_fill_1 FILLER_73_483 ();
 sg13g2_fill_2 FILLER_73_563 ();
 sg13g2_fill_2 FILLER_73_580 ();
 sg13g2_fill_1 FILLER_73_582 ();
 sg13g2_fill_2 FILLER_73_644 ();
 sg13g2_fill_1 FILLER_73_655 ();
 sg13g2_fill_2 FILLER_73_665 ();
 sg13g2_decap_4 FILLER_73_677 ();
 sg13g2_fill_1 FILLER_73_681 ();
 sg13g2_decap_4 FILLER_73_687 ();
 sg13g2_decap_8 FILLER_73_695 ();
 sg13g2_fill_2 FILLER_73_702 ();
 sg13g2_fill_2 FILLER_73_709 ();
 sg13g2_fill_1 FILLER_73_711 ();
 sg13g2_fill_1 FILLER_73_716 ();
 sg13g2_fill_2 FILLER_73_743 ();
 sg13g2_fill_2 FILLER_73_771 ();
 sg13g2_decap_8 FILLER_73_812 ();
 sg13g2_decap_4 FILLER_73_819 ();
 sg13g2_fill_2 FILLER_73_823 ();
 sg13g2_decap_8 FILLER_73_829 ();
 sg13g2_decap_8 FILLER_73_836 ();
 sg13g2_decap_8 FILLER_73_843 ();
 sg13g2_fill_2 FILLER_73_854 ();
 sg13g2_decap_8 FILLER_73_882 ();
 sg13g2_decap_8 FILLER_73_889 ();
 sg13g2_decap_8 FILLER_73_896 ();
 sg13g2_decap_4 FILLER_73_913 ();
 sg13g2_fill_2 FILLER_73_917 ();
 sg13g2_fill_2 FILLER_73_991 ();
 sg13g2_fill_2 FILLER_73_997 ();
 sg13g2_fill_1 FILLER_73_1071 ();
 sg13g2_fill_1 FILLER_73_1076 ();
 sg13g2_fill_1 FILLER_73_1087 ();
 sg13g2_fill_1 FILLER_73_1102 ();
 sg13g2_fill_1 FILLER_73_1107 ();
 sg13g2_fill_1 FILLER_73_1179 ();
 sg13g2_decap_8 FILLER_73_1234 ();
 sg13g2_fill_1 FILLER_73_1241 ();
 sg13g2_fill_1 FILLER_73_1252 ();
 sg13g2_decap_8 FILLER_73_1257 ();
 sg13g2_decap_8 FILLER_73_1264 ();
 sg13g2_fill_1 FILLER_73_1271 ();
 sg13g2_decap_4 FILLER_73_1280 ();
 sg13g2_fill_1 FILLER_73_1342 ();
 sg13g2_fill_1 FILLER_73_1348 ();
 sg13g2_fill_1 FILLER_73_1356 ();
 sg13g2_fill_1 FILLER_73_1388 ();
 sg13g2_decap_4 FILLER_73_1401 ();
 sg13g2_fill_2 FILLER_73_1415 ();
 sg13g2_fill_1 FILLER_73_1417 ();
 sg13g2_fill_2 FILLER_73_1448 ();
 sg13g2_fill_2 FILLER_73_1455 ();
 sg13g2_fill_1 FILLER_73_1457 ();
 sg13g2_fill_1 FILLER_73_1461 ();
 sg13g2_fill_2 FILLER_73_1482 ();
 sg13g2_fill_1 FILLER_73_1484 ();
 sg13g2_fill_2 FILLER_73_1490 ();
 sg13g2_fill_1 FILLER_73_1497 ();
 sg13g2_fill_2 FILLER_73_1524 ();
 sg13g2_fill_1 FILLER_73_1526 ();
 sg13g2_decap_8 FILLER_73_1563 ();
 sg13g2_decap_8 FILLER_73_1570 ();
 sg13g2_fill_2 FILLER_73_1581 ();
 sg13g2_fill_1 FILLER_73_1609 ();
 sg13g2_decap_4 FILLER_73_1614 ();
 sg13g2_fill_2 FILLER_73_1618 ();
 sg13g2_decap_4 FILLER_73_1624 ();
 sg13g2_fill_2 FILLER_73_1632 ();
 sg13g2_fill_2 FILLER_73_1663 ();
 sg13g2_fill_1 FILLER_73_1665 ();
 sg13g2_fill_2 FILLER_73_1670 ();
 sg13g2_fill_2 FILLER_73_1678 ();
 sg13g2_decap_4 FILLER_73_1706 ();
 sg13g2_fill_2 FILLER_73_1710 ();
 sg13g2_decap_8 FILLER_73_1715 ();
 sg13g2_decap_4 FILLER_73_1722 ();
 sg13g2_fill_2 FILLER_73_1743 ();
 sg13g2_fill_1 FILLER_73_1766 ();
 sg13g2_decap_8 FILLER_73_1784 ();
 sg13g2_fill_2 FILLER_73_1791 ();
 sg13g2_fill_1 FILLER_73_1798 ();
 sg13g2_fill_2 FILLER_73_1803 ();
 sg13g2_fill_2 FILLER_73_1810 ();
 sg13g2_fill_2 FILLER_73_1818 ();
 sg13g2_fill_1 FILLER_73_1820 ();
 sg13g2_decap_4 FILLER_73_1826 ();
 sg13g2_decap_4 FILLER_73_1834 ();
 sg13g2_decap_8 FILLER_73_1843 ();
 sg13g2_decap_4 FILLER_73_1850 ();
 sg13g2_fill_1 FILLER_73_1854 ();
 sg13g2_fill_1 FILLER_73_1874 ();
 sg13g2_decap_8 FILLER_73_1879 ();
 sg13g2_decap_4 FILLER_73_1886 ();
 sg13g2_fill_2 FILLER_73_1890 ();
 sg13g2_fill_1 FILLER_73_1926 ();
 sg13g2_decap_8 FILLER_73_1932 ();
 sg13g2_decap_4 FILLER_73_1939 ();
 sg13g2_decap_4 FILLER_73_1954 ();
 sg13g2_fill_2 FILLER_73_1997 ();
 sg13g2_fill_1 FILLER_73_1999 ();
 sg13g2_fill_1 FILLER_73_2015 ();
 sg13g2_fill_1 FILLER_73_2053 ();
 sg13g2_fill_1 FILLER_73_2064 ();
 sg13g2_fill_1 FILLER_73_2070 ();
 sg13g2_fill_1 FILLER_73_2075 ();
 sg13g2_fill_1 FILLER_73_2086 ();
 sg13g2_fill_2 FILLER_73_2099 ();
 sg13g2_fill_1 FILLER_73_2101 ();
 sg13g2_fill_1 FILLER_73_2123 ();
 sg13g2_fill_1 FILLER_73_2137 ();
 sg13g2_fill_2 FILLER_73_2142 ();
 sg13g2_fill_1 FILLER_73_2144 ();
 sg13g2_decap_8 FILLER_73_2150 ();
 sg13g2_fill_1 FILLER_73_2157 ();
 sg13g2_decap_8 FILLER_73_2194 ();
 sg13g2_fill_2 FILLER_73_2201 ();
 sg13g2_fill_2 FILLER_73_2233 ();
 sg13g2_fill_1 FILLER_73_2275 ();
 sg13g2_fill_2 FILLER_73_2336 ();
 sg13g2_fill_1 FILLER_73_2338 ();
 sg13g2_decap_4 FILLER_73_2374 ();
 sg13g2_fill_1 FILLER_73_2378 ();
 sg13g2_decap_4 FILLER_73_2390 ();
 sg13g2_fill_2 FILLER_73_2394 ();
 sg13g2_fill_1 FILLER_73_2402 ();
 sg13g2_decap_4 FILLER_73_2417 ();
 sg13g2_fill_1 FILLER_73_2460 ();
 sg13g2_fill_2 FILLER_73_2466 ();
 sg13g2_fill_1 FILLER_73_2533 ();
 sg13g2_decap_8 FILLER_73_2591 ();
 sg13g2_decap_8 FILLER_73_2598 ();
 sg13g2_decap_8 FILLER_73_2605 ();
 sg13g2_decap_8 FILLER_73_2612 ();
 sg13g2_decap_8 FILLER_73_2619 ();
 sg13g2_decap_8 FILLER_73_2626 ();
 sg13g2_decap_8 FILLER_73_2633 ();
 sg13g2_decap_8 FILLER_73_2640 ();
 sg13g2_decap_8 FILLER_73_2647 ();
 sg13g2_decap_8 FILLER_73_2654 ();
 sg13g2_decap_8 FILLER_73_2661 ();
 sg13g2_fill_2 FILLER_73_2668 ();
 sg13g2_decap_4 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_30 ();
 sg13g2_fill_2 FILLER_74_37 ();
 sg13g2_fill_2 FILLER_74_65 ();
 sg13g2_fill_2 FILLER_74_71 ();
 sg13g2_fill_1 FILLER_74_73 ();
 sg13g2_fill_1 FILLER_74_82 ();
 sg13g2_decap_4 FILLER_74_104 ();
 sg13g2_fill_2 FILLER_74_118 ();
 sg13g2_fill_1 FILLER_74_120 ();
 sg13g2_decap_4 FILLER_74_136 ();
 sg13g2_fill_1 FILLER_74_140 ();
 sg13g2_decap_8 FILLER_74_145 ();
 sg13g2_decap_8 FILLER_74_152 ();
 sg13g2_decap_4 FILLER_74_159 ();
 sg13g2_fill_2 FILLER_74_163 ();
 sg13g2_fill_1 FILLER_74_202 ();
 sg13g2_fill_1 FILLER_74_260 ();
 sg13g2_fill_1 FILLER_74_265 ();
 sg13g2_fill_1 FILLER_74_270 ();
 sg13g2_fill_2 FILLER_74_279 ();
 sg13g2_fill_1 FILLER_74_281 ();
 sg13g2_fill_2 FILLER_74_316 ();
 sg13g2_fill_1 FILLER_74_318 ();
 sg13g2_fill_2 FILLER_74_323 ();
 sg13g2_decap_4 FILLER_74_332 ();
 sg13g2_fill_2 FILLER_74_341 ();
 sg13g2_fill_2 FILLER_74_393 ();
 sg13g2_fill_1 FILLER_74_395 ();
 sg13g2_decap_8 FILLER_74_422 ();
 sg13g2_decap_4 FILLER_74_429 ();
 sg13g2_fill_2 FILLER_74_433 ();
 sg13g2_fill_1 FILLER_74_442 ();
 sg13g2_fill_2 FILLER_74_569 ();
 sg13g2_fill_1 FILLER_74_597 ();
 sg13g2_fill_2 FILLER_74_606 ();
 sg13g2_fill_1 FILLER_74_608 ();
 sg13g2_fill_1 FILLER_74_613 ();
 sg13g2_fill_1 FILLER_74_640 ();
 sg13g2_fill_1 FILLER_74_646 ();
 sg13g2_fill_1 FILLER_74_656 ();
 sg13g2_fill_1 FILLER_74_683 ();
 sg13g2_fill_2 FILLER_74_720 ();
 sg13g2_fill_1 FILLER_74_722 ();
 sg13g2_fill_1 FILLER_74_727 ();
 sg13g2_fill_1 FILLER_74_738 ();
 sg13g2_decap_4 FILLER_74_756 ();
 sg13g2_decap_8 FILLER_74_773 ();
 sg13g2_fill_2 FILLER_74_813 ();
 sg13g2_fill_1 FILLER_74_815 ();
 sg13g2_decap_4 FILLER_74_864 ();
 sg13g2_fill_1 FILLER_74_868 ();
 sg13g2_decap_8 FILLER_74_883 ();
 sg13g2_fill_1 FILLER_74_890 ();
 sg13g2_decap_8 FILLER_74_955 ();
 sg13g2_fill_1 FILLER_74_973 ();
 sg13g2_decap_8 FILLER_74_978 ();
 sg13g2_decap_8 FILLER_74_985 ();
 sg13g2_fill_1 FILLER_74_992 ();
 sg13g2_decap_8 FILLER_74_997 ();
 sg13g2_fill_2 FILLER_74_1004 ();
 sg13g2_fill_1 FILLER_74_1006 ();
 sg13g2_fill_1 FILLER_74_1023 ();
 sg13g2_decap_8 FILLER_74_1034 ();
 sg13g2_decap_4 FILLER_74_1057 ();
 sg13g2_fill_1 FILLER_74_1061 ();
 sg13g2_decap_8 FILLER_74_1078 ();
 sg13g2_decap_4 FILLER_74_1085 ();
 sg13g2_fill_2 FILLER_74_1089 ();
 sg13g2_fill_2 FILLER_74_1126 ();
 sg13g2_fill_2 FILLER_74_1168 ();
 sg13g2_fill_2 FILLER_74_1191 ();
 sg13g2_fill_1 FILLER_74_1193 ();
 sg13g2_decap_8 FILLER_74_1198 ();
 sg13g2_decap_4 FILLER_74_1215 ();
 sg13g2_fill_2 FILLER_74_1219 ();
 sg13g2_fill_2 FILLER_74_1224 ();
 sg13g2_fill_2 FILLER_74_1230 ();
 sg13g2_fill_1 FILLER_74_1232 ();
 sg13g2_decap_4 FILLER_74_1259 ();
 sg13g2_fill_2 FILLER_74_1263 ();
 sg13g2_fill_2 FILLER_74_1301 ();
 sg13g2_fill_2 FILLER_74_1311 ();
 sg13g2_fill_1 FILLER_74_1313 ();
 sg13g2_fill_2 FILLER_74_1333 ();
 sg13g2_fill_1 FILLER_74_1335 ();
 sg13g2_fill_2 FILLER_74_1345 ();
 sg13g2_fill_1 FILLER_74_1377 ();
 sg13g2_fill_2 FILLER_74_1395 ();
 sg13g2_decap_8 FILLER_74_1407 ();
 sg13g2_fill_1 FILLER_74_1414 ();
 sg13g2_fill_2 FILLER_74_1429 ();
 sg13g2_decap_4 FILLER_74_1436 ();
 sg13g2_fill_2 FILLER_74_1447 ();
 sg13g2_fill_1 FILLER_74_1484 ();
 sg13g2_fill_1 FILLER_74_1489 ();
 sg13g2_decap_4 FILLER_74_1495 ();
 sg13g2_fill_1 FILLER_74_1499 ();
 sg13g2_decap_8 FILLER_74_1509 ();
 sg13g2_decap_4 FILLER_74_1516 ();
 sg13g2_fill_1 FILLER_74_1520 ();
 sg13g2_fill_2 FILLER_74_1531 ();
 sg13g2_fill_2 FILLER_74_1559 ();
 sg13g2_fill_1 FILLER_74_1561 ();
 sg13g2_decap_8 FILLER_74_1566 ();
 sg13g2_decap_4 FILLER_74_1573 ();
 sg13g2_fill_2 FILLER_74_1577 ();
 sg13g2_decap_4 FILLER_74_1587 ();
 sg13g2_decap_8 FILLER_74_1595 ();
 sg13g2_decap_8 FILLER_74_1602 ();
 sg13g2_decap_8 FILLER_74_1609 ();
 sg13g2_decap_8 FILLER_74_1616 ();
 sg13g2_decap_4 FILLER_74_1623 ();
 sg13g2_fill_1 FILLER_74_1627 ();
 sg13g2_fill_1 FILLER_74_1649 ();
 sg13g2_fill_1 FILLER_74_1654 ();
 sg13g2_fill_1 FILLER_74_1660 ();
 sg13g2_fill_1 FILLER_74_1666 ();
 sg13g2_fill_1 FILLER_74_1672 ();
 sg13g2_fill_1 FILLER_74_1677 ();
 sg13g2_fill_1 FILLER_74_1683 ();
 sg13g2_decap_4 FILLER_74_1688 ();
 sg13g2_fill_2 FILLER_74_1692 ();
 sg13g2_fill_1 FILLER_74_1697 ();
 sg13g2_fill_1 FILLER_74_1708 ();
 sg13g2_fill_2 FILLER_74_1719 ();
 sg13g2_fill_1 FILLER_74_1721 ();
 sg13g2_decap_8 FILLER_74_1727 ();
 sg13g2_fill_2 FILLER_74_1734 ();
 sg13g2_decap_8 FILLER_74_1746 ();
 sg13g2_fill_1 FILLER_74_1753 ();
 sg13g2_fill_1 FILLER_74_1757 ();
 sg13g2_fill_2 FILLER_74_1778 ();
 sg13g2_fill_1 FILLER_74_1780 ();
 sg13g2_decap_8 FILLER_74_1787 ();
 sg13g2_fill_1 FILLER_74_1794 ();
 sg13g2_fill_1 FILLER_74_1808 ();
 sg13g2_fill_2 FILLER_74_1823 ();
 sg13g2_decap_4 FILLER_74_1847 ();
 sg13g2_fill_2 FILLER_74_1851 ();
 sg13g2_decap_8 FILLER_74_1886 ();
 sg13g2_decap_4 FILLER_74_1898 ();
 sg13g2_decap_8 FILLER_74_1919 ();
 sg13g2_fill_2 FILLER_74_1926 ();
 sg13g2_decap_8 FILLER_74_1933 ();
 sg13g2_decap_4 FILLER_74_1940 ();
 sg13g2_fill_2 FILLER_74_1944 ();
 sg13g2_decap_8 FILLER_74_1949 ();
 sg13g2_decap_4 FILLER_74_1956 ();
 sg13g2_fill_1 FILLER_74_1960 ();
 sg13g2_fill_2 FILLER_74_1966 ();
 sg13g2_fill_1 FILLER_74_1968 ();
 sg13g2_fill_2 FILLER_74_1974 ();
 sg13g2_fill_2 FILLER_74_1988 ();
 sg13g2_fill_1 FILLER_74_1990 ();
 sg13g2_fill_2 FILLER_74_2000 ();
 sg13g2_fill_1 FILLER_74_2006 ();
 sg13g2_fill_2 FILLER_74_2017 ();
 sg13g2_fill_1 FILLER_74_2019 ();
 sg13g2_fill_1 FILLER_74_2040 ();
 sg13g2_decap_4 FILLER_74_2066 ();
 sg13g2_fill_1 FILLER_74_2070 ();
 sg13g2_fill_1 FILLER_74_2080 ();
 sg13g2_fill_1 FILLER_74_2126 ();
 sg13g2_decap_4 FILLER_74_2131 ();
 sg13g2_fill_1 FILLER_74_2135 ();
 sg13g2_fill_1 FILLER_74_2144 ();
 sg13g2_decap_8 FILLER_74_2207 ();
 sg13g2_fill_1 FILLER_74_2214 ();
 sg13g2_fill_1 FILLER_74_2260 ();
 sg13g2_fill_1 FILLER_74_2275 ();
 sg13g2_fill_2 FILLER_74_2304 ();
 sg13g2_fill_2 FILLER_74_2310 ();
 sg13g2_fill_1 FILLER_74_2317 ();
 sg13g2_fill_1 FILLER_74_2326 ();
 sg13g2_fill_1 FILLER_74_2333 ();
 sg13g2_fill_1 FILLER_74_2347 ();
 sg13g2_fill_2 FILLER_74_2383 ();
 sg13g2_fill_1 FILLER_74_2385 ();
 sg13g2_fill_2 FILLER_74_2424 ();
 sg13g2_fill_1 FILLER_74_2426 ();
 sg13g2_decap_4 FILLER_74_2431 ();
 sg13g2_fill_1 FILLER_74_2439 ();
 sg13g2_fill_1 FILLER_74_2455 ();
 sg13g2_fill_2 FILLER_74_2487 ();
 sg13g2_fill_1 FILLER_74_2489 ();
 sg13g2_fill_2 FILLER_74_2496 ();
 sg13g2_fill_1 FILLER_74_2503 ();
 sg13g2_fill_2 FILLER_74_2530 ();
 sg13g2_fill_2 FILLER_74_2560 ();
 sg13g2_decap_8 FILLER_74_2596 ();
 sg13g2_decap_8 FILLER_74_2603 ();
 sg13g2_decap_8 FILLER_74_2610 ();
 sg13g2_decap_8 FILLER_74_2617 ();
 sg13g2_decap_8 FILLER_74_2624 ();
 sg13g2_decap_8 FILLER_74_2631 ();
 sg13g2_decap_8 FILLER_74_2638 ();
 sg13g2_decap_8 FILLER_74_2645 ();
 sg13g2_decap_8 FILLER_74_2652 ();
 sg13g2_decap_8 FILLER_74_2659 ();
 sg13g2_decap_4 FILLER_74_2666 ();
 sg13g2_fill_2 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_38 ();
 sg13g2_fill_1 FILLER_75_45 ();
 sg13g2_decap_8 FILLER_75_59 ();
 sg13g2_fill_2 FILLER_75_66 ();
 sg13g2_decap_4 FILLER_75_78 ();
 sg13g2_fill_1 FILLER_75_82 ();
 sg13g2_fill_2 FILLER_75_104 ();
 sg13g2_fill_1 FILLER_75_106 ();
 sg13g2_decap_4 FILLER_75_112 ();
 sg13g2_fill_1 FILLER_75_147 ();
 sg13g2_decap_8 FILLER_75_157 ();
 sg13g2_decap_8 FILLER_75_164 ();
 sg13g2_fill_2 FILLER_75_171 ();
 sg13g2_decap_4 FILLER_75_177 ();
 sg13g2_fill_1 FILLER_75_198 ();
 sg13g2_fill_2 FILLER_75_233 ();
 sg13g2_fill_1 FILLER_75_240 ();
 sg13g2_decap_8 FILLER_75_270 ();
 sg13g2_decap_4 FILLER_75_277 ();
 sg13g2_fill_1 FILLER_75_281 ();
 sg13g2_fill_1 FILLER_75_288 ();
 sg13g2_fill_2 FILLER_75_351 ();
 sg13g2_fill_1 FILLER_75_353 ();
 sg13g2_decap_8 FILLER_75_359 ();
 sg13g2_decap_4 FILLER_75_366 ();
 sg13g2_fill_2 FILLER_75_370 ();
 sg13g2_decap_8 FILLER_75_376 ();
 sg13g2_decap_8 FILLER_75_383 ();
 sg13g2_decap_4 FILLER_75_390 ();
 sg13g2_decap_4 FILLER_75_415 ();
 sg13g2_fill_1 FILLER_75_419 ();
 sg13g2_decap_4 FILLER_75_424 ();
 sg13g2_fill_2 FILLER_75_428 ();
 sg13g2_fill_1 FILLER_75_449 ();
 sg13g2_fill_2 FILLER_75_465 ();
 sg13g2_decap_8 FILLER_75_500 ();
 sg13g2_fill_2 FILLER_75_507 ();
 sg13g2_fill_1 FILLER_75_509 ();
 sg13g2_fill_2 FILLER_75_528 ();
 sg13g2_fill_2 FILLER_75_563 ();
 sg13g2_decap_4 FILLER_75_576 ();
 sg13g2_fill_1 FILLER_75_580 ();
 sg13g2_fill_1 FILLER_75_596 ();
 sg13g2_fill_2 FILLER_75_607 ();
 sg13g2_decap_8 FILLER_75_631 ();
 sg13g2_decap_4 FILLER_75_638 ();
 sg13g2_fill_2 FILLER_75_642 ();
 sg13g2_decap_8 FILLER_75_649 ();
 sg13g2_decap_4 FILLER_75_675 ();
 sg13g2_fill_2 FILLER_75_679 ();
 sg13g2_decap_8 FILLER_75_717 ();
 sg13g2_decap_8 FILLER_75_724 ();
 sg13g2_decap_8 FILLER_75_731 ();
 sg13g2_decap_4 FILLER_75_738 ();
 sg13g2_fill_1 FILLER_75_742 ();
 sg13g2_decap_4 FILLER_75_757 ();
 sg13g2_fill_1 FILLER_75_761 ();
 sg13g2_fill_1 FILLER_75_792 ();
 sg13g2_decap_8 FILLER_75_798 ();
 sg13g2_fill_2 FILLER_75_805 ();
 sg13g2_fill_1 FILLER_75_843 ();
 sg13g2_decap_4 FILLER_75_862 ();
 sg13g2_fill_2 FILLER_75_866 ();
 sg13g2_decap_4 FILLER_75_878 ();
 sg13g2_fill_2 FILLER_75_908 ();
 sg13g2_fill_1 FILLER_75_910 ();
 sg13g2_decap_4 FILLER_75_946 ();
 sg13g2_fill_1 FILLER_75_980 ();
 sg13g2_fill_2 FILLER_75_985 ();
 sg13g2_decap_8 FILLER_75_1013 ();
 sg13g2_fill_2 FILLER_75_1020 ();
 sg13g2_decap_4 FILLER_75_1028 ();
 sg13g2_fill_2 FILLER_75_1032 ();
 sg13g2_fill_2 FILLER_75_1059 ();
 sg13g2_decap_8 FILLER_75_1135 ();
 sg13g2_decap_8 FILLER_75_1142 ();
 sg13g2_decap_8 FILLER_75_1149 ();
 sg13g2_decap_8 FILLER_75_1156 ();
 sg13g2_fill_1 FILLER_75_1163 ();
 sg13g2_decap_8 FILLER_75_1190 ();
 sg13g2_decap_4 FILLER_75_1197 ();
 sg13g2_fill_1 FILLER_75_1201 ();
 sg13g2_fill_2 FILLER_75_1207 ();
 sg13g2_fill_2 FILLER_75_1254 ();
 sg13g2_decap_8 FILLER_75_1299 ();
 sg13g2_fill_2 FILLER_75_1306 ();
 sg13g2_decap_8 FILLER_75_1346 ();
 sg13g2_fill_2 FILLER_75_1353 ();
 sg13g2_fill_1 FILLER_75_1355 ();
 sg13g2_decap_8 FILLER_75_1409 ();
 sg13g2_fill_2 FILLER_75_1416 ();
 sg13g2_fill_1 FILLER_75_1418 ();
 sg13g2_fill_2 FILLER_75_1445 ();
 sg13g2_fill_2 FILLER_75_1473 ();
 sg13g2_fill_2 FILLER_75_1483 ();
 sg13g2_decap_8 FILLER_75_1495 ();
 sg13g2_decap_8 FILLER_75_1502 ();
 sg13g2_fill_1 FILLER_75_1545 ();
 sg13g2_fill_2 FILLER_75_1550 ();
 sg13g2_fill_1 FILLER_75_1552 ();
 sg13g2_fill_2 FILLER_75_1563 ();
 sg13g2_fill_1 FILLER_75_1565 ();
 sg13g2_decap_8 FILLER_75_1605 ();
 sg13g2_fill_1 FILLER_75_1612 ();
 sg13g2_decap_4 FILLER_75_1617 ();
 sg13g2_decap_8 FILLER_75_1625 ();
 sg13g2_decap_4 FILLER_75_1632 ();
 sg13g2_decap_8 FILLER_75_1646 ();
 sg13g2_decap_8 FILLER_75_1653 ();
 sg13g2_decap_4 FILLER_75_1660 ();
 sg13g2_decap_8 FILLER_75_1681 ();
 sg13g2_decap_8 FILLER_75_1688 ();
 sg13g2_decap_4 FILLER_75_1695 ();
 sg13g2_fill_2 FILLER_75_1699 ();
 sg13g2_fill_1 FILLER_75_1726 ();
 sg13g2_fill_2 FILLER_75_1731 ();
 sg13g2_fill_1 FILLER_75_1742 ();
 sg13g2_fill_2 FILLER_75_1749 ();
 sg13g2_fill_2 FILLER_75_1766 ();
 sg13g2_decap_8 FILLER_75_1778 ();
 sg13g2_fill_2 FILLER_75_1785 ();
 sg13g2_fill_2 FILLER_75_1797 ();
 sg13g2_fill_1 FILLER_75_1799 ();
 sg13g2_fill_2 FILLER_75_1827 ();
 sg13g2_fill_1 FILLER_75_1837 ();
 sg13g2_fill_2 FILLER_75_1843 ();
 sg13g2_fill_1 FILLER_75_1849 ();
 sg13g2_fill_1 FILLER_75_1858 ();
 sg13g2_fill_1 FILLER_75_1871 ();
 sg13g2_fill_1 FILLER_75_1877 ();
 sg13g2_fill_1 FILLER_75_1882 ();
 sg13g2_fill_1 FILLER_75_1887 ();
 sg13g2_decap_8 FILLER_75_1899 ();
 sg13g2_fill_2 FILLER_75_1918 ();
 sg13g2_fill_1 FILLER_75_1920 ();
 sg13g2_fill_1 FILLER_75_1925 ();
 sg13g2_fill_1 FILLER_75_1931 ();
 sg13g2_fill_1 FILLER_75_1941 ();
 sg13g2_decap_8 FILLER_75_1954 ();
 sg13g2_decap_8 FILLER_75_1961 ();
 sg13g2_decap_4 FILLER_75_1968 ();
 sg13g2_fill_1 FILLER_75_1972 ();
 sg13g2_decap_4 FILLER_75_2003 ();
 sg13g2_fill_1 FILLER_75_2007 ();
 sg13g2_fill_1 FILLER_75_2016 ();
 sg13g2_fill_1 FILLER_75_2022 ();
 sg13g2_fill_1 FILLER_75_2027 ();
 sg13g2_fill_1 FILLER_75_2036 ();
 sg13g2_fill_1 FILLER_75_2044 ();
 sg13g2_fill_2 FILLER_75_2052 ();
 sg13g2_fill_1 FILLER_75_2080 ();
 sg13g2_fill_1 FILLER_75_2100 ();
 sg13g2_fill_1 FILLER_75_2111 ();
 sg13g2_fill_1 FILLER_75_2117 ();
 sg13g2_fill_1 FILLER_75_2122 ();
 sg13g2_decap_8 FILLER_75_2138 ();
 sg13g2_decap_8 FILLER_75_2145 ();
 sg13g2_decap_8 FILLER_75_2152 ();
 sg13g2_decap_8 FILLER_75_2159 ();
 sg13g2_fill_1 FILLER_75_2166 ();
 sg13g2_fill_2 FILLER_75_2171 ();
 sg13g2_fill_1 FILLER_75_2173 ();
 sg13g2_fill_1 FILLER_75_2198 ();
 sg13g2_fill_1 FILLER_75_2220 ();
 sg13g2_fill_2 FILLER_75_2226 ();
 sg13g2_fill_1 FILLER_75_2228 ();
 sg13g2_fill_1 FILLER_75_2247 ();
 sg13g2_fill_2 FILLER_75_2269 ();
 sg13g2_decap_8 FILLER_75_2309 ();
 sg13g2_fill_1 FILLER_75_2316 ();
 sg13g2_decap_8 FILLER_75_2323 ();
 sg13g2_decap_4 FILLER_75_2330 ();
 sg13g2_decap_8 FILLER_75_2368 ();
 sg13g2_decap_4 FILLER_75_2375 ();
 sg13g2_fill_1 FILLER_75_2379 ();
 sg13g2_fill_1 FILLER_75_2386 ();
 sg13g2_fill_2 FILLER_75_2402 ();
 sg13g2_fill_1 FILLER_75_2404 ();
 sg13g2_decap_4 FILLER_75_2411 ();
 sg13g2_decap_4 FILLER_75_2432 ();
 sg13g2_fill_2 FILLER_75_2445 ();
 sg13g2_fill_2 FILLER_75_2453 ();
 sg13g2_fill_2 FILLER_75_2468 ();
 sg13g2_fill_1 FILLER_75_2477 ();
 sg13g2_decap_4 FILLER_75_2485 ();
 sg13g2_fill_1 FILLER_75_2495 ();
 sg13g2_fill_2 FILLER_75_2527 ();
 sg13g2_fill_1 FILLER_75_2538 ();
 sg13g2_fill_1 FILLER_75_2553 ();
 sg13g2_fill_1 FILLER_75_2584 ();
 sg13g2_decap_8 FILLER_75_2590 ();
 sg13g2_decap_8 FILLER_75_2597 ();
 sg13g2_decap_8 FILLER_75_2604 ();
 sg13g2_decap_8 FILLER_75_2611 ();
 sg13g2_decap_8 FILLER_75_2618 ();
 sg13g2_decap_8 FILLER_75_2625 ();
 sg13g2_decap_8 FILLER_75_2632 ();
 sg13g2_decap_8 FILLER_75_2639 ();
 sg13g2_decap_8 FILLER_75_2646 ();
 sg13g2_decap_8 FILLER_75_2653 ();
 sg13g2_decap_8 FILLER_75_2660 ();
 sg13g2_fill_2 FILLER_75_2667 ();
 sg13g2_fill_1 FILLER_75_2669 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_fill_2 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_13 ();
 sg13g2_fill_2 FILLER_76_20 ();
 sg13g2_fill_1 FILLER_76_22 ();
 sg13g2_decap_4 FILLER_76_28 ();
 sg13g2_fill_1 FILLER_76_32 ();
 sg13g2_decap_4 FILLER_76_43 ();
 sg13g2_fill_2 FILLER_76_57 ();
 sg13g2_fill_1 FILLER_76_59 ();
 sg13g2_fill_2 FILLER_76_121 ();
 sg13g2_fill_2 FILLER_76_144 ();
 sg13g2_fill_2 FILLER_76_176 ();
 sg13g2_fill_2 FILLER_76_184 ();
 sg13g2_fill_2 FILLER_76_200 ();
 sg13g2_fill_2 FILLER_76_235 ();
 sg13g2_decap_4 FILLER_76_255 ();
 sg13g2_fill_2 FILLER_76_259 ();
 sg13g2_decap_4 FILLER_76_279 ();
 sg13g2_fill_1 FILLER_76_283 ();
 sg13g2_decap_8 FILLER_76_287 ();
 sg13g2_fill_1 FILLER_76_294 ();
 sg13g2_decap_8 FILLER_76_317 ();
 sg13g2_decap_8 FILLER_76_324 ();
 sg13g2_fill_1 FILLER_76_331 ();
 sg13g2_fill_1 FILLER_76_353 ();
 sg13g2_decap_8 FILLER_76_384 ();
 sg13g2_fill_1 FILLER_76_422 ();
 sg13g2_fill_2 FILLER_76_488 ();
 sg13g2_decap_8 FILLER_76_495 ();
 sg13g2_decap_4 FILLER_76_502 ();
 sg13g2_fill_1 FILLER_76_533 ();
 sg13g2_fill_1 FILLER_76_545 ();
 sg13g2_fill_1 FILLER_76_560 ();
 sg13g2_decap_8 FILLER_76_567 ();
 sg13g2_decap_4 FILLER_76_574 ();
 sg13g2_decap_4 FILLER_76_582 ();
 sg13g2_fill_1 FILLER_76_586 ();
 sg13g2_decap_4 FILLER_76_597 ();
 sg13g2_fill_1 FILLER_76_601 ();
 sg13g2_decap_4 FILLER_76_608 ();
 sg13g2_fill_1 FILLER_76_612 ();
 sg13g2_decap_4 FILLER_76_624 ();
 sg13g2_fill_2 FILLER_76_673 ();
 sg13g2_fill_1 FILLER_76_675 ();
 sg13g2_decap_8 FILLER_76_716 ();
 sg13g2_fill_2 FILLER_76_723 ();
 sg13g2_fill_1 FILLER_76_760 ();
 sg13g2_fill_2 FILLER_76_771 ();
 sg13g2_fill_1 FILLER_76_788 ();
 sg13g2_decap_4 FILLER_76_803 ();
 sg13g2_fill_2 FILLER_76_871 ();
 sg13g2_fill_1 FILLER_76_873 ();
 sg13g2_fill_1 FILLER_76_906 ();
 sg13g2_decap_8 FILLER_76_912 ();
 sg13g2_decap_8 FILLER_76_945 ();
 sg13g2_fill_2 FILLER_76_952 ();
 sg13g2_decap_4 FILLER_76_983 ();
 sg13g2_fill_2 FILLER_76_987 ();
 sg13g2_fill_2 FILLER_76_1034 ();
 sg13g2_fill_1 FILLER_76_1036 ();
 sg13g2_fill_2 FILLER_76_1053 ();
 sg13g2_decap_8 FILLER_76_1091 ();
 sg13g2_decap_8 FILLER_76_1098 ();
 sg13g2_fill_2 FILLER_76_1105 ();
 sg13g2_decap_4 FILLER_76_1111 ();
 sg13g2_fill_2 FILLER_76_1115 ();
 sg13g2_fill_1 FILLER_76_1164 ();
 sg13g2_fill_2 FILLER_76_1228 ();
 sg13g2_fill_2 FILLER_76_1244 ();
 sg13g2_fill_1 FILLER_76_1246 ();
 sg13g2_fill_2 FILLER_76_1257 ();
 sg13g2_fill_2 FILLER_76_1282 ();
 sg13g2_decap_8 FILLER_76_1328 ();
 sg13g2_decap_8 FILLER_76_1335 ();
 sg13g2_fill_1 FILLER_76_1342 ();
 sg13g2_fill_2 FILLER_76_1374 ();
 sg13g2_fill_1 FILLER_76_1383 ();
 sg13g2_decap_8 FILLER_76_1397 ();
 sg13g2_decap_8 FILLER_76_1404 ();
 sg13g2_fill_1 FILLER_76_1411 ();
 sg13g2_fill_2 FILLER_76_1422 ();
 sg13g2_fill_1 FILLER_76_1424 ();
 sg13g2_decap_8 FILLER_76_1443 ();
 sg13g2_decap_4 FILLER_76_1450 ();
 sg13g2_fill_1 FILLER_76_1454 ();
 sg13g2_decap_4 FILLER_76_1485 ();
 sg13g2_decap_8 FILLER_76_1502 ();
 sg13g2_fill_1 FILLER_76_1509 ();
 sg13g2_decap_8 FILLER_76_1514 ();
 sg13g2_fill_2 FILLER_76_1525 ();
 sg13g2_fill_1 FILLER_76_1527 ();
 sg13g2_fill_2 FILLER_76_1542 ();
 sg13g2_fill_1 FILLER_76_1544 ();
 sg13g2_decap_8 FILLER_76_1583 ();
 sg13g2_decap_8 FILLER_76_1590 ();
 sg13g2_decap_8 FILLER_76_1597 ();
 sg13g2_decap_8 FILLER_76_1604 ();
 sg13g2_fill_2 FILLER_76_1611 ();
 sg13g2_fill_1 FILLER_76_1613 ();
 sg13g2_decap_4 FILLER_76_1644 ();
 sg13g2_fill_1 FILLER_76_1648 ();
 sg13g2_fill_1 FILLER_76_1657 ();
 sg13g2_fill_2 FILLER_76_1689 ();
 sg13g2_fill_1 FILLER_76_1691 ();
 sg13g2_fill_2 FILLER_76_1701 ();
 sg13g2_fill_1 FILLER_76_1703 ();
 sg13g2_fill_1 FILLER_76_1709 ();
 sg13g2_fill_1 FILLER_76_1717 ();
 sg13g2_fill_2 FILLER_76_1734 ();
 sg13g2_fill_1 FILLER_76_1763 ();
 sg13g2_fill_2 FILLER_76_1772 ();
 sg13g2_fill_1 FILLER_76_1774 ();
 sg13g2_fill_1 FILLER_76_1780 ();
 sg13g2_fill_2 FILLER_76_1824 ();
 sg13g2_fill_1 FILLER_76_1826 ();
 sg13g2_fill_1 FILLER_76_1835 ();
 sg13g2_fill_1 FILLER_76_1840 ();
 sg13g2_fill_2 FILLER_76_1855 ();
 sg13g2_fill_1 FILLER_76_1857 ();
 sg13g2_fill_1 FILLER_76_1883 ();
 sg13g2_fill_2 FILLER_76_1894 ();
 sg13g2_fill_1 FILLER_76_1896 ();
 sg13g2_fill_1 FILLER_76_1920 ();
 sg13g2_fill_1 FILLER_76_1940 ();
 sg13g2_decap_8 FILLER_76_1953 ();
 sg13g2_decap_8 FILLER_76_1960 ();
 sg13g2_decap_8 FILLER_76_1967 ();
 sg13g2_fill_2 FILLER_76_1974 ();
 sg13g2_decap_4 FILLER_76_1982 ();
 sg13g2_fill_2 FILLER_76_1999 ();
 sg13g2_fill_1 FILLER_76_2006 ();
 sg13g2_fill_1 FILLER_76_2035 ();
 sg13g2_fill_1 FILLER_76_2043 ();
 sg13g2_fill_1 FILLER_76_2049 ();
 sg13g2_decap_8 FILLER_76_2078 ();
 sg13g2_fill_2 FILLER_76_2085 ();
 sg13g2_fill_2 FILLER_76_2096 ();
 sg13g2_fill_2 FILLER_76_2107 ();
 sg13g2_fill_1 FILLER_76_2109 ();
 sg13g2_decap_4 FILLER_76_2114 ();
 sg13g2_fill_1 FILLER_76_2118 ();
 sg13g2_decap_4 FILLER_76_2128 ();
 sg13g2_decap_4 FILLER_76_2136 ();
 sg13g2_fill_1 FILLER_76_2140 ();
 sg13g2_fill_2 FILLER_76_2172 ();
 sg13g2_fill_1 FILLER_76_2174 ();
 sg13g2_decap_4 FILLER_76_2188 ();
 sg13g2_decap_8 FILLER_76_2222 ();
 sg13g2_decap_8 FILLER_76_2229 ();
 sg13g2_fill_1 FILLER_76_2236 ();
 sg13g2_fill_2 FILLER_76_2244 ();
 sg13g2_fill_1 FILLER_76_2289 ();
 sg13g2_fill_1 FILLER_76_2303 ();
 sg13g2_fill_2 FILLER_76_2373 ();
 sg13g2_fill_1 FILLER_76_2375 ();
 sg13g2_fill_2 FILLER_76_2408 ();
 sg13g2_fill_2 FILLER_76_2427 ();
 sg13g2_fill_1 FILLER_76_2429 ();
 sg13g2_decap_4 FILLER_76_2440 ();
 sg13g2_decap_8 FILLER_76_2475 ();
 sg13g2_fill_1 FILLER_76_2482 ();
 sg13g2_fill_1 FILLER_76_2492 ();
 sg13g2_fill_2 FILLER_76_2507 ();
 sg13g2_fill_2 FILLER_76_2543 ();
 sg13g2_fill_2 FILLER_76_2564 ();
 sg13g2_decap_8 FILLER_76_2586 ();
 sg13g2_fill_2 FILLER_76_2593 ();
 sg13g2_decap_8 FILLER_76_2603 ();
 sg13g2_decap_8 FILLER_76_2610 ();
 sg13g2_decap_8 FILLER_76_2617 ();
 sg13g2_decap_8 FILLER_76_2624 ();
 sg13g2_decap_8 FILLER_76_2631 ();
 sg13g2_decap_8 FILLER_76_2638 ();
 sg13g2_decap_8 FILLER_76_2645 ();
 sg13g2_decap_8 FILLER_76_2652 ();
 sg13g2_decap_8 FILLER_76_2659 ();
 sg13g2_decap_4 FILLER_76_2666 ();
 sg13g2_decap_4 FILLER_77_0 ();
 sg13g2_fill_1 FILLER_77_4 ();
 sg13g2_fill_2 FILLER_77_90 ();
 sg13g2_fill_1 FILLER_77_123 ();
 sg13g2_fill_1 FILLER_77_150 ();
 sg13g2_decap_8 FILLER_77_243 ();
 sg13g2_decap_8 FILLER_77_250 ();
 sg13g2_decap_8 FILLER_77_257 ();
 sg13g2_fill_1 FILLER_77_279 ();
 sg13g2_fill_2 FILLER_77_310 ();
 sg13g2_fill_2 FILLER_77_322 ();
 sg13g2_fill_1 FILLER_77_324 ();
 sg13g2_decap_4 FILLER_77_330 ();
 sg13g2_fill_2 FILLER_77_334 ();
 sg13g2_fill_2 FILLER_77_346 ();
 sg13g2_fill_1 FILLER_77_348 ();
 sg13g2_decap_4 FILLER_77_369 ();
 sg13g2_fill_1 FILLER_77_373 ();
 sg13g2_fill_2 FILLER_77_379 ();
 sg13g2_decap_8 FILLER_77_385 ();
 sg13g2_decap_8 FILLER_77_392 ();
 sg13g2_decap_4 FILLER_77_399 ();
 sg13g2_fill_2 FILLER_77_403 ();
 sg13g2_fill_1 FILLER_77_409 ();
 sg13g2_fill_1 FILLER_77_414 ();
 sg13g2_fill_2 FILLER_77_474 ();
 sg13g2_fill_1 FILLER_77_483 ();
 sg13g2_decap_8 FILLER_77_495 ();
 sg13g2_decap_4 FILLER_77_502 ();
 sg13g2_fill_2 FILLER_77_506 ();
 sg13g2_fill_1 FILLER_77_516 ();
 sg13g2_fill_1 FILLER_77_551 ();
 sg13g2_fill_1 FILLER_77_561 ();
 sg13g2_fill_2 FILLER_77_611 ();
 sg13g2_decap_4 FILLER_77_629 ();
 sg13g2_fill_2 FILLER_77_659 ();
 sg13g2_fill_1 FILLER_77_661 ();
 sg13g2_fill_1 FILLER_77_665 ();
 sg13g2_decap_8 FILLER_77_671 ();
 sg13g2_decap_8 FILLER_77_678 ();
 sg13g2_fill_2 FILLER_77_685 ();
 sg13g2_decap_4 FILLER_77_753 ();
 sg13g2_fill_1 FILLER_77_757 ();
 sg13g2_fill_1 FILLER_77_790 ();
 sg13g2_decap_4 FILLER_77_801 ();
 sg13g2_decap_4 FILLER_77_826 ();
 sg13g2_fill_1 FILLER_77_830 ();
 sg13g2_fill_1 FILLER_77_883 ();
 sg13g2_fill_1 FILLER_77_888 ();
 sg13g2_fill_2 FILLER_77_893 ();
 sg13g2_decap_4 FILLER_77_905 ();
 sg13g2_fill_1 FILLER_77_909 ();
 sg13g2_fill_1 FILLER_77_918 ();
 sg13g2_decap_4 FILLER_77_929 ();
 sg13g2_fill_2 FILLER_77_933 ();
 sg13g2_fill_1 FILLER_77_955 ();
 sg13g2_fill_1 FILLER_77_960 ();
 sg13g2_fill_1 FILLER_77_987 ();
 sg13g2_fill_1 FILLER_77_1014 ();
 sg13g2_fill_2 FILLER_77_1025 ();
 sg13g2_decap_8 FILLER_77_1063 ();
 sg13g2_fill_2 FILLER_77_1070 ();
 sg13g2_fill_1 FILLER_77_1072 ();
 sg13g2_decap_8 FILLER_77_1097 ();
 sg13g2_decap_4 FILLER_77_1104 ();
 sg13g2_decap_4 FILLER_77_1118 ();
 sg13g2_fill_2 FILLER_77_1122 ();
 sg13g2_decap_4 FILLER_77_1134 ();
 sg13g2_fill_2 FILLER_77_1138 ();
 sg13g2_decap_8 FILLER_77_1148 ();
 sg13g2_decap_8 FILLER_77_1155 ();
 sg13g2_decap_4 FILLER_77_1162 ();
 sg13g2_fill_1 FILLER_77_1166 ();
 sg13g2_fill_2 FILLER_77_1181 ();
 sg13g2_fill_2 FILLER_77_1193 ();
 sg13g2_decap_8 FILLER_77_1205 ();
 sg13g2_decap_8 FILLER_77_1286 ();
 sg13g2_decap_8 FILLER_77_1303 ();
 sg13g2_fill_1 FILLER_77_1314 ();
 sg13g2_decap_8 FILLER_77_1319 ();
 sg13g2_decap_8 FILLER_77_1326 ();
 sg13g2_fill_1 FILLER_77_1369 ();
 sg13g2_decap_4 FILLER_77_1406 ();
 sg13g2_fill_2 FILLER_77_1410 ();
 sg13g2_decap_4 FILLER_77_1448 ();
 sg13g2_fill_1 FILLER_77_1452 ();
 sg13g2_decap_8 FILLER_77_1458 ();
 sg13g2_decap_4 FILLER_77_1489 ();
 sg13g2_fill_1 FILLER_77_1493 ();
 sg13g2_fill_2 FILLER_77_1530 ();
 sg13g2_fill_1 FILLER_77_1532 ();
 sg13g2_fill_2 FILLER_77_1543 ();
 sg13g2_fill_1 FILLER_77_1545 ();
 sg13g2_decap_8 FILLER_77_1572 ();
 sg13g2_fill_2 FILLER_77_1579 ();
 sg13g2_fill_1 FILLER_77_1581 ();
 sg13g2_fill_1 FILLER_77_1592 ();
 sg13g2_decap_4 FILLER_77_1597 ();
 sg13g2_fill_1 FILLER_77_1601 ();
 sg13g2_fill_1 FILLER_77_1727 ();
 sg13g2_fill_1 FILLER_77_1738 ();
 sg13g2_fill_1 FILLER_77_1771 ();
 sg13g2_fill_1 FILLER_77_1777 ();
 sg13g2_fill_1 FILLER_77_1801 ();
 sg13g2_fill_2 FILLER_77_1835 ();
 sg13g2_fill_2 FILLER_77_1845 ();
 sg13g2_fill_1 FILLER_77_1869 ();
 sg13g2_fill_1 FILLER_77_1874 ();
 sg13g2_fill_1 FILLER_77_1880 ();
 sg13g2_fill_1 FILLER_77_1891 ();
 sg13g2_decap_4 FILLER_77_1897 ();
 sg13g2_fill_1 FILLER_77_1909 ();
 sg13g2_fill_2 FILLER_77_1913 ();
 sg13g2_fill_1 FILLER_77_1920 ();
 sg13g2_fill_1 FILLER_77_1926 ();
 sg13g2_fill_2 FILLER_77_1931 ();
 sg13g2_fill_2 FILLER_77_1939 ();
 sg13g2_fill_1 FILLER_77_1946 ();
 sg13g2_fill_2 FILLER_77_2009 ();
 sg13g2_fill_1 FILLER_77_2015 ();
 sg13g2_fill_1 FILLER_77_2020 ();
 sg13g2_fill_2 FILLER_77_2031 ();
 sg13g2_fill_1 FILLER_77_2059 ();
 sg13g2_decap_4 FILLER_77_2074 ();
 sg13g2_decap_8 FILLER_77_2086 ();
 sg13g2_decap_4 FILLER_77_2093 ();
 sg13g2_fill_1 FILLER_77_2102 ();
 sg13g2_fill_1 FILLER_77_2108 ();
 sg13g2_decap_4 FILLER_77_2122 ();
 sg13g2_fill_2 FILLER_77_2126 ();
 sg13g2_decap_8 FILLER_77_2138 ();
 sg13g2_fill_2 FILLER_77_2145 ();
 sg13g2_fill_1 FILLER_77_2147 ();
 sg13g2_fill_1 FILLER_77_2184 ();
 sg13g2_decap_4 FILLER_77_2237 ();
 sg13g2_fill_2 FILLER_77_2246 ();
 sg13g2_fill_1 FILLER_77_2314 ();
 sg13g2_fill_1 FILLER_77_2319 ();
 sg13g2_fill_1 FILLER_77_2330 ();
 sg13g2_fill_2 FILLER_77_2336 ();
 sg13g2_fill_2 FILLER_77_2342 ();
 sg13g2_fill_2 FILLER_77_2348 ();
 sg13g2_fill_1 FILLER_77_2350 ();
 sg13g2_fill_1 FILLER_77_2387 ();
 sg13g2_fill_1 FILLER_77_2433 ();
 sg13g2_fill_2 FILLER_77_2439 ();
 sg13g2_fill_1 FILLER_77_2441 ();
 sg13g2_fill_1 FILLER_77_2446 ();
 sg13g2_decap_4 FILLER_77_2476 ();
 sg13g2_fill_2 FILLER_77_2480 ();
 sg13g2_decap_8 FILLER_77_2589 ();
 sg13g2_decap_8 FILLER_77_2596 ();
 sg13g2_decap_8 FILLER_77_2603 ();
 sg13g2_decap_8 FILLER_77_2610 ();
 sg13g2_decap_8 FILLER_77_2617 ();
 sg13g2_decap_8 FILLER_77_2624 ();
 sg13g2_decap_8 FILLER_77_2631 ();
 sg13g2_decap_8 FILLER_77_2638 ();
 sg13g2_decap_8 FILLER_77_2645 ();
 sg13g2_decap_8 FILLER_77_2652 ();
 sg13g2_decap_8 FILLER_77_2659 ();
 sg13g2_decap_4 FILLER_77_2666 ();
 sg13g2_fill_2 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_2 ();
 sg13g2_fill_2 FILLER_78_39 ();
 sg13g2_fill_2 FILLER_78_72 ();
 sg13g2_fill_1 FILLER_78_74 ();
 sg13g2_fill_1 FILLER_78_85 ();
 sg13g2_fill_2 FILLER_78_114 ();
 sg13g2_decap_4 FILLER_78_121 ();
 sg13g2_fill_1 FILLER_78_125 ();
 sg13g2_fill_1 FILLER_78_179 ();
 sg13g2_fill_1 FILLER_78_230 ();
 sg13g2_decap_8 FILLER_78_299 ();
 sg13g2_fill_1 FILLER_78_327 ();
 sg13g2_fill_2 FILLER_78_333 ();
 sg13g2_fill_2 FILLER_78_356 ();
 sg13g2_decap_4 FILLER_78_384 ();
 sg13g2_decap_8 FILLER_78_393 ();
 sg13g2_fill_2 FILLER_78_400 ();
 sg13g2_fill_1 FILLER_78_402 ();
 sg13g2_fill_1 FILLER_78_456 ();
 sg13g2_fill_2 FILLER_78_462 ();
 sg13g2_fill_1 FILLER_78_464 ();
 sg13g2_fill_2 FILLER_78_482 ();
 sg13g2_fill_2 FILLER_78_489 ();
 sg13g2_fill_2 FILLER_78_517 ();
 sg13g2_fill_2 FILLER_78_528 ();
 sg13g2_fill_2 FILLER_78_575 ();
 sg13g2_fill_2 FILLER_78_603 ();
 sg13g2_fill_2 FILLER_78_667 ();
 sg13g2_fill_1 FILLER_78_669 ();
 sg13g2_fill_1 FILLER_78_712 ();
 sg13g2_fill_2 FILLER_78_717 ();
 sg13g2_decap_8 FILLER_78_755 ();
 sg13g2_decap_4 FILLER_78_762 ();
 sg13g2_decap_4 FILLER_78_807 ();
 sg13g2_fill_1 FILLER_78_811 ();
 sg13g2_fill_2 FILLER_78_816 ();
 sg13g2_decap_4 FILLER_78_891 ();
 sg13g2_fill_1 FILLER_78_895 ();
 sg13g2_fill_1 FILLER_78_912 ();
 sg13g2_fill_1 FILLER_78_923 ();
 sg13g2_fill_1 FILLER_78_976 ();
 sg13g2_fill_1 FILLER_78_1042 ();
 sg13g2_decap_4 FILLER_78_1069 ();
 sg13g2_fill_1 FILLER_78_1099 ();
 sg13g2_fill_2 FILLER_78_1120 ();
 sg13g2_fill_1 FILLER_78_1122 ();
 sg13g2_fill_2 FILLER_78_1133 ();
 sg13g2_decap_4 FILLER_78_1161 ();
 sg13g2_fill_1 FILLER_78_1165 ();
 sg13g2_decap_4 FILLER_78_1189 ();
 sg13g2_fill_1 FILLER_78_1253 ();
 sg13g2_fill_1 FILLER_78_1264 ();
 sg13g2_fill_1 FILLER_78_1317 ();
 sg13g2_decap_8 FILLER_78_1328 ();
 sg13g2_decap_4 FILLER_78_1335 ();
 sg13g2_fill_1 FILLER_78_1339 ();
 sg13g2_decap_4 FILLER_78_1344 ();
 sg13g2_decap_4 FILLER_78_1352 ();
 sg13g2_fill_1 FILLER_78_1356 ();
 sg13g2_decap_4 FILLER_78_1409 ();
 sg13g2_decap_4 FILLER_78_1465 ();
 sg13g2_fill_1 FILLER_78_1499 ();
 sg13g2_fill_1 FILLER_78_1549 ();
 sg13g2_decap_4 FILLER_78_1576 ();
 sg13g2_fill_2 FILLER_78_1590 ();
 sg13g2_decap_8 FILLER_78_1626 ();
 sg13g2_decap_4 FILLER_78_1650 ();
 sg13g2_fill_2 FILLER_78_1654 ();
 sg13g2_decap_4 FILLER_78_1691 ();
 sg13g2_fill_2 FILLER_78_1704 ();
 sg13g2_fill_2 FILLER_78_1711 ();
 sg13g2_fill_1 FILLER_78_1713 ();
 sg13g2_decap_8 FILLER_78_1719 ();
 sg13g2_decap_8 FILLER_78_1773 ();
 sg13g2_fill_2 FILLER_78_1780 ();
 sg13g2_fill_1 FILLER_78_1789 ();
 sg13g2_fill_1 FILLER_78_1799 ();
 sg13g2_fill_1 FILLER_78_1812 ();
 sg13g2_fill_1 FILLER_78_1821 ();
 sg13g2_fill_2 FILLER_78_1843 ();
 sg13g2_fill_1 FILLER_78_1845 ();
 sg13g2_fill_1 FILLER_78_1851 ();
 sg13g2_decap_4 FILLER_78_1862 ();
 sg13g2_fill_2 FILLER_78_1899 ();
 sg13g2_fill_2 FILLER_78_1911 ();
 sg13g2_fill_1 FILLER_78_1913 ();
 sg13g2_decap_4 FILLER_78_1971 ();
 sg13g2_decap_4 FILLER_78_1996 ();
 sg13g2_fill_2 FILLER_78_2000 ();
 sg13g2_decap_4 FILLER_78_2020 ();
 sg13g2_fill_2 FILLER_78_2064 ();
 sg13g2_fill_1 FILLER_78_2066 ();
 sg13g2_fill_2 FILLER_78_2080 ();
 sg13g2_fill_2 FILLER_78_2087 ();
 sg13g2_fill_1 FILLER_78_2089 ();
 sg13g2_fill_1 FILLER_78_2109 ();
 sg13g2_fill_1 FILLER_78_2115 ();
 sg13g2_decap_4 FILLER_78_2121 ();
 sg13g2_fill_2 FILLER_78_2161 ();
 sg13g2_fill_2 FILLER_78_2189 ();
 sg13g2_decap_4 FILLER_78_2195 ();
 sg13g2_fill_2 FILLER_78_2209 ();
 sg13g2_decap_8 FILLER_78_2225 ();
 sg13g2_fill_2 FILLER_78_2232 ();
 sg13g2_fill_1 FILLER_78_2234 ();
 sg13g2_fill_1 FILLER_78_2240 ();
 sg13g2_fill_1 FILLER_78_2267 ();
 sg13g2_fill_1 FILLER_78_2294 ();
 sg13g2_fill_2 FILLER_78_2300 ();
 sg13g2_fill_1 FILLER_78_2328 ();
 sg13g2_fill_1 FILLER_78_2334 ();
 sg13g2_fill_2 FILLER_78_2361 ();
 sg13g2_fill_1 FILLER_78_2363 ();
 sg13g2_fill_1 FILLER_78_2438 ();
 sg13g2_fill_1 FILLER_78_2446 ();
 sg13g2_decap_4 FILLER_78_2460 ();
 sg13g2_fill_1 FILLER_78_2464 ();
 sg13g2_decap_4 FILLER_78_2469 ();
 sg13g2_fill_1 FILLER_78_2582 ();
 sg13g2_decap_8 FILLER_78_2588 ();
 sg13g2_decap_8 FILLER_78_2595 ();
 sg13g2_decap_8 FILLER_78_2602 ();
 sg13g2_decap_8 FILLER_78_2609 ();
 sg13g2_decap_8 FILLER_78_2616 ();
 sg13g2_decap_8 FILLER_78_2623 ();
 sg13g2_decap_8 FILLER_78_2630 ();
 sg13g2_decap_8 FILLER_78_2637 ();
 sg13g2_decap_8 FILLER_78_2644 ();
 sg13g2_decap_8 FILLER_78_2651 ();
 sg13g2_decap_8 FILLER_78_2658 ();
 sg13g2_decap_4 FILLER_78_2665 ();
 sg13g2_fill_1 FILLER_78_2669 ();
 sg13g2_decap_4 FILLER_79_0 ();
 sg13g2_fill_1 FILLER_79_4 ();
 sg13g2_fill_2 FILLER_79_9 ();
 sg13g2_fill_1 FILLER_79_11 ();
 sg13g2_fill_1 FILLER_79_42 ();
 sg13g2_fill_2 FILLER_79_47 ();
 sg13g2_fill_1 FILLER_79_75 ();
 sg13g2_fill_2 FILLER_79_102 ();
 sg13g2_fill_2 FILLER_79_109 ();
 sg13g2_fill_1 FILLER_79_111 ();
 sg13g2_fill_2 FILLER_79_116 ();
 sg13g2_fill_1 FILLER_79_118 ();
 sg13g2_fill_2 FILLER_79_124 ();
 sg13g2_fill_2 FILLER_79_136 ();
 sg13g2_fill_1 FILLER_79_154 ();
 sg13g2_fill_2 FILLER_79_184 ();
 sg13g2_fill_1 FILLER_79_212 ();
 sg13g2_decap_4 FILLER_79_247 ();
 sg13g2_fill_2 FILLER_79_281 ();
 sg13g2_fill_1 FILLER_79_283 ();
 sg13g2_fill_2 FILLER_79_289 ();
 sg13g2_fill_1 FILLER_79_291 ();
 sg13g2_decap_8 FILLER_79_328 ();
 sg13g2_decap_8 FILLER_79_335 ();
 sg13g2_fill_2 FILLER_79_342 ();
 sg13g2_fill_1 FILLER_79_344 ();
 sg13g2_decap_4 FILLER_79_358 ();
 sg13g2_fill_1 FILLER_79_362 ();
 sg13g2_fill_1 FILLER_79_372 ();
 sg13g2_decap_8 FILLER_79_399 ();
 sg13g2_fill_2 FILLER_79_489 ();
 sg13g2_fill_1 FILLER_79_525 ();
 sg13g2_fill_1 FILLER_79_552 ();
 sg13g2_fill_1 FILLER_79_579 ();
 sg13g2_fill_2 FILLER_79_584 ();
 sg13g2_decap_8 FILLER_79_638 ();
 sg13g2_decap_8 FILLER_79_645 ();
 sg13g2_decap_4 FILLER_79_652 ();
 sg13g2_fill_1 FILLER_79_656 ();
 sg13g2_decap_8 FILLER_79_661 ();
 sg13g2_decap_4 FILLER_79_668 ();
 sg13g2_fill_2 FILLER_79_672 ();
 sg13g2_decap_8 FILLER_79_704 ();
 sg13g2_decap_4 FILLER_79_711 ();
 sg13g2_fill_2 FILLER_79_782 ();
 sg13g2_fill_1 FILLER_79_784 ();
 sg13g2_fill_1 FILLER_79_837 ();
 sg13g2_fill_1 FILLER_79_868 ();
 sg13g2_decap_8 FILLER_79_905 ();
 sg13g2_decap_4 FILLER_79_912 ();
 sg13g2_fill_1 FILLER_79_916 ();
 sg13g2_decap_4 FILLER_79_921 ();
 sg13g2_decap_4 FILLER_79_929 ();
 sg13g2_fill_2 FILLER_79_933 ();
 sg13g2_decap_4 FILLER_79_939 ();
 sg13g2_fill_2 FILLER_79_983 ();
 sg13g2_fill_1 FILLER_79_985 ();
 sg13g2_decap_8 FILLER_79_1000 ();
 sg13g2_fill_1 FILLER_79_1007 ();
 sg13g2_fill_2 FILLER_79_1012 ();
 sg13g2_fill_2 FILLER_79_1040 ();
 sg13g2_fill_1 FILLER_79_1042 ();
 sg13g2_fill_2 FILLER_79_1079 ();
 sg13g2_fill_1 FILLER_79_1081 ();
 sg13g2_decap_8 FILLER_79_1112 ();
 sg13g2_fill_2 FILLER_79_1119 ();
 sg13g2_fill_2 FILLER_79_1155 ();
 sg13g2_fill_1 FILLER_79_1213 ();
 sg13g2_decap_8 FILLER_79_1244 ();
 sg13g2_decap_8 FILLER_79_1251 ();
 sg13g2_decap_8 FILLER_79_1258 ();
 sg13g2_fill_2 FILLER_79_1282 ();
 sg13g2_fill_2 FILLER_79_1310 ();
 sg13g2_decap_8 FILLER_79_1338 ();
 sg13g2_decap_8 FILLER_79_1345 ();
 sg13g2_fill_1 FILLER_79_1352 ();
 sg13g2_fill_1 FILLER_79_1393 ();
 sg13g2_decap_8 FILLER_79_1454 ();
 sg13g2_fill_1 FILLER_79_1461 ();
 sg13g2_fill_2 FILLER_79_1508 ();
 sg13g2_fill_1 FILLER_79_1510 ();
 sg13g2_decap_4 FILLER_79_1523 ();
 sg13g2_decap_8 FILLER_79_1579 ();
 sg13g2_fill_2 FILLER_79_1586 ();
 sg13g2_decap_8 FILLER_79_1624 ();
 sg13g2_decap_8 FILLER_79_1631 ();
 sg13g2_decap_8 FILLER_79_1638 ();
 sg13g2_decap_8 FILLER_79_1645 ();
 sg13g2_decap_4 FILLER_79_1652 ();
 sg13g2_fill_1 FILLER_79_1656 ();
 sg13g2_decap_8 FILLER_79_1687 ();
 sg13g2_fill_2 FILLER_79_1760 ();
 sg13g2_fill_1 FILLER_79_1762 ();
 sg13g2_decap_8 FILLER_79_1780 ();
 sg13g2_fill_1 FILLER_79_1794 ();
 sg13g2_decap_8 FILLER_79_1799 ();
 sg13g2_fill_1 FILLER_79_1810 ();
 sg13g2_fill_1 FILLER_79_1816 ();
 sg13g2_fill_2 FILLER_79_1821 ();
 sg13g2_fill_1 FILLER_79_1828 ();
 sg13g2_fill_1 FILLER_79_1837 ();
 sg13g2_fill_2 FILLER_79_1851 ();
 sg13g2_decap_8 FILLER_79_1861 ();
 sg13g2_decap_8 FILLER_79_1868 ();
 sg13g2_fill_2 FILLER_79_1875 ();
 sg13g2_fill_1 FILLER_79_1877 ();
 sg13g2_fill_1 FILLER_79_1882 ();
 sg13g2_fill_2 FILLER_79_1887 ();
 sg13g2_fill_1 FILLER_79_1893 ();
 sg13g2_fill_2 FILLER_79_1898 ();
 sg13g2_fill_2 FILLER_79_1904 ();
 sg13g2_fill_2 FILLER_79_1910 ();
 sg13g2_fill_1 FILLER_79_1916 ();
 sg13g2_fill_1 FILLER_79_1921 ();
 sg13g2_fill_1 FILLER_79_1926 ();
 sg13g2_fill_1 FILLER_79_1932 ();
 sg13g2_fill_1 FILLER_79_1938 ();
 sg13g2_fill_1 FILLER_79_1944 ();
 sg13g2_decap_8 FILLER_79_1975 ();
 sg13g2_decap_8 FILLER_79_1982 ();
 sg13g2_decap_8 FILLER_79_1989 ();
 sg13g2_decap_8 FILLER_79_1996 ();
 sg13g2_decap_8 FILLER_79_2003 ();
 sg13g2_decap_8 FILLER_79_2010 ();
 sg13g2_decap_8 FILLER_79_2017 ();
 sg13g2_decap_8 FILLER_79_2024 ();
 sg13g2_fill_2 FILLER_79_2031 ();
 sg13g2_decap_8 FILLER_79_2036 ();
 sg13g2_fill_1 FILLER_79_2043 ();
 sg13g2_fill_2 FILLER_79_2062 ();
 sg13g2_decap_4 FILLER_79_2068 ();
 sg13g2_fill_2 FILLER_79_2072 ();
 sg13g2_decap_4 FILLER_79_2079 ();
 sg13g2_fill_2 FILLER_79_2083 ();
 sg13g2_decap_4 FILLER_79_2093 ();
 sg13g2_decap_8 FILLER_79_2101 ();
 sg13g2_decap_8 FILLER_79_2108 ();
 sg13g2_decap_8 FILLER_79_2115 ();
 sg13g2_decap_8 FILLER_79_2122 ();
 sg13g2_fill_1 FILLER_79_2159 ();
 sg13g2_fill_1 FILLER_79_2170 ();
 sg13g2_fill_1 FILLER_79_2175 ();
 sg13g2_fill_1 FILLER_79_2202 ();
 sg13g2_fill_1 FILLER_79_2229 ();
 sg13g2_fill_2 FILLER_79_2264 ();
 sg13g2_fill_1 FILLER_79_2271 ();
 sg13g2_fill_1 FILLER_79_2332 ();
 sg13g2_decap_4 FILLER_79_2364 ();
 sg13g2_fill_2 FILLER_79_2372 ();
 sg13g2_decap_8 FILLER_79_2378 ();
 sg13g2_decap_8 FILLER_79_2385 ();
 sg13g2_decap_4 FILLER_79_2392 ();
 sg13g2_fill_2 FILLER_79_2396 ();
 sg13g2_fill_2 FILLER_79_2402 ();
 sg13g2_fill_1 FILLER_79_2404 ();
 sg13g2_decap_4 FILLER_79_2444 ();
 sg13g2_decap_8 FILLER_79_2474 ();
 sg13g2_fill_1 FILLER_79_2481 ();
 sg13g2_fill_1 FILLER_79_2517 ();
 sg13g2_fill_2 FILLER_79_2546 ();
 sg13g2_fill_2 FILLER_79_2552 ();
 sg13g2_decap_8 FILLER_79_2558 ();
 sg13g2_fill_2 FILLER_79_2565 ();
 sg13g2_fill_1 FILLER_79_2567 ();
 sg13g2_decap_8 FILLER_79_2572 ();
 sg13g2_decap_8 FILLER_79_2579 ();
 sg13g2_decap_8 FILLER_79_2586 ();
 sg13g2_decap_8 FILLER_79_2593 ();
 sg13g2_decap_8 FILLER_79_2600 ();
 sg13g2_decap_8 FILLER_79_2607 ();
 sg13g2_decap_8 FILLER_79_2614 ();
 sg13g2_decap_8 FILLER_79_2621 ();
 sg13g2_decap_8 FILLER_79_2628 ();
 sg13g2_decap_8 FILLER_79_2635 ();
 sg13g2_decap_8 FILLER_79_2642 ();
 sg13g2_decap_8 FILLER_79_2649 ();
 sg13g2_decap_8 FILLER_79_2656 ();
 sg13g2_decap_8 FILLER_79_2663 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_fill_1 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_12 ();
 sg13g2_decap_8 FILLER_80_23 ();
 sg13g2_decap_8 FILLER_80_30 ();
 sg13g2_decap_4 FILLER_80_47 ();
 sg13g2_fill_1 FILLER_80_51 ();
 sg13g2_decap_8 FILLER_80_73 ();
 sg13g2_fill_2 FILLER_80_84 ();
 sg13g2_fill_1 FILLER_80_86 ();
 sg13g2_fill_2 FILLER_80_91 ();
 sg13g2_decap_4 FILLER_80_97 ();
 sg13g2_fill_1 FILLER_80_105 ();
 sg13g2_fill_1 FILLER_80_124 ();
 sg13g2_fill_1 FILLER_80_129 ();
 sg13g2_fill_2 FILLER_80_134 ();
 sg13g2_fill_1 FILLER_80_164 ();
 sg13g2_fill_1 FILLER_80_192 ();
 sg13g2_fill_1 FILLER_80_201 ();
 sg13g2_fill_1 FILLER_80_213 ();
 sg13g2_fill_1 FILLER_80_247 ();
 sg13g2_fill_1 FILLER_80_252 ();
 sg13g2_decap_8 FILLER_80_265 ();
 sg13g2_decap_8 FILLER_80_272 ();
 sg13g2_fill_2 FILLER_80_283 ();
 sg13g2_fill_1 FILLER_80_290 ();
 sg13g2_fill_1 FILLER_80_295 ();
 sg13g2_fill_1 FILLER_80_311 ();
 sg13g2_decap_8 FILLER_80_316 ();
 sg13g2_decap_8 FILLER_80_323 ();
 sg13g2_fill_2 FILLER_80_330 ();
 sg13g2_fill_1 FILLER_80_332 ();
 sg13g2_fill_1 FILLER_80_338 ();
 sg13g2_fill_2 FILLER_80_344 ();
 sg13g2_decap_4 FILLER_80_369 ();
 sg13g2_fill_1 FILLER_80_373 ();
 sg13g2_fill_2 FILLER_80_379 ();
 sg13g2_fill_1 FILLER_80_381 ();
 sg13g2_decap_8 FILLER_80_386 ();
 sg13g2_decap_8 FILLER_80_393 ();
 sg13g2_decap_4 FILLER_80_400 ();
 sg13g2_fill_2 FILLER_80_404 ();
 sg13g2_decap_8 FILLER_80_418 ();
 sg13g2_fill_1 FILLER_80_425 ();
 sg13g2_fill_2 FILLER_80_430 ();
 sg13g2_decap_4 FILLER_80_436 ();
 sg13g2_decap_4 FILLER_80_448 ();
 sg13g2_decap_4 FILLER_80_456 ();
 sg13g2_fill_2 FILLER_80_460 ();
 sg13g2_decap_8 FILLER_80_466 ();
 sg13g2_decap_8 FILLER_80_473 ();
 sg13g2_decap_4 FILLER_80_480 ();
 sg13g2_fill_1 FILLER_80_510 ();
 sg13g2_decap_8 FILLER_80_515 ();
 sg13g2_decap_8 FILLER_80_522 ();
 sg13g2_fill_2 FILLER_80_529 ();
 sg13g2_fill_1 FILLER_80_531 ();
 sg13g2_decap_4 FILLER_80_543 ();
 sg13g2_fill_2 FILLER_80_547 ();
 sg13g2_decap_8 FILLER_80_553 ();
 sg13g2_fill_2 FILLER_80_560 ();
 sg13g2_decap_8 FILLER_80_566 ();
 sg13g2_decap_8 FILLER_80_573 ();
 sg13g2_decap_4 FILLER_80_580 ();
 sg13g2_fill_2 FILLER_80_584 ();
 sg13g2_decap_4 FILLER_80_590 ();
 sg13g2_fill_2 FILLER_80_598 ();
 sg13g2_fill_1 FILLER_80_600 ();
 sg13g2_decap_4 FILLER_80_614 ();
 sg13g2_fill_1 FILLER_80_618 ();
 sg13g2_decap_8 FILLER_80_627 ();
 sg13g2_decap_8 FILLER_80_634 ();
 sg13g2_decap_8 FILLER_80_644 ();
 sg13g2_fill_1 FILLER_80_655 ();
 sg13g2_decap_4 FILLER_80_682 ();
 sg13g2_decap_8 FILLER_80_690 ();
 sg13g2_decap_8 FILLER_80_697 ();
 sg13g2_decap_8 FILLER_80_704 ();
 sg13g2_decap_8 FILLER_80_711 ();
 sg13g2_decap_4 FILLER_80_718 ();
 sg13g2_fill_2 FILLER_80_756 ();
 sg13g2_fill_2 FILLER_80_762 ();
 sg13g2_fill_1 FILLER_80_764 ();
 sg13g2_decap_8 FILLER_80_769 ();
 sg13g2_decap_8 FILLER_80_776 ();
 sg13g2_decap_8 FILLER_80_783 ();
 sg13g2_fill_1 FILLER_80_790 ();
 sg13g2_decap_8 FILLER_80_795 ();
 sg13g2_fill_2 FILLER_80_802 ();
 sg13g2_decap_8 FILLER_80_809 ();
 sg13g2_fill_2 FILLER_80_816 ();
 sg13g2_decap_8 FILLER_80_822 ();
 sg13g2_decap_8 FILLER_80_829 ();
 sg13g2_decap_4 FILLER_80_836 ();
 sg13g2_fill_2 FILLER_80_840 ();
 sg13g2_fill_2 FILLER_80_850 ();
 sg13g2_decap_8 FILLER_80_858 ();
 sg13g2_decap_8 FILLER_80_865 ();
 sg13g2_fill_2 FILLER_80_872 ();
 sg13g2_fill_1 FILLER_80_874 ();
 sg13g2_fill_1 FILLER_80_883 ();
 sg13g2_decap_8 FILLER_80_936 ();
 sg13g2_decap_8 FILLER_80_943 ();
 sg13g2_decap_8 FILLER_80_950 ();
 sg13g2_decap_8 FILLER_80_957 ();
 sg13g2_fill_2 FILLER_80_964 ();
 sg13g2_decap_8 FILLER_80_970 ();
 sg13g2_decap_8 FILLER_80_977 ();
 sg13g2_decap_8 FILLER_80_984 ();
 sg13g2_decap_8 FILLER_80_991 ();
 sg13g2_decap_8 FILLER_80_998 ();
 sg13g2_decap_8 FILLER_80_1005 ();
 sg13g2_decap_4 FILLER_80_1012 ();
 sg13g2_fill_2 FILLER_80_1016 ();
 sg13g2_decap_8 FILLER_80_1022 ();
 sg13g2_decap_8 FILLER_80_1029 ();
 sg13g2_decap_8 FILLER_80_1036 ();
 sg13g2_decap_8 FILLER_80_1043 ();
 sg13g2_decap_4 FILLER_80_1054 ();
 sg13g2_fill_2 FILLER_80_1058 ();
 sg13g2_decap_8 FILLER_80_1064 ();
 sg13g2_decap_4 FILLER_80_1071 ();
 sg13g2_fill_1 FILLER_80_1075 ();
 sg13g2_decap_4 FILLER_80_1089 ();
 sg13g2_decap_8 FILLER_80_1097 ();
 sg13g2_decap_8 FILLER_80_1104 ();
 sg13g2_fill_2 FILLER_80_1111 ();
 sg13g2_fill_1 FILLER_80_1113 ();
 sg13g2_fill_2 FILLER_80_1140 ();
 sg13g2_decap_8 FILLER_80_1146 ();
 sg13g2_decap_8 FILLER_80_1153 ();
 sg13g2_decap_4 FILLER_80_1160 ();
 sg13g2_fill_2 FILLER_80_1164 ();
 sg13g2_decap_8 FILLER_80_1170 ();
 sg13g2_decap_8 FILLER_80_1177 ();
 sg13g2_decap_4 FILLER_80_1184 ();
 sg13g2_fill_2 FILLER_80_1188 ();
 sg13g2_decap_8 FILLER_80_1194 ();
 sg13g2_decap_8 FILLER_80_1201 ();
 sg13g2_decap_4 FILLER_80_1208 ();
 sg13g2_fill_1 FILLER_80_1212 ();
 sg13g2_fill_2 FILLER_80_1223 ();
 sg13g2_fill_1 FILLER_80_1225 ();
 sg13g2_fill_2 FILLER_80_1230 ();
 sg13g2_fill_1 FILLER_80_1232 ();
 sg13g2_decap_8 FILLER_80_1237 ();
 sg13g2_decap_8 FILLER_80_1244 ();
 sg13g2_fill_2 FILLER_80_1255 ();
 sg13g2_fill_2 FILLER_80_1295 ();
 sg13g2_fill_1 FILLER_80_1297 ();
 sg13g2_decap_4 FILLER_80_1302 ();
 sg13g2_fill_2 FILLER_80_1316 ();
 sg13g2_fill_1 FILLER_80_1318 ();
 sg13g2_decap_8 FILLER_80_1323 ();
 sg13g2_decap_8 FILLER_80_1330 ();
 sg13g2_decap_8 FILLER_80_1337 ();
 sg13g2_decap_8 FILLER_80_1344 ();
 sg13g2_decap_8 FILLER_80_1351 ();
 sg13g2_decap_8 FILLER_80_1358 ();
 sg13g2_decap_8 FILLER_80_1365 ();
 sg13g2_decap_4 FILLER_80_1372 ();
 sg13g2_fill_2 FILLER_80_1390 ();
 sg13g2_decap_8 FILLER_80_1396 ();
 sg13g2_decap_8 FILLER_80_1438 ();
 sg13g2_decap_8 FILLER_80_1445 ();
 sg13g2_decap_8 FILLER_80_1452 ();
 sg13g2_decap_8 FILLER_80_1459 ();
 sg13g2_fill_2 FILLER_80_1466 ();
 sg13g2_fill_1 FILLER_80_1468 ();
 sg13g2_decap_8 FILLER_80_1499 ();
 sg13g2_decap_8 FILLER_80_1506 ();
 sg13g2_decap_8 FILLER_80_1513 ();
 sg13g2_decap_8 FILLER_80_1520 ();
 sg13g2_decap_4 FILLER_80_1527 ();
 sg13g2_fill_2 FILLER_80_1531 ();
 sg13g2_fill_1 FILLER_80_1537 ();
 sg13g2_decap_8 FILLER_80_1570 ();
 sg13g2_decap_8 FILLER_80_1577 ();
 sg13g2_decap_8 FILLER_80_1584 ();
 sg13g2_decap_8 FILLER_80_1591 ();
 sg13g2_fill_1 FILLER_80_1598 ();
 sg13g2_decap_4 FILLER_80_1603 ();
 sg13g2_decap_8 FILLER_80_1615 ();
 sg13g2_decap_8 FILLER_80_1622 ();
 sg13g2_decap_8 FILLER_80_1629 ();
 sg13g2_decap_8 FILLER_80_1636 ();
 sg13g2_decap_8 FILLER_80_1643 ();
 sg13g2_decap_8 FILLER_80_1650 ();
 sg13g2_decap_4 FILLER_80_1657 ();
 sg13g2_fill_2 FILLER_80_1665 ();
 sg13g2_fill_1 FILLER_80_1667 ();
 sg13g2_decap_8 FILLER_80_1672 ();
 sg13g2_decap_8 FILLER_80_1679 ();
 sg13g2_decap_8 FILLER_80_1686 ();
 sg13g2_decap_8 FILLER_80_1693 ();
 sg13g2_decap_8 FILLER_80_1704 ();
 sg13g2_decap_8 FILLER_80_1711 ();
 sg13g2_decap_8 FILLER_80_1718 ();
 sg13g2_decap_4 FILLER_80_1725 ();
 sg13g2_decap_8 FILLER_80_1733 ();
 sg13g2_fill_2 FILLER_80_1740 ();
 sg13g2_fill_1 FILLER_80_1742 ();
 sg13g2_decap_8 FILLER_80_1747 ();
 sg13g2_decap_8 FILLER_80_1754 ();
 sg13g2_decap_8 FILLER_80_1761 ();
 sg13g2_decap_8 FILLER_80_1768 ();
 sg13g2_decap_8 FILLER_80_1775 ();
 sg13g2_decap_8 FILLER_80_1782 ();
 sg13g2_decap_8 FILLER_80_1789 ();
 sg13g2_decap_8 FILLER_80_1796 ();
 sg13g2_decap_8 FILLER_80_1803 ();
 sg13g2_decap_8 FILLER_80_1810 ();
 sg13g2_decap_4 FILLER_80_1817 ();
 sg13g2_fill_1 FILLER_80_1821 ();
 sg13g2_decap_4 FILLER_80_1826 ();
 sg13g2_decap_8 FILLER_80_1834 ();
 sg13g2_fill_1 FILLER_80_1841 ();
 sg13g2_decap_8 FILLER_80_1851 ();
 sg13g2_decap_8 FILLER_80_1858 ();
 sg13g2_decap_8 FILLER_80_1865 ();
 sg13g2_decap_8 FILLER_80_1872 ();
 sg13g2_decap_8 FILLER_80_1879 ();
 sg13g2_decap_8 FILLER_80_1886 ();
 sg13g2_decap_8 FILLER_80_1893 ();
 sg13g2_decap_8 FILLER_80_1900 ();
 sg13g2_decap_4 FILLER_80_1907 ();
 sg13g2_fill_1 FILLER_80_1911 ();
 sg13g2_decap_4 FILLER_80_1917 ();
 sg13g2_fill_2 FILLER_80_1921 ();
 sg13g2_fill_2 FILLER_80_1927 ();
 sg13g2_fill_1 FILLER_80_1929 ();
 sg13g2_decap_8 FILLER_80_1934 ();
 sg13g2_decap_8 FILLER_80_1941 ();
 sg13g2_decap_8 FILLER_80_1948 ();
 sg13g2_fill_2 FILLER_80_1955 ();
 sg13g2_fill_2 FILLER_80_1961 ();
 sg13g2_fill_1 FILLER_80_1963 ();
 sg13g2_decap_8 FILLER_80_1977 ();
 sg13g2_decap_8 FILLER_80_1984 ();
 sg13g2_decap_8 FILLER_80_1991 ();
 sg13g2_decap_8 FILLER_80_1998 ();
 sg13g2_decap_8 FILLER_80_2005 ();
 sg13g2_decap_8 FILLER_80_2012 ();
 sg13g2_decap_8 FILLER_80_2019 ();
 sg13g2_decap_8 FILLER_80_2026 ();
 sg13g2_decap_8 FILLER_80_2033 ();
 sg13g2_decap_8 FILLER_80_2040 ();
 sg13g2_decap_8 FILLER_80_2047 ();
 sg13g2_decap_8 FILLER_80_2054 ();
 sg13g2_decap_8 FILLER_80_2061 ();
 sg13g2_decap_8 FILLER_80_2068 ();
 sg13g2_decap_8 FILLER_80_2075 ();
 sg13g2_decap_8 FILLER_80_2082 ();
 sg13g2_decap_8 FILLER_80_2089 ();
 sg13g2_decap_8 FILLER_80_2096 ();
 sg13g2_decap_8 FILLER_80_2103 ();
 sg13g2_decap_8 FILLER_80_2110 ();
 sg13g2_decap_8 FILLER_80_2117 ();
 sg13g2_decap_8 FILLER_80_2124 ();
 sg13g2_decap_8 FILLER_80_2131 ();
 sg13g2_decap_8 FILLER_80_2146 ();
 sg13g2_decap_8 FILLER_80_2153 ();
 sg13g2_decap_8 FILLER_80_2160 ();
 sg13g2_decap_8 FILLER_80_2167 ();
 sg13g2_decap_8 FILLER_80_2174 ();
 sg13g2_fill_1 FILLER_80_2181 ();
 sg13g2_decap_8 FILLER_80_2186 ();
 sg13g2_decap_8 FILLER_80_2193 ();
 sg13g2_decap_8 FILLER_80_2200 ();
 sg13g2_fill_2 FILLER_80_2207 ();
 sg13g2_fill_1 FILLER_80_2209 ();
 sg13g2_decap_8 FILLER_80_2214 ();
 sg13g2_decap_8 FILLER_80_2221 ();
 sg13g2_decap_8 FILLER_80_2228 ();
 sg13g2_fill_2 FILLER_80_2235 ();
 sg13g2_decap_4 FILLER_80_2241 ();
 sg13g2_fill_1 FILLER_80_2245 ();
 sg13g2_decap_8 FILLER_80_2259 ();
 sg13g2_decap_8 FILLER_80_2266 ();
 sg13g2_fill_1 FILLER_80_2273 ();
 sg13g2_decap_8 FILLER_80_2277 ();
 sg13g2_fill_1 FILLER_80_2284 ();
 sg13g2_decap_8 FILLER_80_2289 ();
 sg13g2_decap_8 FILLER_80_2296 ();
 sg13g2_decap_4 FILLER_80_2303 ();
 sg13g2_fill_1 FILLER_80_2307 ();
 sg13g2_decap_8 FILLER_80_2325 ();
 sg13g2_decap_4 FILLER_80_2332 ();
 sg13g2_fill_2 FILLER_80_2336 ();
 sg13g2_fill_2 FILLER_80_2342 ();
 sg13g2_decap_8 FILLER_80_2348 ();
 sg13g2_decap_8 FILLER_80_2355 ();
 sg13g2_decap_8 FILLER_80_2392 ();
 sg13g2_decap_4 FILLER_80_2399 ();
 sg13g2_fill_2 FILLER_80_2403 ();
 sg13g2_decap_4 FILLER_80_2409 ();
 sg13g2_fill_2 FILLER_80_2413 ();
 sg13g2_decap_4 FILLER_80_2419 ();
 sg13g2_decap_4 FILLER_80_2449 ();
 sg13g2_fill_2 FILLER_80_2453 ();
 sg13g2_decap_8 FILLER_80_2459 ();
 sg13g2_decap_8 FILLER_80_2466 ();
 sg13g2_decap_8 FILLER_80_2473 ();
 sg13g2_decap_8 FILLER_80_2480 ();
 sg13g2_fill_2 FILLER_80_2487 ();
 sg13g2_fill_1 FILLER_80_2506 ();
 sg13g2_decap_8 FILLER_80_2511 ();
 sg13g2_decap_4 FILLER_80_2518 ();
 sg13g2_fill_2 FILLER_80_2522 ();
 sg13g2_decap_8 FILLER_80_2529 ();
 sg13g2_fill_2 FILLER_80_2536 ();
 sg13g2_fill_1 FILLER_80_2538 ();
 sg13g2_fill_1 FILLER_80_2544 ();
 sg13g2_decap_8 FILLER_80_2571 ();
 sg13g2_decap_8 FILLER_80_2578 ();
 sg13g2_decap_8 FILLER_80_2585 ();
 sg13g2_decap_8 FILLER_80_2592 ();
 sg13g2_decap_8 FILLER_80_2599 ();
 sg13g2_decap_8 FILLER_80_2606 ();
 sg13g2_decap_8 FILLER_80_2613 ();
 sg13g2_decap_8 FILLER_80_2620 ();
 sg13g2_decap_8 FILLER_80_2627 ();
 sg13g2_decap_8 FILLER_80_2634 ();
 sg13g2_decap_8 FILLER_80_2641 ();
 sg13g2_decap_8 FILLER_80_2648 ();
 sg13g2_decap_8 FILLER_80_2655 ();
 sg13g2_decap_8 FILLER_80_2662 ();
 sg13g2_fill_1 FILLER_80_2669 ();
endmodule
