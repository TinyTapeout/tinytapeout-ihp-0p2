module tt_um_vc32_cpu (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire clknet_leaf_0_clk;
 wire \cpu.addr[10] ;
 wire \cpu.addr[11] ;
 wire \cpu.addr[12] ;
 wire \cpu.addr[13] ;
 wire \cpu.addr[14] ;
 wire \cpu.addr[15] ;
 wire \cpu.addr[1] ;
 wire \cpu.addr[2] ;
 wire \cpu.addr[3] ;
 wire \cpu.addr[4] ;
 wire \cpu.addr[5] ;
 wire \cpu.addr[6] ;
 wire \cpu.addr[7] ;
 wire \cpu.addr[8] ;
 wire \cpu.addr[9] ;
 wire \cpu.br ;
 wire \cpu.cond[0] ;
 wire \cpu.cond[1] ;
 wire \cpu.cond[2] ;
 wire \cpu.d_flush_all ;
 wire \cpu.d_rstrobe_d ;
 wire \cpu.d_wstrobe_d ;
 wire \cpu.dcache.flush_write ;
 wire \cpu.dcache.r_data[0][0] ;
 wire \cpu.dcache.r_data[0][10] ;
 wire \cpu.dcache.r_data[0][11] ;
 wire \cpu.dcache.r_data[0][12] ;
 wire \cpu.dcache.r_data[0][13] ;
 wire \cpu.dcache.r_data[0][14] ;
 wire \cpu.dcache.r_data[0][15] ;
 wire \cpu.dcache.r_data[0][16] ;
 wire \cpu.dcache.r_data[0][17] ;
 wire \cpu.dcache.r_data[0][18] ;
 wire \cpu.dcache.r_data[0][19] ;
 wire \cpu.dcache.r_data[0][1] ;
 wire \cpu.dcache.r_data[0][20] ;
 wire \cpu.dcache.r_data[0][21] ;
 wire \cpu.dcache.r_data[0][22] ;
 wire \cpu.dcache.r_data[0][23] ;
 wire \cpu.dcache.r_data[0][24] ;
 wire \cpu.dcache.r_data[0][25] ;
 wire \cpu.dcache.r_data[0][26] ;
 wire \cpu.dcache.r_data[0][27] ;
 wire \cpu.dcache.r_data[0][28] ;
 wire \cpu.dcache.r_data[0][29] ;
 wire \cpu.dcache.r_data[0][2] ;
 wire \cpu.dcache.r_data[0][30] ;
 wire \cpu.dcache.r_data[0][31] ;
 wire \cpu.dcache.r_data[0][3] ;
 wire \cpu.dcache.r_data[0][4] ;
 wire \cpu.dcache.r_data[0][5] ;
 wire \cpu.dcache.r_data[0][6] ;
 wire \cpu.dcache.r_data[0][7] ;
 wire \cpu.dcache.r_data[0][8] ;
 wire \cpu.dcache.r_data[0][9] ;
 wire \cpu.dcache.r_data[1][0] ;
 wire \cpu.dcache.r_data[1][10] ;
 wire \cpu.dcache.r_data[1][11] ;
 wire \cpu.dcache.r_data[1][12] ;
 wire \cpu.dcache.r_data[1][13] ;
 wire \cpu.dcache.r_data[1][14] ;
 wire \cpu.dcache.r_data[1][15] ;
 wire \cpu.dcache.r_data[1][16] ;
 wire \cpu.dcache.r_data[1][17] ;
 wire \cpu.dcache.r_data[1][18] ;
 wire \cpu.dcache.r_data[1][19] ;
 wire \cpu.dcache.r_data[1][1] ;
 wire \cpu.dcache.r_data[1][20] ;
 wire \cpu.dcache.r_data[1][21] ;
 wire \cpu.dcache.r_data[1][22] ;
 wire \cpu.dcache.r_data[1][23] ;
 wire \cpu.dcache.r_data[1][24] ;
 wire \cpu.dcache.r_data[1][25] ;
 wire \cpu.dcache.r_data[1][26] ;
 wire \cpu.dcache.r_data[1][27] ;
 wire \cpu.dcache.r_data[1][28] ;
 wire \cpu.dcache.r_data[1][29] ;
 wire \cpu.dcache.r_data[1][2] ;
 wire \cpu.dcache.r_data[1][30] ;
 wire \cpu.dcache.r_data[1][31] ;
 wire \cpu.dcache.r_data[1][3] ;
 wire \cpu.dcache.r_data[1][4] ;
 wire \cpu.dcache.r_data[1][5] ;
 wire \cpu.dcache.r_data[1][6] ;
 wire \cpu.dcache.r_data[1][7] ;
 wire \cpu.dcache.r_data[1][8] ;
 wire \cpu.dcache.r_data[1][9] ;
 wire \cpu.dcache.r_data[2][0] ;
 wire \cpu.dcache.r_data[2][10] ;
 wire \cpu.dcache.r_data[2][11] ;
 wire \cpu.dcache.r_data[2][12] ;
 wire \cpu.dcache.r_data[2][13] ;
 wire \cpu.dcache.r_data[2][14] ;
 wire \cpu.dcache.r_data[2][15] ;
 wire \cpu.dcache.r_data[2][16] ;
 wire \cpu.dcache.r_data[2][17] ;
 wire \cpu.dcache.r_data[2][18] ;
 wire \cpu.dcache.r_data[2][19] ;
 wire \cpu.dcache.r_data[2][1] ;
 wire \cpu.dcache.r_data[2][20] ;
 wire \cpu.dcache.r_data[2][21] ;
 wire \cpu.dcache.r_data[2][22] ;
 wire \cpu.dcache.r_data[2][23] ;
 wire \cpu.dcache.r_data[2][24] ;
 wire \cpu.dcache.r_data[2][25] ;
 wire \cpu.dcache.r_data[2][26] ;
 wire \cpu.dcache.r_data[2][27] ;
 wire \cpu.dcache.r_data[2][28] ;
 wire \cpu.dcache.r_data[2][29] ;
 wire \cpu.dcache.r_data[2][2] ;
 wire \cpu.dcache.r_data[2][30] ;
 wire \cpu.dcache.r_data[2][31] ;
 wire \cpu.dcache.r_data[2][3] ;
 wire \cpu.dcache.r_data[2][4] ;
 wire \cpu.dcache.r_data[2][5] ;
 wire \cpu.dcache.r_data[2][6] ;
 wire \cpu.dcache.r_data[2][7] ;
 wire \cpu.dcache.r_data[2][8] ;
 wire \cpu.dcache.r_data[2][9] ;
 wire \cpu.dcache.r_data[3][0] ;
 wire \cpu.dcache.r_data[3][10] ;
 wire \cpu.dcache.r_data[3][11] ;
 wire \cpu.dcache.r_data[3][12] ;
 wire \cpu.dcache.r_data[3][13] ;
 wire \cpu.dcache.r_data[3][14] ;
 wire \cpu.dcache.r_data[3][15] ;
 wire \cpu.dcache.r_data[3][16] ;
 wire \cpu.dcache.r_data[3][17] ;
 wire \cpu.dcache.r_data[3][18] ;
 wire \cpu.dcache.r_data[3][19] ;
 wire \cpu.dcache.r_data[3][1] ;
 wire \cpu.dcache.r_data[3][20] ;
 wire \cpu.dcache.r_data[3][21] ;
 wire \cpu.dcache.r_data[3][22] ;
 wire \cpu.dcache.r_data[3][23] ;
 wire \cpu.dcache.r_data[3][24] ;
 wire \cpu.dcache.r_data[3][25] ;
 wire \cpu.dcache.r_data[3][26] ;
 wire \cpu.dcache.r_data[3][27] ;
 wire \cpu.dcache.r_data[3][28] ;
 wire \cpu.dcache.r_data[3][29] ;
 wire \cpu.dcache.r_data[3][2] ;
 wire \cpu.dcache.r_data[3][30] ;
 wire \cpu.dcache.r_data[3][31] ;
 wire \cpu.dcache.r_data[3][3] ;
 wire \cpu.dcache.r_data[3][4] ;
 wire \cpu.dcache.r_data[3][5] ;
 wire \cpu.dcache.r_data[3][6] ;
 wire \cpu.dcache.r_data[3][7] ;
 wire \cpu.dcache.r_data[3][8] ;
 wire \cpu.dcache.r_data[3][9] ;
 wire \cpu.dcache.r_data[4][0] ;
 wire \cpu.dcache.r_data[4][10] ;
 wire \cpu.dcache.r_data[4][11] ;
 wire \cpu.dcache.r_data[4][12] ;
 wire \cpu.dcache.r_data[4][13] ;
 wire \cpu.dcache.r_data[4][14] ;
 wire \cpu.dcache.r_data[4][15] ;
 wire \cpu.dcache.r_data[4][16] ;
 wire \cpu.dcache.r_data[4][17] ;
 wire \cpu.dcache.r_data[4][18] ;
 wire \cpu.dcache.r_data[4][19] ;
 wire \cpu.dcache.r_data[4][1] ;
 wire \cpu.dcache.r_data[4][20] ;
 wire \cpu.dcache.r_data[4][21] ;
 wire \cpu.dcache.r_data[4][22] ;
 wire \cpu.dcache.r_data[4][23] ;
 wire \cpu.dcache.r_data[4][24] ;
 wire \cpu.dcache.r_data[4][25] ;
 wire \cpu.dcache.r_data[4][26] ;
 wire \cpu.dcache.r_data[4][27] ;
 wire \cpu.dcache.r_data[4][28] ;
 wire \cpu.dcache.r_data[4][29] ;
 wire \cpu.dcache.r_data[4][2] ;
 wire \cpu.dcache.r_data[4][30] ;
 wire \cpu.dcache.r_data[4][31] ;
 wire \cpu.dcache.r_data[4][3] ;
 wire \cpu.dcache.r_data[4][4] ;
 wire \cpu.dcache.r_data[4][5] ;
 wire \cpu.dcache.r_data[4][6] ;
 wire \cpu.dcache.r_data[4][7] ;
 wire \cpu.dcache.r_data[4][8] ;
 wire \cpu.dcache.r_data[4][9] ;
 wire \cpu.dcache.r_data[5][0] ;
 wire \cpu.dcache.r_data[5][10] ;
 wire \cpu.dcache.r_data[5][11] ;
 wire \cpu.dcache.r_data[5][12] ;
 wire \cpu.dcache.r_data[5][13] ;
 wire \cpu.dcache.r_data[5][14] ;
 wire \cpu.dcache.r_data[5][15] ;
 wire \cpu.dcache.r_data[5][16] ;
 wire \cpu.dcache.r_data[5][17] ;
 wire \cpu.dcache.r_data[5][18] ;
 wire \cpu.dcache.r_data[5][19] ;
 wire \cpu.dcache.r_data[5][1] ;
 wire \cpu.dcache.r_data[5][20] ;
 wire \cpu.dcache.r_data[5][21] ;
 wire \cpu.dcache.r_data[5][22] ;
 wire \cpu.dcache.r_data[5][23] ;
 wire \cpu.dcache.r_data[5][24] ;
 wire \cpu.dcache.r_data[5][25] ;
 wire \cpu.dcache.r_data[5][26] ;
 wire \cpu.dcache.r_data[5][27] ;
 wire \cpu.dcache.r_data[5][28] ;
 wire \cpu.dcache.r_data[5][29] ;
 wire \cpu.dcache.r_data[5][2] ;
 wire \cpu.dcache.r_data[5][30] ;
 wire \cpu.dcache.r_data[5][31] ;
 wire \cpu.dcache.r_data[5][3] ;
 wire \cpu.dcache.r_data[5][4] ;
 wire \cpu.dcache.r_data[5][5] ;
 wire \cpu.dcache.r_data[5][6] ;
 wire \cpu.dcache.r_data[5][7] ;
 wire \cpu.dcache.r_data[5][8] ;
 wire \cpu.dcache.r_data[5][9] ;
 wire \cpu.dcache.r_data[6][0] ;
 wire \cpu.dcache.r_data[6][10] ;
 wire \cpu.dcache.r_data[6][11] ;
 wire \cpu.dcache.r_data[6][12] ;
 wire \cpu.dcache.r_data[6][13] ;
 wire \cpu.dcache.r_data[6][14] ;
 wire \cpu.dcache.r_data[6][15] ;
 wire \cpu.dcache.r_data[6][16] ;
 wire \cpu.dcache.r_data[6][17] ;
 wire \cpu.dcache.r_data[6][18] ;
 wire \cpu.dcache.r_data[6][19] ;
 wire \cpu.dcache.r_data[6][1] ;
 wire \cpu.dcache.r_data[6][20] ;
 wire \cpu.dcache.r_data[6][21] ;
 wire \cpu.dcache.r_data[6][22] ;
 wire \cpu.dcache.r_data[6][23] ;
 wire \cpu.dcache.r_data[6][24] ;
 wire \cpu.dcache.r_data[6][25] ;
 wire \cpu.dcache.r_data[6][26] ;
 wire \cpu.dcache.r_data[6][27] ;
 wire \cpu.dcache.r_data[6][28] ;
 wire \cpu.dcache.r_data[6][29] ;
 wire \cpu.dcache.r_data[6][2] ;
 wire \cpu.dcache.r_data[6][30] ;
 wire \cpu.dcache.r_data[6][31] ;
 wire \cpu.dcache.r_data[6][3] ;
 wire \cpu.dcache.r_data[6][4] ;
 wire \cpu.dcache.r_data[6][5] ;
 wire \cpu.dcache.r_data[6][6] ;
 wire \cpu.dcache.r_data[6][7] ;
 wire \cpu.dcache.r_data[6][8] ;
 wire \cpu.dcache.r_data[6][9] ;
 wire \cpu.dcache.r_data[7][0] ;
 wire \cpu.dcache.r_data[7][10] ;
 wire \cpu.dcache.r_data[7][11] ;
 wire \cpu.dcache.r_data[7][12] ;
 wire \cpu.dcache.r_data[7][13] ;
 wire \cpu.dcache.r_data[7][14] ;
 wire \cpu.dcache.r_data[7][15] ;
 wire \cpu.dcache.r_data[7][16] ;
 wire \cpu.dcache.r_data[7][17] ;
 wire \cpu.dcache.r_data[7][18] ;
 wire \cpu.dcache.r_data[7][19] ;
 wire \cpu.dcache.r_data[7][1] ;
 wire \cpu.dcache.r_data[7][20] ;
 wire \cpu.dcache.r_data[7][21] ;
 wire \cpu.dcache.r_data[7][22] ;
 wire \cpu.dcache.r_data[7][23] ;
 wire \cpu.dcache.r_data[7][24] ;
 wire \cpu.dcache.r_data[7][25] ;
 wire \cpu.dcache.r_data[7][26] ;
 wire \cpu.dcache.r_data[7][27] ;
 wire \cpu.dcache.r_data[7][28] ;
 wire \cpu.dcache.r_data[7][29] ;
 wire \cpu.dcache.r_data[7][2] ;
 wire \cpu.dcache.r_data[7][30] ;
 wire \cpu.dcache.r_data[7][31] ;
 wire \cpu.dcache.r_data[7][3] ;
 wire \cpu.dcache.r_data[7][4] ;
 wire \cpu.dcache.r_data[7][5] ;
 wire \cpu.dcache.r_data[7][6] ;
 wire \cpu.dcache.r_data[7][7] ;
 wire \cpu.dcache.r_data[7][8] ;
 wire \cpu.dcache.r_data[7][9] ;
 wire \cpu.dcache.r_dirty[0] ;
 wire \cpu.dcache.r_dirty[1] ;
 wire \cpu.dcache.r_dirty[2] ;
 wire \cpu.dcache.r_dirty[3] ;
 wire \cpu.dcache.r_dirty[4] ;
 wire \cpu.dcache.r_dirty[5] ;
 wire \cpu.dcache.r_dirty[6] ;
 wire \cpu.dcache.r_dirty[7] ;
 wire \cpu.dcache.r_offset[0] ;
 wire \cpu.dcache.r_offset[1] ;
 wire \cpu.dcache.r_offset[2] ;
 wire \cpu.dcache.r_tag[0][10] ;
 wire \cpu.dcache.r_tag[0][11] ;
 wire \cpu.dcache.r_tag[0][12] ;
 wire \cpu.dcache.r_tag[0][13] ;
 wire \cpu.dcache.r_tag[0][14] ;
 wire \cpu.dcache.r_tag[0][15] ;
 wire \cpu.dcache.r_tag[0][16] ;
 wire \cpu.dcache.r_tag[0][17] ;
 wire \cpu.dcache.r_tag[0][18] ;
 wire \cpu.dcache.r_tag[0][19] ;
 wire \cpu.dcache.r_tag[0][20] ;
 wire \cpu.dcache.r_tag[0][21] ;
 wire \cpu.dcache.r_tag[0][22] ;
 wire \cpu.dcache.r_tag[0][23] ;
 wire \cpu.dcache.r_tag[0][5] ;
 wire \cpu.dcache.r_tag[0][6] ;
 wire \cpu.dcache.r_tag[0][7] ;
 wire \cpu.dcache.r_tag[0][8] ;
 wire \cpu.dcache.r_tag[0][9] ;
 wire \cpu.dcache.r_tag[1][10] ;
 wire \cpu.dcache.r_tag[1][11] ;
 wire \cpu.dcache.r_tag[1][12] ;
 wire \cpu.dcache.r_tag[1][13] ;
 wire \cpu.dcache.r_tag[1][14] ;
 wire \cpu.dcache.r_tag[1][15] ;
 wire \cpu.dcache.r_tag[1][16] ;
 wire \cpu.dcache.r_tag[1][17] ;
 wire \cpu.dcache.r_tag[1][18] ;
 wire \cpu.dcache.r_tag[1][19] ;
 wire \cpu.dcache.r_tag[1][20] ;
 wire \cpu.dcache.r_tag[1][21] ;
 wire \cpu.dcache.r_tag[1][22] ;
 wire \cpu.dcache.r_tag[1][23] ;
 wire \cpu.dcache.r_tag[1][5] ;
 wire \cpu.dcache.r_tag[1][6] ;
 wire \cpu.dcache.r_tag[1][7] ;
 wire \cpu.dcache.r_tag[1][8] ;
 wire \cpu.dcache.r_tag[1][9] ;
 wire \cpu.dcache.r_tag[2][10] ;
 wire \cpu.dcache.r_tag[2][11] ;
 wire \cpu.dcache.r_tag[2][12] ;
 wire \cpu.dcache.r_tag[2][13] ;
 wire \cpu.dcache.r_tag[2][14] ;
 wire \cpu.dcache.r_tag[2][15] ;
 wire \cpu.dcache.r_tag[2][16] ;
 wire \cpu.dcache.r_tag[2][17] ;
 wire \cpu.dcache.r_tag[2][18] ;
 wire \cpu.dcache.r_tag[2][19] ;
 wire \cpu.dcache.r_tag[2][20] ;
 wire \cpu.dcache.r_tag[2][21] ;
 wire \cpu.dcache.r_tag[2][22] ;
 wire \cpu.dcache.r_tag[2][23] ;
 wire \cpu.dcache.r_tag[2][5] ;
 wire \cpu.dcache.r_tag[2][6] ;
 wire \cpu.dcache.r_tag[2][7] ;
 wire \cpu.dcache.r_tag[2][8] ;
 wire \cpu.dcache.r_tag[2][9] ;
 wire \cpu.dcache.r_tag[3][10] ;
 wire \cpu.dcache.r_tag[3][11] ;
 wire \cpu.dcache.r_tag[3][12] ;
 wire \cpu.dcache.r_tag[3][13] ;
 wire \cpu.dcache.r_tag[3][14] ;
 wire \cpu.dcache.r_tag[3][15] ;
 wire \cpu.dcache.r_tag[3][16] ;
 wire \cpu.dcache.r_tag[3][17] ;
 wire \cpu.dcache.r_tag[3][18] ;
 wire \cpu.dcache.r_tag[3][19] ;
 wire \cpu.dcache.r_tag[3][20] ;
 wire \cpu.dcache.r_tag[3][21] ;
 wire \cpu.dcache.r_tag[3][22] ;
 wire \cpu.dcache.r_tag[3][23] ;
 wire \cpu.dcache.r_tag[3][5] ;
 wire \cpu.dcache.r_tag[3][6] ;
 wire \cpu.dcache.r_tag[3][7] ;
 wire \cpu.dcache.r_tag[3][8] ;
 wire \cpu.dcache.r_tag[3][9] ;
 wire \cpu.dcache.r_tag[4][10] ;
 wire \cpu.dcache.r_tag[4][11] ;
 wire \cpu.dcache.r_tag[4][12] ;
 wire \cpu.dcache.r_tag[4][13] ;
 wire \cpu.dcache.r_tag[4][14] ;
 wire \cpu.dcache.r_tag[4][15] ;
 wire \cpu.dcache.r_tag[4][16] ;
 wire \cpu.dcache.r_tag[4][17] ;
 wire \cpu.dcache.r_tag[4][18] ;
 wire \cpu.dcache.r_tag[4][19] ;
 wire \cpu.dcache.r_tag[4][20] ;
 wire \cpu.dcache.r_tag[4][21] ;
 wire \cpu.dcache.r_tag[4][22] ;
 wire \cpu.dcache.r_tag[4][23] ;
 wire \cpu.dcache.r_tag[4][5] ;
 wire \cpu.dcache.r_tag[4][6] ;
 wire \cpu.dcache.r_tag[4][7] ;
 wire \cpu.dcache.r_tag[4][8] ;
 wire \cpu.dcache.r_tag[4][9] ;
 wire \cpu.dcache.r_tag[5][10] ;
 wire \cpu.dcache.r_tag[5][11] ;
 wire \cpu.dcache.r_tag[5][12] ;
 wire \cpu.dcache.r_tag[5][13] ;
 wire \cpu.dcache.r_tag[5][14] ;
 wire \cpu.dcache.r_tag[5][15] ;
 wire \cpu.dcache.r_tag[5][16] ;
 wire \cpu.dcache.r_tag[5][17] ;
 wire \cpu.dcache.r_tag[5][18] ;
 wire \cpu.dcache.r_tag[5][19] ;
 wire \cpu.dcache.r_tag[5][20] ;
 wire \cpu.dcache.r_tag[5][21] ;
 wire \cpu.dcache.r_tag[5][22] ;
 wire \cpu.dcache.r_tag[5][23] ;
 wire \cpu.dcache.r_tag[5][5] ;
 wire \cpu.dcache.r_tag[5][6] ;
 wire \cpu.dcache.r_tag[5][7] ;
 wire \cpu.dcache.r_tag[5][8] ;
 wire \cpu.dcache.r_tag[5][9] ;
 wire \cpu.dcache.r_tag[6][10] ;
 wire \cpu.dcache.r_tag[6][11] ;
 wire \cpu.dcache.r_tag[6][12] ;
 wire \cpu.dcache.r_tag[6][13] ;
 wire \cpu.dcache.r_tag[6][14] ;
 wire \cpu.dcache.r_tag[6][15] ;
 wire \cpu.dcache.r_tag[6][16] ;
 wire \cpu.dcache.r_tag[6][17] ;
 wire \cpu.dcache.r_tag[6][18] ;
 wire \cpu.dcache.r_tag[6][19] ;
 wire \cpu.dcache.r_tag[6][20] ;
 wire \cpu.dcache.r_tag[6][21] ;
 wire \cpu.dcache.r_tag[6][22] ;
 wire \cpu.dcache.r_tag[6][23] ;
 wire \cpu.dcache.r_tag[6][5] ;
 wire \cpu.dcache.r_tag[6][6] ;
 wire \cpu.dcache.r_tag[6][7] ;
 wire \cpu.dcache.r_tag[6][8] ;
 wire \cpu.dcache.r_tag[6][9] ;
 wire \cpu.dcache.r_tag[7][10] ;
 wire \cpu.dcache.r_tag[7][11] ;
 wire \cpu.dcache.r_tag[7][12] ;
 wire \cpu.dcache.r_tag[7][13] ;
 wire \cpu.dcache.r_tag[7][14] ;
 wire \cpu.dcache.r_tag[7][15] ;
 wire \cpu.dcache.r_tag[7][16] ;
 wire \cpu.dcache.r_tag[7][17] ;
 wire \cpu.dcache.r_tag[7][18] ;
 wire \cpu.dcache.r_tag[7][19] ;
 wire \cpu.dcache.r_tag[7][20] ;
 wire \cpu.dcache.r_tag[7][21] ;
 wire \cpu.dcache.r_tag[7][22] ;
 wire \cpu.dcache.r_tag[7][23] ;
 wire \cpu.dcache.r_tag[7][5] ;
 wire \cpu.dcache.r_tag[7][6] ;
 wire \cpu.dcache.r_tag[7][7] ;
 wire \cpu.dcache.r_tag[7][8] ;
 wire \cpu.dcache.r_tag[7][9] ;
 wire \cpu.dcache.r_valid[0] ;
 wire \cpu.dcache.r_valid[1] ;
 wire \cpu.dcache.r_valid[2] ;
 wire \cpu.dcache.r_valid[3] ;
 wire \cpu.dcache.r_valid[4] ;
 wire \cpu.dcache.r_valid[5] ;
 wire \cpu.dcache.r_valid[6] ;
 wire \cpu.dcache.r_valid[7] ;
 wire \cpu.dcache.wdata[0] ;
 wire \cpu.dcache.wdata[10] ;
 wire \cpu.dcache.wdata[11] ;
 wire \cpu.dcache.wdata[12] ;
 wire \cpu.dcache.wdata[13] ;
 wire \cpu.dcache.wdata[14] ;
 wire \cpu.dcache.wdata[15] ;
 wire \cpu.dcache.wdata[1] ;
 wire \cpu.dcache.wdata[2] ;
 wire \cpu.dcache.wdata[3] ;
 wire \cpu.dcache.wdata[4] ;
 wire \cpu.dcache.wdata[5] ;
 wire \cpu.dcache.wdata[6] ;
 wire \cpu.dcache.wdata[7] ;
 wire \cpu.dcache.wdata[8] ;
 wire \cpu.dcache.wdata[9] ;
 wire \cpu.dec.div ;
 wire \cpu.dec.do_flush_all ;
 wire \cpu.dec.do_flush_write ;
 wire \cpu.dec.do_inv_mmu ;
 wire \cpu.dec.imm[0] ;
 wire \cpu.dec.imm[10] ;
 wire \cpu.dec.imm[11] ;
 wire \cpu.dec.imm[12] ;
 wire \cpu.dec.imm[13] ;
 wire \cpu.dec.imm[14] ;
 wire \cpu.dec.imm[15] ;
 wire \cpu.dec.imm[1] ;
 wire \cpu.dec.imm[2] ;
 wire \cpu.dec.imm[3] ;
 wire \cpu.dec.imm[4] ;
 wire \cpu.dec.imm[5] ;
 wire \cpu.dec.imm[6] ;
 wire \cpu.dec.imm[7] ;
 wire \cpu.dec.imm[8] ;
 wire \cpu.dec.imm[9] ;
 wire \cpu.dec.io ;
 wire \cpu.dec.iready ;
 wire \cpu.dec.jmp ;
 wire \cpu.dec.load ;
 wire \cpu.dec.mult ;
 wire \cpu.dec.needs_rs2 ;
 wire \cpu.dec.r_op[10] ;
 wire \cpu.dec.r_op[1] ;
 wire \cpu.dec.r_op[2] ;
 wire \cpu.dec.r_op[3] ;
 wire \cpu.dec.r_op[4] ;
 wire \cpu.dec.r_op[5] ;
 wire \cpu.dec.r_op[6] ;
 wire \cpu.dec.r_op[7] ;
 wire \cpu.dec.r_op[8] ;
 wire \cpu.dec.r_op[9] ;
 wire \cpu.dec.r_rd[0] ;
 wire \cpu.dec.r_rd[1] ;
 wire \cpu.dec.r_rd[2] ;
 wire \cpu.dec.r_rd[3] ;
 wire \cpu.dec.r_rs1[0] ;
 wire \cpu.dec.r_rs1[1] ;
 wire \cpu.dec.r_rs1[2] ;
 wire \cpu.dec.r_rs1[3] ;
 wire \cpu.dec.r_rs2[0] ;
 wire \cpu.dec.r_rs2[1] ;
 wire \cpu.dec.r_rs2[2] ;
 wire \cpu.dec.r_rs2[3] ;
 wire \cpu.dec.r_rs2_pc ;
 wire \cpu.dec.r_set_cc ;
 wire \cpu.dec.r_store ;
 wire \cpu.dec.r_swapsp ;
 wire \cpu.dec.r_sys_call ;
 wire \cpu.dec.r_trap ;
 wire \cpu.dec.supmode ;
 wire \cpu.dec.user_io ;
 wire \cpu.ex.c_div_running ;
 wire \cpu.ex.c_mult[0] ;
 wire \cpu.ex.c_mult[10] ;
 wire \cpu.ex.c_mult[11] ;
 wire \cpu.ex.c_mult[12] ;
 wire \cpu.ex.c_mult[13] ;
 wire \cpu.ex.c_mult[14] ;
 wire \cpu.ex.c_mult[15] ;
 wire \cpu.ex.c_mult[1] ;
 wire \cpu.ex.c_mult[2] ;
 wire \cpu.ex.c_mult[3] ;
 wire \cpu.ex.c_mult[4] ;
 wire \cpu.ex.c_mult[5] ;
 wire \cpu.ex.c_mult[6] ;
 wire \cpu.ex.c_mult[7] ;
 wire \cpu.ex.c_mult[8] ;
 wire \cpu.ex.c_mult[9] ;
 wire \cpu.ex.c_mult_off[0] ;
 wire \cpu.ex.c_mult_off[1] ;
 wire \cpu.ex.c_mult_off[2] ;
 wire \cpu.ex.c_mult_off[3] ;
 wire \cpu.ex.c_mult_running ;
 wire \cpu.ex.genblk3.c_supmode ;
 wire \cpu.ex.genblk3.r_mmu_d_proxy ;
 wire \cpu.ex.genblk3.r_mmu_enable ;
 wire \cpu.ex.genblk3.r_prev_supmode ;
 wire \cpu.ex.i_flush_all ;
 wire \cpu.ex.ifetch ;
 wire \cpu.ex.io_access ;
 wire \cpu.ex.mmu_read[12] ;
 wire \cpu.ex.mmu_read[13] ;
 wire \cpu.ex.mmu_read[14] ;
 wire \cpu.ex.mmu_read[15] ;
 wire \cpu.ex.mmu_read[1] ;
 wire \cpu.ex.mmu_read[2] ;
 wire \cpu.ex.mmu_read[3] ;
 wire \cpu.ex.mmu_reg_data[0] ;
 wire \cpu.ex.pc[10] ;
 wire \cpu.ex.pc[11] ;
 wire \cpu.ex.pc[12] ;
 wire \cpu.ex.pc[13] ;
 wire \cpu.ex.pc[14] ;
 wire \cpu.ex.pc[15] ;
 wire \cpu.ex.pc[1] ;
 wire \cpu.ex.pc[2] ;
 wire \cpu.ex.pc[3] ;
 wire \cpu.ex.pc[4] ;
 wire \cpu.ex.pc[5] ;
 wire \cpu.ex.pc[6] ;
 wire \cpu.ex.pc[7] ;
 wire \cpu.ex.pc[8] ;
 wire \cpu.ex.pc[9] ;
 wire \cpu.ex.r_10[0] ;
 wire \cpu.ex.r_10[10] ;
 wire \cpu.ex.r_10[11] ;
 wire \cpu.ex.r_10[12] ;
 wire \cpu.ex.r_10[13] ;
 wire \cpu.ex.r_10[14] ;
 wire \cpu.ex.r_10[15] ;
 wire \cpu.ex.r_10[1] ;
 wire \cpu.ex.r_10[2] ;
 wire \cpu.ex.r_10[3] ;
 wire \cpu.ex.r_10[4] ;
 wire \cpu.ex.r_10[5] ;
 wire \cpu.ex.r_10[6] ;
 wire \cpu.ex.r_10[7] ;
 wire \cpu.ex.r_10[8] ;
 wire \cpu.ex.r_10[9] ;
 wire \cpu.ex.r_11[0] ;
 wire \cpu.ex.r_11[10] ;
 wire \cpu.ex.r_11[11] ;
 wire \cpu.ex.r_11[12] ;
 wire \cpu.ex.r_11[13] ;
 wire \cpu.ex.r_11[14] ;
 wire \cpu.ex.r_11[15] ;
 wire \cpu.ex.r_11[1] ;
 wire \cpu.ex.r_11[2] ;
 wire \cpu.ex.r_11[3] ;
 wire \cpu.ex.r_11[4] ;
 wire \cpu.ex.r_11[5] ;
 wire \cpu.ex.r_11[6] ;
 wire \cpu.ex.r_11[7] ;
 wire \cpu.ex.r_11[8] ;
 wire \cpu.ex.r_11[9] ;
 wire \cpu.ex.r_12[0] ;
 wire \cpu.ex.r_12[10] ;
 wire \cpu.ex.r_12[11] ;
 wire \cpu.ex.r_12[12] ;
 wire \cpu.ex.r_12[13] ;
 wire \cpu.ex.r_12[14] ;
 wire \cpu.ex.r_12[15] ;
 wire \cpu.ex.r_12[1] ;
 wire \cpu.ex.r_12[2] ;
 wire \cpu.ex.r_12[3] ;
 wire \cpu.ex.r_12[4] ;
 wire \cpu.ex.r_12[5] ;
 wire \cpu.ex.r_12[6] ;
 wire \cpu.ex.r_12[7] ;
 wire \cpu.ex.r_12[8] ;
 wire \cpu.ex.r_12[9] ;
 wire \cpu.ex.r_13[0] ;
 wire \cpu.ex.r_13[10] ;
 wire \cpu.ex.r_13[11] ;
 wire \cpu.ex.r_13[12] ;
 wire \cpu.ex.r_13[13] ;
 wire \cpu.ex.r_13[14] ;
 wire \cpu.ex.r_13[15] ;
 wire \cpu.ex.r_13[1] ;
 wire \cpu.ex.r_13[2] ;
 wire \cpu.ex.r_13[3] ;
 wire \cpu.ex.r_13[4] ;
 wire \cpu.ex.r_13[5] ;
 wire \cpu.ex.r_13[6] ;
 wire \cpu.ex.r_13[7] ;
 wire \cpu.ex.r_13[8] ;
 wire \cpu.ex.r_13[9] ;
 wire \cpu.ex.r_14[0] ;
 wire \cpu.ex.r_14[10] ;
 wire \cpu.ex.r_14[11] ;
 wire \cpu.ex.r_14[12] ;
 wire \cpu.ex.r_14[13] ;
 wire \cpu.ex.r_14[14] ;
 wire \cpu.ex.r_14[15] ;
 wire \cpu.ex.r_14[1] ;
 wire \cpu.ex.r_14[2] ;
 wire \cpu.ex.r_14[3] ;
 wire \cpu.ex.r_14[4] ;
 wire \cpu.ex.r_14[5] ;
 wire \cpu.ex.r_14[6] ;
 wire \cpu.ex.r_14[7] ;
 wire \cpu.ex.r_14[8] ;
 wire \cpu.ex.r_14[9] ;
 wire \cpu.ex.r_15[0] ;
 wire \cpu.ex.r_15[10] ;
 wire \cpu.ex.r_15[11] ;
 wire \cpu.ex.r_15[12] ;
 wire \cpu.ex.r_15[13] ;
 wire \cpu.ex.r_15[14] ;
 wire \cpu.ex.r_15[15] ;
 wire \cpu.ex.r_15[1] ;
 wire \cpu.ex.r_15[2] ;
 wire \cpu.ex.r_15[3] ;
 wire \cpu.ex.r_15[4] ;
 wire \cpu.ex.r_15[5] ;
 wire \cpu.ex.r_15[6] ;
 wire \cpu.ex.r_15[7] ;
 wire \cpu.ex.r_15[8] ;
 wire \cpu.ex.r_15[9] ;
 wire \cpu.ex.r_8[0] ;
 wire \cpu.ex.r_8[10] ;
 wire \cpu.ex.r_8[11] ;
 wire \cpu.ex.r_8[12] ;
 wire \cpu.ex.r_8[13] ;
 wire \cpu.ex.r_8[14] ;
 wire \cpu.ex.r_8[15] ;
 wire \cpu.ex.r_8[1] ;
 wire \cpu.ex.r_8[2] ;
 wire \cpu.ex.r_8[3] ;
 wire \cpu.ex.r_8[4] ;
 wire \cpu.ex.r_8[5] ;
 wire \cpu.ex.r_8[6] ;
 wire \cpu.ex.r_8[7] ;
 wire \cpu.ex.r_8[8] ;
 wire \cpu.ex.r_8[9] ;
 wire \cpu.ex.r_9[0] ;
 wire \cpu.ex.r_9[10] ;
 wire \cpu.ex.r_9[11] ;
 wire \cpu.ex.r_9[12] ;
 wire \cpu.ex.r_9[13] ;
 wire \cpu.ex.r_9[14] ;
 wire \cpu.ex.r_9[15] ;
 wire \cpu.ex.r_9[1] ;
 wire \cpu.ex.r_9[2] ;
 wire \cpu.ex.r_9[3] ;
 wire \cpu.ex.r_9[4] ;
 wire \cpu.ex.r_9[5] ;
 wire \cpu.ex.r_9[6] ;
 wire \cpu.ex.r_9[7] ;
 wire \cpu.ex.r_9[8] ;
 wire \cpu.ex.r_9[9] ;
 wire \cpu.ex.r_branch_stall ;
 wire \cpu.ex.r_div_running ;
 wire \cpu.ex.r_epc[10] ;
 wire \cpu.ex.r_epc[11] ;
 wire \cpu.ex.r_epc[12] ;
 wire \cpu.ex.r_epc[13] ;
 wire \cpu.ex.r_epc[14] ;
 wire \cpu.ex.r_epc[15] ;
 wire \cpu.ex.r_epc[1] ;
 wire \cpu.ex.r_epc[2] ;
 wire \cpu.ex.r_epc[3] ;
 wire \cpu.ex.r_epc[4] ;
 wire \cpu.ex.r_epc[5] ;
 wire \cpu.ex.r_epc[6] ;
 wire \cpu.ex.r_epc[7] ;
 wire \cpu.ex.r_epc[8] ;
 wire \cpu.ex.r_epc[9] ;
 wire \cpu.ex.r_ie ;
 wire \cpu.ex.r_lr[10] ;
 wire \cpu.ex.r_lr[11] ;
 wire \cpu.ex.r_lr[12] ;
 wire \cpu.ex.r_lr[13] ;
 wire \cpu.ex.r_lr[14] ;
 wire \cpu.ex.r_lr[15] ;
 wire \cpu.ex.r_lr[1] ;
 wire \cpu.ex.r_lr[2] ;
 wire \cpu.ex.r_lr[3] ;
 wire \cpu.ex.r_lr[4] ;
 wire \cpu.ex.r_lr[5] ;
 wire \cpu.ex.r_lr[6] ;
 wire \cpu.ex.r_lr[7] ;
 wire \cpu.ex.r_lr[8] ;
 wire \cpu.ex.r_lr[9] ;
 wire \cpu.ex.r_mult[0] ;
 wire \cpu.ex.r_mult[10] ;
 wire \cpu.ex.r_mult[11] ;
 wire \cpu.ex.r_mult[12] ;
 wire \cpu.ex.r_mult[13] ;
 wire \cpu.ex.r_mult[14] ;
 wire \cpu.ex.r_mult[15] ;
 wire \cpu.ex.r_mult[16] ;
 wire \cpu.ex.r_mult[17] ;
 wire \cpu.ex.r_mult[18] ;
 wire \cpu.ex.r_mult[19] ;
 wire \cpu.ex.r_mult[1] ;
 wire \cpu.ex.r_mult[20] ;
 wire \cpu.ex.r_mult[21] ;
 wire \cpu.ex.r_mult[22] ;
 wire \cpu.ex.r_mult[23] ;
 wire \cpu.ex.r_mult[24] ;
 wire \cpu.ex.r_mult[25] ;
 wire \cpu.ex.r_mult[26] ;
 wire \cpu.ex.r_mult[27] ;
 wire \cpu.ex.r_mult[28] ;
 wire \cpu.ex.r_mult[29] ;
 wire \cpu.ex.r_mult[2] ;
 wire \cpu.ex.r_mult[30] ;
 wire \cpu.ex.r_mult[31] ;
 wire \cpu.ex.r_mult[3] ;
 wire \cpu.ex.r_mult[4] ;
 wire \cpu.ex.r_mult[5] ;
 wire \cpu.ex.r_mult[6] ;
 wire \cpu.ex.r_mult[7] ;
 wire \cpu.ex.r_mult[8] ;
 wire \cpu.ex.r_mult[9] ;
 wire \cpu.ex.r_mult_off[0] ;
 wire \cpu.ex.r_mult_off[1] ;
 wire \cpu.ex.r_mult_off[2] ;
 wire \cpu.ex.r_mult_off[3] ;
 wire \cpu.ex.r_mult_running ;
 wire \cpu.ex.r_prev_ie ;
 wire \cpu.ex.r_read_stall ;
 wire \cpu.ex.r_sp[10] ;
 wire \cpu.ex.r_sp[11] ;
 wire \cpu.ex.r_sp[12] ;
 wire \cpu.ex.r_sp[13] ;
 wire \cpu.ex.r_sp[14] ;
 wire \cpu.ex.r_sp[15] ;
 wire \cpu.ex.r_sp[1] ;
 wire \cpu.ex.r_sp[2] ;
 wire \cpu.ex.r_sp[3] ;
 wire \cpu.ex.r_sp[4] ;
 wire \cpu.ex.r_sp[5] ;
 wire \cpu.ex.r_sp[6] ;
 wire \cpu.ex.r_sp[7] ;
 wire \cpu.ex.r_sp[8] ;
 wire \cpu.ex.r_sp[9] ;
 wire \cpu.ex.r_stmp[0] ;
 wire \cpu.ex.r_stmp[10] ;
 wire \cpu.ex.r_stmp[11] ;
 wire \cpu.ex.r_stmp[12] ;
 wire \cpu.ex.r_stmp[13] ;
 wire \cpu.ex.r_stmp[14] ;
 wire \cpu.ex.r_stmp[15] ;
 wire \cpu.ex.r_stmp[1] ;
 wire \cpu.ex.r_stmp[2] ;
 wire \cpu.ex.r_stmp[3] ;
 wire \cpu.ex.r_stmp[4] ;
 wire \cpu.ex.r_stmp[5] ;
 wire \cpu.ex.r_stmp[6] ;
 wire \cpu.ex.r_stmp[7] ;
 wire \cpu.ex.r_stmp[8] ;
 wire \cpu.ex.r_stmp[9] ;
 wire \cpu.ex.r_wb_addr[0] ;
 wire \cpu.ex.r_wb_addr[1] ;
 wire \cpu.ex.r_wb_addr[2] ;
 wire \cpu.ex.r_wb_addr[3] ;
 wire \cpu.ex.r_wb_swapsp ;
 wire \cpu.ex.r_wb_valid ;
 wire \cpu.ex.r_wmask[0] ;
 wire \cpu.ex.r_wmask[1] ;
 wire \cpu.genblk1.mmu.r_valid_d[0] ;
 wire \cpu.genblk1.mmu.r_valid_d[10] ;
 wire \cpu.genblk1.mmu.r_valid_d[11] ;
 wire \cpu.genblk1.mmu.r_valid_d[12] ;
 wire \cpu.genblk1.mmu.r_valid_d[13] ;
 wire \cpu.genblk1.mmu.r_valid_d[14] ;
 wire \cpu.genblk1.mmu.r_valid_d[15] ;
 wire \cpu.genblk1.mmu.r_valid_d[16] ;
 wire \cpu.genblk1.mmu.r_valid_d[17] ;
 wire \cpu.genblk1.mmu.r_valid_d[18] ;
 wire \cpu.genblk1.mmu.r_valid_d[19] ;
 wire \cpu.genblk1.mmu.r_valid_d[1] ;
 wire \cpu.genblk1.mmu.r_valid_d[20] ;
 wire \cpu.genblk1.mmu.r_valid_d[21] ;
 wire \cpu.genblk1.mmu.r_valid_d[22] ;
 wire \cpu.genblk1.mmu.r_valid_d[23] ;
 wire \cpu.genblk1.mmu.r_valid_d[24] ;
 wire \cpu.genblk1.mmu.r_valid_d[25] ;
 wire \cpu.genblk1.mmu.r_valid_d[26] ;
 wire \cpu.genblk1.mmu.r_valid_d[27] ;
 wire \cpu.genblk1.mmu.r_valid_d[28] ;
 wire \cpu.genblk1.mmu.r_valid_d[29] ;
 wire \cpu.genblk1.mmu.r_valid_d[2] ;
 wire \cpu.genblk1.mmu.r_valid_d[30] ;
 wire \cpu.genblk1.mmu.r_valid_d[31] ;
 wire \cpu.genblk1.mmu.r_valid_d[3] ;
 wire \cpu.genblk1.mmu.r_valid_d[4] ;
 wire \cpu.genblk1.mmu.r_valid_d[5] ;
 wire \cpu.genblk1.mmu.r_valid_d[6] ;
 wire \cpu.genblk1.mmu.r_valid_d[7] ;
 wire \cpu.genblk1.mmu.r_valid_d[8] ;
 wire \cpu.genblk1.mmu.r_valid_d[9] ;
 wire \cpu.genblk1.mmu.r_valid_i[0] ;
 wire \cpu.genblk1.mmu.r_valid_i[10] ;
 wire \cpu.genblk1.mmu.r_valid_i[11] ;
 wire \cpu.genblk1.mmu.r_valid_i[12] ;
 wire \cpu.genblk1.mmu.r_valid_i[13] ;
 wire \cpu.genblk1.mmu.r_valid_i[14] ;
 wire \cpu.genblk1.mmu.r_valid_i[15] ;
 wire \cpu.genblk1.mmu.r_valid_i[16] ;
 wire \cpu.genblk1.mmu.r_valid_i[17] ;
 wire \cpu.genblk1.mmu.r_valid_i[18] ;
 wire \cpu.genblk1.mmu.r_valid_i[19] ;
 wire \cpu.genblk1.mmu.r_valid_i[1] ;
 wire \cpu.genblk1.mmu.r_valid_i[20] ;
 wire \cpu.genblk1.mmu.r_valid_i[21] ;
 wire \cpu.genblk1.mmu.r_valid_i[22] ;
 wire \cpu.genblk1.mmu.r_valid_i[23] ;
 wire \cpu.genblk1.mmu.r_valid_i[24] ;
 wire \cpu.genblk1.mmu.r_valid_i[25] ;
 wire \cpu.genblk1.mmu.r_valid_i[26] ;
 wire \cpu.genblk1.mmu.r_valid_i[27] ;
 wire \cpu.genblk1.mmu.r_valid_i[28] ;
 wire \cpu.genblk1.mmu.r_valid_i[29] ;
 wire \cpu.genblk1.mmu.r_valid_i[2] ;
 wire \cpu.genblk1.mmu.r_valid_i[30] ;
 wire \cpu.genblk1.mmu.r_valid_i[31] ;
 wire \cpu.genblk1.mmu.r_valid_i[3] ;
 wire \cpu.genblk1.mmu.r_valid_i[4] ;
 wire \cpu.genblk1.mmu.r_valid_i[5] ;
 wire \cpu.genblk1.mmu.r_valid_i[6] ;
 wire \cpu.genblk1.mmu.r_valid_i[7] ;
 wire \cpu.genblk1.mmu.r_valid_i[8] ;
 wire \cpu.genblk1.mmu.r_valid_i[9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][9] ;
 wire \cpu.genblk1.mmu.r_writeable_d[0] ;
 wire \cpu.genblk1.mmu.r_writeable_d[10] ;
 wire \cpu.genblk1.mmu.r_writeable_d[11] ;
 wire \cpu.genblk1.mmu.r_writeable_d[12] ;
 wire \cpu.genblk1.mmu.r_writeable_d[13] ;
 wire \cpu.genblk1.mmu.r_writeable_d[14] ;
 wire \cpu.genblk1.mmu.r_writeable_d[15] ;
 wire \cpu.genblk1.mmu.r_writeable_d[16] ;
 wire \cpu.genblk1.mmu.r_writeable_d[17] ;
 wire \cpu.genblk1.mmu.r_writeable_d[18] ;
 wire \cpu.genblk1.mmu.r_writeable_d[19] ;
 wire \cpu.genblk1.mmu.r_writeable_d[1] ;
 wire \cpu.genblk1.mmu.r_writeable_d[20] ;
 wire \cpu.genblk1.mmu.r_writeable_d[21] ;
 wire \cpu.genblk1.mmu.r_writeable_d[22] ;
 wire \cpu.genblk1.mmu.r_writeable_d[23] ;
 wire \cpu.genblk1.mmu.r_writeable_d[24] ;
 wire \cpu.genblk1.mmu.r_writeable_d[25] ;
 wire \cpu.genblk1.mmu.r_writeable_d[26] ;
 wire \cpu.genblk1.mmu.r_writeable_d[27] ;
 wire \cpu.genblk1.mmu.r_writeable_d[28] ;
 wire \cpu.genblk1.mmu.r_writeable_d[29] ;
 wire \cpu.genblk1.mmu.r_writeable_d[2] ;
 wire \cpu.genblk1.mmu.r_writeable_d[30] ;
 wire \cpu.genblk1.mmu.r_writeable_d[31] ;
 wire \cpu.genblk1.mmu.r_writeable_d[3] ;
 wire \cpu.genblk1.mmu.r_writeable_d[4] ;
 wire \cpu.genblk1.mmu.r_writeable_d[5] ;
 wire \cpu.genblk1.mmu.r_writeable_d[6] ;
 wire \cpu.genblk1.mmu.r_writeable_d[7] ;
 wire \cpu.genblk1.mmu.r_writeable_d[8] ;
 wire \cpu.genblk1.mmu.r_writeable_d[9] ;
 wire \cpu.gpio.genblk1[3].srcs_o[0] ;
 wire \cpu.gpio.genblk1[3].srcs_o[11] ;
 wire \cpu.gpio.genblk1[3].srcs_o[1] ;
 wire \cpu.gpio.genblk1[3].srcs_o[2] ;
 wire \cpu.gpio.genblk1[3].srcs_o[3] ;
 wire \cpu.gpio.genblk1[3].srcs_o[4] ;
 wire \cpu.gpio.genblk1[3].srcs_o[5] ;
 wire \cpu.gpio.genblk1[3].srcs_o[6] ;
 wire \cpu.gpio.genblk1[3].srcs_o[7] ;
 wire \cpu.gpio.genblk1[3].srcs_o[8] ;
 wire \cpu.gpio.genblk1[4].srcs_o[0] ;
 wire \cpu.gpio.genblk1[5].srcs_o[0] ;
 wire \cpu.gpio.genblk1[6].srcs_o[0] ;
 wire \cpu.gpio.genblk1[7].srcs_o[0] ;
 wire \cpu.gpio.genblk2[4].srcs_io[0] ;
 wire \cpu.gpio.genblk2[5].srcs_io[0] ;
 wire \cpu.gpio.genblk2[6].srcs_io[0] ;
 wire \cpu.gpio.genblk2[7].srcs_io[0] ;
 wire \cpu.gpio.r_enable_in[0] ;
 wire \cpu.gpio.r_enable_in[1] ;
 wire \cpu.gpio.r_enable_in[2] ;
 wire \cpu.gpio.r_enable_in[3] ;
 wire \cpu.gpio.r_enable_in[4] ;
 wire \cpu.gpio.r_enable_in[5] ;
 wire \cpu.gpio.r_enable_in[6] ;
 wire \cpu.gpio.r_enable_in[7] ;
 wire \cpu.gpio.r_enable_io[4] ;
 wire \cpu.gpio.r_enable_io[5] ;
 wire \cpu.gpio.r_enable_io[6] ;
 wire \cpu.gpio.r_enable_io[7] ;
 wire \cpu.gpio.r_spi_miso_src[0][0] ;
 wire \cpu.gpio.r_spi_miso_src[0][1] ;
 wire \cpu.gpio.r_spi_miso_src[0][2] ;
 wire \cpu.gpio.r_spi_miso_src[0][3] ;
 wire \cpu.gpio.r_spi_miso_src[1][0] ;
 wire \cpu.gpio.r_spi_miso_src[1][1] ;
 wire \cpu.gpio.r_spi_miso_src[1][2] ;
 wire \cpu.gpio.r_spi_miso_src[1][3] ;
 wire \cpu.gpio.r_src_io[4][0] ;
 wire \cpu.gpio.r_src_io[4][1] ;
 wire \cpu.gpio.r_src_io[4][2] ;
 wire \cpu.gpio.r_src_io[4][3] ;
 wire \cpu.gpio.r_src_io[5][0] ;
 wire \cpu.gpio.r_src_io[5][1] ;
 wire \cpu.gpio.r_src_io[5][2] ;
 wire \cpu.gpio.r_src_io[5][3] ;
 wire \cpu.gpio.r_src_io[6][0] ;
 wire \cpu.gpio.r_src_io[6][1] ;
 wire \cpu.gpio.r_src_io[6][2] ;
 wire \cpu.gpio.r_src_io[6][3] ;
 wire \cpu.gpio.r_src_io[7][0] ;
 wire \cpu.gpio.r_src_io[7][1] ;
 wire \cpu.gpio.r_src_io[7][2] ;
 wire \cpu.gpio.r_src_io[7][3] ;
 wire \cpu.gpio.r_src_o[3][0] ;
 wire \cpu.gpio.r_src_o[3][1] ;
 wire \cpu.gpio.r_src_o[3][2] ;
 wire \cpu.gpio.r_src_o[3][3] ;
 wire \cpu.gpio.r_src_o[4][0] ;
 wire \cpu.gpio.r_src_o[4][1] ;
 wire \cpu.gpio.r_src_o[4][2] ;
 wire \cpu.gpio.r_src_o[4][3] ;
 wire \cpu.gpio.r_src_o[5][0] ;
 wire \cpu.gpio.r_src_o[5][1] ;
 wire \cpu.gpio.r_src_o[5][2] ;
 wire \cpu.gpio.r_src_o[5][3] ;
 wire \cpu.gpio.r_src_o[6][0] ;
 wire \cpu.gpio.r_src_o[6][1] ;
 wire \cpu.gpio.r_src_o[6][2] ;
 wire \cpu.gpio.r_src_o[6][3] ;
 wire \cpu.gpio.r_src_o[7][0] ;
 wire \cpu.gpio.r_src_o[7][1] ;
 wire \cpu.gpio.r_src_o[7][2] ;
 wire \cpu.gpio.r_src_o[7][3] ;
 wire \cpu.gpio.r_uart_rx_src[0] ;
 wire \cpu.gpio.r_uart_rx_src[1] ;
 wire \cpu.gpio.r_uart_rx_src[2] ;
 wire \cpu.gpio.uart_rx ;
 wire \cpu.i_wstrobe_d ;
 wire \cpu.icache.r_data[0][0] ;
 wire \cpu.icache.r_data[0][10] ;
 wire \cpu.icache.r_data[0][11] ;
 wire \cpu.icache.r_data[0][12] ;
 wire \cpu.icache.r_data[0][13] ;
 wire \cpu.icache.r_data[0][14] ;
 wire \cpu.icache.r_data[0][15] ;
 wire \cpu.icache.r_data[0][16] ;
 wire \cpu.icache.r_data[0][17] ;
 wire \cpu.icache.r_data[0][18] ;
 wire \cpu.icache.r_data[0][19] ;
 wire \cpu.icache.r_data[0][1] ;
 wire \cpu.icache.r_data[0][20] ;
 wire \cpu.icache.r_data[0][21] ;
 wire \cpu.icache.r_data[0][22] ;
 wire \cpu.icache.r_data[0][23] ;
 wire \cpu.icache.r_data[0][24] ;
 wire \cpu.icache.r_data[0][25] ;
 wire \cpu.icache.r_data[0][26] ;
 wire \cpu.icache.r_data[0][27] ;
 wire \cpu.icache.r_data[0][28] ;
 wire \cpu.icache.r_data[0][29] ;
 wire \cpu.icache.r_data[0][2] ;
 wire \cpu.icache.r_data[0][30] ;
 wire \cpu.icache.r_data[0][31] ;
 wire \cpu.icache.r_data[0][3] ;
 wire \cpu.icache.r_data[0][4] ;
 wire \cpu.icache.r_data[0][5] ;
 wire \cpu.icache.r_data[0][6] ;
 wire \cpu.icache.r_data[0][7] ;
 wire \cpu.icache.r_data[0][8] ;
 wire \cpu.icache.r_data[0][9] ;
 wire \cpu.icache.r_data[1][0] ;
 wire \cpu.icache.r_data[1][10] ;
 wire \cpu.icache.r_data[1][11] ;
 wire \cpu.icache.r_data[1][12] ;
 wire \cpu.icache.r_data[1][13] ;
 wire \cpu.icache.r_data[1][14] ;
 wire \cpu.icache.r_data[1][15] ;
 wire \cpu.icache.r_data[1][16] ;
 wire \cpu.icache.r_data[1][17] ;
 wire \cpu.icache.r_data[1][18] ;
 wire \cpu.icache.r_data[1][19] ;
 wire \cpu.icache.r_data[1][1] ;
 wire \cpu.icache.r_data[1][20] ;
 wire \cpu.icache.r_data[1][21] ;
 wire \cpu.icache.r_data[1][22] ;
 wire \cpu.icache.r_data[1][23] ;
 wire \cpu.icache.r_data[1][24] ;
 wire \cpu.icache.r_data[1][25] ;
 wire \cpu.icache.r_data[1][26] ;
 wire \cpu.icache.r_data[1][27] ;
 wire \cpu.icache.r_data[1][28] ;
 wire \cpu.icache.r_data[1][29] ;
 wire \cpu.icache.r_data[1][2] ;
 wire \cpu.icache.r_data[1][30] ;
 wire \cpu.icache.r_data[1][31] ;
 wire \cpu.icache.r_data[1][3] ;
 wire \cpu.icache.r_data[1][4] ;
 wire \cpu.icache.r_data[1][5] ;
 wire \cpu.icache.r_data[1][6] ;
 wire \cpu.icache.r_data[1][7] ;
 wire \cpu.icache.r_data[1][8] ;
 wire \cpu.icache.r_data[1][9] ;
 wire \cpu.icache.r_data[2][0] ;
 wire \cpu.icache.r_data[2][10] ;
 wire \cpu.icache.r_data[2][11] ;
 wire \cpu.icache.r_data[2][12] ;
 wire \cpu.icache.r_data[2][13] ;
 wire \cpu.icache.r_data[2][14] ;
 wire \cpu.icache.r_data[2][15] ;
 wire \cpu.icache.r_data[2][16] ;
 wire \cpu.icache.r_data[2][17] ;
 wire \cpu.icache.r_data[2][18] ;
 wire \cpu.icache.r_data[2][19] ;
 wire \cpu.icache.r_data[2][1] ;
 wire \cpu.icache.r_data[2][20] ;
 wire \cpu.icache.r_data[2][21] ;
 wire \cpu.icache.r_data[2][22] ;
 wire \cpu.icache.r_data[2][23] ;
 wire \cpu.icache.r_data[2][24] ;
 wire \cpu.icache.r_data[2][25] ;
 wire \cpu.icache.r_data[2][26] ;
 wire \cpu.icache.r_data[2][27] ;
 wire \cpu.icache.r_data[2][28] ;
 wire \cpu.icache.r_data[2][29] ;
 wire \cpu.icache.r_data[2][2] ;
 wire \cpu.icache.r_data[2][30] ;
 wire \cpu.icache.r_data[2][31] ;
 wire \cpu.icache.r_data[2][3] ;
 wire \cpu.icache.r_data[2][4] ;
 wire \cpu.icache.r_data[2][5] ;
 wire \cpu.icache.r_data[2][6] ;
 wire \cpu.icache.r_data[2][7] ;
 wire \cpu.icache.r_data[2][8] ;
 wire \cpu.icache.r_data[2][9] ;
 wire \cpu.icache.r_data[3][0] ;
 wire \cpu.icache.r_data[3][10] ;
 wire \cpu.icache.r_data[3][11] ;
 wire \cpu.icache.r_data[3][12] ;
 wire \cpu.icache.r_data[3][13] ;
 wire \cpu.icache.r_data[3][14] ;
 wire \cpu.icache.r_data[3][15] ;
 wire \cpu.icache.r_data[3][16] ;
 wire \cpu.icache.r_data[3][17] ;
 wire \cpu.icache.r_data[3][18] ;
 wire \cpu.icache.r_data[3][19] ;
 wire \cpu.icache.r_data[3][1] ;
 wire \cpu.icache.r_data[3][20] ;
 wire \cpu.icache.r_data[3][21] ;
 wire \cpu.icache.r_data[3][22] ;
 wire \cpu.icache.r_data[3][23] ;
 wire \cpu.icache.r_data[3][24] ;
 wire \cpu.icache.r_data[3][25] ;
 wire \cpu.icache.r_data[3][26] ;
 wire \cpu.icache.r_data[3][27] ;
 wire \cpu.icache.r_data[3][28] ;
 wire \cpu.icache.r_data[3][29] ;
 wire \cpu.icache.r_data[3][2] ;
 wire \cpu.icache.r_data[3][30] ;
 wire \cpu.icache.r_data[3][31] ;
 wire \cpu.icache.r_data[3][3] ;
 wire \cpu.icache.r_data[3][4] ;
 wire \cpu.icache.r_data[3][5] ;
 wire \cpu.icache.r_data[3][6] ;
 wire \cpu.icache.r_data[3][7] ;
 wire \cpu.icache.r_data[3][8] ;
 wire \cpu.icache.r_data[3][9] ;
 wire \cpu.icache.r_data[4][0] ;
 wire \cpu.icache.r_data[4][10] ;
 wire \cpu.icache.r_data[4][11] ;
 wire \cpu.icache.r_data[4][12] ;
 wire \cpu.icache.r_data[4][13] ;
 wire \cpu.icache.r_data[4][14] ;
 wire \cpu.icache.r_data[4][15] ;
 wire \cpu.icache.r_data[4][16] ;
 wire \cpu.icache.r_data[4][17] ;
 wire \cpu.icache.r_data[4][18] ;
 wire \cpu.icache.r_data[4][19] ;
 wire \cpu.icache.r_data[4][1] ;
 wire \cpu.icache.r_data[4][20] ;
 wire \cpu.icache.r_data[4][21] ;
 wire \cpu.icache.r_data[4][22] ;
 wire \cpu.icache.r_data[4][23] ;
 wire \cpu.icache.r_data[4][24] ;
 wire \cpu.icache.r_data[4][25] ;
 wire \cpu.icache.r_data[4][26] ;
 wire \cpu.icache.r_data[4][27] ;
 wire \cpu.icache.r_data[4][28] ;
 wire \cpu.icache.r_data[4][29] ;
 wire \cpu.icache.r_data[4][2] ;
 wire \cpu.icache.r_data[4][30] ;
 wire \cpu.icache.r_data[4][31] ;
 wire \cpu.icache.r_data[4][3] ;
 wire \cpu.icache.r_data[4][4] ;
 wire \cpu.icache.r_data[4][5] ;
 wire \cpu.icache.r_data[4][6] ;
 wire \cpu.icache.r_data[4][7] ;
 wire \cpu.icache.r_data[4][8] ;
 wire \cpu.icache.r_data[4][9] ;
 wire \cpu.icache.r_data[5][0] ;
 wire \cpu.icache.r_data[5][10] ;
 wire \cpu.icache.r_data[5][11] ;
 wire \cpu.icache.r_data[5][12] ;
 wire \cpu.icache.r_data[5][13] ;
 wire \cpu.icache.r_data[5][14] ;
 wire \cpu.icache.r_data[5][15] ;
 wire \cpu.icache.r_data[5][16] ;
 wire \cpu.icache.r_data[5][17] ;
 wire \cpu.icache.r_data[5][18] ;
 wire \cpu.icache.r_data[5][19] ;
 wire \cpu.icache.r_data[5][1] ;
 wire \cpu.icache.r_data[5][20] ;
 wire \cpu.icache.r_data[5][21] ;
 wire \cpu.icache.r_data[5][22] ;
 wire \cpu.icache.r_data[5][23] ;
 wire \cpu.icache.r_data[5][24] ;
 wire \cpu.icache.r_data[5][25] ;
 wire \cpu.icache.r_data[5][26] ;
 wire \cpu.icache.r_data[5][27] ;
 wire \cpu.icache.r_data[5][28] ;
 wire \cpu.icache.r_data[5][29] ;
 wire \cpu.icache.r_data[5][2] ;
 wire \cpu.icache.r_data[5][30] ;
 wire \cpu.icache.r_data[5][31] ;
 wire \cpu.icache.r_data[5][3] ;
 wire \cpu.icache.r_data[5][4] ;
 wire \cpu.icache.r_data[5][5] ;
 wire \cpu.icache.r_data[5][6] ;
 wire \cpu.icache.r_data[5][7] ;
 wire \cpu.icache.r_data[5][8] ;
 wire \cpu.icache.r_data[5][9] ;
 wire \cpu.icache.r_data[6][0] ;
 wire \cpu.icache.r_data[6][10] ;
 wire \cpu.icache.r_data[6][11] ;
 wire \cpu.icache.r_data[6][12] ;
 wire \cpu.icache.r_data[6][13] ;
 wire \cpu.icache.r_data[6][14] ;
 wire \cpu.icache.r_data[6][15] ;
 wire \cpu.icache.r_data[6][16] ;
 wire \cpu.icache.r_data[6][17] ;
 wire \cpu.icache.r_data[6][18] ;
 wire \cpu.icache.r_data[6][19] ;
 wire \cpu.icache.r_data[6][1] ;
 wire \cpu.icache.r_data[6][20] ;
 wire \cpu.icache.r_data[6][21] ;
 wire \cpu.icache.r_data[6][22] ;
 wire \cpu.icache.r_data[6][23] ;
 wire \cpu.icache.r_data[6][24] ;
 wire \cpu.icache.r_data[6][25] ;
 wire \cpu.icache.r_data[6][26] ;
 wire \cpu.icache.r_data[6][27] ;
 wire \cpu.icache.r_data[6][28] ;
 wire \cpu.icache.r_data[6][29] ;
 wire \cpu.icache.r_data[6][2] ;
 wire \cpu.icache.r_data[6][30] ;
 wire \cpu.icache.r_data[6][31] ;
 wire \cpu.icache.r_data[6][3] ;
 wire \cpu.icache.r_data[6][4] ;
 wire \cpu.icache.r_data[6][5] ;
 wire \cpu.icache.r_data[6][6] ;
 wire \cpu.icache.r_data[6][7] ;
 wire \cpu.icache.r_data[6][8] ;
 wire \cpu.icache.r_data[6][9] ;
 wire \cpu.icache.r_data[7][0] ;
 wire \cpu.icache.r_data[7][10] ;
 wire \cpu.icache.r_data[7][11] ;
 wire \cpu.icache.r_data[7][12] ;
 wire \cpu.icache.r_data[7][13] ;
 wire \cpu.icache.r_data[7][14] ;
 wire \cpu.icache.r_data[7][15] ;
 wire \cpu.icache.r_data[7][16] ;
 wire \cpu.icache.r_data[7][17] ;
 wire \cpu.icache.r_data[7][18] ;
 wire \cpu.icache.r_data[7][19] ;
 wire \cpu.icache.r_data[7][1] ;
 wire \cpu.icache.r_data[7][20] ;
 wire \cpu.icache.r_data[7][21] ;
 wire \cpu.icache.r_data[7][22] ;
 wire \cpu.icache.r_data[7][23] ;
 wire \cpu.icache.r_data[7][24] ;
 wire \cpu.icache.r_data[7][25] ;
 wire \cpu.icache.r_data[7][26] ;
 wire \cpu.icache.r_data[7][27] ;
 wire \cpu.icache.r_data[7][28] ;
 wire \cpu.icache.r_data[7][29] ;
 wire \cpu.icache.r_data[7][2] ;
 wire \cpu.icache.r_data[7][30] ;
 wire \cpu.icache.r_data[7][31] ;
 wire \cpu.icache.r_data[7][3] ;
 wire \cpu.icache.r_data[7][4] ;
 wire \cpu.icache.r_data[7][5] ;
 wire \cpu.icache.r_data[7][6] ;
 wire \cpu.icache.r_data[7][7] ;
 wire \cpu.icache.r_data[7][8] ;
 wire \cpu.icache.r_data[7][9] ;
 wire \cpu.icache.r_offset[0] ;
 wire \cpu.icache.r_offset[1] ;
 wire \cpu.icache.r_offset[2] ;
 wire \cpu.icache.r_tag[0][10] ;
 wire \cpu.icache.r_tag[0][11] ;
 wire \cpu.icache.r_tag[0][12] ;
 wire \cpu.icache.r_tag[0][13] ;
 wire \cpu.icache.r_tag[0][14] ;
 wire \cpu.icache.r_tag[0][15] ;
 wire \cpu.icache.r_tag[0][16] ;
 wire \cpu.icache.r_tag[0][17] ;
 wire \cpu.icache.r_tag[0][18] ;
 wire \cpu.icache.r_tag[0][19] ;
 wire \cpu.icache.r_tag[0][20] ;
 wire \cpu.icache.r_tag[0][21] ;
 wire \cpu.icache.r_tag[0][22] ;
 wire \cpu.icache.r_tag[0][23] ;
 wire \cpu.icache.r_tag[0][5] ;
 wire \cpu.icache.r_tag[0][6] ;
 wire \cpu.icache.r_tag[0][7] ;
 wire \cpu.icache.r_tag[0][8] ;
 wire \cpu.icache.r_tag[0][9] ;
 wire \cpu.icache.r_tag[1][10] ;
 wire \cpu.icache.r_tag[1][11] ;
 wire \cpu.icache.r_tag[1][12] ;
 wire \cpu.icache.r_tag[1][13] ;
 wire \cpu.icache.r_tag[1][14] ;
 wire \cpu.icache.r_tag[1][15] ;
 wire \cpu.icache.r_tag[1][16] ;
 wire \cpu.icache.r_tag[1][17] ;
 wire \cpu.icache.r_tag[1][18] ;
 wire \cpu.icache.r_tag[1][19] ;
 wire \cpu.icache.r_tag[1][20] ;
 wire \cpu.icache.r_tag[1][21] ;
 wire \cpu.icache.r_tag[1][22] ;
 wire \cpu.icache.r_tag[1][23] ;
 wire \cpu.icache.r_tag[1][5] ;
 wire \cpu.icache.r_tag[1][6] ;
 wire \cpu.icache.r_tag[1][7] ;
 wire \cpu.icache.r_tag[1][8] ;
 wire \cpu.icache.r_tag[1][9] ;
 wire \cpu.icache.r_tag[2][10] ;
 wire \cpu.icache.r_tag[2][11] ;
 wire \cpu.icache.r_tag[2][12] ;
 wire \cpu.icache.r_tag[2][13] ;
 wire \cpu.icache.r_tag[2][14] ;
 wire \cpu.icache.r_tag[2][15] ;
 wire \cpu.icache.r_tag[2][16] ;
 wire \cpu.icache.r_tag[2][17] ;
 wire \cpu.icache.r_tag[2][18] ;
 wire \cpu.icache.r_tag[2][19] ;
 wire \cpu.icache.r_tag[2][20] ;
 wire \cpu.icache.r_tag[2][21] ;
 wire \cpu.icache.r_tag[2][22] ;
 wire \cpu.icache.r_tag[2][23] ;
 wire \cpu.icache.r_tag[2][5] ;
 wire \cpu.icache.r_tag[2][6] ;
 wire \cpu.icache.r_tag[2][7] ;
 wire \cpu.icache.r_tag[2][8] ;
 wire \cpu.icache.r_tag[2][9] ;
 wire \cpu.icache.r_tag[3][10] ;
 wire \cpu.icache.r_tag[3][11] ;
 wire \cpu.icache.r_tag[3][12] ;
 wire \cpu.icache.r_tag[3][13] ;
 wire \cpu.icache.r_tag[3][14] ;
 wire \cpu.icache.r_tag[3][15] ;
 wire \cpu.icache.r_tag[3][16] ;
 wire \cpu.icache.r_tag[3][17] ;
 wire \cpu.icache.r_tag[3][18] ;
 wire \cpu.icache.r_tag[3][19] ;
 wire \cpu.icache.r_tag[3][20] ;
 wire \cpu.icache.r_tag[3][21] ;
 wire \cpu.icache.r_tag[3][22] ;
 wire \cpu.icache.r_tag[3][23] ;
 wire \cpu.icache.r_tag[3][5] ;
 wire \cpu.icache.r_tag[3][6] ;
 wire \cpu.icache.r_tag[3][7] ;
 wire \cpu.icache.r_tag[3][8] ;
 wire \cpu.icache.r_tag[3][9] ;
 wire \cpu.icache.r_tag[4][10] ;
 wire \cpu.icache.r_tag[4][11] ;
 wire \cpu.icache.r_tag[4][12] ;
 wire \cpu.icache.r_tag[4][13] ;
 wire \cpu.icache.r_tag[4][14] ;
 wire \cpu.icache.r_tag[4][15] ;
 wire \cpu.icache.r_tag[4][16] ;
 wire \cpu.icache.r_tag[4][17] ;
 wire \cpu.icache.r_tag[4][18] ;
 wire \cpu.icache.r_tag[4][19] ;
 wire \cpu.icache.r_tag[4][20] ;
 wire \cpu.icache.r_tag[4][21] ;
 wire \cpu.icache.r_tag[4][22] ;
 wire \cpu.icache.r_tag[4][23] ;
 wire \cpu.icache.r_tag[4][5] ;
 wire \cpu.icache.r_tag[4][6] ;
 wire \cpu.icache.r_tag[4][7] ;
 wire \cpu.icache.r_tag[4][8] ;
 wire \cpu.icache.r_tag[4][9] ;
 wire \cpu.icache.r_tag[5][10] ;
 wire \cpu.icache.r_tag[5][11] ;
 wire \cpu.icache.r_tag[5][12] ;
 wire \cpu.icache.r_tag[5][13] ;
 wire \cpu.icache.r_tag[5][14] ;
 wire \cpu.icache.r_tag[5][15] ;
 wire \cpu.icache.r_tag[5][16] ;
 wire \cpu.icache.r_tag[5][17] ;
 wire \cpu.icache.r_tag[5][18] ;
 wire \cpu.icache.r_tag[5][19] ;
 wire \cpu.icache.r_tag[5][20] ;
 wire \cpu.icache.r_tag[5][21] ;
 wire \cpu.icache.r_tag[5][22] ;
 wire \cpu.icache.r_tag[5][23] ;
 wire \cpu.icache.r_tag[5][5] ;
 wire \cpu.icache.r_tag[5][6] ;
 wire \cpu.icache.r_tag[5][7] ;
 wire \cpu.icache.r_tag[5][8] ;
 wire \cpu.icache.r_tag[5][9] ;
 wire \cpu.icache.r_tag[6][10] ;
 wire \cpu.icache.r_tag[6][11] ;
 wire \cpu.icache.r_tag[6][12] ;
 wire \cpu.icache.r_tag[6][13] ;
 wire \cpu.icache.r_tag[6][14] ;
 wire \cpu.icache.r_tag[6][15] ;
 wire \cpu.icache.r_tag[6][16] ;
 wire \cpu.icache.r_tag[6][17] ;
 wire \cpu.icache.r_tag[6][18] ;
 wire \cpu.icache.r_tag[6][19] ;
 wire \cpu.icache.r_tag[6][20] ;
 wire \cpu.icache.r_tag[6][21] ;
 wire \cpu.icache.r_tag[6][22] ;
 wire \cpu.icache.r_tag[6][23] ;
 wire \cpu.icache.r_tag[6][5] ;
 wire \cpu.icache.r_tag[6][6] ;
 wire \cpu.icache.r_tag[6][7] ;
 wire \cpu.icache.r_tag[6][8] ;
 wire \cpu.icache.r_tag[6][9] ;
 wire \cpu.icache.r_tag[7][10] ;
 wire \cpu.icache.r_tag[7][11] ;
 wire \cpu.icache.r_tag[7][12] ;
 wire \cpu.icache.r_tag[7][13] ;
 wire \cpu.icache.r_tag[7][14] ;
 wire \cpu.icache.r_tag[7][15] ;
 wire \cpu.icache.r_tag[7][16] ;
 wire \cpu.icache.r_tag[7][17] ;
 wire \cpu.icache.r_tag[7][18] ;
 wire \cpu.icache.r_tag[7][19] ;
 wire \cpu.icache.r_tag[7][20] ;
 wire \cpu.icache.r_tag[7][21] ;
 wire \cpu.icache.r_tag[7][22] ;
 wire \cpu.icache.r_tag[7][23] ;
 wire \cpu.icache.r_tag[7][5] ;
 wire \cpu.icache.r_tag[7][6] ;
 wire \cpu.icache.r_tag[7][7] ;
 wire \cpu.icache.r_tag[7][8] ;
 wire \cpu.icache.r_tag[7][9] ;
 wire \cpu.icache.r_valid[0] ;
 wire \cpu.icache.r_valid[1] ;
 wire \cpu.icache.r_valid[2] ;
 wire \cpu.icache.r_valid[3] ;
 wire \cpu.icache.r_valid[4] ;
 wire \cpu.icache.r_valid[5] ;
 wire \cpu.icache.r_valid[6] ;
 wire \cpu.icache.r_valid[7] ;
 wire \cpu.intr.r_clock ;
 wire \cpu.intr.r_clock_cmp[0] ;
 wire \cpu.intr.r_clock_cmp[10] ;
 wire \cpu.intr.r_clock_cmp[11] ;
 wire \cpu.intr.r_clock_cmp[12] ;
 wire \cpu.intr.r_clock_cmp[13] ;
 wire \cpu.intr.r_clock_cmp[14] ;
 wire \cpu.intr.r_clock_cmp[15] ;
 wire \cpu.intr.r_clock_cmp[16] ;
 wire \cpu.intr.r_clock_cmp[17] ;
 wire \cpu.intr.r_clock_cmp[18] ;
 wire \cpu.intr.r_clock_cmp[19] ;
 wire \cpu.intr.r_clock_cmp[1] ;
 wire \cpu.intr.r_clock_cmp[20] ;
 wire \cpu.intr.r_clock_cmp[21] ;
 wire \cpu.intr.r_clock_cmp[22] ;
 wire \cpu.intr.r_clock_cmp[23] ;
 wire \cpu.intr.r_clock_cmp[24] ;
 wire \cpu.intr.r_clock_cmp[25] ;
 wire \cpu.intr.r_clock_cmp[26] ;
 wire \cpu.intr.r_clock_cmp[27] ;
 wire \cpu.intr.r_clock_cmp[28] ;
 wire \cpu.intr.r_clock_cmp[29] ;
 wire \cpu.intr.r_clock_cmp[2] ;
 wire \cpu.intr.r_clock_cmp[30] ;
 wire \cpu.intr.r_clock_cmp[31] ;
 wire \cpu.intr.r_clock_cmp[3] ;
 wire \cpu.intr.r_clock_cmp[4] ;
 wire \cpu.intr.r_clock_cmp[5] ;
 wire \cpu.intr.r_clock_cmp[6] ;
 wire \cpu.intr.r_clock_cmp[7] ;
 wire \cpu.intr.r_clock_cmp[8] ;
 wire \cpu.intr.r_clock_cmp[9] ;
 wire \cpu.intr.r_clock_count[0] ;
 wire \cpu.intr.r_clock_count[10] ;
 wire \cpu.intr.r_clock_count[11] ;
 wire \cpu.intr.r_clock_count[12] ;
 wire \cpu.intr.r_clock_count[13] ;
 wire \cpu.intr.r_clock_count[14] ;
 wire \cpu.intr.r_clock_count[15] ;
 wire \cpu.intr.r_clock_count[16] ;
 wire \cpu.intr.r_clock_count[17] ;
 wire \cpu.intr.r_clock_count[18] ;
 wire \cpu.intr.r_clock_count[19] ;
 wire \cpu.intr.r_clock_count[1] ;
 wire \cpu.intr.r_clock_count[20] ;
 wire \cpu.intr.r_clock_count[21] ;
 wire \cpu.intr.r_clock_count[22] ;
 wire \cpu.intr.r_clock_count[23] ;
 wire \cpu.intr.r_clock_count[24] ;
 wire \cpu.intr.r_clock_count[25] ;
 wire \cpu.intr.r_clock_count[26] ;
 wire \cpu.intr.r_clock_count[27] ;
 wire \cpu.intr.r_clock_count[28] ;
 wire \cpu.intr.r_clock_count[29] ;
 wire \cpu.intr.r_clock_count[2] ;
 wire \cpu.intr.r_clock_count[30] ;
 wire \cpu.intr.r_clock_count[31] ;
 wire \cpu.intr.r_clock_count[3] ;
 wire \cpu.intr.r_clock_count[4] ;
 wire \cpu.intr.r_clock_count[5] ;
 wire \cpu.intr.r_clock_count[6] ;
 wire \cpu.intr.r_clock_count[7] ;
 wire \cpu.intr.r_clock_count[8] ;
 wire \cpu.intr.r_clock_count[9] ;
 wire \cpu.intr.r_enable[0] ;
 wire \cpu.intr.r_enable[1] ;
 wire \cpu.intr.r_enable[2] ;
 wire \cpu.intr.r_enable[3] ;
 wire \cpu.intr.r_enable[4] ;
 wire \cpu.intr.r_enable[5] ;
 wire \cpu.intr.r_swi ;
 wire \cpu.intr.r_timer ;
 wire \cpu.intr.r_timer_count[0] ;
 wire \cpu.intr.r_timer_count[10] ;
 wire \cpu.intr.r_timer_count[11] ;
 wire \cpu.intr.r_timer_count[12] ;
 wire \cpu.intr.r_timer_count[13] ;
 wire \cpu.intr.r_timer_count[14] ;
 wire \cpu.intr.r_timer_count[15] ;
 wire \cpu.intr.r_timer_count[16] ;
 wire \cpu.intr.r_timer_count[17] ;
 wire \cpu.intr.r_timer_count[18] ;
 wire \cpu.intr.r_timer_count[19] ;
 wire \cpu.intr.r_timer_count[1] ;
 wire \cpu.intr.r_timer_count[20] ;
 wire \cpu.intr.r_timer_count[21] ;
 wire \cpu.intr.r_timer_count[22] ;
 wire \cpu.intr.r_timer_count[23] ;
 wire \cpu.intr.r_timer_count[2] ;
 wire \cpu.intr.r_timer_count[3] ;
 wire \cpu.intr.r_timer_count[4] ;
 wire \cpu.intr.r_timer_count[5] ;
 wire \cpu.intr.r_timer_count[6] ;
 wire \cpu.intr.r_timer_count[7] ;
 wire \cpu.intr.r_timer_count[8] ;
 wire \cpu.intr.r_timer_count[9] ;
 wire \cpu.intr.r_timer_reload[0] ;
 wire \cpu.intr.r_timer_reload[10] ;
 wire \cpu.intr.r_timer_reload[11] ;
 wire \cpu.intr.r_timer_reload[12] ;
 wire \cpu.intr.r_timer_reload[13] ;
 wire \cpu.intr.r_timer_reload[14] ;
 wire \cpu.intr.r_timer_reload[15] ;
 wire \cpu.intr.r_timer_reload[16] ;
 wire \cpu.intr.r_timer_reload[17] ;
 wire \cpu.intr.r_timer_reload[18] ;
 wire \cpu.intr.r_timer_reload[19] ;
 wire \cpu.intr.r_timer_reload[1] ;
 wire \cpu.intr.r_timer_reload[20] ;
 wire \cpu.intr.r_timer_reload[21] ;
 wire \cpu.intr.r_timer_reload[22] ;
 wire \cpu.intr.r_timer_reload[23] ;
 wire \cpu.intr.r_timer_reload[2] ;
 wire \cpu.intr.r_timer_reload[3] ;
 wire \cpu.intr.r_timer_reload[4] ;
 wire \cpu.intr.r_timer_reload[5] ;
 wire \cpu.intr.r_timer_reload[6] ;
 wire \cpu.intr.r_timer_reload[7] ;
 wire \cpu.intr.r_timer_reload[8] ;
 wire \cpu.intr.r_timer_reload[9] ;
 wire \cpu.intr.spi_intr ;
 wire \cpu.qspi.c_rstrobe_d ;
 wire \cpu.qspi.c_wstrobe_d ;
 wire \cpu.qspi.c_wstrobe_i ;
 wire \cpu.qspi.r_count[0] ;
 wire \cpu.qspi.r_count[1] ;
 wire \cpu.qspi.r_count[2] ;
 wire \cpu.qspi.r_count[3] ;
 wire \cpu.qspi.r_count[4] ;
 wire \cpu.qspi.r_ind ;
 wire \cpu.qspi.r_mask[0] ;
 wire \cpu.qspi.r_mask[1] ;
 wire \cpu.qspi.r_mask[2] ;
 wire \cpu.qspi.r_quad[0] ;
 wire \cpu.qspi.r_quad[1] ;
 wire \cpu.qspi.r_quad[2] ;
 wire \cpu.qspi.r_read_delay[0][0] ;
 wire \cpu.qspi.r_read_delay[0][1] ;
 wire \cpu.qspi.r_read_delay[0][2] ;
 wire \cpu.qspi.r_read_delay[0][3] ;
 wire \cpu.qspi.r_read_delay[1][0] ;
 wire \cpu.qspi.r_read_delay[1][1] ;
 wire \cpu.qspi.r_read_delay[1][2] ;
 wire \cpu.qspi.r_read_delay[1][3] ;
 wire \cpu.qspi.r_read_delay[2][0] ;
 wire \cpu.qspi.r_read_delay[2][1] ;
 wire \cpu.qspi.r_read_delay[2][2] ;
 wire \cpu.qspi.r_read_delay[2][3] ;
 wire \cpu.qspi.r_rom_mode[0] ;
 wire \cpu.qspi.r_rom_mode[1] ;
 wire \cpu.qspi.r_state[0] ;
 wire \cpu.qspi.r_state[10] ;
 wire \cpu.qspi.r_state[11] ;
 wire \cpu.qspi.r_state[12] ;
 wire \cpu.qspi.r_state[13] ;
 wire \cpu.qspi.r_state[14] ;
 wire \cpu.qspi.r_state[15] ;
 wire \cpu.qspi.r_state[16] ;
 wire \cpu.qspi.r_state[17] ;
 wire \cpu.qspi.r_state[1] ;
 wire \cpu.qspi.r_state[2] ;
 wire \cpu.qspi.r_state[3] ;
 wire \cpu.qspi.r_state[4] ;
 wire \cpu.qspi.r_state[5] ;
 wire \cpu.qspi.r_state[6] ;
 wire \cpu.qspi.r_state[7] ;
 wire \cpu.qspi.r_state[8] ;
 wire \cpu.qspi.r_state[9] ;
 wire \cpu.r_clk_invert ;
 wire \cpu.spi.r_bits[0] ;
 wire \cpu.spi.r_bits[1] ;
 wire \cpu.spi.r_bits[2] ;
 wire \cpu.spi.r_clk_count[0][0] ;
 wire \cpu.spi.r_clk_count[0][1] ;
 wire \cpu.spi.r_clk_count[0][2] ;
 wire \cpu.spi.r_clk_count[0][3] ;
 wire \cpu.spi.r_clk_count[0][4] ;
 wire \cpu.spi.r_clk_count[0][5] ;
 wire \cpu.spi.r_clk_count[0][6] ;
 wire \cpu.spi.r_clk_count[0][7] ;
 wire \cpu.spi.r_clk_count[1][0] ;
 wire \cpu.spi.r_clk_count[1][1] ;
 wire \cpu.spi.r_clk_count[1][2] ;
 wire \cpu.spi.r_clk_count[1][3] ;
 wire \cpu.spi.r_clk_count[1][4] ;
 wire \cpu.spi.r_clk_count[1][5] ;
 wire \cpu.spi.r_clk_count[1][6] ;
 wire \cpu.spi.r_clk_count[1][7] ;
 wire \cpu.spi.r_clk_count[2][0] ;
 wire \cpu.spi.r_clk_count[2][1] ;
 wire \cpu.spi.r_clk_count[2][2] ;
 wire \cpu.spi.r_clk_count[2][3] ;
 wire \cpu.spi.r_clk_count[2][4] ;
 wire \cpu.spi.r_clk_count[2][5] ;
 wire \cpu.spi.r_clk_count[2][6] ;
 wire \cpu.spi.r_clk_count[2][7] ;
 wire \cpu.spi.r_count[0] ;
 wire \cpu.spi.r_count[1] ;
 wire \cpu.spi.r_count[2] ;
 wire \cpu.spi.r_count[3] ;
 wire \cpu.spi.r_count[4] ;
 wire \cpu.spi.r_count[5] ;
 wire \cpu.spi.r_count[6] ;
 wire \cpu.spi.r_count[7] ;
 wire \cpu.spi.r_in[0] ;
 wire \cpu.spi.r_in[1] ;
 wire \cpu.spi.r_in[2] ;
 wire \cpu.spi.r_in[3] ;
 wire \cpu.spi.r_in[4] ;
 wire \cpu.spi.r_in[5] ;
 wire \cpu.spi.r_in[6] ;
 wire \cpu.spi.r_in[7] ;
 wire \cpu.spi.r_mode[0][0] ;
 wire \cpu.spi.r_mode[0][1] ;
 wire \cpu.spi.r_mode[1][0] ;
 wire \cpu.spi.r_mode[1][1] ;
 wire \cpu.spi.r_mode[2][0] ;
 wire \cpu.spi.r_mode[2][1] ;
 wire \cpu.spi.r_out[0] ;
 wire \cpu.spi.r_out[1] ;
 wire \cpu.spi.r_out[2] ;
 wire \cpu.spi.r_out[3] ;
 wire \cpu.spi.r_out[4] ;
 wire \cpu.spi.r_out[5] ;
 wire \cpu.spi.r_out[6] ;
 wire \cpu.spi.r_out[7] ;
 wire \cpu.spi.r_ready ;
 wire \cpu.spi.r_searching ;
 wire \cpu.spi.r_sel[0] ;
 wire \cpu.spi.r_sel[1] ;
 wire \cpu.spi.r_src[0] ;
 wire \cpu.spi.r_src[1] ;
 wire \cpu.spi.r_src[2] ;
 wire \cpu.spi.r_state[0] ;
 wire \cpu.spi.r_state[1] ;
 wire \cpu.spi.r_state[2] ;
 wire \cpu.spi.r_state[3] ;
 wire \cpu.spi.r_state[4] ;
 wire \cpu.spi.r_state[5] ;
 wire \cpu.spi.r_state[6] ;
 wire \cpu.spi.r_timeout[0] ;
 wire \cpu.spi.r_timeout[1] ;
 wire \cpu.spi.r_timeout[2] ;
 wire \cpu.spi.r_timeout[3] ;
 wire \cpu.spi.r_timeout[4] ;
 wire \cpu.spi.r_timeout[5] ;
 wire \cpu.spi.r_timeout[6] ;
 wire \cpu.spi.r_timeout[7] ;
 wire \cpu.spi.r_timeout_count[0] ;
 wire \cpu.spi.r_timeout_count[1] ;
 wire \cpu.spi.r_timeout_count[2] ;
 wire \cpu.spi.r_timeout_count[3] ;
 wire \cpu.spi.r_timeout_count[4] ;
 wire \cpu.spi.r_timeout_count[5] ;
 wire \cpu.spi.r_timeout_count[6] ;
 wire \cpu.spi.r_timeout_count[7] ;
 wire \cpu.uart.r_div[0] ;
 wire \cpu.uart.r_div[10] ;
 wire \cpu.uart.r_div[11] ;
 wire \cpu.uart.r_div[1] ;
 wire \cpu.uart.r_div[2] ;
 wire \cpu.uart.r_div[3] ;
 wire \cpu.uart.r_div[4] ;
 wire \cpu.uart.r_div[5] ;
 wire \cpu.uart.r_div[6] ;
 wire \cpu.uart.r_div[7] ;
 wire \cpu.uart.r_div[8] ;
 wire \cpu.uart.r_div[9] ;
 wire \cpu.uart.r_div_value[0] ;
 wire \cpu.uart.r_div_value[10] ;
 wire \cpu.uart.r_div_value[11] ;
 wire \cpu.uart.r_div_value[1] ;
 wire \cpu.uart.r_div_value[2] ;
 wire \cpu.uart.r_div_value[3] ;
 wire \cpu.uart.r_div_value[4] ;
 wire \cpu.uart.r_div_value[5] ;
 wire \cpu.uart.r_div_value[6] ;
 wire \cpu.uart.r_div_value[7] ;
 wire \cpu.uart.r_div_value[8] ;
 wire \cpu.uart.r_div_value[9] ;
 wire \cpu.uart.r_ib[0] ;
 wire \cpu.uart.r_ib[1] ;
 wire \cpu.uart.r_ib[2] ;
 wire \cpu.uart.r_ib[3] ;
 wire \cpu.uart.r_ib[4] ;
 wire \cpu.uart.r_ib[5] ;
 wire \cpu.uart.r_ib[6] ;
 wire \cpu.uart.r_in[0] ;
 wire \cpu.uart.r_in[1] ;
 wire \cpu.uart.r_in[2] ;
 wire \cpu.uart.r_in[3] ;
 wire \cpu.uart.r_in[4] ;
 wire \cpu.uart.r_in[5] ;
 wire \cpu.uart.r_in[6] ;
 wire \cpu.uart.r_in[7] ;
 wire \cpu.uart.r_out[0] ;
 wire \cpu.uart.r_out[1] ;
 wire \cpu.uart.r_out[2] ;
 wire \cpu.uart.r_out[3] ;
 wire \cpu.uart.r_out[4] ;
 wire \cpu.uart.r_out[5] ;
 wire \cpu.uart.r_out[6] ;
 wire \cpu.uart.r_out[7] ;
 wire \cpu.uart.r_r ;
 wire \cpu.uart.r_r_int ;
 wire \cpu.uart.r_r_invert ;
 wire \cpu.uart.r_rcnt[0] ;
 wire \cpu.uart.r_rcnt[1] ;
 wire \cpu.uart.r_rstate[0] ;
 wire \cpu.uart.r_rstate[1] ;
 wire \cpu.uart.r_rstate[2] ;
 wire \cpu.uart.r_rstate[3] ;
 wire \cpu.uart.r_x_int ;
 wire \cpu.uart.r_x_invert ;
 wire \cpu.uart.r_xcnt[0] ;
 wire \cpu.uart.r_xcnt[1] ;
 wire \cpu.uart.r_xstate[0] ;
 wire \cpu.uart.r_xstate[1] ;
 wire \cpu.uart.r_xstate[2] ;
 wire \cpu.uart.r_xstate[3] ;
 wire r_reset;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_253_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_257_clk;
 wire clknet_leaf_258_clk;
 wire clknet_leaf_259_clk;
 wire clknet_leaf_260_clk;
 wire clknet_leaf_261_clk;
 wire clknet_leaf_262_clk;
 wire clknet_leaf_263_clk;
 wire clknet_leaf_264_clk;
 wire clknet_leaf_265_clk;
 wire clknet_leaf_266_clk;
 wire clknet_leaf_267_clk;
 wire clknet_leaf_268_clk;
 wire clknet_leaf_269_clk;
 wire clknet_leaf_270_clk;
 wire clknet_leaf_271_clk;
 wire clknet_leaf_272_clk;
 wire clknet_leaf_273_clk;
 wire clknet_leaf_274_clk;
 wire clknet_leaf_275_clk;
 wire clknet_leaf_276_clk;
 wire clknet_leaf_277_clk;
 wire clknet_leaf_278_clk;
 wire clknet_leaf_279_clk;
 wire clknet_leaf_280_clk;
 wire clknet_leaf_281_clk;
 wire clknet_leaf_282_clk;
 wire clknet_leaf_283_clk;
 wire clknet_leaf_284_clk;
 wire clknet_leaf_285_clk;
 wire clknet_leaf_286_clk;
 wire clknet_leaf_287_clk;
 wire clknet_leaf_288_clk;
 wire clknet_leaf_289_clk;
 wire clknet_leaf_290_clk;
 wire clknet_leaf_291_clk;
 wire clknet_leaf_292_clk;
 wire clknet_leaf_293_clk;
 wire clknet_leaf_294_clk;
 wire clknet_leaf_295_clk;
 wire clknet_leaf_296_clk;
 wire clknet_leaf_297_clk;
 wire clknet_leaf_298_clk;
 wire clknet_leaf_299_clk;
 wire clknet_leaf_300_clk;
 wire clknet_leaf_301_clk;
 wire clknet_leaf_302_clk;
 wire clknet_leaf_303_clk;
 wire clknet_leaf_304_clk;
 wire clknet_leaf_305_clk;
 wire clknet_leaf_306_clk;
 wire clknet_leaf_307_clk;
 wire clknet_leaf_308_clk;
 wire clknet_leaf_309_clk;
 wire clknet_leaf_310_clk;
 wire clknet_leaf_311_clk;
 wire clknet_leaf_312_clk;
 wire clknet_leaf_313_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_6_0__leaf_clk;
 wire clknet_6_1__leaf_clk;
 wire clknet_6_2__leaf_clk;
 wire clknet_6_3__leaf_clk;
 wire clknet_6_4__leaf_clk;
 wire clknet_6_5__leaf_clk;
 wire clknet_6_6__leaf_clk;
 wire clknet_6_7__leaf_clk;
 wire clknet_6_8__leaf_clk;
 wire clknet_6_9__leaf_clk;
 wire clknet_6_10__leaf_clk;
 wire clknet_6_11__leaf_clk;
 wire clknet_6_12__leaf_clk;
 wire clknet_6_13__leaf_clk;
 wire clknet_6_14__leaf_clk;
 wire clknet_6_15__leaf_clk;
 wire clknet_6_16__leaf_clk;
 wire clknet_6_17__leaf_clk;
 wire clknet_6_18__leaf_clk;
 wire clknet_6_19__leaf_clk;
 wire clknet_6_20__leaf_clk;
 wire clknet_6_21__leaf_clk;
 wire clknet_6_22__leaf_clk;
 wire clknet_6_23__leaf_clk;
 wire clknet_6_24__leaf_clk;
 wire clknet_6_25__leaf_clk;
 wire clknet_6_26__leaf_clk;
 wire clknet_6_27__leaf_clk;
 wire clknet_6_28__leaf_clk;
 wire clknet_6_29__leaf_clk;
 wire clknet_6_30__leaf_clk;
 wire clknet_6_31__leaf_clk;
 wire clknet_6_32__leaf_clk;
 wire clknet_6_33__leaf_clk;
 wire clknet_6_34__leaf_clk;
 wire clknet_6_35__leaf_clk;
 wire clknet_6_36__leaf_clk;
 wire clknet_6_37__leaf_clk;
 wire clknet_6_38__leaf_clk;
 wire clknet_6_39__leaf_clk;
 wire clknet_6_40__leaf_clk;
 wire clknet_6_41__leaf_clk;
 wire clknet_6_42__leaf_clk;
 wire clknet_6_43__leaf_clk;
 wire clknet_6_44__leaf_clk;
 wire clknet_6_45__leaf_clk;
 wire clknet_6_46__leaf_clk;
 wire clknet_6_47__leaf_clk;
 wire clknet_6_48__leaf_clk;
 wire clknet_6_49__leaf_clk;
 wire clknet_6_50__leaf_clk;
 wire clknet_6_51__leaf_clk;
 wire clknet_6_52__leaf_clk;
 wire clknet_6_53__leaf_clk;
 wire clknet_6_54__leaf_clk;
 wire clknet_6_55__leaf_clk;
 wire clknet_6_56__leaf_clk;
 wire clknet_6_57__leaf_clk;
 wire clknet_6_58__leaf_clk;
 wire clknet_6_59__leaf_clk;
 wire clknet_6_60__leaf_clk;
 wire clknet_6_61__leaf_clk;
 wire clknet_6_62__leaf_clk;
 wire clknet_6_63__leaf_clk;

 sg13g2_buf_1 _14932_ (.A(\cpu.dec.r_op[6] ),
    .X(_08121_));
 sg13g2_buf_1 _14933_ (.A(net1123),
    .X(_08122_));
 sg13g2_inv_1 _14934_ (.Y(_08123_),
    .A(_00173_));
 sg13g2_buf_1 _14935_ (.A(\cpu.ex.r_read_stall ),
    .X(_08124_));
 sg13g2_buf_2 _14936_ (.A(\cpu.ex.r_wmask[1] ),
    .X(_08125_));
 sg13g2_inv_2 _14937_ (.Y(_08126_),
    .A(_08125_));
 sg13g2_buf_2 _14938_ (.A(\cpu.ex.r_wmask[0] ),
    .X(_08127_));
 sg13g2_inv_2 _14939_ (.Y(_08128_),
    .A(_08127_));
 sg13g2_nand2_1 _14940_ (.Y(_08129_),
    .A(_08126_),
    .B(_08128_));
 sg13g2_nor3_1 _14941_ (.A(_08123_),
    .B(_08124_),
    .C(_08129_),
    .Y(_08130_));
 sg13g2_buf_2 _14942_ (.A(_08130_),
    .X(_08131_));
 sg13g2_buf_2 _14943_ (.A(_00177_),
    .X(_08132_));
 sg13g2_buf_2 _14944_ (.A(\cpu.ex.ifetch ),
    .X(_08133_));
 sg13g2_buf_2 _14945_ (.A(\cpu.ex.genblk3.r_mmu_d_proxy ),
    .X(_08134_));
 sg13g2_nor2b_1 _14946_ (.A(_08133_),
    .B_N(_08134_),
    .Y(_08135_));
 sg13g2_nor2_1 _14947_ (.A(_08132_),
    .B(_08135_),
    .Y(_08136_));
 sg13g2_buf_8 _14948_ (.A(\cpu.addr[12] ),
    .X(_08137_));
 sg13g2_buf_8 _14949_ (.A(_08137_),
    .X(_08138_));
 sg13g2_buf_8 _14950_ (.A(\cpu.addr[13] ),
    .X(_08139_));
 sg13g2_buf_8 _14951_ (.A(\cpu.addr[15] ),
    .X(_08140_));
 sg13g2_nor3_1 _14952_ (.A(net1062),
    .B(_08139_),
    .C(net1121),
    .Y(_08141_));
 sg13g2_buf_8 _14953_ (.A(\cpu.addr[14] ),
    .X(_08142_));
 sg13g2_buf_8 _14954_ (.A(net1120),
    .X(_08143_));
 sg13g2_mux2_1 _14955_ (.A0(\cpu.genblk1.mmu.r_valid_d[16] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[20] ),
    .S(net1061),
    .X(_08144_));
 sg13g2_nand2_1 _14956_ (.Y(_08145_),
    .A(_08141_),
    .B(_08144_));
 sg13g2_nor2_1 _14957_ (.A(_08139_),
    .B(net1121),
    .Y(_08146_));
 sg13g2_mux2_1 _14958_ (.A0(\cpu.genblk1.mmu.r_valid_d[17] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[21] ),
    .S(_08142_),
    .X(_08147_));
 sg13g2_nand3_1 _14959_ (.B(_08146_),
    .C(_08147_),
    .A(net1062),
    .Y(_08148_));
 sg13g2_nor2b_1 _14960_ (.A(net1121),
    .B_N(_08139_),
    .Y(_08149_));
 sg13g2_buf_8 _14961_ (.A(_08137_),
    .X(_08150_));
 sg13g2_mux4_1 _14962_ (.S0(net1060),
    .A0(\cpu.genblk1.mmu.r_valid_d[18] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[19] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[22] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[23] ),
    .S1(net1061),
    .X(_08151_));
 sg13g2_nand2_1 _14963_ (.Y(_08152_),
    .A(_08149_),
    .B(_08151_));
 sg13g2_nand4_1 _14964_ (.B(_08145_),
    .C(_08148_),
    .A(_08136_),
    .Y(_08153_),
    .D(_08152_));
 sg13g2_buf_8 _14965_ (.A(_08139_),
    .X(_08154_));
 sg13g2_mux4_1 _14966_ (.S0(net1060),
    .A0(\cpu.genblk1.mmu.r_valid_d[24] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[25] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[28] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[29] ),
    .S1(net1061),
    .X(_08155_));
 sg13g2_nand2_1 _14967_ (.Y(_08156_),
    .A(net1121),
    .B(_08155_));
 sg13g2_mux4_1 _14968_ (.S0(net1060),
    .A0(\cpu.genblk1.mmu.r_valid_d[26] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[27] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[30] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[31] ),
    .S1(net1061),
    .X(_08157_));
 sg13g2_nand3_1 _14969_ (.B(_08140_),
    .C(_08157_),
    .A(net1059),
    .Y(_08158_));
 sg13g2_o21ai_1 _14970_ (.B1(_08158_),
    .Y(_08159_),
    .A1(net1059),
    .A2(_08156_));
 sg13g2_mux2_1 _14971_ (.A0(\cpu.genblk1.mmu.r_valid_d[1] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[3] ),
    .S(net1059),
    .X(_08160_));
 sg13g2_buf_2 _14972_ (.A(net1120),
    .X(_08161_));
 sg13g2_nor2_1 _14973_ (.A(net1058),
    .B(net1121),
    .Y(_08162_));
 sg13g2_nand3_1 _14974_ (.B(_08160_),
    .C(_08162_),
    .A(net1062),
    .Y(_08163_));
 sg13g2_inv_1 _14975_ (.Y(_08164_),
    .A(_08132_));
 sg13g2_nand2b_1 _14976_ (.Y(_08165_),
    .B(_08134_),
    .A_N(_08133_));
 sg13g2_mux2_1 _14977_ (.A0(\cpu.genblk1.mmu.r_valid_d[0] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[2] ),
    .S(net1059),
    .X(_08166_));
 sg13g2_nor3_1 _14978_ (.A(net1062),
    .B(_08143_),
    .C(net1121),
    .Y(_08167_));
 sg13g2_a22oi_1 _14979_ (.Y(_08168_),
    .B1(_08166_),
    .B2(_08167_),
    .A2(_08165_),
    .A1(_08164_));
 sg13g2_buf_2 _14980_ (.A(net1121),
    .X(_08169_));
 sg13g2_mux4_1 _14981_ (.S0(_08150_),
    .A0(\cpu.genblk1.mmu.r_valid_d[12] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[13] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[14] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[15] ),
    .S1(net1059),
    .X(_08170_));
 sg13g2_nand3_1 _14982_ (.B(net1057),
    .C(_08170_),
    .A(net1058),
    .Y(_08171_));
 sg13g2_mux4_1 _14983_ (.S0(_08150_),
    .A0(\cpu.genblk1.mmu.r_valid_d[8] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[9] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[10] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[11] ),
    .S1(_08139_),
    .X(_08172_));
 sg13g2_nor2b_1 _14984_ (.A(net1058),
    .B_N(net1121),
    .Y(_08173_));
 sg13g2_mux4_1 _14985_ (.S0(net1062),
    .A0(\cpu.genblk1.mmu.r_valid_d[4] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[5] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[6] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[7] ),
    .S1(net1059),
    .X(_08174_));
 sg13g2_nor2b_1 _14986_ (.A(_08140_),
    .B_N(_08143_),
    .Y(_08175_));
 sg13g2_a22oi_1 _14987_ (.Y(_08176_),
    .B1(_08174_),
    .B2(_08175_),
    .A2(_08173_),
    .A1(_08172_));
 sg13g2_nand4_1 _14988_ (.B(_08168_),
    .C(_08171_),
    .A(_08163_),
    .Y(_08177_),
    .D(_08176_));
 sg13g2_o21ai_1 _14989_ (.B1(_08177_),
    .Y(_08178_),
    .A1(_08153_),
    .A2(_08159_));
 sg13g2_nor2_1 _14990_ (.A(_08125_),
    .B(_08127_),
    .Y(_08179_));
 sg13g2_buf_2 _14991_ (.A(_08179_),
    .X(_08180_));
 sg13g2_buf_2 _14992_ (.A(\cpu.ex.io_access ),
    .X(_08181_));
 sg13g2_buf_1 _14993_ (.A(\cpu.ex.genblk3.r_mmu_enable ),
    .X(_08182_));
 sg13g2_nand2b_1 _14994_ (.Y(_08183_),
    .B(_08182_),
    .A_N(_08181_));
 sg13g2_buf_2 _14995_ (.A(_08182_),
    .X(_08184_));
 sg13g2_buf_1 _14996_ (.A(\cpu.cond[0] ),
    .X(_08185_));
 sg13g2_buf_1 _14997_ (.A(_00182_),
    .X(_08186_));
 sg13g2_a21oi_2 _14998_ (.B1(net1119),
    .Y(_08187_),
    .A2(_08185_),
    .A1(\cpu.ex.mmu_reg_data[0] ));
 sg13g2_or2_1 _14999_ (.X(_08188_),
    .B(_08187_),
    .A(\cpu.ex.r_read_stall ));
 sg13g2_buf_1 _15000_ (.A(\cpu.ex.mmu_reg_data[0] ),
    .X(_08189_));
 sg13g2_inv_2 _15001_ (.Y(_08190_),
    .A(net1118));
 sg13g2_nand3_1 _15002_ (.B(_08185_),
    .C(net1119),
    .A(_08190_),
    .Y(_08191_));
 sg13g2_nand4_1 _15003_ (.B(_00181_),
    .C(_08188_),
    .A(net1056),
    .Y(_08192_),
    .D(_08191_));
 sg13g2_o21ai_1 _15004_ (.B1(_08192_),
    .Y(_08193_),
    .A1(_08180_),
    .A2(_08183_));
 sg13g2_nand2_1 _15005_ (.Y(_08194_),
    .A(_08178_),
    .B(_08193_));
 sg13g2_mux4_1 _15006_ (.S0(_08137_),
    .A0(\cpu.genblk1.mmu.r_writeable_d[2] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[3] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[6] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[7] ),
    .S1(net1120),
    .X(_08195_));
 sg13g2_nand2_1 _15007_ (.Y(_08196_),
    .A(_08149_),
    .B(_08195_));
 sg13g2_mux2_1 _15008_ (.A0(\cpu.genblk1.mmu.r_writeable_d[0] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[4] ),
    .S(net1120),
    .X(_08197_));
 sg13g2_nand2_1 _15009_ (.Y(_08198_),
    .A(_08141_),
    .B(_08197_));
 sg13g2_mux2_1 _15010_ (.A0(\cpu.genblk1.mmu.r_writeable_d[1] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[5] ),
    .S(net1120),
    .X(_08199_));
 sg13g2_nand3_1 _15011_ (.B(_08146_),
    .C(_08199_),
    .A(net1062),
    .Y(_08200_));
 sg13g2_a221oi_1 _15012_ (.B2(_08165_),
    .C1(_08183_),
    .B1(_08164_),
    .A1(_08126_),
    .Y(_08201_),
    .A2(_08128_));
 sg13g2_and4_1 _15013_ (.A(_08196_),
    .B(_08198_),
    .C(_08200_),
    .D(_08201_),
    .X(_08202_));
 sg13g2_mux4_1 _15014_ (.S0(net1060),
    .A0(\cpu.genblk1.mmu.r_writeable_d[8] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[9] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[12] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[13] ),
    .S1(net1061),
    .X(_08203_));
 sg13g2_mux4_1 _15015_ (.S0(net1060),
    .A0(\cpu.genblk1.mmu.r_writeable_d[10] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[11] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[14] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[15] ),
    .S1(net1061),
    .X(_08204_));
 sg13g2_mux2_1 _15016_ (.A0(_08203_),
    .A1(_08204_),
    .S(net1059),
    .X(_08205_));
 sg13g2_nand2_1 _15017_ (.Y(_08206_),
    .A(net1057),
    .B(_08205_));
 sg13g2_mux4_1 _15018_ (.S0(net1060),
    .A0(\cpu.genblk1.mmu.r_writeable_d[24] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[25] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[28] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[29] ),
    .S1(net1061),
    .X(_08207_));
 sg13g2_mux4_1 _15019_ (.S0(net1060),
    .A0(\cpu.genblk1.mmu.r_writeable_d[26] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[27] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[30] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[31] ),
    .S1(net1061),
    .X(_08208_));
 sg13g2_mux2_1 _15020_ (.A0(_08207_),
    .A1(_08208_),
    .S(net1059),
    .X(_08209_));
 sg13g2_nand2_1 _15021_ (.Y(_08210_),
    .A(net1057),
    .B(_08209_));
 sg13g2_mux4_1 _15022_ (.S0(net1060),
    .A0(\cpu.genblk1.mmu.r_writeable_d[18] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[19] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[22] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[23] ),
    .S1(net1120),
    .X(_08211_));
 sg13g2_nand2_1 _15023_ (.Y(_08212_),
    .A(_08149_),
    .B(_08211_));
 sg13g2_mux2_1 _15024_ (.A0(\cpu.genblk1.mmu.r_writeable_d[16] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[20] ),
    .S(net1120),
    .X(_08213_));
 sg13g2_nand2_1 _15025_ (.Y(_08214_),
    .A(_08141_),
    .B(_08213_));
 sg13g2_mux2_1 _15026_ (.A0(\cpu.genblk1.mmu.r_writeable_d[17] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[21] ),
    .S(net1120),
    .X(_08215_));
 sg13g2_nand3_1 _15027_ (.B(_08146_),
    .C(_08215_),
    .A(net1062),
    .Y(_08216_));
 sg13g2_nor4_1 _15028_ (.A(_08132_),
    .B(_08180_),
    .C(_08183_),
    .D(_08135_),
    .Y(_08217_));
 sg13g2_and4_1 _15029_ (.A(_08212_),
    .B(_08214_),
    .C(_08216_),
    .D(_08217_),
    .X(_08218_));
 sg13g2_a22oi_1 _15030_ (.Y(_08219_),
    .B1(_08210_),
    .B2(_08218_),
    .A2(_08206_),
    .A1(_08202_));
 sg13g2_buf_2 _15031_ (.A(_08219_),
    .X(_08220_));
 sg13g2_o21ai_1 _15032_ (.B1(_08220_),
    .Y(_08221_),
    .A1(_08131_),
    .A2(_08194_));
 sg13g2_buf_2 _15033_ (.A(\cpu.dec.supmode ),
    .X(_08222_));
 sg13g2_nand3_1 _15034_ (.B(net1056),
    .C(_08133_),
    .A(_08222_),
    .Y(_08223_));
 sg13g2_buf_8 _15035_ (.A(\cpu.ex.pc[13] ),
    .X(_08224_));
 sg13g2_buf_8 _15036_ (.A(\cpu.ex.pc[14] ),
    .X(_08225_));
 sg13g2_mux4_1 _15037_ (.S0(_08224_),
    .A0(\cpu.genblk1.mmu.r_valid_i[17] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[19] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[21] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[23] ),
    .S1(net1117),
    .X(_08226_));
 sg13g2_mux4_1 _15038_ (.S0(_08224_),
    .A0(\cpu.genblk1.mmu.r_valid_i[16] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[18] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[20] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[22] ),
    .S1(net1117),
    .X(_08227_));
 sg13g2_buf_8 _15039_ (.A(\cpu.ex.pc[12] ),
    .X(_08228_));
 sg13g2_inv_2 _15040_ (.Y(_08229_),
    .A(_08228_));
 sg13g2_mux2_1 _15041_ (.A0(_08226_),
    .A1(_08227_),
    .S(_08229_),
    .X(_08230_));
 sg13g2_buf_2 _15042_ (.A(\cpu.ex.pc[15] ),
    .X(_08231_));
 sg13g2_inv_1 _15043_ (.Y(_08232_),
    .A(_08231_));
 sg13g2_buf_4 _15044_ (.X(_08233_),
    .A(_08232_));
 sg13g2_o21ai_1 _15045_ (.B1(_08233_),
    .Y(_08234_),
    .A1(_08223_),
    .A2(_08230_));
 sg13g2_mux4_1 _15046_ (.S0(_08224_),
    .A0(\cpu.genblk1.mmu.r_valid_i[25] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[27] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[29] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[31] ),
    .S1(_08225_),
    .X(_08235_));
 sg13g2_nor2_1 _15047_ (.A(_08229_),
    .B(_08235_),
    .Y(_08236_));
 sg13g2_buf_2 _15048_ (.A(_08224_),
    .X(_08237_));
 sg13g2_nand2b_1 _15049_ (.Y(_08238_),
    .B(\cpu.genblk1.mmu.r_valid_i[26] ),
    .A_N(\cpu.ex.pc[14] ));
 sg13g2_nand2_1 _15050_ (.Y(_08239_),
    .A(net1117),
    .B(\cpu.genblk1.mmu.r_valid_i[30] ));
 sg13g2_and4_1 _15051_ (.A(_08229_),
    .B(net1055),
    .C(_08238_),
    .D(_08239_),
    .X(_08240_));
 sg13g2_mux2_1 _15052_ (.A0(\cpu.genblk1.mmu.r_valid_i[24] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[28] ),
    .S(net1117),
    .X(_08241_));
 sg13g2_nor3_1 _15053_ (.A(_08228_),
    .B(net1055),
    .C(_08241_),
    .Y(_08242_));
 sg13g2_nor4_1 _15054_ (.A(_08233_),
    .B(_08236_),
    .C(_08240_),
    .D(_08242_),
    .Y(_08243_));
 sg13g2_inv_1 _15055_ (.Y(_08244_),
    .A(_08222_));
 sg13g2_nand3_1 _15056_ (.B(net1056),
    .C(_08133_),
    .A(_08244_),
    .Y(_08245_));
 sg13g2_mux4_1 _15057_ (.S0(_08228_),
    .A0(\cpu.genblk1.mmu.r_valid_i[8] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[9] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[12] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[13] ),
    .S1(net1117),
    .X(_08246_));
 sg13g2_mux4_1 _15058_ (.S0(_08228_),
    .A0(\cpu.genblk1.mmu.r_valid_i[10] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[11] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[14] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[15] ),
    .S1(_08225_),
    .X(_08247_));
 sg13g2_mux2_1 _15059_ (.A0(_08246_),
    .A1(_08247_),
    .S(_08237_),
    .X(_08248_));
 sg13g2_or2_1 _15060_ (.X(_08249_),
    .B(_08248_),
    .A(_08245_));
 sg13g2_o21ai_1 _15061_ (.B1(_08249_),
    .Y(_08250_),
    .A1(_08223_),
    .A2(_08243_));
 sg13g2_mux4_1 _15062_ (.S0(_08237_),
    .A0(\cpu.genblk1.mmu.r_valid_i[1] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[3] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[5] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[7] ),
    .S1(net1117),
    .X(_08251_));
 sg13g2_mux4_1 _15063_ (.S0(_08224_),
    .A0(\cpu.genblk1.mmu.r_valid_i[0] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[2] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[4] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[6] ),
    .S1(net1117),
    .X(_08252_));
 sg13g2_mux2_1 _15064_ (.A0(_08251_),
    .A1(_08252_),
    .S(_08229_),
    .X(_08253_));
 sg13g2_nor3_1 _15065_ (.A(_08231_),
    .B(_08245_),
    .C(_08253_),
    .Y(_08254_));
 sg13g2_a21oi_1 _15066_ (.A1(_08234_),
    .A2(_08250_),
    .Y(_08255_),
    .B1(_08254_));
 sg13g2_buf_2 _15067_ (.A(_08255_),
    .X(_08256_));
 sg13g2_nor2_1 _15068_ (.A(_08131_),
    .B(_08256_),
    .Y(_08257_));
 sg13g2_nor2_2 _15069_ (.A(_08221_),
    .B(_08257_),
    .Y(_08258_));
 sg13g2_buf_1 _15070_ (.A(_08258_),
    .X(_08259_));
 sg13g2_nand2_2 _15071_ (.Y(_08260_),
    .A(_08123_),
    .B(net387));
 sg13g2_buf_1 _15072_ (.A(net1056),
    .X(_08261_));
 sg13g2_buf_2 _15073_ (.A(_08228_),
    .X(_08262_));
 sg13g2_buf_2 _15074_ (.A(_08262_),
    .X(_08263_));
 sg13g2_buf_2 _15075_ (.A(net1055),
    .X(_08264_));
 sg13g2_buf_1 _15076_ (.A(_08264_),
    .X(_08265_));
 sg13g2_mux4_1 _15077_ (.S0(net919),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][0] ),
    .S1(_08265_),
    .X(_08266_));
 sg13g2_mux4_1 _15078_ (.S0(net919),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][0] ),
    .S1(net798),
    .X(_08267_));
 sg13g2_buf_2 _15079_ (.A(_08262_),
    .X(_08268_));
 sg13g2_buf_1 _15080_ (.A(_08264_),
    .X(_08269_));
 sg13g2_mux4_1 _15081_ (.S0(net918),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][0] ),
    .S1(net797),
    .X(_08270_));
 sg13g2_mux4_1 _15082_ (.S0(net918),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][0] ),
    .S1(_08265_),
    .X(_08271_));
 sg13g2_buf_2 _15083_ (.A(_08233_),
    .X(_08272_));
 sg13g2_buf_1 _15084_ (.A(net1117),
    .X(_08273_));
 sg13g2_buf_1 _15085_ (.A(_08273_),
    .X(_08274_));
 sg13g2_mux4_1 _15086_ (.S0(net796),
    .A0(_08266_),
    .A1(_08267_),
    .A2(_08270_),
    .A3(_08271_),
    .S1(net917),
    .X(_08275_));
 sg13g2_mux4_1 _15087_ (.S0(net918),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][0] ),
    .S1(net798),
    .X(_08276_));
 sg13g2_mux4_1 _15088_ (.S0(net918),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][0] ),
    .S1(net798),
    .X(_08277_));
 sg13g2_mux4_1 _15089_ (.S0(net918),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][0] ),
    .S1(net797),
    .X(_08278_));
 sg13g2_mux4_1 _15090_ (.S0(net918),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][0] ),
    .S1(net797),
    .X(_08279_));
 sg13g2_mux4_1 _15091_ (.S0(net796),
    .A0(_08276_),
    .A1(_08277_),
    .A2(_08278_),
    .A3(_08279_),
    .S1(net917),
    .X(_08280_));
 sg13g2_buf_1 _15092_ (.A(_08244_),
    .X(_08281_));
 sg13g2_mux2_1 _15093_ (.A0(_08275_),
    .A1(_08280_),
    .S(_08281_),
    .X(_08282_));
 sg13g2_nor2_1 _15094_ (.A(_08229_),
    .B(_08261_),
    .Y(_08283_));
 sg13g2_a21oi_1 _15095_ (.A1(_08261_),
    .A2(_08282_),
    .Y(_08284_),
    .B1(_08283_));
 sg13g2_buf_2 _15096_ (.A(_08284_),
    .X(_08285_));
 sg13g2_buf_1 _15097_ (.A(_00174_),
    .X(_08286_));
 sg13g2_buf_2 _15098_ (.A(net1116),
    .X(_08287_));
 sg13g2_buf_2 _15099_ (.A(\cpu.ex.pc[2] ),
    .X(_08288_));
 sg13g2_buf_1 _15100_ (.A(\cpu.ex.pc[4] ),
    .X(_08289_));
 sg13g2_buf_1 _15101_ (.A(\cpu.ex.pc[3] ),
    .X(_08290_));
 sg13g2_nor2b_1 _15102_ (.A(_08289_),
    .B_N(net1115),
    .Y(_08291_));
 sg13g2_nand2b_1 _15103_ (.Y(_08292_),
    .B(_08289_),
    .A_N(net1115));
 sg13g2_o21ai_1 _15104_ (.B1(_08292_),
    .Y(_08293_),
    .A1(_08288_),
    .A2(_08291_));
 sg13g2_nand2_1 _15105_ (.Y(_08294_),
    .A(net1053),
    .B(_08293_));
 sg13g2_buf_2 _15106_ (.A(_08294_),
    .X(_08295_));
 sg13g2_buf_1 _15107_ (.A(_08295_),
    .X(_08296_));
 sg13g2_buf_1 _15108_ (.A(_08296_),
    .X(_08297_));
 sg13g2_buf_1 _15109_ (.A(net541),
    .X(_08298_));
 sg13g2_buf_1 _15110_ (.A(_08295_),
    .X(_08299_));
 sg13g2_buf_1 _15111_ (.A(net620),
    .X(_08300_));
 sg13g2_inv_1 _15112_ (.Y(_08301_),
    .A(_08288_));
 sg13g2_buf_2 _15113_ (.A(_08301_),
    .X(_08302_));
 sg13g2_and2_1 _15114_ (.A(net915),
    .B(_08291_),
    .X(_08303_));
 sg13g2_buf_2 _15115_ (.A(_08303_),
    .X(_08304_));
 sg13g2_buf_1 _15116_ (.A(_08304_),
    .X(_08305_));
 sg13g2_buf_1 _15117_ (.A(_08305_),
    .X(_08306_));
 sg13g2_nor3_1 _15118_ (.A(_08288_),
    .B(net1115),
    .C(net1116),
    .Y(_08307_));
 sg13g2_buf_2 _15119_ (.A(_08307_),
    .X(_08308_));
 sg13g2_buf_1 _15120_ (.A(_08308_),
    .X(_08309_));
 sg13g2_buf_1 _15121_ (.A(_08309_),
    .X(_08310_));
 sg13g2_a22oi_1 _15122_ (.Y(_08311_),
    .B1(net699),
    .B2(\cpu.icache.r_tag[4][12] ),
    .A2(net539),
    .A1(\cpu.icache.r_tag[2][12] ));
 sg13g2_nor3_1 _15123_ (.A(_08301_),
    .B(net1115),
    .C(_08289_),
    .Y(_08312_));
 sg13g2_buf_2 _15124_ (.A(_08312_),
    .X(_08313_));
 sg13g2_buf_1 _15125_ (.A(_08313_),
    .X(_08314_));
 sg13g2_buf_1 _15126_ (.A(net698),
    .X(_08315_));
 sg13g2_nor2_1 _15127_ (.A(_08288_),
    .B(net1116),
    .Y(_08316_));
 sg13g2_buf_2 _15128_ (.A(_08316_),
    .X(_08317_));
 sg13g2_and2_1 _15129_ (.A(net1115),
    .B(_08317_),
    .X(_08318_));
 sg13g2_buf_2 _15130_ (.A(_08318_),
    .X(_08319_));
 sg13g2_buf_1 _15131_ (.A(_08319_),
    .X(_08320_));
 sg13g2_buf_1 _15132_ (.A(_08320_),
    .X(_08321_));
 sg13g2_a22oi_1 _15133_ (.Y(_08322_),
    .B1(net538),
    .B2(\cpu.icache.r_tag[6][12] ),
    .A2(net618),
    .A1(\cpu.icache.r_tag[1][12] ));
 sg13g2_buf_1 _15134_ (.A(_08290_),
    .X(_08323_));
 sg13g2_buf_2 _15135_ (.A(_08323_),
    .X(_08324_));
 sg13g2_buf_1 _15136_ (.A(net914),
    .X(_08325_));
 sg13g2_mux2_1 _15137_ (.A0(\cpu.icache.r_tag[7][12] ),
    .A1(\cpu.icache.r_tag[3][12] ),
    .S(net1053),
    .X(_08326_));
 sg13g2_nor2_1 _15138_ (.A(net1115),
    .B(net1116),
    .Y(_08327_));
 sg13g2_buf_1 _15139_ (.A(_08327_),
    .X(_08328_));
 sg13g2_a22oi_1 _15140_ (.Y(_08329_),
    .B1(net913),
    .B2(\cpu.icache.r_tag[5][12] ),
    .A2(_08326_),
    .A1(net794));
 sg13g2_buf_2 _15141_ (.A(_08288_),
    .X(_08330_));
 sg13g2_buf_1 _15142_ (.A(net1051),
    .X(_08331_));
 sg13g2_buf_1 _15143_ (.A(net912),
    .X(_08332_));
 sg13g2_nand2b_1 _15144_ (.Y(_08333_),
    .B(net793),
    .A_N(_08329_));
 sg13g2_nand4_1 _15145_ (.B(_08311_),
    .C(_08322_),
    .A(net540),
    .Y(_08334_),
    .D(_08333_));
 sg13g2_o21ai_1 _15146_ (.B1(_08334_),
    .Y(_08335_),
    .A1(\cpu.icache.r_tag[0][12] ),
    .A2(net471));
 sg13g2_xnor2_1 _15147_ (.Y(_08336_),
    .A(net438),
    .B(_08335_));
 sg13g2_buf_1 _15148_ (.A(_08264_),
    .X(_08337_));
 sg13g2_buf_2 _15149_ (.A(net792),
    .X(_08338_));
 sg13g2_buf_1 _15150_ (.A(net697),
    .X(_08339_));
 sg13g2_mux4_1 _15151_ (.S0(_08268_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][1] ),
    .S1(net797),
    .X(_08340_));
 sg13g2_mux4_1 _15152_ (.S0(_08268_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][1] ),
    .S1(_08269_),
    .X(_08341_));
 sg13g2_buf_2 _15153_ (.A(_08262_),
    .X(_08342_));
 sg13g2_mux4_1 _15154_ (.S0(net911),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][1] ),
    .S1(net797),
    .X(_08343_));
 sg13g2_mux4_1 _15155_ (.S0(net911),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][1] ),
    .S1(_08269_),
    .X(_08344_));
 sg13g2_mux4_1 _15156_ (.S0(_08272_),
    .A0(_08340_),
    .A1(_08341_),
    .A2(_08343_),
    .A3(_08344_),
    .S1(net917),
    .X(_08345_));
 sg13g2_nand2_1 _15157_ (.Y(_08346_),
    .A(_08222_),
    .B(_08345_));
 sg13g2_mux4_1 _15158_ (.S0(net911),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][1] ),
    .S1(net797),
    .X(_08347_));
 sg13g2_mux4_1 _15159_ (.S0(net911),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][1] ),
    .S1(net797),
    .X(_08348_));
 sg13g2_buf_1 _15160_ (.A(_08264_),
    .X(_08349_));
 sg13g2_mux4_1 _15161_ (.S0(_08342_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][1] ),
    .S1(_08349_),
    .X(_08350_));
 sg13g2_mux4_1 _15162_ (.S0(_08342_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][1] ),
    .S1(net797),
    .X(_08351_));
 sg13g2_mux4_1 _15163_ (.S0(_08272_),
    .A0(_08347_),
    .A1(_08348_),
    .A2(_08350_),
    .A3(_08351_),
    .S1(net917),
    .X(_08352_));
 sg13g2_nand2_1 _15164_ (.Y(_08353_),
    .A(_08281_),
    .B(_08352_));
 sg13g2_nand3_1 _15165_ (.B(_08346_),
    .C(_08353_),
    .A(net920),
    .Y(_08354_));
 sg13g2_o21ai_1 _15166_ (.B1(_08354_),
    .Y(_08355_),
    .A1(net616),
    .A2(net920));
 sg13g2_buf_1 _15167_ (.A(_08355_),
    .X(_08356_));
 sg13g2_buf_1 _15168_ (.A(_08297_),
    .X(_08357_));
 sg13g2_buf_1 _15169_ (.A(_08305_),
    .X(_08358_));
 sg13g2_nor3_1 _15170_ (.A(_08301_),
    .B(net1115),
    .C(_08286_),
    .Y(_08359_));
 sg13g2_buf_2 _15171_ (.A(_08359_),
    .X(_08360_));
 sg13g2_buf_1 _15172_ (.A(_08360_),
    .X(_08361_));
 sg13g2_inv_1 _15173_ (.Y(_08362_),
    .A(net1116));
 sg13g2_and2_1 _15174_ (.A(_08288_),
    .B(\cpu.ex.pc[3] ),
    .X(_08363_));
 sg13g2_buf_2 _15175_ (.A(_08363_),
    .X(_08364_));
 sg13g2_and2_1 _15176_ (.A(net1050),
    .B(_08364_),
    .X(_08365_));
 sg13g2_buf_1 _15177_ (.A(_08365_),
    .X(_08366_));
 sg13g2_buf_1 _15178_ (.A(_08366_),
    .X(_08367_));
 sg13g2_and2_1 _15179_ (.A(\cpu.icache.r_tag[7][13] ),
    .B(net615),
    .X(_08368_));
 sg13g2_a221oi_1 _15180_ (.B2(\cpu.icache.r_tag[5][13] ),
    .C1(_08368_),
    .B1(net696),
    .A1(\cpu.icache.r_tag[2][13] ),
    .Y(_08369_),
    .A2(net537));
 sg13g2_a22oi_1 _15181_ (.Y(_08370_),
    .B1(net618),
    .B2(\cpu.icache.r_tag[1][13] ),
    .A2(net699),
    .A1(\cpu.icache.r_tag[4][13] ));
 sg13g2_and2_1 _15182_ (.A(_08286_),
    .B(_08364_),
    .X(_08371_));
 sg13g2_buf_1 _15183_ (.A(_08371_),
    .X(_08372_));
 sg13g2_buf_2 _15184_ (.A(_08372_),
    .X(_08373_));
 sg13g2_buf_2 _15185_ (.A(net614),
    .X(_08374_));
 sg13g2_a22oi_1 _15186_ (.Y(_08375_),
    .B1(net536),
    .B2(\cpu.icache.r_tag[3][13] ),
    .A2(net538),
    .A1(\cpu.icache.r_tag[6][13] ));
 sg13g2_nand4_1 _15187_ (.B(_08369_),
    .C(_08370_),
    .A(net540),
    .Y(_08376_),
    .D(_08375_));
 sg13g2_o21ai_1 _15188_ (.B1(_08376_),
    .Y(_08377_),
    .A1(\cpu.icache.r_tag[0][13] ),
    .A2(net470));
 sg13g2_xnor2_1 _15189_ (.Y(_08378_),
    .A(net386),
    .B(_08377_));
 sg13g2_nand2_1 _15190_ (.Y(_08379_),
    .A(_08336_),
    .B(_08378_));
 sg13g2_buf_2 _15191_ (.A(_00176_),
    .X(_08380_));
 sg13g2_buf_1 _15192_ (.A(_08380_),
    .X(_08381_));
 sg13g2_buf_2 _15193_ (.A(_08262_),
    .X(_08382_));
 sg13g2_buf_1 _15194_ (.A(net792),
    .X(_08383_));
 sg13g2_mux4_1 _15195_ (.S0(_08382_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][8] ),
    .S1(_08383_),
    .X(_08384_));
 sg13g2_mux4_1 _15196_ (.S0(_08382_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][8] ),
    .S1(_08383_),
    .X(_08385_));
 sg13g2_buf_2 _15197_ (.A(_08262_),
    .X(_08386_));
 sg13g2_mux4_1 _15198_ (.S0(net909),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][8] ),
    .S1(net697),
    .X(_08387_));
 sg13g2_mux4_1 _15199_ (.S0(net909),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][8] ),
    .S1(net697),
    .X(_08388_));
 sg13g2_buf_1 _15200_ (.A(_08233_),
    .X(_08389_));
 sg13g2_mux4_1 _15201_ (.S0(net790),
    .A0(_08384_),
    .A1(_08385_),
    .A2(_08387_),
    .A3(_08388_),
    .S1(net917),
    .X(_08390_));
 sg13g2_mux4_1 _15202_ (.S0(net910),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][8] ),
    .S1(net697),
    .X(_08391_));
 sg13g2_mux4_1 _15203_ (.S0(net910),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][8] ),
    .S1(net697),
    .X(_08392_));
 sg13g2_buf_2 _15204_ (.A(net792),
    .X(_08393_));
 sg13g2_mux4_1 _15205_ (.S0(net909),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][8] ),
    .S1(net694),
    .X(_08394_));
 sg13g2_mux4_1 _15206_ (.S0(net909),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][8] ),
    .S1(net697),
    .X(_08395_));
 sg13g2_mux4_1 _15207_ (.S0(net790),
    .A0(_08391_),
    .A1(_08392_),
    .A2(_08394_),
    .A3(_08395_),
    .S1(net917),
    .X(_08396_));
 sg13g2_buf_1 _15208_ (.A(net916),
    .X(_08397_));
 sg13g2_mux2_1 _15209_ (.A0(_08390_),
    .A1(_08396_),
    .S(net789),
    .X(_08398_));
 sg13g2_nand2b_1 _15210_ (.Y(_08399_),
    .B(_08398_),
    .A_N(net1049));
 sg13g2_buf_1 _15211_ (.A(_08399_),
    .X(_08400_));
 sg13g2_a22oi_1 _15212_ (.Y(_08401_),
    .B1(net699),
    .B2(\cpu.icache.r_tag[4][20] ),
    .A2(net539),
    .A1(\cpu.icache.r_tag[2][20] ));
 sg13g2_buf_1 _15213_ (.A(net698),
    .X(_08402_));
 sg13g2_a22oi_1 _15214_ (.Y(_08403_),
    .B1(net538),
    .B2(\cpu.icache.r_tag[6][20] ),
    .A2(net613),
    .A1(\cpu.icache.r_tag[1][20] ));
 sg13g2_mux2_1 _15215_ (.A0(\cpu.icache.r_tag[7][20] ),
    .A1(\cpu.icache.r_tag[3][20] ),
    .S(net1053),
    .X(_08404_));
 sg13g2_a22oi_1 _15216_ (.Y(_08405_),
    .B1(_08404_),
    .B2(net794),
    .A2(net913),
    .A1(\cpu.icache.r_tag[5][20] ));
 sg13g2_nand2b_1 _15217_ (.Y(_08406_),
    .B(net793),
    .A_N(_08405_));
 sg13g2_nand4_1 _15218_ (.B(_08401_),
    .C(_08403_),
    .A(net540),
    .Y(_08407_),
    .D(_08406_));
 sg13g2_o21ai_1 _15219_ (.B1(_08407_),
    .Y(_08408_),
    .A1(\cpu.icache.r_tag[0][20] ),
    .A2(net470));
 sg13g2_xnor2_1 _15220_ (.Y(_08409_),
    .A(net385),
    .B(_08408_));
 sg13g2_mux4_1 _15221_ (.S0(net909),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][9] ),
    .S1(_08338_),
    .X(_08410_));
 sg13g2_mux4_1 _15222_ (.S0(net909),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][9] ),
    .S1(_08338_),
    .X(_08411_));
 sg13g2_mux4_1 _15223_ (.S0(_08386_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][9] ),
    .S1(net694),
    .X(_08412_));
 sg13g2_mux4_1 _15224_ (.S0(net909),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][9] ),
    .S1(net694),
    .X(_08413_));
 sg13g2_mux4_1 _15225_ (.S0(net790),
    .A0(_08410_),
    .A1(_08411_),
    .A2(_08412_),
    .A3(_08413_),
    .S1(_08274_),
    .X(_08414_));
 sg13g2_mux4_1 _15226_ (.S0(net909),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][9] ),
    .S1(net694),
    .X(_08415_));
 sg13g2_mux4_1 _15227_ (.S0(_08386_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][9] ),
    .S1(net694),
    .X(_08416_));
 sg13g2_mux4_1 _15228_ (.S0(_08263_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][9] ),
    .S1(_08393_),
    .X(_08417_));
 sg13g2_mux4_1 _15229_ (.S0(_08263_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][9] ),
    .S1(_08393_),
    .X(_08418_));
 sg13g2_mux4_1 _15230_ (.S0(_08389_),
    .A0(_08415_),
    .A1(_08416_),
    .A2(_08417_),
    .A3(_08418_),
    .S1(_08274_),
    .X(_08419_));
 sg13g2_mux2_1 _15231_ (.A0(_08414_),
    .A1(_08419_),
    .S(net789),
    .X(_08420_));
 sg13g2_nand2b_1 _15232_ (.Y(_08421_),
    .B(_08420_),
    .A_N(net1049));
 sg13g2_buf_1 _15233_ (.A(_08421_),
    .X(_08422_));
 sg13g2_a22oi_1 _15234_ (.Y(_08423_),
    .B1(_08361_),
    .B2(\cpu.icache.r_tag[5][21] ),
    .A2(net617),
    .A1(\cpu.icache.r_tag[6][21] ));
 sg13g2_buf_1 _15235_ (.A(_08364_),
    .X(_08424_));
 sg13g2_buf_1 _15236_ (.A(net1053),
    .X(_08425_));
 sg13g2_mux2_1 _15237_ (.A0(\cpu.icache.r_tag[7][21] ),
    .A1(\cpu.icache.r_tag[3][21] ),
    .S(net908),
    .X(_08426_));
 sg13g2_a22oi_1 _15238_ (.Y(_08427_),
    .B1(net788),
    .B2(_08426_),
    .A2(net613),
    .A1(\cpu.icache.r_tag[1][21] ));
 sg13g2_a22oi_1 _15239_ (.Y(_08428_),
    .B1(net699),
    .B2(\cpu.icache.r_tag[4][21] ),
    .A2(net537),
    .A1(\cpu.icache.r_tag[2][21] ));
 sg13g2_nand4_1 _15240_ (.B(_08423_),
    .C(_08427_),
    .A(net541),
    .Y(_08429_),
    .D(_08428_));
 sg13g2_o21ai_1 _15241_ (.B1(_08429_),
    .Y(_08430_),
    .A1(\cpu.icache.r_tag[0][21] ),
    .A2(net470));
 sg13g2_xnor2_1 _15242_ (.Y(_08431_),
    .A(net384),
    .B(_08430_));
 sg13g2_buf_2 _15243_ (.A(_08262_),
    .X(_08432_));
 sg13g2_buf_1 _15244_ (.A(net792),
    .X(_08433_));
 sg13g2_mux4_1 _15245_ (.S0(net907),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][4] ),
    .S1(net693),
    .X(_08434_));
 sg13g2_mux4_1 _15246_ (.S0(net907),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][4] ),
    .S1(net693),
    .X(_08435_));
 sg13g2_mux4_1 _15247_ (.S0(net907),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][4] ),
    .S1(net695),
    .X(_08436_));
 sg13g2_mux4_1 _15248_ (.S0(net907),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][4] ),
    .S1(net695),
    .X(_08437_));
 sg13g2_buf_1 _15249_ (.A(_08273_),
    .X(_08438_));
 sg13g2_mux4_1 _15250_ (.S0(net790),
    .A0(_08434_),
    .A1(_08435_),
    .A2(_08436_),
    .A3(_08437_),
    .S1(net906),
    .X(_08439_));
 sg13g2_mux4_1 _15251_ (.S0(_08432_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][4] ),
    .S1(net695),
    .X(_08440_));
 sg13g2_mux4_1 _15252_ (.S0(_08432_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][4] ),
    .S1(net695),
    .X(_08441_));
 sg13g2_mux4_1 _15253_ (.S0(net910),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][4] ),
    .S1(net695),
    .X(_08442_));
 sg13g2_mux4_1 _15254_ (.S0(net910),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][4] ),
    .S1(net695),
    .X(_08443_));
 sg13g2_mux4_1 _15255_ (.S0(net790),
    .A0(_08440_),
    .A1(_08441_),
    .A2(_08442_),
    .A3(_08443_),
    .S1(net906),
    .X(_08444_));
 sg13g2_mux2_1 _15256_ (.A0(_08439_),
    .A1(_08444_),
    .S(net789),
    .X(_08445_));
 sg13g2_nand2b_1 _15257_ (.Y(_08446_),
    .B(_08445_),
    .A_N(net1049));
 sg13g2_buf_2 _15258_ (.A(_08446_),
    .X(_08447_));
 sg13g2_a22oi_1 _15259_ (.Y(_08448_),
    .B1(net699),
    .B2(\cpu.icache.r_tag[4][16] ),
    .A2(net539),
    .A1(\cpu.icache.r_tag[2][16] ));
 sg13g2_a22oi_1 _15260_ (.Y(_08449_),
    .B1(net538),
    .B2(\cpu.icache.r_tag[6][16] ),
    .A2(net618),
    .A1(\cpu.icache.r_tag[1][16] ));
 sg13g2_mux2_1 _15261_ (.A0(\cpu.icache.r_tag[7][16] ),
    .A1(\cpu.icache.r_tag[3][16] ),
    .S(net908),
    .X(_08450_));
 sg13g2_a22oi_1 _15262_ (.Y(_08451_),
    .B1(_08450_),
    .B2(net794),
    .A2(net913),
    .A1(\cpu.icache.r_tag[5][16] ));
 sg13g2_nand2b_1 _15263_ (.Y(_08452_),
    .B(net793),
    .A_N(_08451_));
 sg13g2_nand4_1 _15264_ (.B(_08448_),
    .C(_08449_),
    .A(net540),
    .Y(_08453_),
    .D(_08452_));
 sg13g2_o21ai_1 _15265_ (.B1(_08453_),
    .Y(_08454_),
    .A1(\cpu.icache.r_tag[0][16] ),
    .A2(net471));
 sg13g2_xnor2_1 _15266_ (.Y(_08455_),
    .A(_08447_),
    .B(_08454_));
 sg13g2_mux4_1 _15267_ (.S0(net910),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][2] ),
    .S1(net695),
    .X(_08456_));
 sg13g2_mux4_1 _15268_ (.S0(net910),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][2] ),
    .S1(net695),
    .X(_08457_));
 sg13g2_mux4_1 _15269_ (.S0(net910),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][2] ),
    .S1(net697),
    .X(_08458_));
 sg13g2_mux4_1 _15270_ (.S0(net910),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][2] ),
    .S1(net697),
    .X(_08459_));
 sg13g2_mux4_1 _15271_ (.S0(net916),
    .A0(_08456_),
    .A1(_08457_),
    .A2(_08458_),
    .A3(_08459_),
    .S1(_08231_),
    .X(_08460_));
 sg13g2_nand2b_1 _15272_ (.Y(_08461_),
    .B(net920),
    .A_N(_08460_));
 sg13g2_buf_2 _15273_ (.A(_08228_),
    .X(_08462_));
 sg13g2_buf_2 _15274_ (.A(net1048),
    .X(_08463_));
 sg13g2_buf_2 _15275_ (.A(net905),
    .X(_08464_));
 sg13g2_mux4_1 _15276_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][2] ),
    .S1(net616),
    .X(_08465_));
 sg13g2_mux4_1 _15277_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][2] ),
    .S1(net616),
    .X(_08466_));
 sg13g2_mux4_1 _15278_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][2] ),
    .S1(net616),
    .X(_08467_));
 sg13g2_mux4_1 _15279_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][2] ),
    .S1(net616),
    .X(_08468_));
 sg13g2_mux4_1 _15280_ (.S0(net916),
    .A0(_08465_),
    .A1(_08466_),
    .A2(_08467_),
    .A3(_08468_),
    .S1(_08231_),
    .X(_08469_));
 sg13g2_inv_2 _15281_ (.Y(_08470_),
    .A(_08184_));
 sg13g2_nor2_1 _15282_ (.A(net906),
    .B(_08470_),
    .Y(_08471_));
 sg13g2_a22oi_1 _15283_ (.Y(_08472_),
    .B1(_08469_),
    .B2(_08471_),
    .A2(_08461_),
    .A1(net906));
 sg13g2_buf_2 _15284_ (.A(_08472_),
    .X(_08473_));
 sg13g2_mux2_1 _15285_ (.A0(\cpu.icache.r_tag[7][14] ),
    .A1(\cpu.icache.r_tag[3][14] ),
    .S(net908),
    .X(_08474_));
 sg13g2_a22oi_1 _15286_ (.Y(_08475_),
    .B1(net788),
    .B2(_08474_),
    .A2(net539),
    .A1(\cpu.icache.r_tag[2][14] ));
 sg13g2_a22oi_1 _15287_ (.Y(_08476_),
    .B1(net696),
    .B2(\cpu.icache.r_tag[5][14] ),
    .A2(net618),
    .A1(\cpu.icache.r_tag[1][14] ));
 sg13g2_a22oi_1 _15288_ (.Y(_08477_),
    .B1(net538),
    .B2(\cpu.icache.r_tag[6][14] ),
    .A2(net699),
    .A1(\cpu.icache.r_tag[4][14] ));
 sg13g2_nand4_1 _15289_ (.B(_08475_),
    .C(_08476_),
    .A(net540),
    .Y(_08478_),
    .D(_08477_));
 sg13g2_o21ai_1 _15290_ (.B1(_08478_),
    .Y(_08479_),
    .A1(\cpu.icache.r_tag[0][14] ),
    .A2(net471));
 sg13g2_xnor2_1 _15291_ (.Y(_08480_),
    .A(net382),
    .B(_08479_));
 sg13g2_nand4_1 _15292_ (.B(_08431_),
    .C(_08455_),
    .A(_08409_),
    .Y(_08481_),
    .D(_08480_));
 sg13g2_mux4_1 _15293_ (.S0(net919),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][7] ),
    .S1(net694),
    .X(_08482_));
 sg13g2_mux4_1 _15294_ (.S0(net919),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][7] ),
    .S1(net694),
    .X(_08483_));
 sg13g2_mux4_1 _15295_ (.S0(net919),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][7] ),
    .S1(net798),
    .X(_08484_));
 sg13g2_mux4_1 _15296_ (.S0(net919),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][7] ),
    .S1(net798),
    .X(_08485_));
 sg13g2_mux4_1 _15297_ (.S0(net790),
    .A0(_08482_),
    .A1(_08483_),
    .A2(_08484_),
    .A3(_08485_),
    .S1(net917),
    .X(_08486_));
 sg13g2_mux4_1 _15298_ (.S0(net919),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][7] ),
    .S1(net798),
    .X(_08487_));
 sg13g2_mux4_1 _15299_ (.S0(net919),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][7] ),
    .S1(net694),
    .X(_08488_));
 sg13g2_mux4_1 _15300_ (.S0(net918),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][7] ),
    .S1(net798),
    .X(_08489_));
 sg13g2_mux4_1 _15301_ (.S0(net918),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][7] ),
    .S1(net798),
    .X(_08490_));
 sg13g2_mux4_1 _15302_ (.S0(net796),
    .A0(_08487_),
    .A1(_08488_),
    .A2(_08489_),
    .A3(_08490_),
    .S1(net917),
    .X(_08491_));
 sg13g2_mux2_1 _15303_ (.A0(_08486_),
    .A1(_08491_),
    .S(net789),
    .X(_08492_));
 sg13g2_nand2b_1 _15304_ (.Y(_08493_),
    .B(_08492_),
    .A_N(net1049));
 sg13g2_buf_1 _15305_ (.A(_08493_),
    .X(_08494_));
 sg13g2_mux2_1 _15306_ (.A0(\cpu.icache.r_tag[7][19] ),
    .A1(\cpu.icache.r_tag[3][19] ),
    .S(net908),
    .X(_08495_));
 sg13g2_a22oi_1 _15307_ (.Y(_08496_),
    .B1(net788),
    .B2(_08495_),
    .A2(net537),
    .A1(\cpu.icache.r_tag[2][19] ));
 sg13g2_a22oi_1 _15308_ (.Y(_08497_),
    .B1(net696),
    .B2(\cpu.icache.r_tag[5][19] ),
    .A2(net795),
    .A1(\cpu.icache.r_tag[4][19] ));
 sg13g2_a22oi_1 _15309_ (.Y(_08498_),
    .B1(net617),
    .B2(\cpu.icache.r_tag[6][19] ),
    .A2(net613),
    .A1(\cpu.icache.r_tag[1][19] ));
 sg13g2_nand4_1 _15310_ (.B(_08496_),
    .C(_08497_),
    .A(net541),
    .Y(_08499_),
    .D(_08498_));
 sg13g2_o21ai_1 _15311_ (.B1(_08499_),
    .Y(_08500_),
    .A1(\cpu.icache.r_tag[0][19] ),
    .A2(net470));
 sg13g2_xnor2_1 _15312_ (.Y(_08501_),
    .A(net381),
    .B(_08500_));
 sg13g2_mux4_1 _15313_ (.S0(net907),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][3] ),
    .S1(net693),
    .X(_08502_));
 sg13g2_mux4_1 _15314_ (.S0(net907),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][3] ),
    .S1(_08433_),
    .X(_08503_));
 sg13g2_mux4_1 _15315_ (.S0(net907),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][3] ),
    .S1(net693),
    .X(_08504_));
 sg13g2_mux4_1 _15316_ (.S0(net907),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][3] ),
    .S1(_08433_),
    .X(_08505_));
 sg13g2_mux4_1 _15317_ (.S0(net916),
    .A0(_08502_),
    .A1(_08503_),
    .A2(_08504_),
    .A3(_08505_),
    .S1(net906),
    .X(_08506_));
 sg13g2_a21oi_1 _15318_ (.A1(net920),
    .A2(_08506_),
    .Y(_08507_),
    .B1(_08231_));
 sg13g2_mux4_1 _15319_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][3] ),
    .S1(net693),
    .X(_08508_));
 sg13g2_mux4_1 _15320_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][3] ),
    .S1(net693),
    .X(_08509_));
 sg13g2_mux4_1 _15321_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][3] ),
    .S1(net693),
    .X(_08510_));
 sg13g2_mux4_1 _15322_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][3] ),
    .S1(net693),
    .X(_08511_));
 sg13g2_mux4_1 _15323_ (.S0(net916),
    .A0(_08508_),
    .A1(_08509_),
    .A2(_08510_),
    .A3(_08511_),
    .S1(net906),
    .X(_08512_));
 sg13g2_nor3_1 _15324_ (.A(net790),
    .B(_08470_),
    .C(_08512_),
    .Y(_08513_));
 sg13g2_or2_1 _15325_ (.X(_08514_),
    .B(_08513_),
    .A(_08507_));
 sg13g2_buf_1 _15326_ (.A(_08514_),
    .X(_08515_));
 sg13g2_mux2_1 _15327_ (.A0(\cpu.icache.r_tag[7][15] ),
    .A1(\cpu.icache.r_tag[3][15] ),
    .S(net908),
    .X(_08516_));
 sg13g2_a22oi_1 _15328_ (.Y(_08517_),
    .B1(net788),
    .B2(_08516_),
    .A2(net618),
    .A1(\cpu.icache.r_tag[1][15] ));
 sg13g2_a22oi_1 _15329_ (.Y(_08518_),
    .B1(net699),
    .B2(\cpu.icache.r_tag[4][15] ),
    .A2(net539),
    .A1(\cpu.icache.r_tag[2][15] ));
 sg13g2_a22oi_1 _15330_ (.Y(_08519_),
    .B1(_08361_),
    .B2(\cpu.icache.r_tag[5][15] ),
    .A2(net538),
    .A1(\cpu.icache.r_tag[6][15] ));
 sg13g2_nand4_1 _15331_ (.B(_08517_),
    .C(_08518_),
    .A(net540),
    .Y(_08520_),
    .D(_08519_));
 sg13g2_o21ai_1 _15332_ (.B1(_08520_),
    .Y(_08521_),
    .A1(\cpu.icache.r_tag[0][15] ),
    .A2(net471));
 sg13g2_xnor2_1 _15333_ (.Y(_08522_),
    .A(net380),
    .B(_08521_));
 sg13g2_mux4_1 _15334_ (.S0(_08462_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][11] ),
    .S1(_08264_),
    .X(_08523_));
 sg13g2_mux4_1 _15335_ (.S0(net1048),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][11] ),
    .S1(_08264_),
    .X(_08524_));
 sg13g2_mux4_1 _15336_ (.S0(net1048),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][11] ),
    .S1(net1055),
    .X(_08525_));
 sg13g2_mux4_1 _15337_ (.S0(net1048),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][11] ),
    .S1(net1055),
    .X(_08526_));
 sg13g2_mux4_1 _15338_ (.S0(_08233_),
    .A0(_08523_),
    .A1(_08524_),
    .A2(_08525_),
    .A3(_08526_),
    .S1(net1054),
    .X(_08527_));
 sg13g2_mux4_1 _15339_ (.S0(net1048),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][11] ),
    .S1(net1055),
    .X(_08528_));
 sg13g2_mux4_1 _15340_ (.S0(net1048),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][11] ),
    .S1(_08264_),
    .X(_08529_));
 sg13g2_mux4_1 _15341_ (.S0(_08228_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][11] ),
    .S1(net1055),
    .X(_08530_));
 sg13g2_mux4_1 _15342_ (.S0(net1048),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][11] ),
    .S1(net1055),
    .X(_08531_));
 sg13g2_mux4_1 _15343_ (.S0(_08233_),
    .A0(_08528_),
    .A1(_08529_),
    .A2(_08530_),
    .A3(_08531_),
    .S1(net1054),
    .X(_08532_));
 sg13g2_mux2_1 _15344_ (.A0(_08527_),
    .A1(_08532_),
    .S(_08244_),
    .X(_08533_));
 sg13g2_nand2b_1 _15345_ (.Y(_08534_),
    .B(_08533_),
    .A_N(net1049));
 sg13g2_buf_1 _15346_ (.A(_08534_),
    .X(_08535_));
 sg13g2_and2_1 _15347_ (.A(\cpu.icache.r_tag[7][23] ),
    .B(net615),
    .X(_08536_));
 sg13g2_a221oi_1 _15348_ (.B2(\cpu.icache.r_tag[5][23] ),
    .C1(_08536_),
    .B1(net696),
    .A1(\cpu.icache.r_tag[2][23] ),
    .Y(_08537_),
    .A2(net619));
 sg13g2_a22oi_1 _15349_ (.Y(_08538_),
    .B1(net613),
    .B2(\cpu.icache.r_tag[1][23] ),
    .A2(net795),
    .A1(\cpu.icache.r_tag[4][23] ));
 sg13g2_a22oi_1 _15350_ (.Y(_08539_),
    .B1(net614),
    .B2(\cpu.icache.r_tag[3][23] ),
    .A2(net617),
    .A1(\cpu.icache.r_tag[6][23] ));
 sg13g2_nand4_1 _15351_ (.B(_08537_),
    .C(_08538_),
    .A(net620),
    .Y(_08540_),
    .D(_08539_));
 sg13g2_o21ai_1 _15352_ (.B1(_08540_),
    .Y(_08541_),
    .A1(\cpu.icache.r_tag[0][23] ),
    .A2(net541));
 sg13g2_xor2_1 _15353_ (.B(_08541_),
    .A(net469),
    .X(_08542_));
 sg13g2_mux4_1 _15354_ (.S0(net911),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][5] ),
    .S1(net791),
    .X(_08543_));
 sg13g2_mux4_1 _15355_ (.S0(net911),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][5] ),
    .S1(net791),
    .X(_08544_));
 sg13g2_buf_1 _15356_ (.A(_08264_),
    .X(_08545_));
 sg13g2_mux4_1 _15357_ (.S0(net905),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][5] ),
    .S1(net786),
    .X(_08546_));
 sg13g2_mux4_1 _15358_ (.S0(net905),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][5] ),
    .S1(net791),
    .X(_08547_));
 sg13g2_mux4_1 _15359_ (.S0(net796),
    .A0(_08543_),
    .A1(_08544_),
    .A2(_08546_),
    .A3(_08547_),
    .S1(net1054),
    .X(_08548_));
 sg13g2_mux4_1 _15360_ (.S0(net911),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][5] ),
    .S1(net791),
    .X(_08549_));
 sg13g2_mux4_1 _15361_ (.S0(net911),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][5] ),
    .S1(net791),
    .X(_08550_));
 sg13g2_buf_2 _15362_ (.A(net1048),
    .X(_08551_));
 sg13g2_mux4_1 _15363_ (.S0(net904),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][5] ),
    .S1(_08545_),
    .X(_08552_));
 sg13g2_mux4_1 _15364_ (.S0(_08551_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][5] ),
    .S1(net786),
    .X(_08553_));
 sg13g2_mux4_1 _15365_ (.S0(net796),
    .A0(_08549_),
    .A1(_08550_),
    .A2(_08552_),
    .A3(_08553_),
    .S1(net1054),
    .X(_08554_));
 sg13g2_mux2_1 _15366_ (.A0(_08548_),
    .A1(_08554_),
    .S(net916),
    .X(_08555_));
 sg13g2_nand2b_1 _15367_ (.Y(_08556_),
    .B(_08555_),
    .A_N(net1049));
 sg13g2_buf_1 _15368_ (.A(_08556_),
    .X(_08557_));
 sg13g2_and2_1 _15369_ (.A(\cpu.icache.r_tag[3][17] ),
    .B(net614),
    .X(_08558_));
 sg13g2_a221oi_1 _15370_ (.B2(\cpu.icache.r_tag[5][17] ),
    .C1(_08558_),
    .B1(net696),
    .A1(\cpu.icache.r_tag[2][17] ),
    .Y(_08559_),
    .A2(net619));
 sg13g2_a22oi_1 _15371_ (.Y(_08560_),
    .B1(net613),
    .B2(\cpu.icache.r_tag[1][17] ),
    .A2(net795),
    .A1(\cpu.icache.r_tag[4][17] ));
 sg13g2_a22oi_1 _15372_ (.Y(_08561_),
    .B1(net615),
    .B2(\cpu.icache.r_tag[7][17] ),
    .A2(net617),
    .A1(\cpu.icache.r_tag[6][17] ));
 sg13g2_nand4_1 _15373_ (.B(_08559_),
    .C(_08560_),
    .A(net541),
    .Y(_08562_),
    .D(_08561_));
 sg13g2_o21ai_1 _15374_ (.B1(_08562_),
    .Y(_08563_),
    .A1(\cpu.icache.r_tag[0][17] ),
    .A2(net540));
 sg13g2_xor2_1 _15375_ (.B(_08563_),
    .A(net437),
    .X(_08564_));
 sg13g2_mux4_1 _15376_ (.S0(net905),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][6] ),
    .S1(net791),
    .X(_08565_));
 sg13g2_mux4_1 _15377_ (.S0(net905),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][6] ),
    .S1(net791),
    .X(_08566_));
 sg13g2_mux4_1 _15378_ (.S0(net904),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][6] ),
    .S1(net786),
    .X(_08567_));
 sg13g2_mux4_1 _15379_ (.S0(net904),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][6] ),
    .S1(net786),
    .X(_08568_));
 sg13g2_mux4_1 _15380_ (.S0(net796),
    .A0(_08565_),
    .A1(_08566_),
    .A2(_08567_),
    .A3(_08568_),
    .S1(net1054),
    .X(_08569_));
 sg13g2_mux4_1 _15381_ (.S0(net905),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][6] ),
    .S1(net786),
    .X(_08570_));
 sg13g2_mux4_1 _15382_ (.S0(net905),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][6] ),
    .S1(net786),
    .X(_08571_));
 sg13g2_mux4_1 _15383_ (.S0(net904),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][6] ),
    .S1(net792),
    .X(_08572_));
 sg13g2_mux4_1 _15384_ (.S0(_08551_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][6] ),
    .S1(net792),
    .X(_08573_));
 sg13g2_mux4_1 _15385_ (.S0(net796),
    .A0(_08570_),
    .A1(_08571_),
    .A2(_08572_),
    .A3(_08573_),
    .S1(net1054),
    .X(_08574_));
 sg13g2_mux2_1 _15386_ (.A0(_08569_),
    .A1(_08574_),
    .S(net916),
    .X(_08575_));
 sg13g2_nand2b_1 _15387_ (.Y(_08576_),
    .B(_08575_),
    .A_N(net1049));
 sg13g2_buf_2 _15388_ (.A(_08576_),
    .X(_08577_));
 sg13g2_a22oi_1 _15389_ (.Y(_08578_),
    .B1(net613),
    .B2(\cpu.icache.r_tag[1][18] ),
    .A2(net795),
    .A1(\cpu.icache.r_tag[4][18] ));
 sg13g2_a22oi_1 _15390_ (.Y(_08579_),
    .B1(net614),
    .B2(\cpu.icache.r_tag[3][18] ),
    .A2(net537),
    .A1(\cpu.icache.r_tag[2][18] ));
 sg13g2_mux2_1 _15391_ (.A0(\cpu.icache.r_tag[5][18] ),
    .A1(\cpu.icache.r_tag[7][18] ),
    .S(net1052),
    .X(_08580_));
 sg13g2_nor2b_1 _15392_ (.A(_08288_),
    .B_N(net1052),
    .Y(_08581_));
 sg13g2_buf_2 _15393_ (.A(_08581_),
    .X(_08582_));
 sg13g2_a22oi_1 _15394_ (.Y(_08583_),
    .B1(_08582_),
    .B2(\cpu.icache.r_tag[6][18] ),
    .A2(_08580_),
    .A1(net1051));
 sg13g2_or2_1 _15395_ (.X(_08584_),
    .B(_08583_),
    .A(net908));
 sg13g2_nand4_1 _15396_ (.B(_08578_),
    .C(_08579_),
    .A(net620),
    .Y(_08585_),
    .D(_08584_));
 sg13g2_o21ai_1 _15397_ (.B1(_08585_),
    .Y(_08586_),
    .A1(\cpu.icache.r_tag[0][18] ),
    .A2(net540));
 sg13g2_xor2_1 _15398_ (.B(_08586_),
    .A(net436),
    .X(_08587_));
 sg13g2_nor3_1 _15399_ (.A(_08542_),
    .B(_08564_),
    .C(_08587_),
    .Y(_08588_));
 sg13g2_mux4_1 _15400_ (.S0(_08463_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][10] ),
    .S1(net791),
    .X(_08589_));
 sg13g2_mux4_1 _15401_ (.S0(_08463_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][10] ),
    .S1(_08349_),
    .X(_08590_));
 sg13g2_mux4_1 _15402_ (.S0(net904),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][10] ),
    .S1(net792),
    .X(_08591_));
 sg13g2_mux4_1 _15403_ (.S0(net904),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][10] ),
    .S1(net786),
    .X(_08592_));
 sg13g2_mux4_1 _15404_ (.S0(net796),
    .A0(_08589_),
    .A1(_08590_),
    .A2(_08591_),
    .A3(_08592_),
    .S1(net1054),
    .X(_08593_));
 sg13g2_mux4_1 _15405_ (.S0(net904),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][10] ),
    .S1(_08545_),
    .X(_08594_));
 sg13g2_mux4_1 _15406_ (.S0(net905),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][10] ),
    .S1(net786),
    .X(_08595_));
 sg13g2_mux4_1 _15407_ (.S0(_08262_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][10] ),
    .S1(net792),
    .X(_08596_));
 sg13g2_mux4_1 _15408_ (.S0(net904),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][10] ),
    .S1(_08337_),
    .X(_08597_));
 sg13g2_mux4_1 _15409_ (.S0(_08233_),
    .A0(_08594_),
    .A1(_08595_),
    .A2(_08596_),
    .A3(_08597_),
    .S1(net1054),
    .X(_08598_));
 sg13g2_mux2_1 _15410_ (.A0(_08593_),
    .A1(_08598_),
    .S(net916),
    .X(_08599_));
 sg13g2_nand2b_1 _15411_ (.Y(_08600_),
    .B(_08599_),
    .A_N(_08381_));
 sg13g2_buf_1 _15412_ (.A(_08600_),
    .X(_08601_));
 sg13g2_a22oi_1 _15413_ (.Y(_08602_),
    .B1(net795),
    .B2(\cpu.icache.r_tag[4][22] ),
    .A2(net537),
    .A1(\cpu.icache.r_tag[2][22] ));
 sg13g2_a22oi_1 _15414_ (.Y(_08603_),
    .B1(net617),
    .B2(\cpu.icache.r_tag[6][22] ),
    .A2(net698),
    .A1(\cpu.icache.r_tag[1][22] ));
 sg13g2_mux2_1 _15415_ (.A0(\cpu.icache.r_tag[7][22] ),
    .A1(\cpu.icache.r_tag[3][22] ),
    .S(net1053),
    .X(_08604_));
 sg13g2_buf_1 _15416_ (.A(net1052),
    .X(_08605_));
 sg13g2_a22oi_1 _15417_ (.Y(_08606_),
    .B1(_08604_),
    .B2(net903),
    .A2(net913),
    .A1(\cpu.icache.r_tag[5][22] ));
 sg13g2_nand2b_1 _15418_ (.Y(_08607_),
    .B(net912),
    .A_N(_08606_));
 sg13g2_nand4_1 _15419_ (.B(_08602_),
    .C(_08603_),
    .A(net620),
    .Y(_08608_),
    .D(_08607_));
 sg13g2_o21ai_1 _15420_ (.B1(_08608_),
    .Y(_08609_),
    .A1(\cpu.icache.r_tag[0][22] ),
    .A2(net541));
 sg13g2_xor2_1 _15421_ (.B(_08609_),
    .A(net435),
    .X(_08610_));
 sg13g2_buf_1 _15422_ (.A(\cpu.ex.pc[7] ),
    .X(_08611_));
 sg13g2_a22oi_1 _15423_ (.Y(_08612_),
    .B1(_08360_),
    .B2(\cpu.icache.r_tag[5][7] ),
    .A2(_08304_),
    .A1(\cpu.icache.r_tag[2][7] ));
 sg13g2_a22oi_1 _15424_ (.Y(_08613_),
    .B1(_08313_),
    .B2(\cpu.icache.r_tag[1][7] ),
    .A2(_08308_),
    .A1(\cpu.icache.r_tag[4][7] ));
 sg13g2_mux2_1 _15425_ (.A0(\cpu.icache.r_tag[7][7] ),
    .A1(\cpu.icache.r_tag[3][7] ),
    .S(net1116),
    .X(_08614_));
 sg13g2_a22oi_1 _15426_ (.Y(_08615_),
    .B1(_08614_),
    .B2(net1051),
    .A2(_08317_),
    .A1(\cpu.icache.r_tag[6][7] ));
 sg13g2_nand2b_1 _15427_ (.Y(_08616_),
    .B(net914),
    .A_N(_08615_));
 sg13g2_nand4_1 _15428_ (.B(_08612_),
    .C(_08613_),
    .A(_08295_),
    .Y(_08617_),
    .D(_08616_));
 sg13g2_o21ai_1 _15429_ (.B1(_08617_),
    .Y(_08618_),
    .A1(\cpu.icache.r_tag[0][7] ),
    .A2(net621));
 sg13g2_xor2_1 _15430_ (.B(_08618_),
    .A(_08611_),
    .X(_08619_));
 sg13g2_buf_1 _15431_ (.A(\cpu.ex.pc[8] ),
    .X(_08620_));
 sg13g2_a22oi_1 _15432_ (.Y(_08621_),
    .B1(net696),
    .B2(\cpu.icache.r_tag[5][8] ),
    .A2(net619),
    .A1(\cpu.icache.r_tag[2][8] ));
 sg13g2_a22oi_1 _15433_ (.Y(_08622_),
    .B1(net698),
    .B2(\cpu.icache.r_tag[1][8] ),
    .A2(_08308_),
    .A1(\cpu.icache.r_tag[4][8] ));
 sg13g2_mux2_1 _15434_ (.A0(\cpu.icache.r_tag[7][8] ),
    .A1(\cpu.icache.r_tag[3][8] ),
    .S(net1053),
    .X(_08623_));
 sg13g2_a22oi_1 _15435_ (.Y(_08624_),
    .B1(_08623_),
    .B2(net1051),
    .A2(_08317_),
    .A1(\cpu.icache.r_tag[6][8] ));
 sg13g2_nand2b_1 _15436_ (.Y(_08625_),
    .B(net903),
    .A_N(_08624_));
 sg13g2_nand4_1 _15437_ (.B(_08621_),
    .C(_08622_),
    .A(net621),
    .Y(_08626_),
    .D(_08625_));
 sg13g2_o21ai_1 _15438_ (.B1(_08626_),
    .Y(_08627_),
    .A1(\cpu.icache.r_tag[0][8] ),
    .A2(net620));
 sg13g2_xor2_1 _15439_ (.B(_08627_),
    .A(_08620_),
    .X(_08628_));
 sg13g2_buf_1 _15440_ (.A(\cpu.ex.pc[11] ),
    .X(_08629_));
 sg13g2_a22oi_1 _15441_ (.Y(_08630_),
    .B1(_08360_),
    .B2(\cpu.icache.r_tag[5][11] ),
    .A2(net619),
    .A1(\cpu.icache.r_tag[2][11] ));
 sg13g2_a22oi_1 _15442_ (.Y(_08631_),
    .B1(net698),
    .B2(\cpu.icache.r_tag[1][11] ),
    .A2(_08308_),
    .A1(\cpu.icache.r_tag[4][11] ));
 sg13g2_mux2_1 _15443_ (.A0(\cpu.icache.r_tag[7][11] ),
    .A1(\cpu.icache.r_tag[3][11] ),
    .S(net1053),
    .X(_08632_));
 sg13g2_a22oi_1 _15444_ (.Y(_08633_),
    .B1(_08632_),
    .B2(net1051),
    .A2(_08317_),
    .A1(\cpu.icache.r_tag[6][11] ));
 sg13g2_nand2b_1 _15445_ (.Y(_08634_),
    .B(net903),
    .A_N(_08633_));
 sg13g2_nand4_1 _15446_ (.B(_08630_),
    .C(_08631_),
    .A(net621),
    .Y(_08635_),
    .D(_08634_));
 sg13g2_o21ai_1 _15447_ (.B1(_08635_),
    .Y(_08636_),
    .A1(\cpu.icache.r_tag[0][11] ),
    .A2(net620));
 sg13g2_xor2_1 _15448_ (.B(_08636_),
    .A(_08629_),
    .X(_08637_));
 sg13g2_nand3_1 _15449_ (.B(_08628_),
    .C(_08637_),
    .A(_08619_),
    .Y(_08638_));
 sg13g2_buf_1 _15450_ (.A(\cpu.ex.pc[10] ),
    .X(_08639_));
 sg13g2_mux2_1 _15451_ (.A0(\cpu.icache.r_tag[4][10] ),
    .A1(\cpu.icache.r_tag[6][10] ),
    .S(net1052),
    .X(_08640_));
 sg13g2_a22oi_1 _15452_ (.Y(_08641_),
    .B1(_08640_),
    .B2(_08317_),
    .A2(_08372_),
    .A1(\cpu.icache.r_tag[3][10] ));
 sg13g2_a22oi_1 _15453_ (.Y(_08642_),
    .B1(_08360_),
    .B2(\cpu.icache.r_tag[5][10] ),
    .A2(_08304_),
    .A1(\cpu.icache.r_tag[2][10] ));
 sg13g2_a22oi_1 _15454_ (.Y(_08643_),
    .B1(_08366_),
    .B2(\cpu.icache.r_tag[7][10] ),
    .A2(_08313_),
    .A1(\cpu.icache.r_tag[1][10] ));
 sg13g2_nand4_1 _15455_ (.B(_08641_),
    .C(_08642_),
    .A(_08295_),
    .Y(_08644_),
    .D(_08643_));
 sg13g2_o21ai_1 _15456_ (.B1(_08644_),
    .Y(_08645_),
    .A1(\cpu.icache.r_tag[0][10] ),
    .A2(net621));
 sg13g2_xor2_1 _15457_ (.B(_08645_),
    .A(_08639_),
    .X(_08646_));
 sg13g2_inv_1 _15458_ (.Y(_08647_),
    .A(\cpu.ex.pc[6] ));
 sg13g2_buf_1 _15459_ (.A(_08647_),
    .X(_08648_));
 sg13g2_mux2_1 _15460_ (.A0(\cpu.icache.r_tag[4][6] ),
    .A1(\cpu.icache.r_tag[6][6] ),
    .S(_08323_),
    .X(_08649_));
 sg13g2_a22oi_1 _15461_ (.Y(_08650_),
    .B1(_08649_),
    .B2(_08317_),
    .A2(_08372_),
    .A1(\cpu.icache.r_tag[3][6] ));
 sg13g2_a22oi_1 _15462_ (.Y(_08651_),
    .B1(_08360_),
    .B2(\cpu.icache.r_tag[5][6] ),
    .A2(_08304_),
    .A1(\cpu.icache.r_tag[2][6] ));
 sg13g2_a22oi_1 _15463_ (.Y(_08652_),
    .B1(_08366_),
    .B2(\cpu.icache.r_tag[7][6] ),
    .A2(_08313_),
    .A1(\cpu.icache.r_tag[1][6] ));
 sg13g2_nand4_1 _15464_ (.B(_08650_),
    .C(_08651_),
    .A(_08295_),
    .Y(_08653_),
    .D(_08652_));
 sg13g2_o21ai_1 _15465_ (.B1(_08653_),
    .Y(_08654_),
    .A1(\cpu.icache.r_tag[0][6] ),
    .A2(net621));
 sg13g2_xnor2_1 _15466_ (.Y(_08655_),
    .A(net1047),
    .B(_08654_));
 sg13g2_buf_2 _15467_ (.A(\cpu.ex.pc[9] ),
    .X(_08656_));
 sg13g2_and2_1 _15468_ (.A(net1116),
    .B(_08293_),
    .X(_08657_));
 sg13g2_buf_1 _15469_ (.A(_08657_),
    .X(_08658_));
 sg13g2_mux2_1 _15470_ (.A0(\cpu.icache.r_tag[7][9] ),
    .A1(\cpu.icache.r_tag[3][9] ),
    .S(net1116),
    .X(_08659_));
 sg13g2_a22oi_1 _15471_ (.Y(_08660_),
    .B1(_08659_),
    .B2(net1052),
    .A2(_08327_),
    .A1(\cpu.icache.r_tag[5][9] ));
 sg13g2_nor2b_1 _15472_ (.A(_08289_),
    .B_N(\cpu.icache.r_tag[2][9] ),
    .Y(_08661_));
 sg13g2_a21o_1 _15473_ (.A2(\cpu.icache.r_tag[6][9] ),
    .A1(_08362_),
    .B1(_08661_),
    .X(_08662_));
 sg13g2_a221oi_1 _15474_ (.B2(net1052),
    .C1(net1051),
    .B1(_08662_),
    .A1(\cpu.icache.r_tag[4][9] ),
    .Y(_08663_),
    .A2(_08327_));
 sg13g2_a21oi_1 _15475_ (.A1(net1051),
    .A2(_08660_),
    .Y(_08664_),
    .B1(_08663_));
 sg13g2_a221oi_1 _15476_ (.B2(\cpu.icache.r_tag[1][9] ),
    .C1(_08664_),
    .B1(_08313_),
    .A1(\cpu.icache.r_tag[0][9] ),
    .Y(_08665_),
    .A2(_08658_));
 sg13g2_xnor2_1 _15477_ (.Y(_08666_),
    .A(_08656_),
    .B(_08665_));
 sg13g2_buf_1 _15478_ (.A(_08289_),
    .X(_08667_));
 sg13g2_mux4_1 _15479_ (.S0(net1051),
    .A0(\cpu.icache.r_valid[4] ),
    .A1(\cpu.icache.r_valid[5] ),
    .A2(\cpu.icache.r_valid[6] ),
    .A3(\cpu.icache.r_valid[7] ),
    .S1(_08605_),
    .X(_08668_));
 sg13g2_mux4_1 _15480_ (.S0(_08330_),
    .A0(\cpu.icache.r_valid[0] ),
    .A1(\cpu.icache.r_valid[1] ),
    .A2(\cpu.icache.r_valid[2] ),
    .A3(\cpu.icache.r_valid[3] ),
    .S1(_08324_),
    .X(_08669_));
 sg13g2_nor2b_1 _15481_ (.A(net1046),
    .B_N(_08669_),
    .Y(_08670_));
 sg13g2_a21oi_1 _15482_ (.A1(_08667_),
    .A2(_08668_),
    .Y(_08671_),
    .B1(_08670_));
 sg13g2_nor2_1 _15483_ (.A(_08666_),
    .B(_08671_),
    .Y(_08672_));
 sg13g2_buf_1 _15484_ (.A(\cpu.ex.pc[5] ),
    .X(_08673_));
 sg13g2_a22oi_1 _15485_ (.Y(_08674_),
    .B1(net795),
    .B2(\cpu.icache.r_tag[4][5] ),
    .A2(net619),
    .A1(\cpu.icache.r_tag[2][5] ));
 sg13g2_a22oi_1 _15486_ (.Y(_08675_),
    .B1(_08319_),
    .B2(\cpu.icache.r_tag[6][5] ),
    .A2(net698),
    .A1(\cpu.icache.r_tag[1][5] ));
 sg13g2_mux2_1 _15487_ (.A0(\cpu.icache.r_tag[7][5] ),
    .A1(\cpu.icache.r_tag[3][5] ),
    .S(net1053),
    .X(_08676_));
 sg13g2_a22oi_1 _15488_ (.Y(_08677_),
    .B1(_08676_),
    .B2(net914),
    .A2(_08327_),
    .A1(\cpu.icache.r_tag[5][5] ));
 sg13g2_nand2b_1 _15489_ (.Y(_08678_),
    .B(net912),
    .A_N(_08677_));
 sg13g2_nand4_1 _15490_ (.B(_08674_),
    .C(_08675_),
    .A(net621),
    .Y(_08679_),
    .D(_08678_));
 sg13g2_o21ai_1 _15491_ (.B1(_08679_),
    .Y(_08680_),
    .A1(\cpu.icache.r_tag[0][5] ),
    .A2(net620));
 sg13g2_xor2_1 _15492_ (.B(_08680_),
    .A(_08673_),
    .X(_08681_));
 sg13g2_nand4_1 _15493_ (.B(_08655_),
    .C(_08672_),
    .A(_08646_),
    .Y(_08682_),
    .D(_08681_));
 sg13g2_nor3_1 _15494_ (.A(_08610_),
    .B(_08638_),
    .C(_08682_),
    .Y(_08683_));
 sg13g2_nand4_1 _15495_ (.B(_08522_),
    .C(_08588_),
    .A(_08501_),
    .Y(_08684_),
    .D(_08683_));
 sg13g2_or4_1 _15496_ (.A(_08260_),
    .B(_08379_),
    .C(_08481_),
    .D(_08684_),
    .X(_08685_));
 sg13g2_buf_1 _15497_ (.A(_08685_),
    .X(_08686_));
 sg13g2_buf_1 _15498_ (.A(_08686_),
    .X(_08687_));
 sg13g2_buf_1 _15499_ (.A(net152),
    .X(_08688_));
 sg13g2_buf_1 _15500_ (.A(net470),
    .X(_08689_));
 sg13g2_nor2_1 _15501_ (.A(_00192_),
    .B(net434),
    .Y(_08690_));
 sg13g2_buf_1 _15502_ (.A(_08425_),
    .X(_08691_));
 sg13g2_mux2_1 _15503_ (.A0(\cpu.icache.r_data[7][31] ),
    .A1(\cpu.icache.r_data[3][31] ),
    .S(net785),
    .X(_08692_));
 sg13g2_buf_1 _15504_ (.A(_08325_),
    .X(_08693_));
 sg13g2_a22oi_1 _15505_ (.Y(_08694_),
    .B1(_08692_),
    .B2(net692),
    .A2(net913),
    .A1(\cpu.icache.r_data[5][31] ));
 sg13g2_buf_1 _15506_ (.A(_08332_),
    .X(_08695_));
 sg13g2_nand2b_1 _15507_ (.Y(_08696_),
    .B(net691),
    .A_N(_08694_));
 sg13g2_buf_1 _15508_ (.A(net618),
    .X(_08697_));
 sg13g2_buf_1 _15509_ (.A(net617),
    .X(_08698_));
 sg13g2_a22oi_1 _15510_ (.Y(_08699_),
    .B1(net534),
    .B2(\cpu.icache.r_data[6][31] ),
    .A2(net535),
    .A1(\cpu.icache.r_data[1][31] ));
 sg13g2_buf_1 _15511_ (.A(net539),
    .X(_08700_));
 sg13g2_buf_1 _15512_ (.A(net795),
    .X(_08701_));
 sg13g2_a22oi_1 _15513_ (.Y(_08702_),
    .B1(net690),
    .B2(\cpu.icache.r_data[4][31] ),
    .A2(net468),
    .A1(\cpu.icache.r_data[2][31] ));
 sg13g2_nand3_1 _15514_ (.B(_08699_),
    .C(_08702_),
    .A(_08696_),
    .Y(_08703_));
 sg13g2_buf_1 _15515_ (.A(\cpu.ex.pc[1] ),
    .X(_08704_));
 sg13g2_buf_1 _15516_ (.A(_08704_),
    .X(_08705_));
 sg13g2_buf_1 _15517_ (.A(net1045),
    .X(_08706_));
 sg13g2_buf_1 _15518_ (.A(_08706_),
    .X(_08707_));
 sg13g2_o21ai_1 _15519_ (.B1(net784),
    .Y(_08708_),
    .A1(_08690_),
    .A2(_08703_));
 sg13g2_inv_1 _15520_ (.Y(_08709_),
    .A(_08704_));
 sg13g2_buf_1 _15521_ (.A(_08658_),
    .X(_08710_));
 sg13g2_nand2_1 _15522_ (.Y(_08711_),
    .A(_00191_),
    .B(net612));
 sg13g2_buf_1 _15523_ (.A(net696),
    .X(_08712_));
 sg13g2_and2_1 _15524_ (.A(\cpu.icache.r_data[4][15] ),
    .B(net690),
    .X(_08713_));
 sg13g2_a221oi_1 _15525_ (.B2(\cpu.icache.r_data[5][15] ),
    .C1(_08713_),
    .B1(net611),
    .A1(\cpu.icache.r_data[1][15] ),
    .Y(_08714_),
    .A2(_08697_));
 sg13g2_a22oi_1 _15526_ (.Y(_08715_),
    .B1(net615),
    .B2(\cpu.icache.r_data[7][15] ),
    .A2(net468),
    .A1(\cpu.icache.r_data[2][15] ));
 sg13g2_buf_1 _15527_ (.A(net536),
    .X(_08716_));
 sg13g2_a22oi_1 _15528_ (.Y(_08717_),
    .B1(net467),
    .B2(\cpu.icache.r_data[3][15] ),
    .A2(net534),
    .A1(\cpu.icache.r_data[6][15] ));
 sg13g2_nand4_1 _15529_ (.B(_08714_),
    .C(_08715_),
    .A(net434),
    .Y(_08718_),
    .D(_08717_));
 sg13g2_nand3_1 _15530_ (.B(_08711_),
    .C(_08718_),
    .A(net1044),
    .Y(_08719_));
 sg13g2_and2_1 _15531_ (.A(_08708_),
    .B(_08719_),
    .X(_08720_));
 sg13g2_buf_1 _15532_ (.A(_08720_),
    .X(_08721_));
 sg13g2_nand2_1 _15533_ (.Y(_08722_),
    .A(\cpu.icache.r_data[4][13] ),
    .B(_08308_));
 sg13g2_a22oi_1 _15534_ (.Y(_08723_),
    .B1(_08360_),
    .B2(\cpu.icache.r_data[5][13] ),
    .A2(_08313_),
    .A1(\cpu.icache.r_data[1][13] ));
 sg13g2_a22oi_1 _15535_ (.Y(_08724_),
    .B1(_08366_),
    .B2(\cpu.icache.r_data[7][13] ),
    .A2(_08304_),
    .A1(\cpu.icache.r_data[2][13] ));
 sg13g2_a22oi_1 _15536_ (.Y(_08725_),
    .B1(net614),
    .B2(\cpu.icache.r_data[3][13] ),
    .A2(_08319_),
    .A1(\cpu.icache.r_data[6][13] ));
 sg13g2_nand4_1 _15537_ (.B(_08723_),
    .C(_08724_),
    .A(_08722_),
    .Y(_08726_),
    .D(_08725_));
 sg13g2_mux2_1 _15538_ (.A0(\cpu.icache.r_data[0][13] ),
    .A1(_08726_),
    .S(net621),
    .X(_08727_));
 sg13g2_mux2_1 _15539_ (.A0(\cpu.icache.r_data[7][29] ),
    .A1(\cpu.icache.r_data[3][29] ),
    .S(_08287_),
    .X(_08728_));
 sg13g2_a22oi_1 _15540_ (.Y(_08729_),
    .B1(_08728_),
    .B2(net903),
    .A2(net913),
    .A1(\cpu.icache.r_data[5][29] ));
 sg13g2_nand2b_1 _15541_ (.Y(_08730_),
    .B(net912),
    .A_N(_08729_));
 sg13g2_a22oi_1 _15542_ (.Y(_08731_),
    .B1(_08319_),
    .B2(\cpu.icache.r_data[6][29] ),
    .A2(_08304_),
    .A1(\cpu.icache.r_data[2][29] ));
 sg13g2_a22oi_1 _15543_ (.Y(_08732_),
    .B1(_08313_),
    .B2(\cpu.icache.r_data[1][29] ),
    .A2(_08308_),
    .A1(\cpu.icache.r_data[4][29] ));
 sg13g2_nand2_1 _15544_ (.Y(_08733_),
    .A(_08731_),
    .B(_08732_));
 sg13g2_a21oi_1 _15545_ (.A1(\cpu.icache.r_data[0][29] ),
    .A2(_08658_),
    .Y(_08734_),
    .B1(_08733_));
 sg13g2_nand3_1 _15546_ (.B(_08730_),
    .C(_08734_),
    .A(net1045),
    .Y(_08735_));
 sg13g2_o21ai_1 _15547_ (.B1(_08735_),
    .Y(_08736_),
    .A1(net1045),
    .A2(_08727_));
 sg13g2_buf_1 _15548_ (.A(_08736_),
    .X(_08737_));
 sg13g2_nor2_1 _15549_ (.A(_00190_),
    .B(net541),
    .Y(_08738_));
 sg13g2_buf_1 _15550_ (.A(net785),
    .X(_08739_));
 sg13g2_mux2_1 _15551_ (.A0(\cpu.icache.r_data[5][30] ),
    .A1(\cpu.icache.r_data[7][30] ),
    .S(net914),
    .X(_08740_));
 sg13g2_nor2_1 _15552_ (.A(_08288_),
    .B(net1115),
    .Y(_08741_));
 sg13g2_buf_2 _15553_ (.A(_08741_),
    .X(_08742_));
 sg13g2_a22oi_1 _15554_ (.Y(_08743_),
    .B1(_08742_),
    .B2(\cpu.icache.r_data[4][30] ),
    .A2(_08740_),
    .A1(net912));
 sg13g2_nor2_1 _15555_ (.A(net689),
    .B(_08743_),
    .Y(_08744_));
 sg13g2_a22oi_1 _15556_ (.Y(_08745_),
    .B1(net614),
    .B2(\cpu.icache.r_data[3][30] ),
    .A2(net617),
    .A1(\cpu.icache.r_data[6][30] ));
 sg13g2_a22oi_1 _15557_ (.Y(_08746_),
    .B1(net613),
    .B2(\cpu.icache.r_data[1][30] ),
    .A2(net537),
    .A1(\cpu.icache.r_data[2][30] ));
 sg13g2_nand2_1 _15558_ (.Y(_08747_),
    .A(_08745_),
    .B(_08746_));
 sg13g2_nor3_1 _15559_ (.A(_08738_),
    .B(_08744_),
    .C(_08747_),
    .Y(_08748_));
 sg13g2_nand2_1 _15560_ (.Y(_08749_),
    .A(_00189_),
    .B(_08658_));
 sg13g2_nor2b_1 _15561_ (.A(net914),
    .B_N(\cpu.icache.r_data[4][14] ),
    .Y(_08750_));
 sg13g2_a21oi_1 _15562_ (.A1(net914),
    .A2(\cpu.icache.r_data[6][14] ),
    .Y(_08751_),
    .B1(_08750_));
 sg13g2_nor2_2 _15563_ (.A(net915),
    .B(net1052),
    .Y(_08752_));
 sg13g2_a22oi_1 _15564_ (.Y(_08753_),
    .B1(_08364_),
    .B2(\cpu.icache.r_data[7][14] ),
    .A2(_08752_),
    .A1(\cpu.icache.r_data[5][14] ));
 sg13g2_o21ai_1 _15565_ (.B1(_08753_),
    .Y(_08754_),
    .A1(net912),
    .A2(_08751_));
 sg13g2_nand2_1 _15566_ (.Y(_08755_),
    .A(net1050),
    .B(_08754_));
 sg13g2_nand2_1 _15567_ (.Y(_08756_),
    .A(\cpu.icache.r_data[1][14] ),
    .B(_08402_));
 sg13g2_a22oi_1 _15568_ (.Y(_08757_),
    .B1(net614),
    .B2(\cpu.icache.r_data[3][14] ),
    .A2(net537),
    .A1(\cpu.icache.r_data[2][14] ));
 sg13g2_nand4_1 _15569_ (.B(_08755_),
    .C(_08756_),
    .A(net541),
    .Y(_08758_),
    .D(_08757_));
 sg13g2_a21oi_1 _15570_ (.A1(_08749_),
    .A2(_08758_),
    .Y(_08759_),
    .B1(net1045));
 sg13g2_a21o_1 _15571_ (.A2(_08748_),
    .A1(net784),
    .B1(_08759_),
    .X(_08760_));
 sg13g2_buf_1 _15572_ (.A(_08760_),
    .X(_08761_));
 sg13g2_nand2_2 _15573_ (.Y(_08762_),
    .A(net305),
    .B(_08761_));
 sg13g2_nor2_1 _15574_ (.A(_08721_),
    .B(_08762_),
    .Y(_08763_));
 sg13g2_buf_1 _15575_ (.A(_08763_),
    .X(_08764_));
 sg13g2_buf_1 _15576_ (.A(_08764_),
    .X(_08765_));
 sg13g2_buf_1 _15577_ (.A(net784),
    .X(_08766_));
 sg13g2_mux2_1 _15578_ (.A0(\cpu.icache.r_data[7][16] ),
    .A1(\cpu.icache.r_data[3][16] ),
    .S(net785),
    .X(_08767_));
 sg13g2_a22oi_1 _15579_ (.Y(_08768_),
    .B1(_08767_),
    .B2(net692),
    .A2(net913),
    .A1(\cpu.icache.r_data[5][16] ));
 sg13g2_nand2b_1 _15580_ (.Y(_08769_),
    .B(net691),
    .A_N(_08768_));
 sg13g2_buf_1 _15581_ (.A(_08698_),
    .X(_08770_));
 sg13g2_a22oi_1 _15582_ (.Y(_08771_),
    .B1(net466),
    .B2(\cpu.icache.r_data[6][16] ),
    .A2(net690),
    .A1(\cpu.icache.r_data[4][16] ));
 sg13g2_a22oi_1 _15583_ (.Y(_08772_),
    .B1(net535),
    .B2(\cpu.icache.r_data[1][16] ),
    .A2(net468),
    .A1(\cpu.icache.r_data[2][16] ));
 sg13g2_nand3_1 _15584_ (.B(_08771_),
    .C(_08772_),
    .A(_08769_),
    .Y(_08773_));
 sg13g2_a21oi_1 _15585_ (.A1(\cpu.icache.r_data[0][16] ),
    .A2(net612),
    .Y(_08774_),
    .B1(_08773_));
 sg13g2_mux2_1 _15586_ (.A0(\cpu.icache.r_data[4][0] ),
    .A1(\cpu.icache.r_data[6][0] ),
    .S(net794),
    .X(_08775_));
 sg13g2_a22oi_1 _15587_ (.Y(_08776_),
    .B1(_08775_),
    .B2(_08317_),
    .A2(net467),
    .A1(\cpu.icache.r_data[3][0] ));
 sg13g2_a22oi_1 _15588_ (.Y(_08777_),
    .B1(net535),
    .B2(\cpu.icache.r_data[1][0] ),
    .A2(net468),
    .A1(\cpu.icache.r_data[2][0] ));
 sg13g2_a22oi_1 _15589_ (.Y(_08778_),
    .B1(net615),
    .B2(\cpu.icache.r_data[7][0] ),
    .A2(net611),
    .A1(\cpu.icache.r_data[5][0] ));
 sg13g2_nand4_1 _15590_ (.B(_08776_),
    .C(_08777_),
    .A(net434),
    .Y(_08779_),
    .D(_08778_));
 sg13g2_o21ai_1 _15591_ (.B1(_08779_),
    .Y(_08780_),
    .A1(\cpu.icache.r_data[0][0] ),
    .A2(net434));
 sg13g2_and2_1 _15592_ (.A(net1044),
    .B(_08780_),
    .X(_08781_));
 sg13g2_a21o_1 _15593_ (.A2(_08774_),
    .A1(_08766_),
    .B1(_08781_),
    .X(_08782_));
 sg13g2_buf_1 _15594_ (.A(_08782_),
    .X(_08783_));
 sg13g2_buf_1 _15595_ (.A(_08358_),
    .X(_08784_));
 sg13g2_buf_1 _15596_ (.A(_08402_),
    .X(_08785_));
 sg13g2_a22oi_1 _15597_ (.Y(_08786_),
    .B1(net533),
    .B2(\cpu.icache.r_data[1][1] ),
    .A2(_08784_),
    .A1(\cpu.icache.r_data[2][1] ));
 sg13g2_a22oi_1 _15598_ (.Y(_08787_),
    .B1(net467),
    .B2(\cpu.icache.r_data[3][1] ),
    .A2(_08321_),
    .A1(\cpu.icache.r_data[6][1] ));
 sg13g2_mux2_1 _15599_ (.A0(\cpu.icache.r_data[5][1] ),
    .A1(\cpu.icache.r_data[7][1] ),
    .S(net903),
    .X(_08788_));
 sg13g2_a22oi_1 _15600_ (.Y(_08789_),
    .B1(_08788_),
    .B2(net793),
    .A2(_08742_),
    .A1(\cpu.icache.r_data[4][1] ));
 sg13g2_or2_1 _15601_ (.X(_08790_),
    .B(_08789_),
    .A(net689));
 sg13g2_nand3_1 _15602_ (.B(_08787_),
    .C(_08790_),
    .A(_08786_),
    .Y(_08791_));
 sg13g2_mux2_1 _15603_ (.A0(\cpu.icache.r_data[0][1] ),
    .A1(_08791_),
    .S(net471),
    .X(_08792_));
 sg13g2_mux2_1 _15604_ (.A0(\cpu.icache.r_data[7][17] ),
    .A1(\cpu.icache.r_data[3][17] ),
    .S(_08691_),
    .X(_08793_));
 sg13g2_a22oi_1 _15605_ (.Y(_08794_),
    .B1(_08793_),
    .B2(net692),
    .A2(net913),
    .A1(\cpu.icache.r_data[5][17] ));
 sg13g2_nand2b_1 _15606_ (.Y(_08795_),
    .B(_08695_),
    .A_N(_08794_));
 sg13g2_a22oi_1 _15607_ (.Y(_08796_),
    .B1(_08698_),
    .B2(\cpu.icache.r_data[6][17] ),
    .A2(net465),
    .A1(\cpu.icache.r_data[2][17] ));
 sg13g2_a22oi_1 _15608_ (.Y(_08797_),
    .B1(net533),
    .B2(\cpu.icache.r_data[1][17] ),
    .A2(net690),
    .A1(\cpu.icache.r_data[4][17] ));
 sg13g2_nand2_1 _15609_ (.Y(_08798_),
    .A(_08796_),
    .B(_08797_));
 sg13g2_a21oi_1 _15610_ (.A1(\cpu.icache.r_data[0][17] ),
    .A2(net612),
    .Y(_08799_),
    .B1(_08798_));
 sg13g2_nand3_1 _15611_ (.B(_08795_),
    .C(_08799_),
    .A(net902),
    .Y(_08800_));
 sg13g2_o21ai_1 _15612_ (.B1(_08800_),
    .Y(_08801_),
    .A1(net902),
    .A2(_08792_));
 sg13g2_buf_1 _15613_ (.A(_08801_),
    .X(_08802_));
 sg13g2_inv_1 _15614_ (.Y(_08803_),
    .A(_08802_));
 sg13g2_buf_1 _15615_ (.A(_08803_),
    .X(_08804_));
 sg13g2_nor2_1 _15616_ (.A(net212),
    .B(net150),
    .Y(_08805_));
 sg13g2_buf_1 _15617_ (.A(_08805_),
    .X(_08806_));
 sg13g2_nand2_2 _15618_ (.Y(_08807_),
    .A(net151),
    .B(_08806_));
 sg13g2_a22oi_1 _15619_ (.Y(_08808_),
    .B1(_08320_),
    .B2(\cpu.icache.r_data[6][6] ),
    .A2(net698),
    .A1(\cpu.icache.r_data[1][6] ));
 sg13g2_a22oi_1 _15620_ (.Y(_08809_),
    .B1(net614),
    .B2(\cpu.icache.r_data[3][6] ),
    .A2(net619),
    .A1(\cpu.icache.r_data[2][6] ));
 sg13g2_mux2_1 _15621_ (.A0(\cpu.icache.r_data[5][6] ),
    .A1(\cpu.icache.r_data[7][6] ),
    .S(net1052),
    .X(_08810_));
 sg13g2_a22oi_1 _15622_ (.Y(_08811_),
    .B1(_08810_),
    .B2(_08330_),
    .A2(_08742_),
    .A1(\cpu.icache.r_data[4][6] ));
 sg13g2_or2_1 _15623_ (.X(_08812_),
    .B(_08811_),
    .A(net908));
 sg13g2_and4_1 _15624_ (.A(_08299_),
    .B(_08808_),
    .C(_08809_),
    .D(_08812_),
    .X(_08813_));
 sg13g2_a21oi_1 _15625_ (.A1(_00195_),
    .A2(_08658_),
    .Y(_08814_),
    .B1(_08813_));
 sg13g2_nor2_1 _15626_ (.A(_00196_),
    .B(net620),
    .Y(_08815_));
 sg13g2_mux2_1 _15627_ (.A0(\cpu.icache.r_data[5][22] ),
    .A1(\cpu.icache.r_data[7][22] ),
    .S(_08324_),
    .X(_08816_));
 sg13g2_a22oi_1 _15628_ (.Y(_08817_),
    .B1(_08816_),
    .B2(net912),
    .A2(_08742_),
    .A1(\cpu.icache.r_data[4][22] ));
 sg13g2_nor2_1 _15629_ (.A(net785),
    .B(_08817_),
    .Y(_08818_));
 sg13g2_a22oi_1 _15630_ (.Y(_08819_),
    .B1(net617),
    .B2(\cpu.icache.r_data[6][22] ),
    .A2(net537),
    .A1(\cpu.icache.r_data[2][22] ));
 sg13g2_a22oi_1 _15631_ (.Y(_08820_),
    .B1(_08373_),
    .B2(\cpu.icache.r_data[3][22] ),
    .A2(net698),
    .A1(\cpu.icache.r_data[1][22] ));
 sg13g2_nand2_1 _15632_ (.Y(_08821_),
    .A(_08819_),
    .B(_08820_));
 sg13g2_or4_1 _15633_ (.A(net1044),
    .B(_08815_),
    .C(_08818_),
    .D(_08821_),
    .X(_08822_));
 sg13g2_o21ai_1 _15634_ (.B1(_08822_),
    .Y(_08823_),
    .A1(net1045),
    .A2(_08814_));
 sg13g2_buf_1 _15635_ (.A(_08823_),
    .X(_08824_));
 sg13g2_inv_1 _15636_ (.Y(_08825_),
    .A(_00193_));
 sg13g2_a22oi_1 _15637_ (.Y(_08826_),
    .B1(_08360_),
    .B2(\cpu.icache.r_data[5][5] ),
    .A2(_08314_),
    .A1(\cpu.icache.r_data[1][5] ));
 sg13g2_a22oi_1 _15638_ (.Y(_08827_),
    .B1(_08373_),
    .B2(\cpu.icache.r_data[3][5] ),
    .A2(net619),
    .A1(\cpu.icache.r_data[2][5] ));
 sg13g2_mux2_1 _15639_ (.A0(\cpu.icache.r_data[4][5] ),
    .A1(\cpu.icache.r_data[6][5] ),
    .S(_08290_),
    .X(_08828_));
 sg13g2_a22oi_1 _15640_ (.Y(_08829_),
    .B1(_08828_),
    .B2(net915),
    .A2(_08364_),
    .A1(\cpu.icache.r_data[7][5] ));
 sg13g2_or2_1 _15641_ (.X(_08830_),
    .B(_08829_),
    .A(net908));
 sg13g2_nand4_1 _15642_ (.B(_08826_),
    .C(_08827_),
    .A(net621),
    .Y(_08831_),
    .D(_08830_));
 sg13g2_o21ai_1 _15643_ (.B1(_08831_),
    .Y(_08832_),
    .A1(_08825_),
    .A2(_08299_));
 sg13g2_mux2_1 _15644_ (.A0(\cpu.icache.r_data[7][21] ),
    .A1(\cpu.icache.r_data[3][21] ),
    .S(_08287_),
    .X(_08833_));
 sg13g2_a22oi_1 _15645_ (.Y(_08834_),
    .B1(_08364_),
    .B2(_08833_),
    .A2(_08319_),
    .A1(\cpu.icache.r_data[6][21] ));
 sg13g2_a22oi_1 _15646_ (.Y(_08835_),
    .B1(_08309_),
    .B2(\cpu.icache.r_data[4][21] ),
    .A2(net619),
    .A1(\cpu.icache.r_data[2][21] ));
 sg13g2_a22oi_1 _15647_ (.Y(_08836_),
    .B1(_08360_),
    .B2(\cpu.icache.r_data[5][21] ),
    .A2(_08314_),
    .A1(\cpu.icache.r_data[1][21] ));
 sg13g2_nand3_1 _15648_ (.B(_08835_),
    .C(_08836_),
    .A(_08834_),
    .Y(_08837_));
 sg13g2_nor2_1 _15649_ (.A(_00194_),
    .B(_08296_),
    .Y(_08838_));
 sg13g2_o21ai_1 _15650_ (.B1(net1045),
    .Y(_08839_),
    .A1(_08837_),
    .A2(_08838_));
 sg13g2_o21ai_1 _15651_ (.B1(_08839_),
    .Y(_08840_),
    .A1(net1045),
    .A2(_08832_));
 sg13g2_buf_1 _15652_ (.A(_08840_),
    .X(_08841_));
 sg13g2_inv_1 _15653_ (.Y(_08842_),
    .A(_08841_));
 sg13g2_nand2_2 _15654_ (.Y(_08843_),
    .A(_08824_),
    .B(_08842_));
 sg13g2_inv_1 _15655_ (.Y(_08844_),
    .A(_00187_));
 sg13g2_a22oi_1 _15656_ (.Y(_08845_),
    .B1(net611),
    .B2(\cpu.icache.r_data[5][11] ),
    .A2(net533),
    .A1(\cpu.icache.r_data[1][11] ));
 sg13g2_a22oi_1 _15657_ (.Y(_08846_),
    .B1(net467),
    .B2(\cpu.icache.r_data[3][11] ),
    .A2(net465),
    .A1(\cpu.icache.r_data[2][11] ));
 sg13g2_mux2_1 _15658_ (.A0(\cpu.icache.r_data[4][11] ),
    .A1(\cpu.icache.r_data[6][11] ),
    .S(net903),
    .X(_08847_));
 sg13g2_a22oi_1 _15659_ (.Y(_08848_),
    .B1(_08847_),
    .B2(net915),
    .A2(net788),
    .A1(\cpu.icache.r_data[7][11] ));
 sg13g2_or2_1 _15660_ (.X(_08849_),
    .B(_08848_),
    .A(_08739_));
 sg13g2_nand4_1 _15661_ (.B(_08845_),
    .C(_08846_),
    .A(net471),
    .Y(_08850_),
    .D(_08849_));
 sg13g2_o21ai_1 _15662_ (.B1(_08850_),
    .Y(_08851_),
    .A1(_08844_),
    .A2(net434));
 sg13g2_nand2_1 _15663_ (.Y(_08852_),
    .A(\cpu.icache.r_data[2][27] ),
    .B(net465));
 sg13g2_a22oi_1 _15664_ (.Y(_08853_),
    .B1(net533),
    .B2(\cpu.icache.r_data[1][27] ),
    .A2(_08701_),
    .A1(\cpu.icache.r_data[4][27] ));
 sg13g2_a22oi_1 _15665_ (.Y(_08854_),
    .B1(net615),
    .B2(\cpu.icache.r_data[7][27] ),
    .A2(_08712_),
    .A1(\cpu.icache.r_data[5][27] ));
 sg13g2_a22oi_1 _15666_ (.Y(_08855_),
    .B1(net467),
    .B2(\cpu.icache.r_data[3][27] ),
    .A2(net534),
    .A1(\cpu.icache.r_data[6][27] ));
 sg13g2_nand4_1 _15667_ (.B(_08853_),
    .C(_08854_),
    .A(_08852_),
    .Y(_08856_),
    .D(_08855_));
 sg13g2_nor2_1 _15668_ (.A(_00188_),
    .B(net471),
    .Y(_08857_));
 sg13g2_o21ai_1 _15669_ (.B1(net902),
    .Y(_08858_),
    .A1(_08856_),
    .A2(_08857_));
 sg13g2_o21ai_1 _15670_ (.B1(_08858_),
    .Y(_08859_),
    .A1(net784),
    .A2(_08851_));
 sg13g2_buf_1 _15671_ (.A(_08859_),
    .X(_08860_));
 sg13g2_nor2_1 _15672_ (.A(_00186_),
    .B(net471),
    .Y(_08861_));
 sg13g2_mux2_1 _15673_ (.A0(\cpu.icache.r_data[4][26] ),
    .A1(\cpu.icache.r_data[6][26] ),
    .S(net794),
    .X(_08862_));
 sg13g2_a22oi_1 _15674_ (.Y(_08863_),
    .B1(_08862_),
    .B2(net915),
    .A2(net788),
    .A1(\cpu.icache.r_data[7][26] ));
 sg13g2_nor2_1 _15675_ (.A(net689),
    .B(_08863_),
    .Y(_08864_));
 sg13g2_a22oi_1 _15676_ (.Y(_08865_),
    .B1(_08716_),
    .B2(\cpu.icache.r_data[3][26] ),
    .A2(net468),
    .A1(\cpu.icache.r_data[2][26] ));
 sg13g2_a22oi_1 _15677_ (.Y(_08866_),
    .B1(net611),
    .B2(\cpu.icache.r_data[5][26] ),
    .A2(net535),
    .A1(\cpu.icache.r_data[1][26] ));
 sg13g2_nand2_1 _15678_ (.Y(_08867_),
    .A(_08865_),
    .B(_08866_));
 sg13g2_nor3_1 _15679_ (.A(_08861_),
    .B(_08864_),
    .C(_08867_),
    .Y(_08868_));
 sg13g2_nand2_1 _15680_ (.Y(_08869_),
    .A(_00185_),
    .B(net612));
 sg13g2_a22oi_1 _15681_ (.Y(_08870_),
    .B1(net534),
    .B2(\cpu.icache.r_data[6][10] ),
    .A2(net533),
    .A1(\cpu.icache.r_data[1][10] ));
 sg13g2_a22oi_1 _15682_ (.Y(_08871_),
    .B1(_08701_),
    .B2(\cpu.icache.r_data[4][10] ),
    .A2(net465),
    .A1(\cpu.icache.r_data[2][10] ));
 sg13g2_mux2_1 _15683_ (.A0(\cpu.icache.r_data[7][10] ),
    .A1(\cpu.icache.r_data[3][10] ),
    .S(_08425_),
    .X(_08872_));
 sg13g2_a22oi_1 _15684_ (.Y(_08873_),
    .B1(_08872_),
    .B2(net692),
    .A2(_08328_),
    .A1(\cpu.icache.r_data[5][10] ));
 sg13g2_nand2b_1 _15685_ (.Y(_08874_),
    .B(net793),
    .A_N(_08873_));
 sg13g2_nand4_1 _15686_ (.B(_08870_),
    .C(_08871_),
    .A(_08689_),
    .Y(_08875_),
    .D(_08874_));
 sg13g2_a21oi_1 _15687_ (.A1(_08869_),
    .A2(_08875_),
    .Y(_08876_),
    .B1(net902));
 sg13g2_a21oi_1 _15688_ (.A1(net784),
    .A2(_08868_),
    .Y(_08877_),
    .B1(_08876_));
 sg13g2_buf_1 _15689_ (.A(_08877_),
    .X(_08878_));
 sg13g2_nand2_1 _15690_ (.Y(_08879_),
    .A(_08860_),
    .B(_08878_));
 sg13g2_nor4_1 _15691_ (.A(_08687_),
    .B(_08807_),
    .C(_08843_),
    .D(_08879_),
    .Y(_08880_));
 sg13g2_a21o_1 _15692_ (.A2(_08688_),
    .A1(_08122_),
    .B1(_08880_),
    .X(_00017_));
 sg13g2_buf_1 _15693_ (.A(\cpu.dec.r_op[4] ),
    .X(_08881_));
 sg13g2_buf_1 _15694_ (.A(net1114),
    .X(_08882_));
 sg13g2_buf_1 _15695_ (.A(net152),
    .X(_08883_));
 sg13g2_nor2_1 _15696_ (.A(_00198_),
    .B(net434),
    .Y(_08884_));
 sg13g2_mux2_1 _15697_ (.A0(\cpu.icache.r_data[5][28] ),
    .A1(\cpu.icache.r_data[7][28] ),
    .S(net692),
    .X(_08885_));
 sg13g2_a22oi_1 _15698_ (.Y(_08886_),
    .B1(_08885_),
    .B2(_08695_),
    .A2(_08582_),
    .A1(\cpu.icache.r_data[6][28] ));
 sg13g2_nor2_1 _15699_ (.A(net689),
    .B(_08886_),
    .Y(_08887_));
 sg13g2_buf_1 _15700_ (.A(net690),
    .X(_08888_));
 sg13g2_buf_2 _15701_ (.A(net467),
    .X(_08889_));
 sg13g2_a22oi_1 _15702_ (.Y(_08890_),
    .B1(net433),
    .B2(\cpu.icache.r_data[3][28] ),
    .A2(net610),
    .A1(\cpu.icache.r_data[4][28] ));
 sg13g2_a22oi_1 _15703_ (.Y(_08891_),
    .B1(net535),
    .B2(\cpu.icache.r_data[1][28] ),
    .A2(net468),
    .A1(\cpu.icache.r_data[2][28] ));
 sg13g2_nand2_1 _15704_ (.Y(_08892_),
    .A(_08890_),
    .B(_08891_));
 sg13g2_nor3_1 _15705_ (.A(_08884_),
    .B(_08887_),
    .C(_08892_),
    .Y(_08893_));
 sg13g2_nand2_1 _15706_ (.Y(_08894_),
    .A(_00197_),
    .B(_08710_));
 sg13g2_and2_1 _15707_ (.A(\cpu.icache.r_data[4][12] ),
    .B(net690),
    .X(_08895_));
 sg13g2_a221oi_1 _15708_ (.B2(\cpu.icache.r_data[5][12] ),
    .C1(_08895_),
    .B1(net611),
    .A1(\cpu.icache.r_data[1][12] ),
    .Y(_08896_),
    .A2(_08697_));
 sg13g2_a22oi_1 _15709_ (.Y(_08897_),
    .B1(net615),
    .B2(\cpu.icache.r_data[7][12] ),
    .A2(_08700_),
    .A1(\cpu.icache.r_data[2][12] ));
 sg13g2_a22oi_1 _15710_ (.Y(_08898_),
    .B1(_08889_),
    .B2(\cpu.icache.r_data[3][12] ),
    .A2(net534),
    .A1(\cpu.icache.r_data[6][12] ));
 sg13g2_nand4_1 _15711_ (.B(_08896_),
    .C(_08897_),
    .A(net434),
    .Y(_08899_),
    .D(_08898_));
 sg13g2_a21oi_1 _15712_ (.A1(_08894_),
    .A2(_08899_),
    .Y(_08900_),
    .B1(_08707_));
 sg13g2_a21oi_2 _15713_ (.B1(_08900_),
    .Y(_08901_),
    .A2(_08893_),
    .A1(net784));
 sg13g2_buf_1 _15714_ (.A(_08901_),
    .X(_08902_));
 sg13g2_nand3_1 _15715_ (.B(net234),
    .C(net211),
    .A(_08860_),
    .Y(_08903_));
 sg13g2_buf_1 _15716_ (.A(_08903_),
    .X(_08904_));
 sg13g2_buf_1 _15717_ (.A(_08802_),
    .X(_08905_));
 sg13g2_nor2_1 _15718_ (.A(net212),
    .B(net186),
    .Y(_08906_));
 sg13g2_nand2_1 _15719_ (.Y(_08907_),
    .A(_08764_),
    .B(_08906_));
 sg13g2_buf_1 _15720_ (.A(_08907_),
    .X(_08908_));
 sg13g2_nor4_1 _15721_ (.A(net187),
    .B(_08843_),
    .C(_08904_),
    .D(_08908_),
    .Y(_08909_));
 sg13g2_a21o_1 _15722_ (.A2(_08883_),
    .A1(net1043),
    .B1(_08909_),
    .X(_00015_));
 sg13g2_buf_1 _15723_ (.A(\cpu.dec.r_op[5] ),
    .X(_08910_));
 sg13g2_buf_1 _15724_ (.A(_08910_),
    .X(_08911_));
 sg13g2_buf_1 _15725_ (.A(_08860_),
    .X(_08912_));
 sg13g2_inv_2 _15726_ (.Y(_08913_),
    .A(_08878_));
 sg13g2_nor4_1 _15727_ (.A(net187),
    .B(_08807_),
    .C(net210),
    .D(_08913_),
    .Y(_08914_));
 sg13g2_a21o_1 _15728_ (.A2(net122),
    .A1(_08911_),
    .B1(_08914_),
    .X(_00016_));
 sg13g2_inv_1 _15729_ (.Y(_08915_),
    .A(\cpu.dec.r_op[7] ));
 sg13g2_and4_1 _15730_ (.A(_08646_),
    .B(_08655_),
    .C(_08619_),
    .D(_08672_),
    .X(_08916_));
 sg13g2_nand4_1 _15731_ (.B(_08628_),
    .C(_08637_),
    .A(_08916_),
    .Y(_08917_),
    .D(_08681_));
 sg13g2_or4_1 _15732_ (.A(_08542_),
    .B(_08610_),
    .C(_08564_),
    .D(_08917_),
    .X(_08918_));
 sg13g2_inv_1 _15733_ (.Y(_08919_),
    .A(_08587_));
 sg13g2_nand4_1 _15734_ (.B(_08431_),
    .C(_08919_),
    .A(_08409_),
    .Y(_08920_),
    .D(_08501_));
 sg13g2_nand3_1 _15735_ (.B(_08455_),
    .C(_08480_),
    .A(_08522_),
    .Y(_08921_));
 sg13g2_nor4_1 _15736_ (.A(_08379_),
    .B(_08918_),
    .C(_08920_),
    .D(_08921_),
    .Y(_08922_));
 sg13g2_inv_2 _15737_ (.Y(_08923_),
    .A(_08922_));
 sg13g2_nor2_1 _15738_ (.A(_08260_),
    .B(_08923_),
    .Y(_08924_));
 sg13g2_buf_1 _15739_ (.A(_08924_),
    .X(_08925_));
 sg13g2_buf_1 _15740_ (.A(net121),
    .X(_08926_));
 sg13g2_buf_1 _15741_ (.A(net121),
    .X(_08927_));
 sg13g2_buf_1 _15742_ (.A(_08841_),
    .X(_08928_));
 sg13g2_buf_1 _15743_ (.A(_08824_),
    .X(_08929_));
 sg13g2_nor3_1 _15744_ (.A(net233),
    .B(_08879_),
    .C(_08908_),
    .Y(_08930_));
 sg13g2_nand3_1 _15745_ (.B(net254),
    .C(_08930_),
    .A(_08927_),
    .Y(_08931_));
 sg13g2_o21ai_1 _15746_ (.B1(_08931_),
    .Y(_00018_),
    .A1(_08915_),
    .A2(net105));
 sg13g2_buf_2 _15747_ (.A(\cpu.dec.r_op[3] ),
    .X(_08932_));
 sg13g2_buf_1 _15748_ (.A(_08932_),
    .X(_08933_));
 sg13g2_inv_1 _15749_ (.Y(_08934_),
    .A(net1041));
 sg13g2_nand2_1 _15750_ (.Y(_08935_),
    .A(_08708_),
    .B(_08719_));
 sg13g2_inv_1 _15751_ (.Y(_08936_),
    .A(net305));
 sg13g2_buf_1 _15752_ (.A(_08936_),
    .X(_08937_));
 sg13g2_a21oi_1 _15753_ (.A1(net1045),
    .A2(_08748_),
    .Y(_08938_),
    .B1(_08759_));
 sg13g2_buf_1 _15754_ (.A(_08938_),
    .X(_08939_));
 sg13g2_nor2_1 _15755_ (.A(net232),
    .B(net253),
    .Y(_08940_));
 sg13g2_buf_1 _15756_ (.A(_08940_),
    .X(_08941_));
 sg13g2_nand2_1 _15757_ (.Y(_08942_),
    .A(_08935_),
    .B(net185));
 sg13g2_buf_1 _15758_ (.A(_08942_),
    .X(_08943_));
 sg13g2_a21oi_1 _15759_ (.A1(_08766_),
    .A2(_08774_),
    .Y(_08944_),
    .B1(_08781_));
 sg13g2_buf_1 _15760_ (.A(_08944_),
    .X(_08945_));
 sg13g2_nand2_1 _15761_ (.Y(_08946_),
    .A(_08945_),
    .B(_08802_));
 sg13g2_buf_2 _15762_ (.A(_08946_),
    .X(_08947_));
 sg13g2_nor2_1 _15763_ (.A(net120),
    .B(_08947_),
    .Y(_08948_));
 sg13g2_inv_2 _15764_ (.Y(_08949_),
    .A(_08901_));
 sg13g2_nand2b_1 _15765_ (.Y(_08950_),
    .B(_08949_),
    .A_N(_08879_));
 sg13g2_nand2_1 _15766_ (.Y(_08951_),
    .A(net233),
    .B(net254));
 sg13g2_nor2_1 _15767_ (.A(_08950_),
    .B(_08951_),
    .Y(_08952_));
 sg13g2_nand3_1 _15768_ (.B(_08948_),
    .C(_08952_),
    .A(_08927_),
    .Y(_08953_));
 sg13g2_o21ai_1 _15769_ (.B1(_08953_),
    .Y(_00014_),
    .A1(_08934_),
    .A2(net105));
 sg13g2_nand2_1 _15770_ (.Y(_08954_),
    .A(net210),
    .B(_08913_));
 sg13g2_nor2_1 _15771_ (.A(net233),
    .B(_08950_),
    .Y(_08955_));
 sg13g2_nand2_1 _15772_ (.Y(_08956_),
    .A(net254),
    .B(_08955_));
 sg13g2_a21oi_1 _15773_ (.A1(_08954_),
    .A2(_08956_),
    .Y(_08957_),
    .B1(_08807_));
 sg13g2_buf_1 _15774_ (.A(\cpu.dec.r_op[2] ),
    .X(_08958_));
 sg13g2_buf_1 _15775_ (.A(net1113),
    .X(_08959_));
 sg13g2_buf_1 _15776_ (.A(net187),
    .X(_08960_));
 sg13g2_mux2_1 _15777_ (.A0(_08957_),
    .A1(net1040),
    .S(net149),
    .X(_00013_));
 sg13g2_nor2b_1 _15778_ (.A(r_reset),
    .B_N(net1),
    .Y(_08961_));
 sg13g2_buf_1 _15779_ (.A(_08961_),
    .X(_08962_));
 sg13g2_buf_1 _15780_ (.A(net1039),
    .X(_08963_));
 sg13g2_buf_1 _15781_ (.A(net901),
    .X(_08964_));
 sg13g2_buf_1 _15782_ (.A(net783),
    .X(_08965_));
 sg13g2_buf_2 _15783_ (.A(\cpu.ex.r_ie ),
    .X(_08966_));
 sg13g2_inv_1 _15784_ (.Y(_08967_),
    .A(_08966_));
 sg13g2_buf_1 _15785_ (.A(\cpu.intr.r_clock ),
    .X(_08968_));
 sg13g2_buf_1 _15786_ (.A(\cpu.intr.r_timer ),
    .X(_08969_));
 sg13g2_buf_1 _15787_ (.A(\cpu.intr.r_enable[2] ),
    .X(_08970_));
 sg13g2_a22oi_1 _15788_ (.Y(_08971_),
    .B1(_08969_),
    .B2(_08970_),
    .A2(\cpu.intr.r_enable[1] ),
    .A1(_08968_));
 sg13g2_buf_1 _15789_ (.A(\cpu.uart.r_x_int ),
    .X(_08972_));
 sg13g2_buf_2 _15790_ (.A(\cpu.uart.r_r_int ),
    .X(_08973_));
 sg13g2_o21ai_1 _15791_ (.B1(\cpu.intr.r_enable[0] ),
    .Y(_08974_),
    .A1(_08972_),
    .A2(_08973_));
 sg13g2_buf_1 _15792_ (.A(\cpu.intr.r_swi ),
    .X(_08975_));
 sg13g2_buf_2 _15793_ (.A(\cpu.intr.spi_intr ),
    .X(_08976_));
 sg13g2_a22oi_1 _15794_ (.Y(_08977_),
    .B1(_08976_),
    .B2(\cpu.intr.r_enable[5] ),
    .A2(_08975_),
    .A1(\cpu.intr.r_enable[3] ));
 sg13g2_nand3_1 _15795_ (.B(_08974_),
    .C(_08977_),
    .A(_08971_),
    .Y(_08978_));
 sg13g2_buf_2 _15796_ (.A(_08978_),
    .X(_08979_));
 sg13g2_buf_1 _15797_ (.A(ui_in[3]),
    .X(_08980_));
 sg13g2_nand2_1 _15798_ (.Y(_08981_),
    .A(\cpu.gpio.r_enable_in[3] ),
    .B(_08980_));
 sg13g2_buf_2 _15799_ (.A(uio_in[4]),
    .X(_08982_));
 sg13g2_nand2_1 _15800_ (.Y(_08983_),
    .A(\cpu.gpio.r_enable_io[4] ),
    .B(_08982_));
 sg13g2_buf_1 _15801_ (.A(\cpu.gpio.r_enable_io[5] ),
    .X(_08984_));
 sg13g2_buf_1 _15802_ (.A(uio_in[5]),
    .X(_08985_));
 sg13g2_nand2_1 _15803_ (.Y(_08986_),
    .A(_08984_),
    .B(_08985_));
 sg13g2_buf_2 _15804_ (.A(ui_in[7]),
    .X(_08987_));
 sg13g2_nand2_1 _15805_ (.Y(_08988_),
    .A(\cpu.gpio.r_enable_in[7] ),
    .B(_08987_));
 sg13g2_and4_1 _15806_ (.A(_08981_),
    .B(_08983_),
    .C(_08986_),
    .D(_08988_),
    .X(_08989_));
 sg13g2_buf_1 _15807_ (.A(\cpu.gpio.r_enable_in[0] ),
    .X(_08990_));
 sg13g2_buf_2 _15808_ (.A(ui_in[0]),
    .X(_08991_));
 sg13g2_buf_2 _15809_ (.A(\cpu.gpio.r_enable_io[7] ),
    .X(_08992_));
 sg13g2_buf_1 _15810_ (.A(uio_in[7]),
    .X(_08993_));
 sg13g2_a22oi_1 _15811_ (.Y(_08994_),
    .B1(_08992_),
    .B2(_08993_),
    .A2(_08991_),
    .A1(_08990_));
 sg13g2_buf_1 _15812_ (.A(\cpu.gpio.r_enable_in[4] ),
    .X(_08995_));
 sg13g2_buf_8 _15813_ (.A(ui_in[4]),
    .X(_08996_));
 sg13g2_buf_2 _15814_ (.A(\cpu.gpio.r_enable_in[6] ),
    .X(_08997_));
 sg13g2_buf_2 _15815_ (.A(ui_in[6]),
    .X(_08998_));
 sg13g2_a22oi_1 _15816_ (.Y(_08999_),
    .B1(_08997_),
    .B2(_08998_),
    .A2(_08996_),
    .A1(_08995_));
 sg13g2_buf_8 _15817_ (.A(ui_in[2]),
    .X(_09000_));
 sg13g2_buf_1 _15818_ (.A(\cpu.gpio.r_enable_in[5] ),
    .X(_09001_));
 sg13g2_buf_2 _15819_ (.A(ui_in[5]),
    .X(_09002_));
 sg13g2_a22oi_1 _15820_ (.Y(_09003_),
    .B1(_09001_),
    .B2(_09002_),
    .A2(_09000_),
    .A1(\cpu.gpio.r_enable_in[2] ));
 sg13g2_buf_8 _15821_ (.A(ui_in[1]),
    .X(_09004_));
 sg13g2_buf_2 _15822_ (.A(uio_in[6]),
    .X(_09005_));
 sg13g2_a22oi_1 _15823_ (.Y(_09006_),
    .B1(\cpu.gpio.r_enable_io[6] ),
    .B2(_09005_),
    .A2(_09004_),
    .A1(\cpu.gpio.r_enable_in[1] ));
 sg13g2_and4_1 _15824_ (.A(_08994_),
    .B(_08999_),
    .C(_09003_),
    .D(_09006_),
    .X(_09007_));
 sg13g2_buf_2 _15825_ (.A(\cpu.intr.r_enable[4] ),
    .X(_09008_));
 sg13g2_inv_1 _15826_ (.Y(_09009_),
    .A(_09008_));
 sg13g2_a21oi_2 _15827_ (.B1(_09009_),
    .Y(_09010_),
    .A2(_09007_),
    .A1(_08989_));
 sg13g2_nor2_1 _15828_ (.A(_08979_),
    .B(_09010_),
    .Y(_09011_));
 sg13g2_nor2_1 _15829_ (.A(_08967_),
    .B(_09011_),
    .Y(_09012_));
 sg13g2_buf_1 _15830_ (.A(\cpu.dec.r_trap ),
    .X(_09013_));
 sg13g2_a21oi_1 _15831_ (.A1(_08222_),
    .A2(_09012_),
    .Y(_09014_),
    .B1(_09013_));
 sg13g2_and2_1 _15832_ (.A(_08258_),
    .B(_09014_),
    .X(_09015_));
 sg13g2_buf_1 _15833_ (.A(_09015_),
    .X(_09016_));
 sg13g2_nor2b_1 _15834_ (.A(_00181_),
    .B_N(_09016_),
    .Y(_09017_));
 sg13g2_inv_1 _15835_ (.Y(_09018_),
    .A(net1122));
 sg13g2_nor2_1 _15836_ (.A(net1118),
    .B(net1119),
    .Y(_09019_));
 sg13g2_a21oi_1 _15837_ (.A1(net1118),
    .A2(_08124_),
    .Y(_09020_),
    .B1(_09019_));
 sg13g2_buf_1 _15838_ (.A(_08185_),
    .X(_09021_));
 sg13g2_a22oi_1 _15839_ (.Y(_09022_),
    .B1(_09020_),
    .B2(_09021_),
    .A2(_09018_),
    .A1(_08186_));
 sg13g2_buf_2 _15840_ (.A(\cpu.addr[6] ),
    .X(_09023_));
 sg13g2_buf_1 _15841_ (.A(\cpu.addr[8] ),
    .X(_09024_));
 sg13g2_buf_2 _15842_ (.A(_09024_),
    .X(_09025_));
 sg13g2_buf_2 _15843_ (.A(\cpu.addr[7] ),
    .X(_09026_));
 sg13g2_nor2b_1 _15844_ (.A(net1037),
    .B_N(_09026_),
    .Y(_09027_));
 sg13g2_buf_1 _15845_ (.A(_09027_),
    .X(_09028_));
 sg13g2_nand2_1 _15846_ (.Y(_09029_),
    .A(_09023_),
    .B(_09028_));
 sg13g2_buf_1 _15847_ (.A(_09029_),
    .X(_09030_));
 sg13g2_buf_1 _15848_ (.A(_00201_),
    .X(_09031_));
 sg13g2_buf_1 _15849_ (.A(\cpu.addr[2] ),
    .X(_09032_));
 sg13g2_buf_1 _15850_ (.A(_09032_),
    .X(_09033_));
 sg13g2_buf_8 _15851_ (.A(net1036),
    .X(_09034_));
 sg13g2_buf_1 _15852_ (.A(_09034_),
    .X(_09035_));
 sg13g2_buf_1 _15853_ (.A(net782),
    .X(_09036_));
 sg13g2_buf_1 _15854_ (.A(net686),
    .X(_09037_));
 sg13g2_buf_1 _15855_ (.A(\cpu.addr[1] ),
    .X(_09038_));
 sg13g2_nor2_1 _15856_ (.A(net609),
    .B(net1111),
    .Y(_09039_));
 sg13g2_nand2_2 _15857_ (.Y(_09040_),
    .A(_09031_),
    .B(_09039_));
 sg13g2_nor2_1 _15858_ (.A(_09030_),
    .B(_09040_),
    .Y(_09041_));
 sg13g2_and3_1 _15859_ (.X(_09042_),
    .A(_09017_),
    .B(_09022_),
    .C(_09041_));
 sg13g2_buf_1 _15860_ (.A(_09042_),
    .X(_09043_));
 sg13g2_buf_2 _15861_ (.A(\cpu.spi.r_state[1] ),
    .X(_09044_));
 sg13g2_nand3_1 _15862_ (.B(_08129_),
    .C(_09016_),
    .A(_08181_),
    .Y(_09045_));
 sg13g2_buf_1 _15863_ (.A(_09045_),
    .X(_09046_));
 sg13g2_or2_1 _15864_ (.X(_09047_),
    .B(_09046_),
    .A(_09030_));
 sg13g2_buf_2 _15865_ (.A(_09047_),
    .X(_09048_));
 sg13g2_buf_2 _15866_ (.A(\cpu.addr[3] ),
    .X(_09049_));
 sg13g2_buf_8 _15867_ (.A(_09049_),
    .X(_09050_));
 sg13g2_inv_2 _15868_ (.Y(_09051_),
    .A(net1035));
 sg13g2_buf_1 _15869_ (.A(_09051_),
    .X(_09052_));
 sg13g2_nand2b_1 _15870_ (.Y(_09053_),
    .B(net781),
    .A_N(_09048_));
 sg13g2_buf_2 _15871_ (.A(_09053_),
    .X(_09054_));
 sg13g2_nand2_1 _15872_ (.Y(_09055_),
    .A(_09044_),
    .B(_09054_));
 sg13g2_buf_2 _15873_ (.A(_09055_),
    .X(_09056_));
 sg13g2_buf_1 _15874_ (.A(\cpu.spi.r_state[6] ),
    .X(_09057_));
 sg13g2_buf_1 _15875_ (.A(_09057_),
    .X(_09058_));
 sg13g2_buf_1 _15876_ (.A(\cpu.spi.r_bits[0] ),
    .X(_09059_));
 sg13g2_buf_1 _15877_ (.A(\cpu.spi.r_bits[1] ),
    .X(_09060_));
 sg13g2_nor3_1 _15878_ (.A(_09059_),
    .B(_09060_),
    .C(\cpu.spi.r_bits[2] ),
    .Y(_09061_));
 sg13g2_nor3_2 _15879_ (.A(\cpu.spi.r_timeout_count[0] ),
    .B(\cpu.spi.r_timeout_count[1] ),
    .C(\cpu.spi.r_timeout_count[2] ),
    .Y(_09062_));
 sg13g2_nor2b_1 _15880_ (.A(\cpu.spi.r_timeout_count[3] ),
    .B_N(_09062_),
    .Y(_09063_));
 sg13g2_nand2b_1 _15881_ (.Y(_09064_),
    .B(_09063_),
    .A_N(\cpu.spi.r_timeout_count[4] ));
 sg13g2_nor2_1 _15882_ (.A(\cpu.spi.r_timeout_count[5] ),
    .B(_09064_),
    .Y(_09065_));
 sg13g2_nand2b_1 _15883_ (.Y(_09066_),
    .B(_09065_),
    .A_N(\cpu.spi.r_timeout_count[6] ));
 sg13g2_buf_1 _15884_ (.A(_09066_),
    .X(_09067_));
 sg13g2_o21ai_1 _15885_ (.B1(\cpu.spi.r_searching ),
    .Y(_09068_),
    .A1(\cpu.spi.r_timeout_count[7] ),
    .A2(_09067_));
 sg13g2_nand2_1 _15886_ (.Y(_09069_),
    .A(_09061_),
    .B(_09068_));
 sg13g2_buf_1 _15887_ (.A(\cpu.spi.r_in[3] ),
    .X(_09070_));
 sg13g2_buf_1 _15888_ (.A(\cpu.spi.r_in[6] ),
    .X(_09071_));
 sg13g2_buf_1 _15889_ (.A(\cpu.spi.r_in[1] ),
    .X(_09072_));
 sg13g2_buf_1 _15890_ (.A(\cpu.spi.r_in[0] ),
    .X(_09073_));
 sg13g2_nand2_1 _15891_ (.Y(_09074_),
    .A(_09072_),
    .B(_09073_));
 sg13g2_nand3_1 _15892_ (.B(_09071_),
    .C(_09074_),
    .A(_09070_),
    .Y(_09075_));
 sg13g2_buf_1 _15893_ (.A(\cpu.spi.r_in[2] ),
    .X(_09076_));
 sg13g2_buf_1 _15894_ (.A(\cpu.spi.r_in[5] ),
    .X(_09077_));
 sg13g2_buf_1 _15895_ (.A(\cpu.spi.r_in[4] ),
    .X(_09078_));
 sg13g2_nand4_1 _15896_ (.B(_09077_),
    .C(_09078_),
    .A(_09076_),
    .Y(_09079_),
    .D(\cpu.spi.r_in[7] ));
 sg13g2_nor2_1 _15897_ (.A(_09075_),
    .B(_09079_),
    .Y(_09080_));
 sg13g2_o21ai_1 _15898_ (.B1(\cpu.spi.r_searching ),
    .Y(_09081_),
    .A1(_00200_),
    .A2(_09080_));
 sg13g2_nand2_2 _15899_ (.Y(_09082_),
    .A(_09069_),
    .B(_09081_));
 sg13g2_buf_1 _15900_ (.A(\cpu.spi.r_count[7] ),
    .X(_09083_));
 sg13g2_buf_1 _15901_ (.A(\cpu.spi.r_count[2] ),
    .X(_09084_));
 sg13g2_buf_1 _15902_ (.A(\cpu.spi.r_count[0] ),
    .X(_09085_));
 sg13g2_or2_1 _15903_ (.X(_09086_),
    .B(\cpu.spi.r_count[1] ),
    .A(_09085_));
 sg13g2_buf_1 _15904_ (.A(_09086_),
    .X(_09087_));
 sg13g2_nor3_1 _15905_ (.A(_09084_),
    .B(\cpu.spi.r_count[3] ),
    .C(_09087_),
    .Y(_09088_));
 sg13g2_nor2b_1 _15906_ (.A(\cpu.spi.r_count[4] ),
    .B_N(_09088_),
    .Y(_09089_));
 sg13g2_nor2b_1 _15907_ (.A(\cpu.spi.r_count[5] ),
    .B_N(_09089_),
    .Y(_09090_));
 sg13g2_nor2b_1 _15908_ (.A(\cpu.spi.r_count[6] ),
    .B_N(_09090_),
    .Y(_09091_));
 sg13g2_buf_1 _15909_ (.A(_09091_),
    .X(_09092_));
 sg13g2_nor2b_1 _15910_ (.A(_09083_),
    .B_N(_09092_),
    .Y(_09093_));
 sg13g2_buf_1 _15911_ (.A(_09093_),
    .X(_09094_));
 sg13g2_buf_1 _15912_ (.A(net379),
    .X(_09095_));
 sg13g2_nand3_1 _15913_ (.B(_09082_),
    .C(net304),
    .A(net1034),
    .Y(_09096_));
 sg13g2_o21ai_1 _15914_ (.B1(_09096_),
    .Y(_09097_),
    .A1(_09043_),
    .A2(_09056_));
 sg13g2_and2_1 _15915_ (.A(net687),
    .B(_09097_),
    .X(_00030_));
 sg13g2_buf_1 _15916_ (.A(_09044_),
    .X(_09098_));
 sg13g2_buf_1 _15917_ (.A(net1033),
    .X(_09099_));
 sg13g2_buf_2 _15918_ (.A(_09049_),
    .X(_09100_));
 sg13g2_buf_1 _15919_ (.A(net1032),
    .X(_09101_));
 sg13g2_buf_8 _15920_ (.A(net898),
    .X(_09102_));
 sg13g2_buf_1 _15921_ (.A(net780),
    .X(_09103_));
 sg13g2_buf_1 _15922_ (.A(net685),
    .X(_09104_));
 sg13g2_buf_1 _15923_ (.A(net608),
    .X(_09105_));
 sg13g2_buf_1 _15924_ (.A(net532),
    .X(_09106_));
 sg13g2_nor2_1 _15925_ (.A(net464),
    .B(_09048_),
    .Y(_09107_));
 sg13g2_buf_2 _15926_ (.A(_09107_),
    .X(_09108_));
 sg13g2_buf_1 _15927_ (.A(_09108_),
    .X(_09109_));
 sg13g2_a21oi_1 _15928_ (.A1(_09099_),
    .A2(_09109_),
    .Y(_09110_),
    .B1(\cpu.spi.r_state[5] ));
 sg13g2_buf_1 _15929_ (.A(\cpu.spi.r_state[4] ),
    .X(_09111_));
 sg13g2_nand2b_1 _15930_ (.Y(_09112_),
    .B(_09092_),
    .A_N(_09083_));
 sg13g2_buf_1 _15931_ (.A(_09112_),
    .X(_09113_));
 sg13g2_inv_2 _15932_ (.Y(_09114_),
    .A(_09057_));
 sg13g2_nor2_1 _15933_ (.A(_09114_),
    .B(_09082_),
    .Y(_09115_));
 sg13g2_nor3_1 _15934_ (.A(net1110),
    .B(net378),
    .C(_09115_),
    .Y(_09116_));
 sg13g2_buf_2 _15935_ (.A(\cpu.spi.r_state[2] ),
    .X(_09117_));
 sg13g2_buf_1 _15936_ (.A(net901),
    .X(_09118_));
 sg13g2_o21ai_1 _15937_ (.B1(net779),
    .Y(_09119_),
    .A1(_09117_),
    .A2(net304));
 sg13g2_a21oi_1 _15938_ (.A1(_09110_),
    .A2(_09116_),
    .Y(_00031_),
    .B1(_09119_));
 sg13g2_nand2b_1 _15939_ (.Y(_09120_),
    .B(net1),
    .A_N(r_reset));
 sg13g2_buf_2 _15940_ (.A(_09120_),
    .X(_09121_));
 sg13g2_buf_1 _15941_ (.A(_09121_),
    .X(_09122_));
 sg13g2_buf_2 _15942_ (.A(net897),
    .X(_09123_));
 sg13g2_buf_2 _15943_ (.A(net778),
    .X(_09124_));
 sg13g2_inv_1 _15944_ (.Y(_09125_),
    .A(_09044_));
 sg13g2_nor2_1 _15945_ (.A(_09125_),
    .B(_09109_),
    .Y(_09126_));
 sg13g2_buf_1 _15946_ (.A(\cpu.spi.r_state[3] ),
    .X(_09127_));
 sg13g2_a21oi_1 _15947_ (.A1(_09043_),
    .A2(_09126_),
    .Y(_09128_),
    .B1(_09127_));
 sg13g2_nor3_1 _15948_ (.A(net684),
    .B(_09095_),
    .C(_09128_),
    .Y(_00032_));
 sg13g2_buf_1 _15949_ (.A(net778),
    .X(_09129_));
 sg13g2_buf_1 _15950_ (.A(_09129_),
    .X(_09130_));
 sg13g2_nor2_1 _15951_ (.A(_09040_),
    .B(_09048_),
    .Y(_09131_));
 sg13g2_buf_1 _15952_ (.A(\cpu.spi.r_state[0] ),
    .X(_09132_));
 sg13g2_a22oi_1 _15953_ (.Y(_09133_),
    .B1(_09131_),
    .B2(_09132_),
    .A2(net378),
    .A1(net1110));
 sg13g2_nor2_1 _15954_ (.A(net607),
    .B(_09133_),
    .Y(_00033_));
 sg13g2_nor3_1 _15955_ (.A(net684),
    .B(net304),
    .C(_09110_),
    .Y(_00034_));
 sg13g2_nand2_1 _15956_ (.Y(_09134_),
    .A(net1034),
    .B(net378));
 sg13g2_nand2_1 _15957_ (.Y(_09135_),
    .A(_09117_),
    .B(net304));
 sg13g2_buf_2 _15958_ (.A(net778),
    .X(_09136_));
 sg13g2_buf_1 _15959_ (.A(_09136_),
    .X(_09137_));
 sg13g2_a21oi_1 _15960_ (.A1(_09134_),
    .A2(_09135_),
    .Y(_00035_),
    .B1(net606));
 sg13g2_buf_1 _15961_ (.A(\cpu.ex.r_div_running ),
    .X(_09138_));
 sg13g2_buf_1 _15962_ (.A(\cpu.ex.r_mult_off[1] ),
    .X(_09139_));
 sg13g2_buf_1 _15963_ (.A(\cpu.ex.r_mult_off[2] ),
    .X(_09140_));
 sg13g2_buf_2 _15964_ (.A(\cpu.ex.r_mult_off[0] ),
    .X(_09141_));
 sg13g2_inv_1 _15965_ (.Y(_09142_),
    .A(\cpu.dec.div ));
 sg13g2_nand3b_1 _15966_ (.B(\cpu.dec.iready ),
    .C(_00183_),
    .Y(_09143_),
    .A_N(\cpu.ex.r_branch_stall ));
 sg13g2_buf_1 _15967_ (.A(_09143_),
    .X(_09144_));
 sg13g2_or3_1 _15968_ (.A(_09142_),
    .B(_09121_),
    .C(net1031),
    .X(_09145_));
 sg13g2_buf_1 _15969_ (.A(_09145_),
    .X(_09146_));
 sg13g2_inv_1 _15970_ (.Y(_09147_),
    .A(\cpu.dec.mult ));
 sg13g2_or3_1 _15971_ (.A(_09147_),
    .B(_09121_),
    .C(net1031),
    .X(_09148_));
 sg13g2_buf_2 _15972_ (.A(_09148_),
    .X(_09149_));
 sg13g2_nand3_1 _15973_ (.B(_09146_),
    .C(_09149_),
    .A(_09141_),
    .Y(_09150_));
 sg13g2_buf_2 _15974_ (.A(_09150_),
    .X(\cpu.ex.c_mult_off[0] ));
 sg13g2_nor4_2 _15975_ (.A(net1109),
    .B(_09140_),
    .C(\cpu.ex.r_mult_off[3] ),
    .Y(_09151_),
    .D(\cpu.ex.c_mult_off[0] ));
 sg13g2_nor3_1 _15976_ (.A(_09142_),
    .B(_09121_),
    .C(net1031),
    .Y(_09152_));
 sg13g2_buf_2 _15977_ (.A(_09152_),
    .X(_09153_));
 sg13g2_o21ai_1 _15978_ (.B1(net1039),
    .Y(_09154_),
    .A1(_09138_),
    .A2(_09153_));
 sg13g2_a21oi_1 _15979_ (.A1(_09138_),
    .A2(_09151_),
    .Y(\cpu.ex.c_div_running ),
    .B1(_09154_));
 sg13g2_buf_1 _15980_ (.A(\cpu.ex.r_mult_running ),
    .X(_09155_));
 sg13g2_inv_1 _15981_ (.Y(_09156_),
    .A(_09155_));
 sg13g2_buf_1 _15982_ (.A(_09149_),
    .X(_09157_));
 sg13g2_nand2_2 _15983_ (.Y(_09158_),
    .A(_09156_),
    .B(net683));
 sg13g2_nand2_1 _15984_ (.Y(_09159_),
    .A(net1039),
    .B(_09158_));
 sg13g2_a21oi_1 _15985_ (.A1(_09155_),
    .A2(_09151_),
    .Y(\cpu.ex.c_mult_running ),
    .B1(_09159_));
 sg13g2_o21ai_1 _15986_ (.B1(_09132_),
    .Y(_09160_),
    .A1(_09040_),
    .A2(_09048_));
 sg13g2_and2_1 _15987_ (.A(net1039),
    .B(_09160_),
    .X(_09161_));
 sg13g2_buf_1 _15988_ (.A(_09161_),
    .X(_09162_));
 sg13g2_o21ai_1 _15989_ (.B1(_09162_),
    .Y(_00029_),
    .A1(net378),
    .A2(_09128_));
 sg13g2_buf_1 _15990_ (.A(\cpu.qspi.r_state[17] ),
    .X(_09163_));
 sg13g2_buf_1 _15991_ (.A(_08133_),
    .X(_09164_));
 sg13g2_inv_1 _15992_ (.Y(_09165_),
    .A(_08181_));
 sg13g2_buf_1 _15993_ (.A(_09165_),
    .X(_09166_));
 sg13g2_and2_1 _15994_ (.A(_09166_),
    .B(_09016_),
    .X(_09167_));
 sg13g2_buf_1 _15995_ (.A(_09167_),
    .X(_09168_));
 sg13g2_mux4_1 _15996_ (.S0(net686),
    .A0(\cpu.dcache.r_valid[4] ),
    .A1(\cpu.dcache.r_valid[5] ),
    .A2(\cpu.dcache.r_valid[6] ),
    .A3(\cpu.dcache.r_valid[7] ),
    .S1(net685),
    .X(_09169_));
 sg13g2_mux4_1 _15997_ (.S0(net686),
    .A0(\cpu.dcache.r_valid[0] ),
    .A1(\cpu.dcache.r_valid[1] ),
    .A2(\cpu.dcache.r_valid[2] ),
    .A3(\cpu.dcache.r_valid[3] ),
    .S1(_09103_),
    .X(_09170_));
 sg13g2_buf_2 _15998_ (.A(\cpu.addr[4] ),
    .X(_09171_));
 sg13g2_inv_1 _15999_ (.Y(_09172_),
    .A(_09171_));
 sg13g2_buf_1 _16000_ (.A(_09172_),
    .X(_09173_));
 sg13g2_buf_1 _16001_ (.A(net895),
    .X(_09174_));
 sg13g2_mux2_1 _16002_ (.A0(_09169_),
    .A1(_09170_),
    .S(net777),
    .X(_09175_));
 sg13g2_mux4_1 _16003_ (.S0(net686),
    .A0(\cpu.dcache.r_dirty[4] ),
    .A1(\cpu.dcache.r_dirty[5] ),
    .A2(\cpu.dcache.r_dirty[6] ),
    .A3(\cpu.dcache.r_dirty[7] ),
    .S1(net685),
    .X(_09176_));
 sg13g2_mux4_1 _16004_ (.S0(net686),
    .A0(\cpu.dcache.r_dirty[0] ),
    .A1(\cpu.dcache.r_dirty[1] ),
    .A2(\cpu.dcache.r_dirty[2] ),
    .A3(\cpu.dcache.r_dirty[3] ),
    .S1(net685),
    .X(_09177_));
 sg13g2_mux2_1 _16005_ (.A0(_09176_),
    .A1(_09177_),
    .S(net777),
    .X(_09178_));
 sg13g2_and4_1 _16006_ (.A(_08258_),
    .B(_09014_),
    .C(_09175_),
    .D(_09178_),
    .X(_09179_));
 sg13g2_buf_1 _16007_ (.A(_09179_),
    .X(_09180_));
 sg13g2_inv_1 _16008_ (.Y(_09181_),
    .A(_09180_));
 sg13g2_buf_1 _16009_ (.A(\cpu.dcache.flush_write ),
    .X(_09182_));
 sg13g2_buf_1 _16010_ (.A(_08136_),
    .X(_09183_));
 sg13g2_buf_8 _16011_ (.A(net1062),
    .X(_09184_));
 sg13g2_buf_8 _16012_ (.A(_09184_),
    .X(_09185_));
 sg13g2_buf_2 _16013_ (.A(_08154_),
    .X(_09186_));
 sg13g2_buf_1 _16014_ (.A(_09186_),
    .X(_09187_));
 sg13g2_mux4_1 _16015_ (.S0(net775),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][4] ),
    .S1(net774),
    .X(_09188_));
 sg13g2_mux4_1 _16016_ (.S0(net775),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][4] ),
    .S1(net774),
    .X(_09189_));
 sg13g2_buf_2 _16017_ (.A(_08138_),
    .X(_09190_));
 sg13g2_buf_1 _16018_ (.A(_09186_),
    .X(_09191_));
 sg13g2_mux4_1 _16019_ (.S0(net894),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][4] ),
    .S1(net773),
    .X(_09192_));
 sg13g2_mux4_1 _16020_ (.S0(net894),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][4] ),
    .S1(net773),
    .X(_09193_));
 sg13g2_mux4_1 _16021_ (.S0(net1058),
    .A0(_09188_),
    .A1(_09189_),
    .A2(_09192_),
    .A3(_09193_),
    .S1(net1057),
    .X(_09194_));
 sg13g2_nand2_1 _16022_ (.Y(_09195_),
    .A(net776),
    .B(_09194_));
 sg13g2_nand2_1 _16023_ (.Y(_09196_),
    .A(_08164_),
    .B(_08165_));
 sg13g2_buf_4 _16024_ (.X(_09197_),
    .A(_09196_));
 sg13g2_buf_1 _16025_ (.A(_09197_),
    .X(_09198_));
 sg13g2_mux4_1 _16026_ (.S0(_09185_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][4] ),
    .S1(_09187_),
    .X(_09199_));
 sg13g2_mux4_1 _16027_ (.S0(net775),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][4] ),
    .S1(net774),
    .X(_09200_));
 sg13g2_buf_2 _16028_ (.A(_08138_),
    .X(_09201_));
 sg13g2_buf_1 _16029_ (.A(_08154_),
    .X(_09202_));
 sg13g2_mux4_1 _16030_ (.S0(net893),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][4] ),
    .S1(net892),
    .X(_09203_));
 sg13g2_mux4_1 _16031_ (.S0(net894),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][4] ),
    .S1(net773),
    .X(_09204_));
 sg13g2_mux4_1 _16032_ (.S0(net1058),
    .A0(_09199_),
    .A1(_09200_),
    .A2(_09203_),
    .A3(_09204_),
    .S1(net1057),
    .X(_09205_));
 sg13g2_nand2_1 _16033_ (.Y(_09206_),
    .A(net682),
    .B(_09205_));
 sg13g2_a21oi_2 _16034_ (.B1(_08380_),
    .Y(_09207_),
    .A2(_09206_),
    .A1(_09195_));
 sg13g2_buf_1 _16035_ (.A(_09207_),
    .X(_09208_));
 sg13g2_buf_1 _16036_ (.A(_00206_),
    .X(_09209_));
 sg13g2_nor2b_1 _16037_ (.A(_09100_),
    .B_N(net1108),
    .Y(_09210_));
 sg13g2_nand2_1 _16038_ (.Y(_09211_),
    .A(_09035_),
    .B(_09210_));
 sg13g2_buf_2 _16039_ (.A(_09211_),
    .X(_09212_));
 sg13g2_nand3b_1 _16040_ (.B(net1035),
    .C(\cpu.dcache.r_tag[6][16] ),
    .Y(_09213_),
    .A_N(net1036));
 sg13g2_nand3b_1 _16041_ (.B(\cpu.dcache.r_tag[5][16] ),
    .C(net1036),
    .Y(_09214_),
    .A_N(_09050_));
 sg13g2_a21o_1 _16042_ (.A2(_09214_),
    .A1(_09213_),
    .B1(net895),
    .X(_09215_));
 sg13g2_inv_1 _16043_ (.Y(_09216_),
    .A(net1112));
 sg13g2_buf_1 _16044_ (.A(_09216_),
    .X(_09217_));
 sg13g2_buf_1 _16045_ (.A(_09171_),
    .X(_09218_));
 sg13g2_nor2b_2 _16046_ (.A(net1035),
    .B_N(net1029),
    .Y(_09219_));
 sg13g2_nand3_1 _16047_ (.B(\cpu.dcache.r_tag[4][16] ),
    .C(_09219_),
    .A(net891),
    .Y(_09220_));
 sg13g2_and3_1 _16048_ (.X(_09221_),
    .A(net1112),
    .B(_09171_),
    .C(_09049_));
 sg13g2_buf_1 _16049_ (.A(_09221_),
    .X(_09222_));
 sg13g2_and2_1 _16050_ (.A(_09049_),
    .B(_00206_),
    .X(_09223_));
 sg13g2_buf_1 _16051_ (.A(_09223_),
    .X(_09224_));
 sg13g2_mux2_1 _16052_ (.A0(\cpu.dcache.r_tag[2][16] ),
    .A1(\cpu.dcache.r_tag[3][16] ),
    .S(_09033_),
    .X(_09225_));
 sg13g2_a22oi_1 _16053_ (.Y(_09226_),
    .B1(net890),
    .B2(_09225_),
    .A2(_09222_),
    .A1(\cpu.dcache.r_tag[7][16] ));
 sg13g2_and3_1 _16054_ (.X(_09227_),
    .A(_09215_),
    .B(_09220_),
    .C(_09226_));
 sg13g2_or2_1 _16055_ (.X(_09228_),
    .B(_09049_),
    .A(_09171_));
 sg13g2_buf_1 _16056_ (.A(_09228_),
    .X(_09229_));
 sg13g2_buf_1 _16057_ (.A(_09229_),
    .X(_09230_));
 sg13g2_mux2_1 _16058_ (.A0(_00225_),
    .A1(_09227_),
    .S(net772),
    .X(_09231_));
 sg13g2_nor2_1 _16059_ (.A(\cpu.dcache.r_tag[1][16] ),
    .B(_09212_),
    .Y(_09232_));
 sg13g2_a22oi_1 _16060_ (.Y(_09233_),
    .B1(_09232_),
    .B2(_09227_),
    .A2(_09231_),
    .A1(_09212_));
 sg13g2_xor2_1 _16061_ (.B(_09233_),
    .A(net432),
    .X(_09234_));
 sg13g2_buf_8 _16062_ (.A(_09184_),
    .X(_09235_));
 sg13g2_buf_2 _16063_ (.A(_09186_),
    .X(_09236_));
 sg13g2_mux4_1 _16064_ (.S0(net771),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][6] ),
    .S1(net770),
    .X(_09237_));
 sg13g2_mux4_1 _16065_ (.S0(net771),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][6] ),
    .S1(net770),
    .X(_09238_));
 sg13g2_mux4_1 _16066_ (.S0(net894),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][6] ),
    .S1(net773),
    .X(_09239_));
 sg13g2_mux4_1 _16067_ (.S0(net894),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][6] ),
    .S1(net773),
    .X(_09240_));
 sg13g2_buf_2 _16068_ (.A(net1058),
    .X(_09241_));
 sg13g2_buf_1 _16069_ (.A(net1057),
    .X(_09242_));
 sg13g2_mux4_1 _16070_ (.S0(net889),
    .A0(_09237_),
    .A1(_09238_),
    .A2(_09239_),
    .A3(_09240_),
    .S1(net888),
    .X(_09243_));
 sg13g2_nand2_1 _16071_ (.Y(_09244_),
    .A(net776),
    .B(_09243_));
 sg13g2_mux4_1 _16072_ (.S0(net775),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][6] ),
    .S1(net774),
    .X(_09245_));
 sg13g2_mux4_1 _16073_ (.S0(net775),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][6] ),
    .S1(_09236_),
    .X(_09246_));
 sg13g2_mux4_1 _16074_ (.S0(net894),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][6] ),
    .S1(net773),
    .X(_09247_));
 sg13g2_mux4_1 _16075_ (.S0(_09190_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][6] ),
    .S1(_09191_),
    .X(_09248_));
 sg13g2_mux4_1 _16076_ (.S0(net1058),
    .A0(_09245_),
    .A1(_09246_),
    .A2(_09247_),
    .A3(_09248_),
    .S1(net1057),
    .X(_09249_));
 sg13g2_nand2_1 _16077_ (.Y(_09250_),
    .A(net682),
    .B(_09249_));
 sg13g2_a21oi_2 _16078_ (.B1(_08380_),
    .Y(_09251_),
    .A2(_09250_),
    .A1(_09244_));
 sg13g2_buf_1 _16079_ (.A(_09251_),
    .X(_09252_));
 sg13g2_and3_1 _16080_ (.X(_09253_),
    .A(net1112),
    .B(net1032),
    .C(net1108));
 sg13g2_buf_2 _16081_ (.A(_09253_),
    .X(_09254_));
 sg13g2_buf_1 _16082_ (.A(_09254_),
    .X(_09255_));
 sg13g2_nand2_1 _16083_ (.Y(_09256_),
    .A(\cpu.dcache.r_tag[3][18] ),
    .B(net681));
 sg13g2_and2_1 _16084_ (.A(_09033_),
    .B(_09210_),
    .X(_09257_));
 sg13g2_buf_1 _16085_ (.A(_09257_),
    .X(_09258_));
 sg13g2_buf_1 _16086_ (.A(_09258_),
    .X(_09259_));
 sg13g2_nor2b_1 _16087_ (.A(net1112),
    .B_N(_09171_),
    .Y(_09260_));
 sg13g2_buf_2 _16088_ (.A(_09260_),
    .X(_09261_));
 sg13g2_and2_1 _16089_ (.A(_09051_),
    .B(_09261_),
    .X(_09262_));
 sg13g2_buf_1 _16090_ (.A(_09262_),
    .X(_09263_));
 sg13g2_a22oi_1 _16091_ (.Y(_09264_),
    .B1(_09263_),
    .B2(\cpu.dcache.r_tag[4][18] ),
    .A2(net605),
    .A1(\cpu.dcache.r_tag[1][18] ));
 sg13g2_buf_1 _16092_ (.A(_09222_),
    .X(_09265_));
 sg13g2_and2_1 _16093_ (.A(_09216_),
    .B(net890),
    .X(_09266_));
 sg13g2_buf_2 _16094_ (.A(_09266_),
    .X(_09267_));
 sg13g2_a22oi_1 _16095_ (.Y(_09268_),
    .B1(_09267_),
    .B2(\cpu.dcache.r_tag[2][18] ),
    .A2(net769),
    .A1(\cpu.dcache.r_tag[7][18] ));
 sg13g2_buf_1 _16096_ (.A(net891),
    .X(_09269_));
 sg13g2_nand3_1 _16097_ (.B(net780),
    .C(\cpu.dcache.r_tag[6][18] ),
    .A(_09218_),
    .Y(_09270_));
 sg13g2_o21ai_1 _16098_ (.B1(_09270_),
    .Y(_09271_),
    .A1(_00227_),
    .A2(net772));
 sg13g2_nor3_1 _16099_ (.A(_09216_),
    .B(net895),
    .C(net1035),
    .Y(_09272_));
 sg13g2_buf_2 _16100_ (.A(_09272_),
    .X(_09273_));
 sg13g2_buf_1 _16101_ (.A(net1108),
    .X(_09274_));
 sg13g2_nor3_1 _16102_ (.A(net1028),
    .B(_00227_),
    .C(net772),
    .Y(_09275_));
 sg13g2_a221oi_1 _16103_ (.B2(\cpu.dcache.r_tag[5][18] ),
    .C1(_09275_),
    .B1(_09273_),
    .A1(net768),
    .Y(_09276_),
    .A2(_09271_));
 sg13g2_nand4_1 _16104_ (.B(_09264_),
    .C(_09268_),
    .A(_09256_),
    .Y(_09277_),
    .D(_09276_));
 sg13g2_xor2_1 _16105_ (.B(_09277_),
    .A(net431),
    .X(_09278_));
 sg13g2_buf_2 _16106_ (.A(_09184_),
    .X(_09279_));
 sg13g2_buf_1 _16107_ (.A(_09186_),
    .X(_09280_));
 sg13g2_mux4_1 _16108_ (.S0(net767),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][10] ),
    .S1(net766),
    .X(_09281_));
 sg13g2_mux4_1 _16109_ (.S0(net767),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][10] ),
    .S1(net766),
    .X(_09282_));
 sg13g2_mux4_1 _16110_ (.S0(net771),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][10] ),
    .S1(net770),
    .X(_09283_));
 sg13g2_mux4_1 _16111_ (.S0(net771),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][10] ),
    .S1(net770),
    .X(_09284_));
 sg13g2_mux4_1 _16112_ (.S0(net889),
    .A0(_09281_),
    .A1(_09282_),
    .A2(_09283_),
    .A3(_09284_),
    .S1(net888),
    .X(_09285_));
 sg13g2_nand2_1 _16113_ (.Y(_09286_),
    .A(net776),
    .B(_09285_));
 sg13g2_mux4_1 _16114_ (.S0(net767),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][10] ),
    .S1(net766),
    .X(_09287_));
 sg13g2_mux4_1 _16115_ (.S0(net767),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][10] ),
    .S1(net766),
    .X(_09288_));
 sg13g2_mux4_1 _16116_ (.S0(net771),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][10] ),
    .S1(net770),
    .X(_09289_));
 sg13g2_mux4_1 _16117_ (.S0(_09235_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][10] ),
    .S1(net770),
    .X(_09290_));
 sg13g2_mux4_1 _16118_ (.S0(_09241_),
    .A0(_09287_),
    .A1(_09288_),
    .A2(_09289_),
    .A3(_09290_),
    .S1(_09242_),
    .X(_09291_));
 sg13g2_nand2_1 _16119_ (.Y(_09292_),
    .A(_09198_),
    .B(_09291_));
 sg13g2_a21oi_2 _16120_ (.B1(_08380_),
    .Y(_09293_),
    .A2(_09292_),
    .A1(_09286_));
 sg13g2_buf_1 _16121_ (.A(_09293_),
    .X(_09294_));
 sg13g2_nor2b_1 _16122_ (.A(net1036),
    .B_N(net1032),
    .Y(_09295_));
 sg13g2_buf_1 _16123_ (.A(_09295_),
    .X(_09296_));
 sg13g2_buf_1 _16124_ (.A(_09296_),
    .X(_09297_));
 sg13g2_mux2_1 _16125_ (.A0(\cpu.dcache.r_tag[5][22] ),
    .A1(\cpu.dcache.r_tag[7][22] ),
    .S(net780),
    .X(_09298_));
 sg13g2_a22oi_1 _16126_ (.Y(_09299_),
    .B1(_09298_),
    .B2(net686),
    .A2(_09297_),
    .A1(\cpu.dcache.r_tag[6][22] ));
 sg13g2_buf_1 _16127_ (.A(_09263_),
    .X(_09300_));
 sg13g2_and2_1 _16128_ (.A(net1112),
    .B(net1108),
    .X(_09301_));
 sg13g2_buf_2 _16129_ (.A(_09301_),
    .X(_09302_));
 sg13g2_nor2_1 _16130_ (.A(_09229_),
    .B(_09302_),
    .Y(_09303_));
 sg13g2_buf_1 _16131_ (.A(_09303_),
    .X(_09304_));
 sg13g2_inv_2 _16132_ (.Y(_09305_),
    .A(net1028));
 sg13g2_buf_1 _16133_ (.A(net1035),
    .X(_09306_));
 sg13g2_mux2_1 _16134_ (.A0(\cpu.dcache.r_tag[1][22] ),
    .A1(\cpu.dcache.r_tag[3][22] ),
    .S(net887),
    .X(_09307_));
 sg13g2_a22oi_1 _16135_ (.Y(_09308_),
    .B1(_09307_),
    .B2(net782),
    .A2(_09296_),
    .A1(\cpu.dcache.r_tag[2][22] ));
 sg13g2_nor2_1 _16136_ (.A(_09305_),
    .B(_09308_),
    .Y(_09309_));
 sg13g2_a221oi_1 _16137_ (.B2(\cpu.dcache.r_tag[0][22] ),
    .C1(_09309_),
    .B1(_09304_),
    .A1(\cpu.dcache.r_tag[4][22] ),
    .Y(_09310_),
    .A2(_09300_));
 sg13g2_o21ai_1 _16138_ (.B1(_09310_),
    .Y(_09311_),
    .A1(net895),
    .A2(_09299_));
 sg13g2_xor2_1 _16139_ (.B(_09311_),
    .A(net430),
    .X(_09312_));
 sg13g2_buf_1 _16140_ (.A(net1058),
    .X(_09313_));
 sg13g2_mux4_1 _16141_ (.S0(net767),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][2] ),
    .S1(_09280_),
    .X(_09314_));
 sg13g2_mux4_1 _16142_ (.S0(net767),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][2] ),
    .S1(net766),
    .X(_09315_));
 sg13g2_mux4_1 _16143_ (.S0(net771),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][2] ),
    .S1(net770),
    .X(_09316_));
 sg13g2_mux4_1 _16144_ (.S0(_09235_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][2] ),
    .S1(_09236_),
    .X(_09317_));
 sg13g2_mux4_1 _16145_ (.S0(_09197_),
    .A0(_09314_),
    .A1(_09315_),
    .A2(_09316_),
    .A3(_09317_),
    .S1(net888),
    .X(_09318_));
 sg13g2_nand2_1 _16146_ (.Y(_09319_),
    .A(_08184_),
    .B(_09318_));
 sg13g2_buf_2 _16147_ (.A(_09186_),
    .X(_09320_));
 sg13g2_mux4_1 _16148_ (.S0(_09279_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][2] ),
    .S1(net765),
    .X(_09321_));
 sg13g2_buf_2 _16149_ (.A(_09184_),
    .X(_09322_));
 sg13g2_mux4_1 _16150_ (.S0(net764),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][2] ),
    .S1(net765),
    .X(_09323_));
 sg13g2_mux4_1 _16151_ (.S0(net771),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][2] ),
    .S1(net770),
    .X(_09324_));
 sg13g2_mux4_1 _16152_ (.S0(_09279_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][2] ),
    .S1(_09280_),
    .X(_09325_));
 sg13g2_mux4_1 _16153_ (.S0(_09197_),
    .A0(_09321_),
    .A1(_09323_),
    .A2(_09324_),
    .A3(_09325_),
    .S1(net888),
    .X(_09326_));
 sg13g2_o21ai_1 _16154_ (.B1(net886),
    .Y(_09327_),
    .A1(_08470_),
    .A2(_09326_));
 sg13g2_o21ai_1 _16155_ (.B1(_09327_),
    .Y(_09328_),
    .A1(_09313_),
    .A2(_09319_));
 sg13g2_buf_1 _16156_ (.A(_09328_),
    .X(_09329_));
 sg13g2_buf_1 _16157_ (.A(_09212_),
    .X(_09330_));
 sg13g2_nor2_1 _16158_ (.A(net891),
    .B(net895),
    .Y(_09331_));
 sg13g2_mux2_1 _16159_ (.A0(\cpu.dcache.r_tag[5][14] ),
    .A1(\cpu.dcache.r_tag[7][14] ),
    .S(net898),
    .X(_09332_));
 sg13g2_inv_1 _16160_ (.Y(_09333_),
    .A(\cpu.dcache.r_tag[4][14] ));
 sg13g2_nand2b_1 _16161_ (.Y(_09334_),
    .B(net1029),
    .A_N(_09100_));
 sg13g2_buf_2 _16162_ (.A(_09334_),
    .X(_09335_));
 sg13g2_nand3_1 _16163_ (.B(net1108),
    .C(\cpu.dcache.r_tag[2][14] ),
    .A(net898),
    .Y(_09336_));
 sg13g2_o21ai_1 _16164_ (.B1(_09336_),
    .Y(_09337_),
    .A1(_09333_),
    .A2(_09335_));
 sg13g2_inv_1 _16165_ (.Y(_09338_),
    .A(\cpu.dcache.r_tag[6][14] ));
 sg13g2_nand3b_1 _16166_ (.B(net1029),
    .C(net1032),
    .Y(_09339_),
    .A_N(net1112));
 sg13g2_buf_1 _16167_ (.A(_09339_),
    .X(_09340_));
 sg13g2_nand4_1 _16168_ (.B(net898),
    .C(net1108),
    .A(net900),
    .Y(_09341_),
    .D(\cpu.dcache.r_tag[3][14] ));
 sg13g2_o21ai_1 _16169_ (.B1(_09341_),
    .Y(_09342_),
    .A1(_09338_),
    .A2(_09340_));
 sg13g2_a221oi_1 _16170_ (.B2(net891),
    .C1(_09342_),
    .B1(_09337_),
    .A1(_09331_),
    .Y(_09343_),
    .A2(_09332_));
 sg13g2_mux2_1 _16171_ (.A0(_00223_),
    .A1(_09343_),
    .S(net772),
    .X(_09344_));
 sg13g2_nor2_1 _16172_ (.A(\cpu.dcache.r_tag[1][14] ),
    .B(_09212_),
    .Y(_09345_));
 sg13g2_a22oi_1 _16173_ (.Y(_09346_),
    .B1(_09345_),
    .B2(_09343_),
    .A2(_09344_),
    .A1(net531));
 sg13g2_xor2_1 _16174_ (.B(_09346_),
    .A(net429),
    .X(_09347_));
 sg13g2_nor4_1 _16175_ (.A(_09234_),
    .B(_09278_),
    .C(_09312_),
    .D(_09347_),
    .Y(_09348_));
 sg13g2_mux4_1 _16176_ (.S0(net775),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][5] ),
    .S1(net774),
    .X(_09349_));
 sg13g2_mux4_1 _16177_ (.S0(net775),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][5] ),
    .S1(net774),
    .X(_09350_));
 sg13g2_mux4_1 _16178_ (.S0(net893),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][5] ),
    .S1(net773),
    .X(_09351_));
 sg13g2_mux4_1 _16179_ (.S0(net894),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][5] ),
    .S1(net773),
    .X(_09352_));
 sg13g2_mux4_1 _16180_ (.S0(_08161_),
    .A0(_09349_),
    .A1(_09350_),
    .A2(_09351_),
    .A3(_09352_),
    .S1(net1057),
    .X(_09353_));
 sg13g2_nand2_1 _16181_ (.Y(_09354_),
    .A(_08136_),
    .B(_09353_));
 sg13g2_mux4_1 _16182_ (.S0(_09190_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][5] ),
    .S1(_09191_),
    .X(_09355_));
 sg13g2_mux4_1 _16183_ (.S0(net775),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][5] ),
    .S1(net774),
    .X(_09356_));
 sg13g2_mux4_1 _16184_ (.S0(net893),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][5] ),
    .S1(net892),
    .X(_09357_));
 sg13g2_mux4_1 _16185_ (.S0(net893),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][5] ),
    .S1(net892),
    .X(_09358_));
 sg13g2_mux4_1 _16186_ (.S0(_08161_),
    .A0(_09355_),
    .A1(_09356_),
    .A2(_09357_),
    .A3(_09358_),
    .S1(_08169_),
    .X(_09359_));
 sg13g2_nand2_1 _16187_ (.Y(_09360_),
    .A(net682),
    .B(_09359_));
 sg13g2_a21oi_2 _16188_ (.B1(_08380_),
    .Y(_09361_),
    .A2(_09360_),
    .A1(_09354_));
 sg13g2_buf_1 _16189_ (.A(_09361_),
    .X(_09362_));
 sg13g2_mux2_1 _16190_ (.A0(\cpu.dcache.r_tag[1][17] ),
    .A1(\cpu.dcache.r_tag[3][17] ),
    .S(net780),
    .X(_09363_));
 sg13g2_a22oi_1 _16191_ (.Y(_09364_),
    .B1(_09363_),
    .B2(net686),
    .A2(_09296_),
    .A1(\cpu.dcache.r_tag[2][17] ));
 sg13g2_inv_1 _16192_ (.Y(_09365_),
    .A(_00226_));
 sg13g2_nor2b_1 _16193_ (.A(net1035),
    .B_N(net1036),
    .Y(_09366_));
 sg13g2_buf_2 _16194_ (.A(_09366_),
    .X(_09367_));
 sg13g2_mux2_1 _16195_ (.A0(\cpu.dcache.r_tag[4][17] ),
    .A1(\cpu.dcache.r_tag[6][17] ),
    .S(net898),
    .X(_09368_));
 sg13g2_a22oi_1 _16196_ (.Y(_09369_),
    .B1(_09368_),
    .B2(net891),
    .A2(_09367_),
    .A1(\cpu.dcache.r_tag[5][17] ));
 sg13g2_nor2_1 _16197_ (.A(net895),
    .B(_09369_),
    .Y(_09370_));
 sg13g2_a221oi_1 _16198_ (.B2(_09365_),
    .C1(_09370_),
    .B1(_09304_),
    .A1(\cpu.dcache.r_tag[7][17] ),
    .Y(_09371_),
    .A2(net769));
 sg13g2_o21ai_1 _16199_ (.B1(_09371_),
    .Y(_09372_),
    .A1(_09305_),
    .A2(_09364_));
 sg13g2_xor2_1 _16200_ (.B(_09372_),
    .A(net428),
    .X(_09373_));
 sg13g2_nand2b_1 _16201_ (.Y(_09374_),
    .B(_09304_),
    .A_N(_00224_));
 sg13g2_a22oi_1 _16202_ (.Y(_09375_),
    .B1(_09273_),
    .B2(\cpu.dcache.r_tag[5][15] ),
    .A2(_09254_),
    .A1(\cpu.dcache.r_tag[3][15] ));
 sg13g2_a22oi_1 _16203_ (.Y(_09376_),
    .B1(_09267_),
    .B2(\cpu.dcache.r_tag[2][15] ),
    .A2(_09258_),
    .A1(\cpu.dcache.r_tag[1][15] ));
 sg13g2_mux2_1 _16204_ (.A0(\cpu.dcache.r_tag[4][15] ),
    .A1(\cpu.dcache.r_tag[6][15] ),
    .S(net887),
    .X(_09377_));
 sg13g2_and2_1 _16205_ (.A(net1112),
    .B(net1032),
    .X(_09378_));
 sg13g2_buf_2 _16206_ (.A(_09378_),
    .X(_09379_));
 sg13g2_a22oi_1 _16207_ (.Y(_09380_),
    .B1(_09379_),
    .B2(\cpu.dcache.r_tag[7][15] ),
    .A2(_09377_),
    .A1(net891));
 sg13g2_buf_1 _16208_ (.A(_09218_),
    .X(_09381_));
 sg13g2_buf_1 _16209_ (.A(net885),
    .X(_09382_));
 sg13g2_nand2b_1 _16210_ (.Y(_09383_),
    .B(net763),
    .A_N(_09380_));
 sg13g2_nand4_1 _16211_ (.B(_09375_),
    .C(_09376_),
    .A(_09374_),
    .Y(_09384_),
    .D(_09383_));
 sg13g2_buf_1 _16212_ (.A(_08169_),
    .X(_09385_));
 sg13g2_mux4_1 _16213_ (.S0(net893),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][3] ),
    .S1(_09202_),
    .X(_09386_));
 sg13g2_mux4_1 _16214_ (.S0(_09201_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][3] ),
    .S1(net892),
    .X(_09387_));
 sg13g2_mux4_1 _16215_ (.S0(net893),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][3] ),
    .S1(_09202_),
    .X(_09388_));
 sg13g2_mux4_1 _16216_ (.S0(net893),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][3] ),
    .S1(net892),
    .X(_09389_));
 sg13g2_mux4_1 _16217_ (.S0(_09197_),
    .A0(_09386_),
    .A1(_09387_),
    .A2(_09388_),
    .A3(_09389_),
    .S1(_09313_),
    .X(_09390_));
 sg13g2_nand2_1 _16218_ (.Y(_09391_),
    .A(net1056),
    .B(_09390_));
 sg13g2_mux4_1 _16219_ (.S0(net894),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][3] ),
    .S1(net774),
    .X(_09392_));
 sg13g2_mux4_1 _16220_ (.S0(_09185_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][3] ),
    .S1(_09187_),
    .X(_09393_));
 sg13g2_mux4_1 _16221_ (.S0(net893),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][3] ),
    .S1(net892),
    .X(_09394_));
 sg13g2_mux4_1 _16222_ (.S0(_09201_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][3] ),
    .S1(net892),
    .X(_09395_));
 sg13g2_mux4_1 _16223_ (.S0(_09197_),
    .A0(_09392_),
    .A1(_09393_),
    .A2(_09394_),
    .A3(_09395_),
    .S1(net886),
    .X(_09396_));
 sg13g2_o21ai_1 _16224_ (.B1(_09385_),
    .Y(_09397_),
    .A1(_08470_),
    .A2(_09396_));
 sg13g2_o21ai_1 _16225_ (.B1(_09397_),
    .Y(_09398_),
    .A1(net884),
    .A2(_09391_));
 sg13g2_buf_1 _16226_ (.A(_09398_),
    .X(_09399_));
 sg13g2_xor2_1 _16227_ (.B(net427),
    .A(_09384_),
    .X(_09400_));
 sg13g2_buf_2 _16228_ (.A(net771),
    .X(_09401_));
 sg13g2_buf_2 _16229_ (.A(net766),
    .X(_09402_));
 sg13g2_mux4_1 _16230_ (.S0(net679),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][11] ),
    .S1(net678),
    .X(_09403_));
 sg13g2_mux4_1 _16231_ (.S0(net679),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][11] ),
    .S1(net678),
    .X(_09404_));
 sg13g2_mux4_1 _16232_ (.S0(net679),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][11] ),
    .S1(net678),
    .X(_09405_));
 sg13g2_mux4_1 _16233_ (.S0(net679),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][11] ),
    .S1(net678),
    .X(_09406_));
 sg13g2_mux4_1 _16234_ (.S0(net886),
    .A0(_09403_),
    .A1(_09404_),
    .A2(_09405_),
    .A3(_09406_),
    .S1(net884),
    .X(_09407_));
 sg13g2_nand2_1 _16235_ (.Y(_09408_),
    .A(net776),
    .B(_09407_));
 sg13g2_mux4_1 _16236_ (.S0(net679),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][11] ),
    .S1(net678),
    .X(_09409_));
 sg13g2_mux4_1 _16237_ (.S0(_09401_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][11] ),
    .S1(net678),
    .X(_09410_));
 sg13g2_buf_2 _16238_ (.A(_09184_),
    .X(_09411_));
 sg13g2_buf_2 _16239_ (.A(net892),
    .X(_09412_));
 sg13g2_mux4_1 _16240_ (.S0(_09411_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][11] ),
    .S1(net761),
    .X(_09413_));
 sg13g2_mux4_1 _16241_ (.S0(net762),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][11] ),
    .S1(net761),
    .X(_09414_));
 sg13g2_mux4_1 _16242_ (.S0(net886),
    .A0(_09409_),
    .A1(_09410_),
    .A2(_09413_),
    .A3(_09414_),
    .S1(net884),
    .X(_09415_));
 sg13g2_nand2_1 _16243_ (.Y(_09416_),
    .A(_09198_),
    .B(_09415_));
 sg13g2_a21oi_2 _16244_ (.B1(_08381_),
    .Y(_09417_),
    .A2(_09416_),
    .A1(_09408_));
 sg13g2_nand2_1 _16245_ (.Y(_09418_),
    .A(\cpu.dcache.r_tag[3][23] ),
    .B(_09255_));
 sg13g2_and2_1 _16246_ (.A(net1035),
    .B(_09261_),
    .X(_09419_));
 sg13g2_buf_1 _16247_ (.A(_09419_),
    .X(_09420_));
 sg13g2_a22oi_1 _16248_ (.Y(_09421_),
    .B1(net677),
    .B2(\cpu.dcache.r_tag[6][23] ),
    .A2(_09259_),
    .A1(\cpu.dcache.r_tag[1][23] ));
 sg13g2_inv_1 _16249_ (.Y(_09422_),
    .A(_00229_));
 sg13g2_a22oi_1 _16250_ (.Y(_09423_),
    .B1(_09304_),
    .B2(_09422_),
    .A2(_09267_),
    .A1(\cpu.dcache.r_tag[2][23] ));
 sg13g2_mux2_1 _16251_ (.A0(\cpu.dcache.r_tag[5][23] ),
    .A1(\cpu.dcache.r_tag[7][23] ),
    .S(net887),
    .X(_09424_));
 sg13g2_nor2_1 _16252_ (.A(net1112),
    .B(net1032),
    .Y(_09425_));
 sg13g2_buf_2 _16253_ (.A(_09425_),
    .X(_09426_));
 sg13g2_a22oi_1 _16254_ (.Y(_09427_),
    .B1(_09426_),
    .B2(\cpu.dcache.r_tag[4][23] ),
    .A2(_09424_),
    .A1(net782));
 sg13g2_nand2b_1 _16255_ (.Y(_09428_),
    .B(net763),
    .A_N(_09427_));
 sg13g2_nand4_1 _16256_ (.B(_09421_),
    .C(_09423_),
    .A(_09418_),
    .Y(_09429_),
    .D(_09428_));
 sg13g2_xor2_1 _16257_ (.B(_09429_),
    .A(_09417_),
    .X(_09430_));
 sg13g2_buf_2 _16258_ (.A(_09184_),
    .X(_09431_));
 sg13g2_buf_2 _16259_ (.A(_09186_),
    .X(_09432_));
 sg13g2_mux4_1 _16260_ (.S0(net760),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][9] ),
    .S1(net759),
    .X(_09433_));
 sg13g2_mux4_1 _16261_ (.S0(net760),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][9] ),
    .S1(net759),
    .X(_09434_));
 sg13g2_mux4_1 _16262_ (.S0(net764),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][9] ),
    .S1(net765),
    .X(_09435_));
 sg13g2_mux4_1 _16263_ (.S0(net764),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][9] ),
    .S1(net765),
    .X(_09436_));
 sg13g2_mux4_1 _16264_ (.S0(net889),
    .A0(_09433_),
    .A1(_09434_),
    .A2(_09435_),
    .A3(_09436_),
    .S1(net888),
    .X(_09437_));
 sg13g2_nand2_1 _16265_ (.Y(_09438_),
    .A(net776),
    .B(_09437_));
 sg13g2_mux4_1 _16266_ (.S0(net764),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][9] ),
    .S1(_09432_),
    .X(_09439_));
 sg13g2_mux4_1 _16267_ (.S0(_09431_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][9] ),
    .S1(_09432_),
    .X(_09440_));
 sg13g2_mux4_1 _16268_ (.S0(net767),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][9] ),
    .S1(net766),
    .X(_09441_));
 sg13g2_mux4_1 _16269_ (.S0(net767),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][9] ),
    .S1(net766),
    .X(_09442_));
 sg13g2_mux4_1 _16270_ (.S0(net889),
    .A0(_09439_),
    .A1(_09440_),
    .A2(_09441_),
    .A3(_09442_),
    .S1(net888),
    .X(_09443_));
 sg13g2_nand2_1 _16271_ (.Y(_09444_),
    .A(net682),
    .B(_09443_));
 sg13g2_a21oi_2 _16272_ (.B1(_08380_),
    .Y(_09445_),
    .A2(_09444_),
    .A1(_09438_));
 sg13g2_buf_1 _16273_ (.A(_09445_),
    .X(_09446_));
 sg13g2_buf_1 _16274_ (.A(_09304_),
    .X(_09447_));
 sg13g2_nand2_1 _16275_ (.Y(_09448_),
    .A(\cpu.dcache.r_tag[0][21] ),
    .B(_09447_));
 sg13g2_buf_1 _16276_ (.A(_09267_),
    .X(_09449_));
 sg13g2_a22oi_1 _16277_ (.Y(_09450_),
    .B1(_09449_),
    .B2(\cpu.dcache.r_tag[2][21] ),
    .A2(_09259_),
    .A1(\cpu.dcache.r_tag[1][21] ));
 sg13g2_a22oi_1 _16278_ (.Y(_09451_),
    .B1(_09255_),
    .B2(\cpu.dcache.r_tag[3][21] ),
    .A2(net769),
    .A1(\cpu.dcache.r_tag[7][21] ));
 sg13g2_mux2_1 _16279_ (.A0(\cpu.dcache.r_tag[4][21] ),
    .A1(\cpu.dcache.r_tag[6][21] ),
    .S(net780),
    .X(_09452_));
 sg13g2_a22oi_1 _16280_ (.Y(_09453_),
    .B1(_09452_),
    .B2(net768),
    .A2(_09367_),
    .A1(\cpu.dcache.r_tag[5][21] ));
 sg13g2_nand2b_1 _16281_ (.Y(_09454_),
    .B(_09382_),
    .A_N(_09453_));
 sg13g2_nand4_1 _16282_ (.B(_09450_),
    .C(_09451_),
    .A(_09448_),
    .Y(_09455_),
    .D(_09454_));
 sg13g2_xor2_1 _16283_ (.B(_09455_),
    .A(net426),
    .X(_09456_));
 sg13g2_nor4_1 _16284_ (.A(_09373_),
    .B(_09400_),
    .C(_09430_),
    .D(_09456_),
    .Y(_09457_));
 sg13g2_nand2_1 _16285_ (.Y(_09458_),
    .A(_09348_),
    .B(_09457_));
 sg13g2_mux2_1 _16286_ (.A0(\cpu.dcache.r_tag[4][13] ),
    .A1(\cpu.dcache.r_tag[6][13] ),
    .S(net780),
    .X(_09459_));
 sg13g2_a22oi_1 _16287_ (.Y(_09460_),
    .B1(_09459_),
    .B2(net768),
    .A2(_09379_),
    .A1(\cpu.dcache.r_tag[7][13] ));
 sg13g2_nor2_1 _16288_ (.A(_09171_),
    .B(net1032),
    .Y(_09461_));
 sg13g2_buf_1 _16289_ (.A(_09461_),
    .X(_09462_));
 sg13g2_nand2b_1 _16290_ (.Y(_09463_),
    .B(net758),
    .A_N(_09302_));
 sg13g2_buf_2 _16291_ (.A(_09463_),
    .X(_09464_));
 sg13g2_a22oi_1 _16292_ (.Y(_09465_),
    .B1(_09273_),
    .B2(\cpu.dcache.r_tag[5][13] ),
    .A2(_09254_),
    .A1(\cpu.dcache.r_tag[3][13] ));
 sg13g2_o21ai_1 _16293_ (.B1(_09465_),
    .Y(_09466_),
    .A1(_00222_),
    .A2(_09464_));
 sg13g2_a221oi_1 _16294_ (.B2(\cpu.dcache.r_tag[2][13] ),
    .C1(_09466_),
    .B1(_09449_),
    .A1(\cpu.dcache.r_tag[1][13] ),
    .Y(_09467_),
    .A2(net605));
 sg13g2_o21ai_1 _16295_ (.B1(_09467_),
    .Y(_09468_),
    .A1(net895),
    .A2(_09460_));
 sg13g2_mux4_1 _16296_ (.S0(net762),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][1] ),
    .S1(_09402_),
    .X(_09469_));
 sg13g2_mux4_1 _16297_ (.S0(_09401_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][1] ),
    .S1(_09402_),
    .X(_09470_));
 sg13g2_mux4_1 _16298_ (.S0(net762),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][1] ),
    .S1(_09412_),
    .X(_09471_));
 sg13g2_mux4_1 _16299_ (.S0(net762),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][1] ),
    .S1(_09412_),
    .X(_09472_));
 sg13g2_mux4_1 _16300_ (.S0(net886),
    .A0(_09469_),
    .A1(_09470_),
    .A2(_09471_),
    .A3(_09472_),
    .S1(net884),
    .X(_09473_));
 sg13g2_buf_2 _16301_ (.A(_09186_),
    .X(_09474_));
 sg13g2_mux4_1 _16302_ (.S0(net760),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][1] ),
    .S1(_09474_),
    .X(_09475_));
 sg13g2_buf_2 _16303_ (.A(_09184_),
    .X(_09476_));
 sg13g2_mux4_1 _16304_ (.S0(net756),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][1] ),
    .S1(net757),
    .X(_09477_));
 sg13g2_mux4_1 _16305_ (.S0(net764),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][1] ),
    .S1(net765),
    .X(_09478_));
 sg13g2_mux4_1 _16306_ (.S0(net764),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][1] ),
    .S1(net765),
    .X(_09479_));
 sg13g2_mux4_1 _16307_ (.S0(_09241_),
    .A0(_09475_),
    .A1(_09477_),
    .A2(_09478_),
    .A3(_09479_),
    .S1(_09242_),
    .X(_09480_));
 sg13g2_and2_1 _16308_ (.A(net776),
    .B(_09480_),
    .X(_09481_));
 sg13g2_a21oi_1 _16309_ (.A1(net682),
    .A2(_09473_),
    .Y(_09482_),
    .B1(_09481_));
 sg13g2_buf_1 _16310_ (.A(net678),
    .X(_09483_));
 sg13g2_nor2_1 _16311_ (.A(net920),
    .B(net601),
    .Y(_09484_));
 sg13g2_a21oi_1 _16312_ (.A1(net920),
    .A2(_09482_),
    .Y(_09485_),
    .B1(_09484_));
 sg13g2_buf_1 _16313_ (.A(_09485_),
    .X(_09486_));
 sg13g2_xnor2_1 _16314_ (.Y(_09487_),
    .A(_09468_),
    .B(_09486_));
 sg13g2_mux4_1 _16315_ (.S0(net762),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][0] ),
    .S1(net761),
    .X(_09488_));
 sg13g2_mux4_1 _16316_ (.S0(_09411_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][0] ),
    .S1(net761),
    .X(_09489_));
 sg13g2_mux4_1 _16317_ (.S0(net762),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][0] ),
    .S1(net761),
    .X(_09490_));
 sg13g2_mux4_1 _16318_ (.S0(net762),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][0] ),
    .S1(net761),
    .X(_09491_));
 sg13g2_mux4_1 _16319_ (.S0(net886),
    .A0(_09488_),
    .A1(_09489_),
    .A2(_09490_),
    .A3(_09491_),
    .S1(net884),
    .X(_09492_));
 sg13g2_mux4_1 _16320_ (.S0(_09431_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][0] ),
    .S1(net759),
    .X(_09493_));
 sg13g2_mux4_1 _16321_ (.S0(net760),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][0] ),
    .S1(net759),
    .X(_09494_));
 sg13g2_mux4_1 _16322_ (.S0(_09322_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][0] ),
    .S1(_09320_),
    .X(_09495_));
 sg13g2_mux4_1 _16323_ (.S0(_09322_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][0] ),
    .S1(_09320_),
    .X(_09496_));
 sg13g2_mux4_1 _16324_ (.S0(net889),
    .A0(_09493_),
    .A1(_09494_),
    .A2(_09495_),
    .A3(_09496_),
    .S1(net888),
    .X(_09497_));
 sg13g2_and2_1 _16325_ (.A(_09183_),
    .B(_09497_),
    .X(_09498_));
 sg13g2_a21oi_1 _16326_ (.A1(net682),
    .A2(_09492_),
    .Y(_09499_),
    .B1(_09498_));
 sg13g2_nor2_1 _16327_ (.A(net1056),
    .B(net679),
    .Y(_09500_));
 sg13g2_a21oi_1 _16328_ (.A1(net920),
    .A2(_09499_),
    .Y(_09501_),
    .B1(_09500_));
 sg13g2_buf_1 _16329_ (.A(_09501_),
    .X(_09502_));
 sg13g2_a22oi_1 _16330_ (.Y(_09503_),
    .B1(net677),
    .B2(\cpu.dcache.r_tag[6][12] ),
    .A2(_09273_),
    .A1(\cpu.dcache.r_tag[5][12] ));
 sg13g2_a22oi_1 _16331_ (.Y(_09504_),
    .B1(_09267_),
    .B2(\cpu.dcache.r_tag[2][12] ),
    .A2(net769),
    .A1(\cpu.dcache.r_tag[7][12] ));
 sg13g2_a22oi_1 _16332_ (.Y(_09505_),
    .B1(_09263_),
    .B2(\cpu.dcache.r_tag[4][12] ),
    .A2(_09254_),
    .A1(\cpu.dcache.r_tag[3][12] ));
 sg13g2_and3_1 _16333_ (.X(_09506_),
    .A(_09503_),
    .B(_09504_),
    .C(_09505_));
 sg13g2_mux2_1 _16334_ (.A0(_00221_),
    .A1(_09506_),
    .S(net772),
    .X(_09507_));
 sg13g2_nor2_1 _16335_ (.A(\cpu.dcache.r_tag[1][12] ),
    .B(net531),
    .Y(_09508_));
 sg13g2_a22oi_1 _16336_ (.Y(_09509_),
    .B1(_09508_),
    .B2(_09506_),
    .A2(_09507_),
    .A1(_09330_));
 sg13g2_xnor2_1 _16337_ (.Y(_09510_),
    .A(net376),
    .B(_09509_));
 sg13g2_nand2_1 _16338_ (.Y(_09511_),
    .A(_09487_),
    .B(_09510_));
 sg13g2_mux2_1 _16339_ (.A0(\cpu.dcache.r_tag[5][9] ),
    .A1(\cpu.dcache.r_tag[7][9] ),
    .S(net780),
    .X(_09512_));
 sg13g2_a22oi_1 _16340_ (.Y(_09513_),
    .B1(_09512_),
    .B2(net782),
    .A2(_09426_),
    .A1(\cpu.dcache.r_tag[4][9] ));
 sg13g2_nor2_1 _16341_ (.A(net895),
    .B(_09513_),
    .Y(_09514_));
 sg13g2_mux2_1 _16342_ (.A0(\cpu.dcache.r_tag[1][9] ),
    .A1(\cpu.dcache.r_tag[3][9] ),
    .S(net887),
    .X(_09515_));
 sg13g2_a22oi_1 _16343_ (.Y(_09516_),
    .B1(_09515_),
    .B2(net782),
    .A2(_09296_),
    .A1(\cpu.dcache.r_tag[2][9] ));
 sg13g2_nand3_1 _16344_ (.B(_09306_),
    .C(\cpu.dcache.r_tag[6][9] ),
    .A(net1029),
    .Y(_09517_));
 sg13g2_o21ai_1 _16345_ (.B1(_09517_),
    .Y(_09518_),
    .A1(_00216_),
    .A2(_09229_));
 sg13g2_nor3_1 _16346_ (.A(net1028),
    .B(_00216_),
    .C(_09229_),
    .Y(_09519_));
 sg13g2_a21oi_1 _16347_ (.A1(_09269_),
    .A2(_09518_),
    .Y(_09520_),
    .B1(_09519_));
 sg13g2_o21ai_1 _16348_ (.B1(_09520_),
    .Y(_09521_),
    .A1(_09305_),
    .A2(_09516_));
 sg13g2_nor2_1 _16349_ (.A(_09514_),
    .B(_09521_),
    .Y(_09522_));
 sg13g2_xor2_1 _16350_ (.B(_09522_),
    .A(_00215_),
    .X(_09523_));
 sg13g2_a22oi_1 _16351_ (.Y(_09524_),
    .B1(_09302_),
    .B2(\cpu.dcache.r_tag[3][8] ),
    .A2(_09261_),
    .A1(\cpu.dcache.r_tag[6][8] ));
 sg13g2_nand2_1 _16352_ (.Y(_09525_),
    .A(net780),
    .B(_09524_));
 sg13g2_a22oi_1 _16353_ (.Y(_09526_),
    .B1(_09302_),
    .B2(\cpu.dcache.r_tag[1][8] ),
    .A2(_09261_),
    .A1(\cpu.dcache.r_tag[4][8] ));
 sg13g2_nand2_1 _16354_ (.Y(_09527_),
    .A(_09051_),
    .B(_09526_));
 sg13g2_and2_1 _16355_ (.A(net900),
    .B(\cpu.dcache.r_tag[5][8] ),
    .X(_09528_));
 sg13g2_a22oi_1 _16356_ (.Y(_09529_),
    .B1(_09528_),
    .B2(_09219_),
    .A2(_09267_),
    .A1(\cpu.dcache.r_tag[2][8] ));
 sg13g2_o21ai_1 _16357_ (.B1(_09529_),
    .Y(_09530_),
    .A1(_00214_),
    .A2(_09464_));
 sg13g2_a221oi_1 _16358_ (.B2(_09527_),
    .C1(_09530_),
    .B1(_09525_),
    .A1(\cpu.dcache.r_tag[7][8] ),
    .Y(_09531_),
    .A2(_09265_));
 sg13g2_xor2_1 _16359_ (.B(_09531_),
    .A(_00213_),
    .X(_09532_));
 sg13g2_a22oi_1 _16360_ (.Y(_09533_),
    .B1(\cpu.dcache.r_tag[3][10] ),
    .B2(net1028),
    .A2(\cpu.dcache.r_tag[7][10] ),
    .A1(net885));
 sg13g2_a221oi_1 _16361_ (.B2(net1028),
    .C1(net782),
    .B1(\cpu.dcache.r_tag[2][10] ),
    .A1(net885),
    .Y(_09534_),
    .A2(\cpu.dcache.r_tag[6][10] ));
 sg13g2_a21oi_1 _16362_ (.A1(_09036_),
    .A2(_09533_),
    .Y(_09535_),
    .B1(_09534_));
 sg13g2_mux2_1 _16363_ (.A0(\cpu.dcache.r_tag[4][10] ),
    .A1(\cpu.dcache.r_tag[5][10] ),
    .S(net900),
    .X(_09536_));
 sg13g2_nor3_1 _16364_ (.A(net885),
    .B(_00218_),
    .C(_09302_),
    .Y(_09537_));
 sg13g2_a221oi_1 _16365_ (.B2(net885),
    .C1(_09537_),
    .B1(_09536_),
    .A1(\cpu.dcache.r_tag[1][10] ),
    .Y(_09538_),
    .A2(_09302_));
 sg13g2_nand2_1 _16366_ (.Y(_09539_),
    .A(_09051_),
    .B(_09538_));
 sg13g2_o21ai_1 _16367_ (.B1(_09539_),
    .Y(_09540_),
    .A1(_09051_),
    .A2(_09535_));
 sg13g2_xor2_1 _16368_ (.B(_09540_),
    .A(_00217_),
    .X(_09541_));
 sg13g2_buf_1 _16369_ (.A(_00207_),
    .X(_09542_));
 sg13g2_inv_1 _16370_ (.Y(_09543_),
    .A(_09542_));
 sg13g2_buf_1 _16371_ (.A(_09543_),
    .X(_09544_));
 sg13g2_a22oi_1 _16372_ (.Y(_09545_),
    .B1(\cpu.dcache.r_tag[3][5] ),
    .B2(_09209_),
    .A2(\cpu.dcache.r_tag[7][5] ),
    .A1(net1029));
 sg13g2_nand3b_1 _16373_ (.B(net1028),
    .C(\cpu.dcache.r_tag[2][5] ),
    .Y(_09546_),
    .A_N(net900));
 sg13g2_o21ai_1 _16374_ (.B1(_09546_),
    .Y(_09547_),
    .A1(_09217_),
    .A2(_09545_));
 sg13g2_nand2_1 _16375_ (.Y(_09548_),
    .A(_09102_),
    .B(_09547_));
 sg13g2_nand3_1 _16376_ (.B(net887),
    .C(\cpu.dcache.r_tag[6][5] ),
    .A(net1029),
    .Y(_09549_));
 sg13g2_o21ai_1 _16377_ (.B1(_09549_),
    .Y(_09550_),
    .A1(_00208_),
    .A2(net772));
 sg13g2_nand2_1 _16378_ (.Y(_09551_),
    .A(_09269_),
    .B(_09550_));
 sg13g2_mux2_1 _16379_ (.A0(\cpu.dcache.r_tag[4][5] ),
    .A1(\cpu.dcache.r_tag[5][5] ),
    .S(net900),
    .X(_09552_));
 sg13g2_nor3_1 _16380_ (.A(_09274_),
    .B(_00208_),
    .C(net772),
    .Y(_09553_));
 sg13g2_a221oi_1 _16381_ (.B2(_09552_),
    .C1(_09553_),
    .B1(_09219_),
    .A1(\cpu.dcache.r_tag[1][5] ),
    .Y(_09554_),
    .A2(_09258_));
 sg13g2_nand3_1 _16382_ (.B(_09551_),
    .C(_09554_),
    .A(_09548_),
    .Y(_09555_));
 sg13g2_xnor2_1 _16383_ (.Y(_09556_),
    .A(_09544_),
    .B(_09555_));
 sg13g2_mux2_1 _16384_ (.A0(\cpu.dcache.r_tag[4][6] ),
    .A1(\cpu.dcache.r_tag[6][6] ),
    .S(net1035),
    .X(_09557_));
 sg13g2_and3_1 _16385_ (.X(_09558_),
    .A(net1036),
    .B(net898),
    .C(\cpu.dcache.r_tag[7][6] ));
 sg13g2_a21o_1 _16386_ (.A2(_09557_),
    .A1(net891),
    .B1(_09558_),
    .X(_09559_));
 sg13g2_nand2_1 _16387_ (.Y(_09560_),
    .A(net887),
    .B(\cpu.dcache.r_tag[2][6] ));
 sg13g2_nand3b_1 _16388_ (.B(\cpu.dcache.r_tag[1][6] ),
    .C(net900),
    .Y(_09561_),
    .A_N(_09306_));
 sg13g2_o21ai_1 _16389_ (.B1(_09561_),
    .Y(_09562_),
    .A1(net782),
    .A2(_09560_));
 sg13g2_nand3_1 _16390_ (.B(net1108),
    .C(\cpu.dcache.r_tag[3][6] ),
    .A(net887),
    .Y(_09563_));
 sg13g2_nand3b_1 _16391_ (.B(\cpu.dcache.r_tag[5][6] ),
    .C(net1029),
    .Y(_09564_),
    .A_N(net887));
 sg13g2_a21oi_1 _16392_ (.A1(_09563_),
    .A2(_09564_),
    .Y(_09565_),
    .B1(net891));
 sg13g2_a221oi_1 _16393_ (.B2(_09274_),
    .C1(_09565_),
    .B1(_09562_),
    .A1(_09381_),
    .Y(_09566_),
    .A2(_09559_));
 sg13g2_o21ai_1 _16394_ (.B1(_09566_),
    .Y(_09567_),
    .A1(_00210_),
    .A2(_09464_));
 sg13g2_xor2_1 _16395_ (.B(_09567_),
    .A(_00209_),
    .X(_09568_));
 sg13g2_nand2_1 _16396_ (.Y(_09569_),
    .A(_09556_),
    .B(_09568_));
 sg13g2_nor4_1 _16397_ (.A(_09523_),
    .B(_09532_),
    .C(_09541_),
    .D(_09569_),
    .Y(_09570_));
 sg13g2_nand2_1 _16398_ (.Y(_09571_),
    .A(\cpu.dcache.r_tag[6][7] ),
    .B(net677));
 sg13g2_a22oi_1 _16399_ (.Y(_09572_),
    .B1(_09426_),
    .B2(\cpu.dcache.r_tag[4][7] ),
    .A2(_09379_),
    .A1(\cpu.dcache.r_tag[7][7] ));
 sg13g2_nand2b_1 _16400_ (.Y(_09573_),
    .B(net885),
    .A_N(_09572_));
 sg13g2_mux2_1 _16401_ (.A0(\cpu.dcache.r_tag[2][7] ),
    .A1(\cpu.dcache.r_tag[3][7] ),
    .S(net900),
    .X(_09574_));
 sg13g2_a22oi_1 _16402_ (.Y(_09575_),
    .B1(_09574_),
    .B2(net890),
    .A2(_09273_),
    .A1(\cpu.dcache.r_tag[5][7] ));
 sg13g2_nand3_1 _16403_ (.B(_09573_),
    .C(_09575_),
    .A(_09571_),
    .Y(_09576_));
 sg13g2_nand2_1 _16404_ (.Y(_09577_),
    .A(_00212_),
    .B(net758));
 sg13g2_o21ai_1 _16405_ (.B1(_09577_),
    .Y(_09578_),
    .A1(net758),
    .A2(_09576_));
 sg13g2_o21ai_1 _16406_ (.B1(net605),
    .Y(_09579_),
    .A1(\cpu.dcache.r_tag[1][7] ),
    .A2(_09576_));
 sg13g2_o21ai_1 _16407_ (.B1(_09579_),
    .Y(_09580_),
    .A1(net605),
    .A2(_09578_));
 sg13g2_xor2_1 _16408_ (.B(_09580_),
    .A(_00211_),
    .X(_09581_));
 sg13g2_buf_2 _16409_ (.A(net772),
    .X(_09582_));
 sg13g2_a22oi_1 _16410_ (.Y(_09583_),
    .B1(_09367_),
    .B2(\cpu.dcache.r_tag[5][11] ),
    .A2(_09296_),
    .A1(\cpu.dcache.r_tag[6][11] ));
 sg13g2_inv_1 _16411_ (.Y(_09584_),
    .A(_09583_));
 sg13g2_a22oi_1 _16412_ (.Y(_09585_),
    .B1(_09224_),
    .B2(\cpu.dcache.r_tag[2][11] ),
    .A2(_09219_),
    .A1(\cpu.dcache.r_tag[4][11] ));
 sg13g2_a22oi_1 _16413_ (.Y(_09586_),
    .B1(_09254_),
    .B2(\cpu.dcache.r_tag[3][11] ),
    .A2(net769),
    .A1(\cpu.dcache.r_tag[7][11] ));
 sg13g2_o21ai_1 _16414_ (.B1(_09586_),
    .Y(_09587_),
    .A1(net782),
    .A2(_09585_));
 sg13g2_a21oi_1 _16415_ (.A1(net885),
    .A2(_09584_),
    .Y(_09588_),
    .B1(_09587_));
 sg13g2_and2_1 _16416_ (.A(_00220_),
    .B(net758),
    .X(_09589_));
 sg13g2_a21oi_1 _16417_ (.A1(_09582_),
    .A2(_09588_),
    .Y(_09590_),
    .B1(_09589_));
 sg13g2_nand3b_1 _16418_ (.B(net605),
    .C(_09588_),
    .Y(_09591_),
    .A_N(\cpu.dcache.r_tag[1][11] ));
 sg13g2_o21ai_1 _16419_ (.B1(_09591_),
    .Y(_09592_),
    .A1(net605),
    .A2(_09590_));
 sg13g2_xnor2_1 _16420_ (.Y(_09593_),
    .A(_00219_),
    .B(_09592_));
 sg13g2_mux4_1 _16421_ (.S0(net756),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][8] ),
    .S1(net757),
    .X(_09594_));
 sg13g2_mux4_1 _16422_ (.S0(net756),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][8] ),
    .S1(net757),
    .X(_09595_));
 sg13g2_mux4_1 _16423_ (.S0(net760),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][8] ),
    .S1(net759),
    .X(_09596_));
 sg13g2_mux4_1 _16424_ (.S0(net760),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][8] ),
    .S1(net759),
    .X(_09597_));
 sg13g2_mux4_1 _16425_ (.S0(net889),
    .A0(_09594_),
    .A1(_09595_),
    .A2(_09596_),
    .A3(_09597_),
    .S1(net884),
    .X(_09598_));
 sg13g2_nand2_1 _16426_ (.Y(_09599_),
    .A(net776),
    .B(_09598_));
 sg13g2_mux4_1 _16427_ (.S0(net756),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][8] ),
    .S1(net757),
    .X(_09600_));
 sg13g2_mux4_1 _16428_ (.S0(net756),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][8] ),
    .S1(net757),
    .X(_09601_));
 sg13g2_mux4_1 _16429_ (.S0(net764),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][8] ),
    .S1(net765),
    .X(_09602_));
 sg13g2_mux4_1 _16430_ (.S0(net764),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][8] ),
    .S1(net765),
    .X(_09603_));
 sg13g2_mux4_1 _16431_ (.S0(net889),
    .A0(_09600_),
    .A1(_09601_),
    .A2(_09602_),
    .A3(_09603_),
    .S1(net888),
    .X(_09604_));
 sg13g2_nand2_1 _16432_ (.Y(_09605_),
    .A(net682),
    .B(_09604_));
 sg13g2_a21oi_2 _16433_ (.B1(_08380_),
    .Y(_09606_),
    .A2(_09605_),
    .A1(_09599_));
 sg13g2_buf_1 _16434_ (.A(_09606_),
    .X(_09607_));
 sg13g2_nand2_1 _16435_ (.Y(_09608_),
    .A(net898),
    .B(\cpu.dcache.r_tag[6][20] ));
 sg13g2_nand3b_1 _16436_ (.B(\cpu.dcache.r_tag[5][20] ),
    .C(net1036),
    .Y(_09609_),
    .A_N(net898));
 sg13g2_o21ai_1 _16437_ (.B1(_09609_),
    .Y(_09610_),
    .A1(net900),
    .A2(_09608_));
 sg13g2_inv_1 _16438_ (.Y(_09611_),
    .A(\cpu.dcache.r_tag[4][20] ));
 sg13g2_nand3_1 _16439_ (.B(net1108),
    .C(\cpu.dcache.r_tag[2][20] ),
    .A(_09101_),
    .Y(_09612_));
 sg13g2_o21ai_1 _16440_ (.B1(_09612_),
    .Y(_09613_),
    .A1(_09611_),
    .A2(_09335_));
 sg13g2_inv_1 _16441_ (.Y(_09614_),
    .A(\cpu.dcache.r_tag[7][20] ));
 sg13g2_nand3_1 _16442_ (.B(net1029),
    .C(net1032),
    .A(net1036),
    .Y(_09615_));
 sg13g2_buf_2 _16443_ (.A(_09615_),
    .X(_09616_));
 sg13g2_nand4_1 _16444_ (.B(_09101_),
    .C(_09209_),
    .A(_09034_),
    .Y(_09617_),
    .D(\cpu.dcache.r_tag[3][20] ));
 sg13g2_o21ai_1 _16445_ (.B1(_09617_),
    .Y(_09618_),
    .A1(_09614_),
    .A2(_09616_));
 sg13g2_a221oi_1 _16446_ (.B2(_09217_),
    .C1(_09618_),
    .B1(_09613_),
    .A1(net885),
    .Y(_09619_),
    .A2(_09610_));
 sg13g2_nor2_1 _16447_ (.A(\cpu.dcache.r_tag[0][20] ),
    .B(_09230_),
    .Y(_09620_));
 sg13g2_a21o_1 _16448_ (.A2(_09619_),
    .A1(_09230_),
    .B1(_09620_),
    .X(_09621_));
 sg13g2_nor2_1 _16449_ (.A(\cpu.dcache.r_tag[1][20] ),
    .B(_09212_),
    .Y(_09622_));
 sg13g2_a22oi_1 _16450_ (.Y(_09623_),
    .B1(_09622_),
    .B2(_09619_),
    .A2(_09621_),
    .A1(_09330_));
 sg13g2_xor2_1 _16451_ (.B(_09623_),
    .A(net425),
    .X(_09624_));
 sg13g2_mux4_1 _16452_ (.S0(_09476_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][7] ),
    .S1(net761),
    .X(_09625_));
 sg13g2_mux4_1 _16453_ (.S0(net762),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][7] ),
    .S1(net761),
    .X(_09626_));
 sg13g2_mux4_1 _16454_ (.S0(net756),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][7] ),
    .S1(net757),
    .X(_09627_));
 sg13g2_mux4_1 _16455_ (.S0(_09476_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][7] ),
    .S1(_09474_),
    .X(_09628_));
 sg13g2_mux4_1 _16456_ (.S0(net886),
    .A0(_09625_),
    .A1(_09626_),
    .A2(_09627_),
    .A3(_09628_),
    .S1(net884),
    .X(_09629_));
 sg13g2_nand2_1 _16457_ (.Y(_09630_),
    .A(net776),
    .B(_09629_));
 sg13g2_mux4_1 _16458_ (.S0(net756),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][7] ),
    .S1(net757),
    .X(_09631_));
 sg13g2_mux4_1 _16459_ (.S0(net756),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][7] ),
    .S1(net757),
    .X(_09632_));
 sg13g2_mux4_1 _16460_ (.S0(net760),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][7] ),
    .S1(net759),
    .X(_09633_));
 sg13g2_mux4_1 _16461_ (.S0(net760),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][7] ),
    .S1(net759),
    .X(_09634_));
 sg13g2_mux4_1 _16462_ (.S0(net889),
    .A0(_09631_),
    .A1(_09632_),
    .A2(_09633_),
    .A3(_09634_),
    .S1(net884),
    .X(_09635_));
 sg13g2_nand2_1 _16463_ (.Y(_09636_),
    .A(net682),
    .B(_09635_));
 sg13g2_a21oi_2 _16464_ (.B1(net1049),
    .Y(_09637_),
    .A2(_09636_),
    .A1(_09630_));
 sg13g2_buf_1 _16465_ (.A(_09637_),
    .X(_09638_));
 sg13g2_nor2_1 _16466_ (.A(_00228_),
    .B(_09464_),
    .Y(_09639_));
 sg13g2_a221oi_1 _16467_ (.B2(\cpu.dcache.r_tag[6][19] ),
    .C1(_09639_),
    .B1(net677),
    .A1(\cpu.dcache.r_tag[3][19] ),
    .Y(_09640_),
    .A2(_09254_));
 sg13g2_a22oi_1 _16468_ (.Y(_09641_),
    .B1(net602),
    .B2(\cpu.dcache.r_tag[2][19] ),
    .A2(net605),
    .A1(\cpu.dcache.r_tag[1][19] ));
 sg13g2_mux2_1 _16469_ (.A0(\cpu.dcache.r_tag[5][19] ),
    .A1(\cpu.dcache.r_tag[7][19] ),
    .S(_09102_),
    .X(_09642_));
 sg13g2_a22oi_1 _16470_ (.Y(_09643_),
    .B1(_09642_),
    .B2(net686),
    .A2(_09426_),
    .A1(\cpu.dcache.r_tag[4][19] ));
 sg13g2_nand2b_1 _16471_ (.Y(_09644_),
    .B(_09382_),
    .A_N(_09643_));
 sg13g2_and3_1 _16472_ (.X(_09645_),
    .A(_09640_),
    .B(_09641_),
    .C(_09644_));
 sg13g2_xnor2_1 _16473_ (.Y(_09646_),
    .A(_09638_),
    .B(_09645_));
 sg13g2_nor2_1 _16474_ (.A(_09624_),
    .B(_09646_),
    .Y(_09647_));
 sg13g2_nand4_1 _16475_ (.B(_09581_),
    .C(_09593_),
    .A(_09570_),
    .Y(_09648_),
    .D(_09647_));
 sg13g2_nor4_1 _16476_ (.A(_09182_),
    .B(_09458_),
    .C(_09511_),
    .D(_09648_),
    .Y(_09649_));
 sg13g2_inv_1 _16477_ (.Y(_09650_),
    .A(_09175_));
 sg13g2_nor4_1 _16478_ (.A(_09650_),
    .B(_09458_),
    .C(_09511_),
    .D(_09648_),
    .Y(_09651_));
 sg13g2_or3_1 _16479_ (.A(_09182_),
    .B(_09180_),
    .C(_09651_),
    .X(_09652_));
 sg13g2_buf_1 _16480_ (.A(_09652_),
    .X(_09653_));
 sg13g2_o21ai_1 _16481_ (.B1(_09653_),
    .Y(_09654_),
    .A1(_09181_),
    .A2(_09649_));
 sg13g2_and2_1 _16482_ (.A(_09168_),
    .B(_09654_),
    .X(_09655_));
 sg13g2_nand2b_1 _16483_ (.Y(_09656_),
    .B(_08180_),
    .A_N(_09022_));
 sg13g2_a22oi_1 _16484_ (.Y(_09657_),
    .B1(_09655_),
    .B2(_09656_),
    .A2(_08923_),
    .A1(net1030));
 sg13g2_nand2_1 _16485_ (.Y(_09658_),
    .A(_09163_),
    .B(_09657_));
 sg13g2_buf_1 _16486_ (.A(\cpu.qspi.r_state[7] ),
    .X(_09659_));
 sg13g2_buf_2 _16487_ (.A(\cpu.qspi.r_ind ),
    .X(_09660_));
 sg13g2_buf_1 _16488_ (.A(_00230_),
    .X(_09661_));
 sg13g2_buf_1 _16489_ (.A(\cpu.qspi.r_count[0] ),
    .X(_09662_));
 sg13g2_buf_2 _16490_ (.A(\cpu.qspi.r_count[1] ),
    .X(_09663_));
 sg13g2_buf_1 _16491_ (.A(\cpu.qspi.r_count[2] ),
    .X(_09664_));
 sg13g2_nor3_1 _16492_ (.A(_09662_),
    .B(_09663_),
    .C(_09664_),
    .Y(_09665_));
 sg13g2_nor2b_1 _16493_ (.A(\cpu.qspi.r_count[3] ),
    .B_N(_09665_),
    .Y(_09666_));
 sg13g2_buf_1 _16494_ (.A(_09666_),
    .X(_09667_));
 sg13g2_and2_1 _16495_ (.A(_09661_),
    .B(_09667_),
    .X(_09668_));
 sg13g2_buf_1 _16496_ (.A(_09668_),
    .X(_09669_));
 sg13g2_buf_1 _16497_ (.A(\cpu.qspi.r_state[2] ),
    .X(_09670_));
 sg13g2_buf_1 _16498_ (.A(\cpu.qspi.r_state[1] ),
    .X(_09671_));
 sg13g2_a221oi_1 _16499_ (.B2(_09670_),
    .C1(_09671_),
    .B1(_09669_),
    .A1(_09659_),
    .Y(_09672_),
    .A2(_09660_));
 sg13g2_a21oi_1 _16500_ (.A1(_09658_),
    .A2(_09672_),
    .Y(_00026_),
    .B1(net606));
 sg13g2_buf_1 _16501_ (.A(\cpu.qspi.r_state[16] ),
    .X(_09673_));
 sg13g2_nand2_1 _16502_ (.Y(_09674_),
    .A(_09661_),
    .B(_09667_));
 sg13g2_buf_1 _16503_ (.A(_09674_),
    .X(_09675_));
 sg13g2_nor3_1 _16504_ (.A(net1030),
    .B(_09181_),
    .C(_09649_),
    .Y(_09676_));
 sg13g2_buf_2 _16505_ (.A(_09676_),
    .X(_09677_));
 sg13g2_buf_2 _16506_ (.A(\cpu.qspi.r_state[8] ),
    .X(_09678_));
 sg13g2_a22oi_1 _16507_ (.Y(_09679_),
    .B1(_09677_),
    .B2(_09678_),
    .A2(net600),
    .A1(_09673_));
 sg13g2_nor2_1 _16508_ (.A(net607),
    .B(_09679_),
    .Y(_00025_));
 sg13g2_buf_1 _16509_ (.A(\cpu.qspi.r_state[4] ),
    .X(_09680_));
 sg13g2_buf_1 _16510_ (.A(\cpu.qspi.r_state[9] ),
    .X(_09681_));
 sg13g2_a21oi_1 _16511_ (.A1(_09680_),
    .A2(_09669_),
    .Y(_09682_),
    .B1(_09681_));
 sg13g2_nor2_1 _16512_ (.A(net607),
    .B(_09682_),
    .Y(_00022_));
 sg13g2_buf_1 _16513_ (.A(\cpu.qspi.r_rom_mode[1] ),
    .X(_09683_));
 sg13g2_buf_1 _16514_ (.A(\cpu.qspi.r_rom_mode[0] ),
    .X(_09684_));
 sg13g2_inv_1 _16515_ (.Y(_09685_),
    .A(_08133_));
 sg13g2_buf_1 _16516_ (.A(_09685_),
    .X(_09686_));
 sg13g2_buf_1 _16517_ (.A(_09417_),
    .X(_09687_));
 sg13g2_nor2_1 _16518_ (.A(net882),
    .B(_08535_),
    .Y(_09688_));
 sg13g2_a21oi_1 _16519_ (.A1(net882),
    .A2(net375),
    .Y(_09689_),
    .B1(_09688_));
 sg13g2_nor2b_1 _16520_ (.A(_09684_),
    .B_N(_09689_),
    .Y(_09690_));
 sg13g2_a21oi_1 _16521_ (.A1(_09684_),
    .A2(_09677_),
    .Y(_09691_),
    .B1(_09690_));
 sg13g2_and2_1 _16522_ (.A(_09683_),
    .B(_09691_),
    .X(_09692_));
 sg13g2_buf_2 _16523_ (.A(_09692_),
    .X(_09693_));
 sg13g2_nor3_1 _16524_ (.A(_09684_),
    .B(_09683_),
    .C(_09689_),
    .Y(_09694_));
 sg13g2_buf_2 _16525_ (.A(_09694_),
    .X(_09695_));
 sg13g2_nor2_1 _16526_ (.A(_09695_),
    .B(_09693_),
    .Y(_09696_));
 sg13g2_buf_2 _16527_ (.A(_09696_),
    .X(_09697_));
 sg13g2_and2_1 _16528_ (.A(\cpu.qspi.r_quad[2] ),
    .B(_09695_),
    .X(_09698_));
 sg13g2_a221oi_1 _16529_ (.B2(\cpu.qspi.r_quad[0] ),
    .C1(_09698_),
    .B1(_09697_),
    .A1(\cpu.qspi.r_quad[1] ),
    .Y(_09699_),
    .A2(_09693_));
 sg13g2_buf_2 _16530_ (.A(_09699_),
    .X(_09700_));
 sg13g2_inv_1 _16531_ (.Y(_09701_),
    .A(_09700_));
 sg13g2_nand3b_1 _16532_ (.B(_08964_),
    .C(_09163_),
    .Y(_09702_),
    .A_N(_09657_));
 sg13g2_nand3_1 _16533_ (.B(_08964_),
    .C(net600),
    .A(_09680_),
    .Y(_09703_));
 sg13g2_o21ai_1 _16534_ (.B1(_09703_),
    .Y(_00028_),
    .A1(_09701_),
    .A2(_09702_));
 sg13g2_nand2_1 _16535_ (.Y(_09704_),
    .A(_09670_),
    .B(_09675_));
 sg13g2_buf_2 _16536_ (.A(\cpu.qspi.r_state[14] ),
    .X(_09705_));
 sg13g2_nand2_1 _16537_ (.Y(_09706_),
    .A(_09705_),
    .B(_09669_));
 sg13g2_a21oi_1 _16538_ (.A1(_09704_),
    .A2(_09706_),
    .Y(_00027_),
    .B1(net606));
 sg13g2_inv_1 _16539_ (.Y(_09707_),
    .A(_09660_));
 sg13g2_a21o_1 _16540_ (.A2(_09707_),
    .A1(_09659_),
    .B1(net684),
    .X(_00021_));
 sg13g2_buf_2 _16541_ (.A(\cpu.dec.r_op[1] ),
    .X(_09708_));
 sg13g2_inv_1 _16542_ (.Y(_09709_),
    .A(_09708_));
 sg13g2_buf_1 _16543_ (.A(_08842_),
    .X(_09710_));
 sg13g2_nand3_1 _16544_ (.B(net231),
    .C(_08930_),
    .A(net121),
    .Y(_09711_));
 sg13g2_o21ai_1 _16545_ (.B1(_09711_),
    .Y(_00012_),
    .A1(_09709_),
    .A2(_08926_));
 sg13g2_buf_2 _16546_ (.A(\cpu.dec.r_op[10] ),
    .X(_09712_));
 sg13g2_inv_1 _16547_ (.Y(_09713_),
    .A(_09712_));
 sg13g2_nor2_1 _16548_ (.A(_08860_),
    .B(_08877_),
    .Y(_09714_));
 sg13g2_nand3_1 _16549_ (.B(_08948_),
    .C(_09714_),
    .A(net121),
    .Y(_09715_));
 sg13g2_o21ai_1 _16550_ (.B1(_09715_),
    .Y(_00011_),
    .A1(_09713_),
    .A2(net105));
 sg13g2_nand3_1 _16551_ (.B(net231),
    .C(_08955_),
    .A(_08948_),
    .Y(_09716_));
 sg13g2_o21ai_1 _16552_ (.B1(_09716_),
    .Y(_09717_),
    .A1(_08908_),
    .A2(_08954_));
 sg13g2_buf_2 _16553_ (.A(\cpu.dec.r_op[9] ),
    .X(_09718_));
 sg13g2_buf_1 _16554_ (.A(_09718_),
    .X(_09719_));
 sg13g2_mux2_1 _16555_ (.A0(_09717_),
    .A1(net1027),
    .S(net149),
    .X(_00020_));
 sg13g2_buf_1 _16556_ (.A(_00257_),
    .X(_09720_));
 sg13g2_buf_1 _16557_ (.A(\cpu.qspi.r_state[12] ),
    .X(_09721_));
 sg13g2_nand2_1 _16558_ (.Y(_09722_),
    .A(_09721_),
    .B(net600));
 sg13g2_a21oi_1 _16559_ (.A1(_09720_),
    .A2(_09722_),
    .Y(_00023_),
    .B1(net606));
 sg13g2_buf_1 _16560_ (.A(\cpu.qspi.r_state[5] ),
    .X(_09723_));
 sg13g2_inv_1 _16561_ (.Y(_09724_),
    .A(_09723_));
 sg13g2_nand2_1 _16562_ (.Y(_09725_),
    .A(_09705_),
    .B(net600));
 sg13g2_a21oi_1 _16563_ (.A1(_09724_),
    .A2(_09725_),
    .Y(_00024_),
    .B1(_09137_));
 sg13g2_buf_1 _16564_ (.A(_08721_),
    .X(_09726_));
 sg13g2_nand2_2 _16565_ (.Y(_09727_),
    .A(net209),
    .B(net185));
 sg13g2_nand2_1 _16566_ (.Y(_09728_),
    .A(_08783_),
    .B(_08804_));
 sg13g2_buf_2 _16567_ (.A(_09728_),
    .X(_09729_));
 sg13g2_nor2_1 _16568_ (.A(_09727_),
    .B(_09729_),
    .Y(_09730_));
 sg13g2_buf_2 _16569_ (.A(\cpu.dec.r_op[8] ),
    .X(_09731_));
 sg13g2_buf_1 _16570_ (.A(_09731_),
    .X(_09732_));
 sg13g2_mux2_1 _16571_ (.A0(_09730_),
    .A1(net1026),
    .S(net149),
    .X(_00019_));
 sg13g2_nor3_1 _16572_ (.A(\cpu.uart.r_div[0] ),
    .B(\cpu.uart.r_div[1] ),
    .C(\cpu.uart.r_div[2] ),
    .Y(_09733_));
 sg13g2_nor2b_1 _16573_ (.A(\cpu.uart.r_div[3] ),
    .B_N(_09733_),
    .Y(_09734_));
 sg13g2_nor2b_1 _16574_ (.A(\cpu.uart.r_div[4] ),
    .B_N(_09734_),
    .Y(_09735_));
 sg13g2_nor2b_1 _16575_ (.A(\cpu.uart.r_div[5] ),
    .B_N(_09735_),
    .Y(_09736_));
 sg13g2_nor2b_1 _16576_ (.A(\cpu.uart.r_div[6] ),
    .B_N(_09736_),
    .Y(_09737_));
 sg13g2_nand2b_1 _16577_ (.Y(_09738_),
    .B(_09737_),
    .A_N(\cpu.uart.r_div[7] ));
 sg13g2_nor2_1 _16578_ (.A(\cpu.uart.r_div[8] ),
    .B(_09738_),
    .Y(_09739_));
 sg13g2_nand2b_1 _16579_ (.Y(_09740_),
    .B(_09739_),
    .A_N(\cpu.uart.r_div[9] ));
 sg13g2_buf_1 _16580_ (.A(_09740_),
    .X(_09741_));
 sg13g2_nor3_1 _16581_ (.A(\cpu.uart.r_div[11] ),
    .B(\cpu.uart.r_div[10] ),
    .C(_09741_),
    .Y(_09742_));
 sg13g2_buf_1 _16582_ (.A(_09742_),
    .X(_09743_));
 sg13g2_buf_1 _16583_ (.A(_09743_),
    .X(_09744_));
 sg13g2_nor2_1 _16584_ (.A(net897),
    .B(_09744_),
    .Y(_09745_));
 sg13g2_buf_1 _16585_ (.A(_09745_),
    .X(_09746_));
 sg13g2_buf_1 _16586_ (.A(net208),
    .X(_09747_));
 sg13g2_mux2_1 _16587_ (.A0(\cpu.uart.r_div_value[0] ),
    .A1(_00258_),
    .S(net184),
    .X(_00079_));
 sg13g2_xnor2_1 _16588_ (.Y(_09748_),
    .A(\cpu.uart.r_div[0] ),
    .B(\cpu.uart.r_div[1] ));
 sg13g2_mux2_1 _16589_ (.A0(\cpu.uart.r_div_value[1] ),
    .A1(_09748_),
    .S(net184),
    .X(_00082_));
 sg13g2_o21ai_1 _16590_ (.B1(\cpu.uart.r_div[2] ),
    .Y(_09749_),
    .A1(\cpu.uart.r_div[0] ),
    .A2(\cpu.uart.r_div[1] ));
 sg13g2_nor2b_1 _16591_ (.A(_09733_),
    .B_N(_09749_),
    .Y(_09750_));
 sg13g2_nor2_1 _16592_ (.A(\cpu.uart.r_div_value[2] ),
    .B(net208),
    .Y(_09751_));
 sg13g2_a21oi_1 _16593_ (.A1(_09747_),
    .A2(_09750_),
    .Y(_00083_),
    .B1(_09751_));
 sg13g2_xnor2_1 _16594_ (.Y(_09752_),
    .A(\cpu.uart.r_div[3] ),
    .B(_09733_));
 sg13g2_nor2_1 _16595_ (.A(\cpu.uart.r_div_value[3] ),
    .B(net208),
    .Y(_09753_));
 sg13g2_a21oi_1 _16596_ (.A1(_09747_),
    .A2(_09752_),
    .Y(_00084_),
    .B1(_09753_));
 sg13g2_xnor2_1 _16597_ (.Y(_09754_),
    .A(\cpu.uart.r_div[4] ),
    .B(_09734_));
 sg13g2_nor2_1 _16598_ (.A(\cpu.uart.r_div_value[4] ),
    .B(net208),
    .Y(_09755_));
 sg13g2_a21oi_1 _16599_ (.A1(net184),
    .A2(_09754_),
    .Y(_00085_),
    .B1(_09755_));
 sg13g2_xnor2_1 _16600_ (.Y(_09756_),
    .A(\cpu.uart.r_div[5] ),
    .B(_09735_));
 sg13g2_nor2_1 _16601_ (.A(\cpu.uart.r_div_value[5] ),
    .B(net208),
    .Y(_09757_));
 sg13g2_a21oi_1 _16602_ (.A1(net184),
    .A2(_09756_),
    .Y(_00086_),
    .B1(_09757_));
 sg13g2_xnor2_1 _16603_ (.Y(_09758_),
    .A(\cpu.uart.r_div[6] ),
    .B(_09736_));
 sg13g2_nor2_1 _16604_ (.A(\cpu.uart.r_div_value[6] ),
    .B(net208),
    .Y(_09759_));
 sg13g2_a21oi_1 _16605_ (.A1(net184),
    .A2(_09758_),
    .Y(_00087_),
    .B1(_09759_));
 sg13g2_xnor2_1 _16606_ (.Y(_09760_),
    .A(\cpu.uart.r_div[7] ),
    .B(_09737_));
 sg13g2_nor2_1 _16607_ (.A(\cpu.uart.r_div_value[7] ),
    .B(_09746_),
    .Y(_09761_));
 sg13g2_a21oi_1 _16608_ (.A1(net184),
    .A2(_09760_),
    .Y(_00088_),
    .B1(_09761_));
 sg13g2_xor2_1 _16609_ (.B(_09738_),
    .A(\cpu.uart.r_div[8] ),
    .X(_09762_));
 sg13g2_nor2_1 _16610_ (.A(\cpu.uart.r_div_value[8] ),
    .B(net208),
    .Y(_09763_));
 sg13g2_a21oi_1 _16611_ (.A1(net184),
    .A2(_09762_),
    .Y(_00089_),
    .B1(_09763_));
 sg13g2_xnor2_1 _16612_ (.Y(_09764_),
    .A(\cpu.uart.r_div[9] ),
    .B(_09739_));
 sg13g2_nor2_1 _16613_ (.A(\cpu.uart.r_div_value[9] ),
    .B(net208),
    .Y(_09765_));
 sg13g2_a21oi_1 _16614_ (.A1(net184),
    .A2(_09764_),
    .Y(_00090_),
    .B1(_09765_));
 sg13g2_buf_1 _16615_ (.A(\cpu.uart.r_div_value[10] ),
    .X(_09766_));
 sg13g2_inv_1 _16616_ (.Y(_09767_),
    .A(_09766_));
 sg13g2_nand2_1 _16617_ (.Y(_09768_),
    .A(net901),
    .B(_09741_));
 sg13g2_o21ai_1 _16618_ (.B1(_09768_),
    .Y(_09769_),
    .A1(\cpu.uart.r_div[11] ),
    .A2(_09766_));
 sg13g2_inv_1 _16619_ (.Y(_09770_),
    .A(\cpu.uart.r_div[10] ));
 sg13g2_nor3_1 _16620_ (.A(_09770_),
    .B(net778),
    .C(_09741_),
    .Y(_09771_));
 sg13g2_a221oi_1 _16621_ (.B2(_09770_),
    .C1(_09771_),
    .B1(_09769_),
    .A1(_09767_),
    .Y(_00080_),
    .A2(net684));
 sg13g2_nor2_1 _16622_ (.A(\cpu.uart.r_div[10] ),
    .B(_09741_),
    .Y(_09772_));
 sg13g2_nand2_1 _16623_ (.Y(_09773_),
    .A(\cpu.uart.r_div[11] ),
    .B(net783));
 sg13g2_o21ai_1 _16624_ (.B1(\cpu.uart.r_div_value[11] ),
    .Y(_09774_),
    .A1(net778),
    .A2(net252));
 sg13g2_o21ai_1 _16625_ (.B1(_09774_),
    .Y(_00081_),
    .A1(_09772_),
    .A2(_09773_));
 sg13g2_buf_1 _16626_ (.A(_09038_),
    .X(_09775_));
 sg13g2_buf_1 _16627_ (.A(net1025),
    .X(_09776_));
 sg13g2_buf_1 _16628_ (.A(net881),
    .X(_09777_));
 sg13g2_buf_1 _16629_ (.A(_09265_),
    .X(_09778_));
 sg13g2_buf_1 _16630_ (.A(net675),
    .X(_09779_));
 sg13g2_buf_1 _16631_ (.A(net599),
    .X(_09780_));
 sg13g2_buf_2 _16632_ (.A(\cpu.addr[5] ),
    .X(_09781_));
 sg13g2_nor3_2 _16633_ (.A(_09781_),
    .B(net1037),
    .C(_09026_),
    .Y(_09782_));
 sg13g2_nand2_1 _16634_ (.Y(_09783_),
    .A(_09023_),
    .B(_09782_));
 sg13g2_buf_1 _16635_ (.A(_09783_),
    .X(_09784_));
 sg13g2_nor2_1 _16636_ (.A(_09046_),
    .B(net674),
    .Y(_09785_));
 sg13g2_buf_2 _16637_ (.A(_09785_),
    .X(_09786_));
 sg13g2_nand3_1 _16638_ (.B(net530),
    .C(_09786_),
    .A(net755),
    .Y(_09787_));
 sg13g2_buf_1 _16639_ (.A(_09787_),
    .X(_09788_));
 sg13g2_buf_1 _16640_ (.A(\cpu.intr.r_timer_count[19] ),
    .X(_09789_));
 sg13g2_buf_1 _16641_ (.A(\cpu.intr.r_timer_count[18] ),
    .X(_09790_));
 sg13g2_buf_1 _16642_ (.A(\cpu.intr.r_timer_count[17] ),
    .X(_09791_));
 sg13g2_buf_1 _16643_ (.A(\cpu.intr.r_timer_count[16] ),
    .X(_09792_));
 sg13g2_buf_1 _16644_ (.A(\cpu.intr.r_timer_count[11] ),
    .X(_09793_));
 sg13g2_buf_1 _16645_ (.A(\cpu.intr.r_timer_count[10] ),
    .X(_09794_));
 sg13g2_buf_1 _16646_ (.A(\cpu.intr.r_timer_count[7] ),
    .X(_09795_));
 sg13g2_buf_1 _16647_ (.A(\cpu.intr.r_timer_count[1] ),
    .X(_09796_));
 sg13g2_nor3_1 _16648_ (.A(_09796_),
    .B(\cpu.intr.r_timer_count[0] ),
    .C(\cpu.intr.r_timer_count[2] ),
    .Y(_09797_));
 sg13g2_nor2b_1 _16649_ (.A(\cpu.intr.r_timer_count[3] ),
    .B_N(_09797_),
    .Y(_09798_));
 sg13g2_nor2b_1 _16650_ (.A(\cpu.intr.r_timer_count[4] ),
    .B_N(_09798_),
    .Y(_09799_));
 sg13g2_nor2b_1 _16651_ (.A(\cpu.intr.r_timer_count[5] ),
    .B_N(_09799_),
    .Y(_09800_));
 sg13g2_nand2b_1 _16652_ (.Y(_09801_),
    .B(_09800_),
    .A_N(\cpu.intr.r_timer_count[6] ));
 sg13g2_nor3_1 _16653_ (.A(_09795_),
    .B(\cpu.intr.r_timer_count[8] ),
    .C(_09801_),
    .Y(_09802_));
 sg13g2_nand2b_1 _16654_ (.Y(_09803_),
    .B(_09802_),
    .A_N(\cpu.intr.r_timer_count[9] ));
 sg13g2_buf_1 _16655_ (.A(_09803_),
    .X(_09804_));
 sg13g2_nor4_1 _16656_ (.A(_09793_),
    .B(_09794_),
    .C(\cpu.intr.r_timer_count[12] ),
    .D(_09804_),
    .Y(_09805_));
 sg13g2_nor2b_1 _16657_ (.A(\cpu.intr.r_timer_count[13] ),
    .B_N(_09805_),
    .Y(_09806_));
 sg13g2_nor2b_1 _16658_ (.A(\cpu.intr.r_timer_count[14] ),
    .B_N(_09806_),
    .Y(_09807_));
 sg13g2_nand2b_2 _16659_ (.Y(_09808_),
    .B(_09807_),
    .A_N(\cpu.intr.r_timer_count[15] ));
 sg13g2_nor3_2 _16660_ (.A(_09791_),
    .B(_09792_),
    .C(_09808_),
    .Y(_09809_));
 sg13g2_nor2b_1 _16661_ (.A(_09790_),
    .B_N(_09809_),
    .Y(_09810_));
 sg13g2_nand2b_1 _16662_ (.Y(_09811_),
    .B(_09810_),
    .A_N(_09789_));
 sg13g2_buf_1 _16663_ (.A(_09811_),
    .X(_09812_));
 sg13g2_buf_1 _16664_ (.A(\cpu.intr.r_timer_count[21] ),
    .X(_09813_));
 sg13g2_buf_2 _16665_ (.A(\cpu.intr.r_timer_count[20] ),
    .X(_09814_));
 sg13g2_buf_1 _16666_ (.A(\cpu.intr.r_timer_count[23] ),
    .X(_09815_));
 sg13g2_buf_1 _16667_ (.A(\cpu.intr.r_timer_count[22] ),
    .X(_09816_));
 sg13g2_nor4_2 _16668_ (.A(_09813_),
    .B(_09814_),
    .C(_09815_),
    .Y(_09817_),
    .D(_09816_));
 sg13g2_nand2b_1 _16669_ (.Y(_09818_),
    .B(_09817_),
    .A_N(_09812_));
 sg13g2_buf_2 _16670_ (.A(_09818_),
    .X(_09819_));
 sg13g2_nand2_1 _16671_ (.Y(_09820_),
    .A(_09788_),
    .B(_09819_));
 sg13g2_buf_2 _16672_ (.A(_09820_),
    .X(_09821_));
 sg13g2_buf_8 _16673_ (.A(_09821_),
    .X(_09822_));
 sg13g2_mux2_1 _16674_ (.A0(_00264_),
    .A1(\cpu.intr.r_timer_reload[0] ),
    .S(net65),
    .X(_00055_));
 sg13g2_buf_8 _16675_ (.A(_09821_),
    .X(_09823_));
 sg13g2_xor2_1 _16676_ (.B(\cpu.intr.r_timer_count[0] ),
    .A(_09796_),
    .X(_09824_));
 sg13g2_nand2_1 _16677_ (.Y(_09825_),
    .A(\cpu.intr.r_timer_reload[1] ),
    .B(net65));
 sg13g2_o21ai_1 _16678_ (.B1(_09825_),
    .Y(_00066_),
    .A1(net64),
    .A2(_09824_));
 sg13g2_o21ai_1 _16679_ (.B1(\cpu.intr.r_timer_count[2] ),
    .Y(_09826_),
    .A1(_09796_),
    .A2(\cpu.intr.r_timer_count[0] ));
 sg13g2_nor2b_1 _16680_ (.A(_09797_),
    .B_N(_09826_),
    .Y(_09827_));
 sg13g2_nand2_1 _16681_ (.Y(_09828_),
    .A(\cpu.intr.r_timer_reload[2] ),
    .B(net65));
 sg13g2_o21ai_1 _16682_ (.B1(_09828_),
    .Y(_00071_),
    .A1(net64),
    .A2(_09827_));
 sg13g2_xnor2_1 _16683_ (.Y(_09829_),
    .A(\cpu.intr.r_timer_count[3] ),
    .B(_09797_));
 sg13g2_nand2_1 _16684_ (.Y(_09830_),
    .A(\cpu.intr.r_timer_reload[3] ),
    .B(_09822_));
 sg13g2_o21ai_1 _16685_ (.B1(_09830_),
    .Y(_00072_),
    .A1(_09823_),
    .A2(_09829_));
 sg13g2_xnor2_1 _16686_ (.Y(_09831_),
    .A(\cpu.intr.r_timer_count[4] ),
    .B(_09798_));
 sg13g2_nand2_1 _16687_ (.Y(_09832_),
    .A(\cpu.intr.r_timer_reload[4] ),
    .B(_09822_));
 sg13g2_o21ai_1 _16688_ (.B1(_09832_),
    .Y(_00073_),
    .A1(net64),
    .A2(_09831_));
 sg13g2_xnor2_1 _16689_ (.Y(_09833_),
    .A(\cpu.intr.r_timer_count[5] ),
    .B(_09799_));
 sg13g2_buf_8 _16690_ (.A(_09821_),
    .X(_09834_));
 sg13g2_nand2_1 _16691_ (.Y(_09835_),
    .A(\cpu.intr.r_timer_reload[5] ),
    .B(net63));
 sg13g2_o21ai_1 _16692_ (.B1(_09835_),
    .Y(_00074_),
    .A1(_09823_),
    .A2(_09833_));
 sg13g2_xnor2_1 _16693_ (.Y(_09836_),
    .A(\cpu.intr.r_timer_count[6] ),
    .B(_09800_));
 sg13g2_nand2_1 _16694_ (.Y(_09837_),
    .A(\cpu.intr.r_timer_reload[6] ),
    .B(net63));
 sg13g2_o21ai_1 _16695_ (.B1(_09837_),
    .Y(_00075_),
    .A1(net64),
    .A2(_09836_));
 sg13g2_xor2_1 _16696_ (.B(_09801_),
    .A(_09795_),
    .X(_09838_));
 sg13g2_nand2_1 _16697_ (.Y(_09839_),
    .A(\cpu.intr.r_timer_reload[7] ),
    .B(net63));
 sg13g2_o21ai_1 _16698_ (.B1(_09839_),
    .Y(_00076_),
    .A1(net64),
    .A2(_09838_));
 sg13g2_nor2_1 _16699_ (.A(_09795_),
    .B(_09801_),
    .Y(_09840_));
 sg13g2_xnor2_1 _16700_ (.Y(_09841_),
    .A(\cpu.intr.r_timer_count[8] ),
    .B(_09840_));
 sg13g2_nand2_1 _16701_ (.Y(_09842_),
    .A(\cpu.intr.r_timer_reload[8] ),
    .B(net63));
 sg13g2_o21ai_1 _16702_ (.B1(_09842_),
    .Y(_00077_),
    .A1(net64),
    .A2(_09841_));
 sg13g2_xnor2_1 _16703_ (.Y(_09843_),
    .A(\cpu.intr.r_timer_count[9] ),
    .B(_09802_));
 sg13g2_nand2_1 _16704_ (.Y(_09844_),
    .A(\cpu.intr.r_timer_reload[9] ),
    .B(net63));
 sg13g2_o21ai_1 _16705_ (.B1(_09844_),
    .Y(_00078_),
    .A1(net64),
    .A2(_09843_));
 sg13g2_xor2_1 _16706_ (.B(_09804_),
    .A(_09794_),
    .X(_09845_));
 sg13g2_nand2_1 _16707_ (.Y(_09846_),
    .A(\cpu.intr.r_timer_reload[10] ),
    .B(net63));
 sg13g2_o21ai_1 _16708_ (.B1(_09846_),
    .Y(_00056_),
    .A1(net64),
    .A2(_09845_));
 sg13g2_nor3_1 _16709_ (.A(_09793_),
    .B(_09794_),
    .C(_09804_),
    .Y(_09847_));
 sg13g2_o21ai_1 _16710_ (.B1(_09793_),
    .Y(_09848_),
    .A1(_09794_),
    .A2(_09804_));
 sg13g2_nor2b_1 _16711_ (.A(_09847_),
    .B_N(_09848_),
    .Y(_09849_));
 sg13g2_nand2_1 _16712_ (.Y(_09850_),
    .A(\cpu.intr.r_timer_reload[11] ),
    .B(_09834_));
 sg13g2_o21ai_1 _16713_ (.B1(_09850_),
    .Y(_00057_),
    .A1(net65),
    .A2(_09849_));
 sg13g2_xnor2_1 _16714_ (.Y(_09851_),
    .A(\cpu.intr.r_timer_count[12] ),
    .B(_09847_));
 sg13g2_nand2_1 _16715_ (.Y(_09852_),
    .A(\cpu.intr.r_timer_reload[12] ),
    .B(net63));
 sg13g2_o21ai_1 _16716_ (.B1(_09852_),
    .Y(_00058_),
    .A1(net65),
    .A2(_09851_));
 sg13g2_xnor2_1 _16717_ (.Y(_09853_),
    .A(\cpu.intr.r_timer_count[13] ),
    .B(_09805_));
 sg13g2_nand2_1 _16718_ (.Y(_09854_),
    .A(\cpu.intr.r_timer_reload[13] ),
    .B(_09834_));
 sg13g2_o21ai_1 _16719_ (.B1(_09854_),
    .Y(_00059_),
    .A1(net65),
    .A2(_09853_));
 sg13g2_xnor2_1 _16720_ (.Y(_09855_),
    .A(\cpu.intr.r_timer_count[14] ),
    .B(_09806_));
 sg13g2_nand2_1 _16721_ (.Y(_09856_),
    .A(\cpu.intr.r_timer_reload[14] ),
    .B(net63));
 sg13g2_o21ai_1 _16722_ (.B1(_09856_),
    .Y(_00060_),
    .A1(net65),
    .A2(_09855_));
 sg13g2_xnor2_1 _16723_ (.Y(_09857_),
    .A(\cpu.intr.r_timer_count[15] ),
    .B(_09807_));
 sg13g2_nand2_1 _16724_ (.Y(_09858_),
    .A(\cpu.intr.r_timer_reload[15] ),
    .B(_09821_));
 sg13g2_o21ai_1 _16725_ (.B1(_09858_),
    .Y(_00061_),
    .A1(net65),
    .A2(_09857_));
 sg13g2_buf_1 _16726_ (.A(\cpu.dcache.wdata[0] ),
    .X(_09859_));
 sg13g2_buf_1 _16727_ (.A(_09859_),
    .X(_09860_));
 sg13g2_buf_1 _16728_ (.A(net1024),
    .X(_09861_));
 sg13g2_nor4_1 _16729_ (.A(_09791_),
    .B(_09789_),
    .C(_09790_),
    .D(\cpu.intr.r_timer_reload[16] ),
    .Y(_09862_));
 sg13g2_a21oi_1 _16730_ (.A1(_09817_),
    .A2(_09862_),
    .Y(_09863_),
    .B1(_09792_));
 sg13g2_mux2_1 _16731_ (.A0(_09863_),
    .A1(_09792_),
    .S(_09808_),
    .X(_09864_));
 sg13g2_buf_1 _16732_ (.A(_09788_),
    .X(_09865_));
 sg13g2_mux2_1 _16733_ (.A0(net880),
    .A1(_09864_),
    .S(net102),
    .X(_00062_));
 sg13g2_nor2_1 _16734_ (.A(\cpu.intr.r_timer_reload[17] ),
    .B(_09819_),
    .Y(_09866_));
 sg13g2_o21ai_1 _16735_ (.B1(_09791_),
    .Y(_09867_),
    .A1(_09792_),
    .A2(_09808_));
 sg13g2_inv_1 _16736_ (.Y(_09868_),
    .A(_09867_));
 sg13g2_o21ai_1 _16737_ (.B1(net102),
    .Y(_09869_),
    .A1(_09809_),
    .A2(_09868_));
 sg13g2_buf_1 _16738_ (.A(\cpu.dcache.wdata[1] ),
    .X(_09870_));
 sg13g2_buf_1 _16739_ (.A(_09870_),
    .X(_09871_));
 sg13g2_inv_2 _16740_ (.Y(_09872_),
    .A(net1111));
 sg13g2_buf_1 _16741_ (.A(_09872_),
    .X(_09873_));
 sg13g2_buf_1 _16742_ (.A(net879),
    .X(_09874_));
 sg13g2_buf_2 _16743_ (.A(net754),
    .X(_09875_));
 sg13g2_buf_1 _16744_ (.A(_09616_),
    .X(_09876_));
 sg13g2_nor4_1 _16745_ (.A(net673),
    .B(_09046_),
    .C(net672),
    .D(_09784_),
    .Y(_09877_));
 sg13g2_buf_1 _16746_ (.A(_09877_),
    .X(_09878_));
 sg13g2_buf_1 _16747_ (.A(_09878_),
    .X(_09879_));
 sg13g2_nand2_1 _16748_ (.Y(_09880_),
    .A(net1023),
    .B(net148));
 sg13g2_o21ai_1 _16749_ (.B1(_09880_),
    .Y(_00063_),
    .A1(_09866_),
    .A2(_09869_));
 sg13g2_buf_1 _16750_ (.A(\cpu.dcache.wdata[2] ),
    .X(_09881_));
 sg13g2_inv_1 _16751_ (.Y(_09882_),
    .A(_09881_));
 sg13g2_buf_1 _16752_ (.A(_09882_),
    .X(_09883_));
 sg13g2_buf_1 _16753_ (.A(net878),
    .X(_09884_));
 sg13g2_xnor2_1 _16754_ (.Y(_09885_),
    .A(_09790_),
    .B(_09809_));
 sg13g2_nor2_1 _16755_ (.A(_09878_),
    .B(_09885_),
    .Y(_09886_));
 sg13g2_o21ai_1 _16756_ (.B1(_09886_),
    .Y(_09887_),
    .A1(\cpu.intr.r_timer_reload[18] ),
    .A2(_09819_));
 sg13g2_o21ai_1 _16757_ (.B1(_09887_),
    .Y(_00064_),
    .A1(net753),
    .A2(net102));
 sg13g2_xor2_1 _16758_ (.B(_09810_),
    .A(_09789_),
    .X(_09888_));
 sg13g2_o21ai_1 _16759_ (.B1(_09888_),
    .Y(_09889_),
    .A1(\cpu.intr.r_timer_reload[19] ),
    .A2(_09819_));
 sg13g2_buf_1 _16760_ (.A(\cpu.dcache.wdata[3] ),
    .X(_09890_));
 sg13g2_nand2_1 _16761_ (.Y(_09891_),
    .A(net1106),
    .B(net148));
 sg13g2_o21ai_1 _16762_ (.B1(_09891_),
    .Y(_00065_),
    .A1(net148),
    .A2(_09889_));
 sg13g2_nor2b_1 _16763_ (.A(\cpu.intr.r_timer_reload[20] ),
    .B_N(_09817_),
    .Y(_09892_));
 sg13g2_nor3_1 _16764_ (.A(_09814_),
    .B(_09812_),
    .C(_09892_),
    .Y(_09893_));
 sg13g2_a21oi_1 _16765_ (.A1(_09814_),
    .A2(_09812_),
    .Y(_09894_),
    .B1(_09893_));
 sg13g2_buf_1 _16766_ (.A(\cpu.dcache.wdata[4] ),
    .X(_09895_));
 sg13g2_buf_1 _16767_ (.A(net1105),
    .X(_09896_));
 sg13g2_nand2_1 _16768_ (.Y(_09897_),
    .A(net1022),
    .B(net148));
 sg13g2_o21ai_1 _16769_ (.B1(_09897_),
    .Y(_00067_),
    .A1(net148),
    .A2(_09894_));
 sg13g2_nor2_1 _16770_ (.A(_09814_),
    .B(_09812_),
    .Y(_09898_));
 sg13g2_xnor2_1 _16771_ (.Y(_09899_),
    .A(_09813_),
    .B(_09898_));
 sg13g2_o21ai_1 _16772_ (.B1(_09788_),
    .Y(_09900_),
    .A1(\cpu.intr.r_timer_reload[21] ),
    .A2(_09819_));
 sg13g2_buf_2 _16773_ (.A(\cpu.dcache.wdata[5] ),
    .X(_09901_));
 sg13g2_buf_1 _16774_ (.A(_09901_),
    .X(_09902_));
 sg13g2_nand2_1 _16775_ (.Y(_09903_),
    .A(net1021),
    .B(_09878_));
 sg13g2_o21ai_1 _16776_ (.B1(_09903_),
    .Y(_00068_),
    .A1(_09899_),
    .A2(_09900_));
 sg13g2_nor3_1 _16777_ (.A(_09813_),
    .B(_09814_),
    .C(_09812_),
    .Y(_09904_));
 sg13g2_xnor2_1 _16778_ (.Y(_09905_),
    .A(_09816_),
    .B(_09904_));
 sg13g2_o21ai_1 _16779_ (.B1(_09788_),
    .Y(_09906_),
    .A1(\cpu.intr.r_timer_reload[22] ),
    .A2(_09819_));
 sg13g2_buf_2 _16780_ (.A(\cpu.dcache.wdata[6] ),
    .X(_09907_));
 sg13g2_buf_1 _16781_ (.A(_09907_),
    .X(_09908_));
 sg13g2_nand2_1 _16782_ (.Y(_09909_),
    .A(net1020),
    .B(_09878_));
 sg13g2_o21ai_1 _16783_ (.B1(_09909_),
    .Y(_00069_),
    .A1(_09905_),
    .A2(_09906_));
 sg13g2_buf_1 _16784_ (.A(\cpu.dcache.wdata[7] ),
    .X(_09910_));
 sg13g2_buf_1 _16785_ (.A(net1104),
    .X(_09911_));
 sg13g2_nor2b_1 _16786_ (.A(_09815_),
    .B_N(\cpu.intr.r_timer_reload[23] ),
    .Y(_09912_));
 sg13g2_nand2b_1 _16787_ (.Y(_09913_),
    .B(_09904_),
    .A_N(_09816_));
 sg13g2_mux2_1 _16788_ (.A0(_09912_),
    .A1(_09815_),
    .S(_09913_),
    .X(_09914_));
 sg13g2_mux2_1 _16789_ (.A0(net1019),
    .A1(_09914_),
    .S(net102),
    .X(_00070_));
 sg13g2_buf_1 _16790_ (.A(net604),
    .X(_09915_));
 sg13g2_buf_1 _16791_ (.A(_09915_),
    .X(_09916_));
 sg13g2_nand2_1 _16792_ (.Y(_09917_),
    .A(net463),
    .B(_09786_));
 sg13g2_buf_1 _16793_ (.A(_09917_),
    .X(_09918_));
 sg13g2_buf_1 _16794_ (.A(_09918_),
    .X(_09919_));
 sg13g2_nand2_1 _16795_ (.Y(_09920_),
    .A(net781),
    .B(_09261_));
 sg13g2_nor2_1 _16796_ (.A(net1025),
    .B(_09920_),
    .Y(_09921_));
 sg13g2_buf_1 _16797_ (.A(_09921_),
    .X(_09922_));
 sg13g2_buf_1 _16798_ (.A(net528),
    .X(_09923_));
 sg13g2_and2_1 _16799_ (.A(_09786_),
    .B(net462),
    .X(_09924_));
 sg13g2_buf_2 _16800_ (.A(_09924_),
    .X(_09925_));
 sg13g2_buf_1 _16801_ (.A(_09925_),
    .X(_09926_));
 sg13g2_buf_1 _16802_ (.A(net1024),
    .X(_09927_));
 sg13g2_a22oi_1 _16803_ (.Y(_09928_),
    .B1(net100),
    .B2(net877),
    .A2(_09919_),
    .A1(_00265_));
 sg13g2_inv_1 _16804_ (.Y(_00036_),
    .A(_09928_));
 sg13g2_buf_1 _16805_ (.A(_09870_),
    .X(_09929_));
 sg13g2_buf_1 _16806_ (.A(\cpu.intr.r_clock_count[0] ),
    .X(_09930_));
 sg13g2_buf_2 _16807_ (.A(\cpu.intr.r_clock_count[1] ),
    .X(_09931_));
 sg13g2_xor2_1 _16808_ (.B(_09931_),
    .A(_09930_),
    .X(_09932_));
 sg13g2_buf_1 _16809_ (.A(_09918_),
    .X(_09933_));
 sg13g2_buf_1 _16810_ (.A(net99),
    .X(_09934_));
 sg13g2_a22oi_1 _16811_ (.Y(_09935_),
    .B1(_09932_),
    .B2(net84),
    .A2(net100),
    .A1(net1018));
 sg13g2_inv_1 _16812_ (.Y(_00043_),
    .A(_09935_));
 sg13g2_buf_1 _16813_ (.A(_09881_),
    .X(_09936_));
 sg13g2_buf_1 _16814_ (.A(net1017),
    .X(_09937_));
 sg13g2_buf_1 _16815_ (.A(\cpu.intr.r_clock_count[2] ),
    .X(_09938_));
 sg13g2_nand2_1 _16816_ (.Y(_09939_),
    .A(_09930_),
    .B(_09931_));
 sg13g2_xnor2_1 _16817_ (.Y(_09940_),
    .A(_09938_),
    .B(_09939_));
 sg13g2_a22oi_1 _16818_ (.Y(_09941_),
    .B1(_09940_),
    .B2(net84),
    .A2(net100),
    .A1(net876));
 sg13g2_inv_1 _16819_ (.Y(_00044_),
    .A(_09941_));
 sg13g2_buf_1 _16820_ (.A(net1106),
    .X(_09942_));
 sg13g2_buf_2 _16821_ (.A(\cpu.intr.r_clock_count[3] ),
    .X(_09943_));
 sg13g2_nand2_1 _16822_ (.Y(_09944_),
    .A(_09931_),
    .B(_09938_));
 sg13g2_nor2_1 _16823_ (.A(_00265_),
    .B(_09944_),
    .Y(_09945_));
 sg13g2_xor2_1 _16824_ (.B(_09945_),
    .A(_09943_),
    .X(_09946_));
 sg13g2_a22oi_1 _16825_ (.Y(_09947_),
    .B1(_09946_),
    .B2(net84),
    .A2(net100),
    .A1(net1016));
 sg13g2_inv_1 _16826_ (.Y(_00045_),
    .A(_09947_));
 sg13g2_buf_2 _16827_ (.A(\cpu.intr.r_clock_count[4] ),
    .X(_09948_));
 sg13g2_and4_1 _16828_ (.A(_09930_),
    .B(_09931_),
    .C(_09938_),
    .D(_09943_),
    .X(_09949_));
 sg13g2_buf_1 _16829_ (.A(_09949_),
    .X(_09950_));
 sg13g2_xor2_1 _16830_ (.B(_09950_),
    .A(_09948_),
    .X(_09951_));
 sg13g2_a22oi_1 _16831_ (.Y(_09952_),
    .B1(_09951_),
    .B2(net84),
    .A2(_09926_),
    .A1(net1022));
 sg13g2_inv_1 _16832_ (.Y(_00046_),
    .A(_09952_));
 sg13g2_buf_2 _16833_ (.A(\cpu.intr.r_clock_count[5] ),
    .X(_09953_));
 sg13g2_nand3_1 _16834_ (.B(_09948_),
    .C(_09945_),
    .A(_09943_),
    .Y(_09954_));
 sg13g2_xnor2_1 _16835_ (.Y(_09955_),
    .A(_09953_),
    .B(_09954_));
 sg13g2_a22oi_1 _16836_ (.Y(_09956_),
    .B1(_09955_),
    .B2(net84),
    .A2(net100),
    .A1(net1021));
 sg13g2_inv_1 _16837_ (.Y(_00047_),
    .A(_09956_));
 sg13g2_buf_1 _16838_ (.A(net1020),
    .X(_09957_));
 sg13g2_buf_1 _16839_ (.A(_09925_),
    .X(_09958_));
 sg13g2_buf_1 _16840_ (.A(\cpu.intr.r_clock_count[6] ),
    .X(_09959_));
 sg13g2_nand3_1 _16841_ (.B(_09953_),
    .C(_09950_),
    .A(_09948_),
    .Y(_09960_));
 sg13g2_xor2_1 _16842_ (.B(_09960_),
    .A(_09959_),
    .X(_09961_));
 sg13g2_nand2_1 _16843_ (.Y(_09962_),
    .A(net768),
    .B(_09038_));
 sg13g2_buf_1 _16844_ (.A(_09962_),
    .X(_09963_));
 sg13g2_nor2_2 _16845_ (.A(_09335_),
    .B(net598),
    .Y(_09964_));
 sg13g2_buf_1 _16846_ (.A(_09964_),
    .X(_09965_));
 sg13g2_buf_1 _16847_ (.A(net461),
    .X(_09966_));
 sg13g2_and2_1 _16848_ (.A(_09786_),
    .B(net423),
    .X(_09967_));
 sg13g2_buf_1 _16849_ (.A(_09967_),
    .X(_09968_));
 sg13g2_nor3_1 _16850_ (.A(net98),
    .B(_09961_),
    .C(_09968_),
    .Y(_09969_));
 sg13g2_a21o_1 _16851_ (.A2(_09926_),
    .A1(net875),
    .B1(_09969_),
    .X(_00048_));
 sg13g2_buf_1 _16852_ (.A(\cpu.intr.r_clock_count[7] ),
    .X(_09970_));
 sg13g2_and3_1 _16853_ (.X(_09971_),
    .A(_09943_),
    .B(_09948_),
    .C(_09945_));
 sg13g2_nand3_1 _16854_ (.B(_09959_),
    .C(_09971_),
    .A(_09953_),
    .Y(_09972_));
 sg13g2_xnor2_1 _16855_ (.Y(_09973_),
    .A(_09970_),
    .B(_09972_));
 sg13g2_a22oi_1 _16856_ (.Y(_09974_),
    .B1(_09973_),
    .B2(net84),
    .A2(net100),
    .A1(net1019));
 sg13g2_inv_1 _16857_ (.Y(_00049_),
    .A(_09974_));
 sg13g2_buf_2 _16858_ (.A(\cpu.dcache.wdata[8] ),
    .X(_09975_));
 sg13g2_buf_2 _16859_ (.A(\cpu.intr.r_clock_count[8] ),
    .X(_09976_));
 sg13g2_nand2_1 _16860_ (.Y(_09977_),
    .A(_09948_),
    .B(_09950_));
 sg13g2_nand3_1 _16861_ (.B(_09959_),
    .C(_09970_),
    .A(_09953_),
    .Y(_09978_));
 sg13g2_nor2_1 _16862_ (.A(_09977_),
    .B(_09978_),
    .Y(_09979_));
 sg13g2_xor2_1 _16863_ (.B(_09979_),
    .A(_09976_),
    .X(_09980_));
 sg13g2_a22oi_1 _16864_ (.Y(_09981_),
    .B1(_09980_),
    .B2(net84),
    .A2(net100),
    .A1(_09975_));
 sg13g2_inv_1 _16865_ (.Y(_00050_),
    .A(_09981_));
 sg13g2_buf_1 _16866_ (.A(\cpu.intr.r_clock_count[9] ),
    .X(_09982_));
 sg13g2_nand2_1 _16867_ (.Y(_09983_),
    .A(_09976_),
    .B(_09979_));
 sg13g2_xnor2_1 _16868_ (.Y(_09984_),
    .A(_09982_),
    .B(_09983_));
 sg13g2_a22oi_1 _16869_ (.Y(_09985_),
    .B1(_09984_),
    .B2(_09934_),
    .A2(net100),
    .A1(\cpu.dcache.wdata[9] ));
 sg13g2_inv_1 _16870_ (.Y(_00051_),
    .A(_09985_));
 sg13g2_buf_2 _16871_ (.A(\cpu.dcache.wdata[10] ),
    .X(_09986_));
 sg13g2_buf_1 _16872_ (.A(\cpu.intr.r_clock_count[10] ),
    .X(_09987_));
 sg13g2_nand3_1 _16873_ (.B(_09982_),
    .C(_09979_),
    .A(_09976_),
    .Y(_09988_));
 sg13g2_xnor2_1 _16874_ (.Y(_09989_),
    .A(_09987_),
    .B(_09988_));
 sg13g2_a22oi_1 _16875_ (.Y(_09990_),
    .B1(_09989_),
    .B2(net84),
    .A2(net98),
    .A1(_09986_));
 sg13g2_inv_1 _16876_ (.Y(_00037_),
    .A(_09990_));
 sg13g2_buf_2 _16877_ (.A(\cpu.dcache.wdata[11] ),
    .X(_09991_));
 sg13g2_buf_2 _16878_ (.A(\cpu.intr.r_clock_count[11] ),
    .X(_09992_));
 sg13g2_nand3_1 _16879_ (.B(_09982_),
    .C(_09987_),
    .A(_09976_),
    .Y(_09993_));
 sg13g2_nor2_1 _16880_ (.A(_09978_),
    .B(_09993_),
    .Y(_09994_));
 sg13g2_nand2_1 _16881_ (.Y(_09995_),
    .A(_09971_),
    .B(_09994_));
 sg13g2_xnor2_1 _16882_ (.Y(_09996_),
    .A(_09992_),
    .B(_09995_));
 sg13g2_a22oi_1 _16883_ (.Y(_09997_),
    .B1(_09996_),
    .B2(net101),
    .A2(net98),
    .A1(_09991_));
 sg13g2_inv_1 _16884_ (.Y(_00038_),
    .A(_09997_));
 sg13g2_buf_1 _16885_ (.A(\cpu.intr.r_clock_count[12] ),
    .X(_09998_));
 sg13g2_nand4_1 _16886_ (.B(_09992_),
    .C(_09950_),
    .A(_09948_),
    .Y(_09999_),
    .D(_09994_));
 sg13g2_xnor2_1 _16887_ (.Y(_10000_),
    .A(_09998_),
    .B(_09999_));
 sg13g2_a22oi_1 _16888_ (.Y(_10001_),
    .B1(_10000_),
    .B2(net101),
    .A2(net98),
    .A1(\cpu.dcache.wdata[12] ));
 sg13g2_inv_1 _16889_ (.Y(_00039_),
    .A(_10001_));
 sg13g2_buf_2 _16890_ (.A(\cpu.intr.r_clock_count[13] ),
    .X(_10002_));
 sg13g2_nand3_1 _16891_ (.B(_09998_),
    .C(_09994_),
    .A(_09992_),
    .Y(_10003_));
 sg13g2_buf_1 _16892_ (.A(_10003_),
    .X(_10004_));
 sg13g2_nor2_1 _16893_ (.A(_09954_),
    .B(_10004_),
    .Y(_10005_));
 sg13g2_xor2_1 _16894_ (.B(_10005_),
    .A(_10002_),
    .X(_10006_));
 sg13g2_a22oi_1 _16895_ (.Y(_10007_),
    .B1(_10006_),
    .B2(net101),
    .A2(net98),
    .A1(\cpu.dcache.wdata[13] ));
 sg13g2_inv_1 _16896_ (.Y(_00040_),
    .A(_10007_));
 sg13g2_buf_2 _16897_ (.A(\cpu.intr.r_clock_count[14] ),
    .X(_10008_));
 sg13g2_nor2_1 _16898_ (.A(_09977_),
    .B(_10004_),
    .Y(_10009_));
 sg13g2_nand2_1 _16899_ (.Y(_10010_),
    .A(_10002_),
    .B(_10009_));
 sg13g2_xnor2_1 _16900_ (.Y(_10011_),
    .A(_10008_),
    .B(_10010_));
 sg13g2_a22oi_1 _16901_ (.Y(_10012_),
    .B1(_10011_),
    .B2(net101),
    .A2(_09958_),
    .A1(\cpu.dcache.wdata[14] ));
 sg13g2_inv_1 _16902_ (.Y(_00041_),
    .A(_10012_));
 sg13g2_buf_1 _16903_ (.A(\cpu.intr.r_clock_count[15] ),
    .X(_10013_));
 sg13g2_nand3_1 _16904_ (.B(_10008_),
    .C(_10005_),
    .A(_10002_),
    .Y(_10014_));
 sg13g2_xnor2_1 _16905_ (.Y(_10015_),
    .A(_10013_),
    .B(_10014_));
 sg13g2_a22oi_1 _16906_ (.Y(_10016_),
    .B1(_10015_),
    .B2(net101),
    .A2(net98),
    .A1(\cpu.dcache.wdata[15] ));
 sg13g2_inv_1 _16907_ (.Y(_00042_),
    .A(_10016_));
 sg13g2_buf_2 _16908_ (.A(\cpu.ex.r_wb_valid ),
    .X(_10017_));
 sg13g2_inv_1 _16909_ (.Y(_10018_),
    .A(_10017_));
 sg13g2_buf_1 _16910_ (.A(\cpu.ex.r_wb_addr[3] ),
    .X(_10019_));
 sg13g2_inv_1 _16911_ (.Y(_10020_),
    .A(_10019_));
 sg13g2_buf_2 _16912_ (.A(\cpu.ex.r_wb_addr[2] ),
    .X(_10021_));
 sg13g2_nand2_1 _16913_ (.Y(_10022_),
    .A(_10020_),
    .B(_10021_));
 sg13g2_buf_8 _16914_ (.A(\cpu.ex.r_wb_addr[1] ),
    .X(_10023_));
 sg13g2_buf_1 _16915_ (.A(\cpu.ex.r_wb_addr[0] ),
    .X(_10024_));
 sg13g2_buf_8 _16916_ (.A(_10024_),
    .X(_10025_));
 sg13g2_nand2_1 _16917_ (.Y(_10026_),
    .A(net1102),
    .B(net1015));
 sg13g2_nor3_1 _16918_ (.A(_10018_),
    .B(_10022_),
    .C(_10026_),
    .Y(_10027_));
 sg13g2_buf_2 _16919_ (.A(_10027_),
    .X(_10028_));
 sg13g2_buf_1 _16920_ (.A(_10028_),
    .X(_10029_));
 sg13g2_nand2_2 _16921_ (.Y(_10030_),
    .A(_10017_),
    .B(\cpu.dec.r_set_cc ));
 sg13g2_nor2_1 _16922_ (.A(_10029_),
    .B(_10030_),
    .Y(_10031_));
 sg13g2_inv_1 _16923_ (.Y(_10032_),
    .A(_00269_));
 sg13g2_nor4_1 _16924_ (.A(\cpu.ex.r_wb_addr[1] ),
    .B(_10024_),
    .C(net1103),
    .D(_10021_),
    .Y(_10033_));
 sg13g2_nor2_1 _16925_ (.A(_10018_),
    .B(_10033_),
    .Y(_10034_));
 sg13g2_buf_1 _16926_ (.A(\cpu.dec.r_rs1[3] ),
    .X(_10035_));
 sg13g2_buf_8 _16927_ (.A(_10035_),
    .X(_10036_));
 sg13g2_xor2_1 _16928_ (.B(_10036_),
    .A(net1103),
    .X(_10037_));
 sg13g2_buf_4 _16929_ (.X(_10038_),
    .A(\cpu.dec.r_rs1[0] ));
 sg13g2_xor2_1 _16930_ (.B(_10038_),
    .A(_10025_),
    .X(_10039_));
 sg13g2_buf_2 _16931_ (.A(\cpu.dec.r_rs1[2] ),
    .X(_10040_));
 sg13g2_xor2_1 _16932_ (.B(_10040_),
    .A(_10021_),
    .X(_10041_));
 sg13g2_buf_2 _16933_ (.A(\cpu.dec.r_rs1[1] ),
    .X(_10042_));
 sg13g2_buf_8 _16934_ (.A(_10042_),
    .X(_10043_));
 sg13g2_xor2_1 _16935_ (.B(_10043_),
    .A(net1102),
    .X(_10044_));
 sg13g2_nor4_1 _16936_ (.A(_10037_),
    .B(_10039_),
    .C(_10041_),
    .D(_10044_),
    .Y(_10045_));
 sg13g2_nand2_1 _16937_ (.Y(_10046_),
    .A(_10034_),
    .B(_10045_));
 sg13g2_buf_1 _16938_ (.A(_10046_),
    .X(_10047_));
 sg13g2_nor2_1 _16939_ (.A(_09036_),
    .B(net596),
    .Y(_10048_));
 sg13g2_buf_2 _16940_ (.A(_10043_),
    .X(_10049_));
 sg13g2_buf_1 _16941_ (.A(_10049_),
    .X(_10050_));
 sg13g2_buf_1 _16942_ (.A(net752),
    .X(_10051_));
 sg13g2_buf_1 _16943_ (.A(net671),
    .X(_10052_));
 sg13g2_buf_8 _16944_ (.A(_10038_),
    .X(_10053_));
 sg13g2_buf_8 _16945_ (.A(net1012),
    .X(_10054_));
 sg13g2_buf_1 _16946_ (.A(net873),
    .X(_10055_));
 sg13g2_buf_1 _16947_ (.A(_10055_),
    .X(_10056_));
 sg13g2_nor2b_1 _16948_ (.A(net1014),
    .B_N(_10040_),
    .Y(_10057_));
 sg13g2_buf_2 _16949_ (.A(_10057_),
    .X(_10058_));
 sg13g2_buf_1 _16950_ (.A(_10058_),
    .X(_10059_));
 sg13g2_buf_8 _16951_ (.A(_10040_),
    .X(_10060_));
 sg13g2_nor2b_1 _16952_ (.A(net1011),
    .B_N(net1014),
    .Y(_10061_));
 sg13g2_buf_1 _16953_ (.A(_10061_),
    .X(_10062_));
 sg13g2_buf_1 _16954_ (.A(_10062_),
    .X(_10063_));
 sg13g2_a22oi_1 _16955_ (.Y(_10064_),
    .B1(net668),
    .B2(\cpu.ex.r_10[2] ),
    .A2(net669),
    .A1(\cpu.ex.r_stmp[2] ));
 sg13g2_buf_8 _16956_ (.A(net1011),
    .X(_10065_));
 sg13g2_buf_2 _16957_ (.A(net872),
    .X(_10066_));
 sg13g2_nor2b_1 _16958_ (.A(_00238_),
    .B_N(net750),
    .Y(_10067_));
 sg13g2_nor2b_1 _16959_ (.A(net750),
    .B_N(\cpu.ex.r_11[2] ),
    .Y(_10068_));
 sg13g2_buf_8 _16960_ (.A(net1014),
    .X(_10069_));
 sg13g2_and2_1 _16961_ (.A(net873),
    .B(_10069_),
    .X(_10070_));
 sg13g2_buf_1 _16962_ (.A(_10070_),
    .X(_10071_));
 sg13g2_o21ai_1 _16963_ (.B1(_10071_),
    .Y(_10072_),
    .A1(_10067_),
    .A2(_10068_));
 sg13g2_o21ai_1 _16964_ (.B1(_10072_),
    .Y(_10073_),
    .A1(net670),
    .A2(_10064_));
 sg13g2_nand2_1 _16965_ (.Y(_10074_),
    .A(net595),
    .B(_10073_));
 sg13g2_buf_1 _16966_ (.A(\cpu.ex.r_mult[18] ),
    .X(_10075_));
 sg13g2_nor2b_1 _16967_ (.A(net871),
    .B_N(net1013),
    .Y(_10076_));
 sg13g2_buf_1 _16968_ (.A(_10076_),
    .X(_10077_));
 sg13g2_buf_1 _16969_ (.A(_10069_),
    .X(_10078_));
 sg13g2_buf_2 _16970_ (.A(\cpu.ex.mmu_read[2] ),
    .X(_10079_));
 sg13g2_inv_2 _16971_ (.Y(_10080_),
    .A(_10079_));
 sg13g2_nand2_1 _16972_ (.Y(_10081_),
    .A(net749),
    .B(\cpu.ex.r_13[2] ));
 sg13g2_o21ai_1 _16973_ (.B1(_10081_),
    .Y(_10082_),
    .A1(net749),
    .A2(_10080_));
 sg13g2_inv_1 _16974_ (.Y(_10083_),
    .A(net874));
 sg13g2_buf_1 _16975_ (.A(_10083_),
    .X(_10084_));
 sg13g2_a22oi_1 _16976_ (.Y(_10085_),
    .B1(_10082_),
    .B2(net666),
    .A2(net667),
    .A1(_10075_));
 sg13g2_mux2_1 _16977_ (.A0(\cpu.ex.r_lr[2] ),
    .A1(\cpu.ex.r_9[2] ),
    .S(net749),
    .X(_10086_));
 sg13g2_a22oi_1 _16978_ (.Y(_10087_),
    .B1(_10086_),
    .B2(net666),
    .A2(net667),
    .A1(\cpu.ex.r_epc[2] ));
 sg13g2_inv_1 _16979_ (.Y(_10088_),
    .A(net871));
 sg13g2_nor2_1 _16980_ (.A(_10083_),
    .B(net748),
    .Y(_10089_));
 sg13g2_nand2_1 _16981_ (.Y(_10090_),
    .A(net749),
    .B(\cpu.ex.r_12[2] ));
 sg13g2_o21ai_1 _16982_ (.B1(_10090_),
    .Y(_10091_),
    .A1(_08244_),
    .A2(net749));
 sg13g2_a22oi_1 _16983_ (.Y(_10092_),
    .B1(_10091_),
    .B2(_10084_),
    .A2(_10089_),
    .A1(\cpu.ex.r_14[2] ));
 sg13g2_buf_1 _16984_ (.A(\cpu.ex.r_sp[2] ),
    .X(_10093_));
 sg13g2_nor2b_1 _16985_ (.A(net1013),
    .B_N(net1014),
    .Y(_10094_));
 sg13g2_buf_1 _16986_ (.A(_10094_),
    .X(_10095_));
 sg13g2_buf_1 _16987_ (.A(_10095_),
    .X(_10096_));
 sg13g2_a22oi_1 _16988_ (.Y(_10097_),
    .B1(net665),
    .B2(\cpu.ex.r_8[2] ),
    .A2(net667),
    .A1(_10093_));
 sg13g2_inv_1 _16989_ (.Y(_10098_),
    .A(net872));
 sg13g2_buf_2 _16990_ (.A(_10098_),
    .X(_10099_));
 sg13g2_inv_1 _16991_ (.Y(_10100_),
    .A(_10038_));
 sg13g2_buf_1 _16992_ (.A(_10100_),
    .X(_10101_));
 sg13g2_mux4_1 _16993_ (.S0(_10099_),
    .A0(_10085_),
    .A1(_10087_),
    .A2(_10092_),
    .A3(_10097_),
    .S1(net870),
    .X(_10102_));
 sg13g2_and3_1 _16994_ (.X(_10103_),
    .A(_10047_),
    .B(_10074_),
    .C(_10102_));
 sg13g2_nor2_1 _16995_ (.A(_10048_),
    .B(_10103_),
    .Y(_10104_));
 sg13g2_nand4_1 _16996_ (.B(_08983_),
    .C(_08986_),
    .A(_08981_),
    .Y(_10105_),
    .D(_08988_));
 sg13g2_nand4_1 _16997_ (.B(_08999_),
    .C(_09003_),
    .A(_08994_),
    .Y(_10106_),
    .D(_09006_));
 sg13g2_buf_1 _16998_ (.A(_00252_),
    .X(_10107_));
 sg13g2_nor4_2 _16999_ (.A(_10042_),
    .B(_10038_),
    .C(_10035_),
    .Y(_10108_),
    .D(_10040_));
 sg13g2_or3_1 _17000_ (.A(_09013_),
    .B(_10107_),
    .C(_10108_),
    .X(_10109_));
 sg13g2_nor4_2 _17001_ (.A(_08979_),
    .B(_10105_),
    .C(_10106_),
    .Y(_10110_),
    .D(_10109_));
 sg13g2_nor4_1 _17002_ (.A(_09013_),
    .B(_09008_),
    .C(_10107_),
    .D(_10108_),
    .Y(_10111_));
 sg13g2_nor2b_1 _17003_ (.A(_08979_),
    .B_N(_10111_),
    .Y(_10112_));
 sg13g2_nor4_1 _17004_ (.A(_09013_),
    .B(_08966_),
    .C(_10107_),
    .D(_10108_),
    .Y(_10113_));
 sg13g2_or3_1 _17005_ (.A(_10110_),
    .B(_10112_),
    .C(_10113_),
    .X(_10114_));
 sg13g2_buf_8 _17006_ (.A(_10114_),
    .X(_10115_));
 sg13g2_and2_1 _17007_ (.A(_08220_),
    .B(_10115_),
    .X(_10116_));
 sg13g2_buf_1 _17008_ (.A(_10116_),
    .X(_10117_));
 sg13g2_a221oi_1 _17009_ (.B2(_08250_),
    .C1(_08254_),
    .B1(_08234_),
    .A1(_08178_),
    .Y(_10118_),
    .A2(_08193_));
 sg13g2_buf_8 _17010_ (.A(_10118_),
    .X(_10119_));
 sg13g2_buf_2 _17011_ (.A(\cpu.br ),
    .X(_10120_));
 sg13g2_inv_1 _17012_ (.Y(_10121_),
    .A(_10120_));
 sg13g2_a21o_1 _17013_ (.A2(_10115_),
    .A1(_08131_),
    .B1(_10121_),
    .X(_10122_));
 sg13g2_buf_1 _17014_ (.A(_10122_),
    .X(_10123_));
 sg13g2_a21o_1 _17015_ (.A2(net460),
    .A1(_10117_),
    .B1(_10123_),
    .X(_10124_));
 sg13g2_buf_8 _17016_ (.A(_10124_),
    .X(_10125_));
 sg13g2_buf_8 _17017_ (.A(_10125_),
    .X(_10126_));
 sg13g2_mux2_1 _17018_ (.A0(_10032_),
    .A1(_10104_),
    .S(net251),
    .X(_10127_));
 sg13g2_buf_2 _17019_ (.A(_10127_),
    .X(_10128_));
 sg13g2_buf_1 _17020_ (.A(\cpu.dec.r_rs2_pc ),
    .X(_10129_));
 sg13g2_buf_2 _17021_ (.A(\cpu.dec.needs_rs2 ),
    .X(_10130_));
 sg13g2_inv_2 _17022_ (.Y(_10131_),
    .A(_10130_));
 sg13g2_nor2_1 _17023_ (.A(net1101),
    .B(_10131_),
    .Y(_10132_));
 sg13g2_buf_2 _17024_ (.A(_10132_),
    .X(_10133_));
 sg13g2_buf_1 _17025_ (.A(\cpu.dec.r_rs2[2] ),
    .X(_10134_));
 sg13g2_xnor2_1 _17026_ (.Y(_10135_),
    .A(_10021_),
    .B(net1100));
 sg13g2_buf_8 _17027_ (.A(\cpu.dec.r_rs2[1] ),
    .X(_10136_));
 sg13g2_xnor2_1 _17028_ (.Y(_10137_),
    .A(_10023_),
    .B(_10136_));
 sg13g2_buf_1 _17029_ (.A(\cpu.dec.r_rs2[3] ),
    .X(_10138_));
 sg13g2_buf_8 _17030_ (.A(net1099),
    .X(_10139_));
 sg13g2_xnor2_1 _17031_ (.Y(_10140_),
    .A(net1103),
    .B(net1010));
 sg13g2_buf_1 _17032_ (.A(\cpu.dec.r_rs2[0] ),
    .X(_10141_));
 sg13g2_xnor2_1 _17033_ (.Y(_10142_),
    .A(_10024_),
    .B(net1098));
 sg13g2_and4_1 _17034_ (.A(_10135_),
    .B(_10137_),
    .C(_10140_),
    .D(_10142_),
    .X(_10143_));
 sg13g2_buf_8 _17035_ (.A(_10136_),
    .X(_10144_));
 sg13g2_nor2_2 _17036_ (.A(net1098),
    .B(net1009),
    .Y(_10145_));
 sg13g2_nor2_1 _17037_ (.A(net1010),
    .B(net1100),
    .Y(_10146_));
 sg13g2_buf_1 _17038_ (.A(_10146_),
    .X(_10147_));
 sg13g2_a22oi_1 _17039_ (.Y(_10148_),
    .B1(_10145_),
    .B2(_10147_),
    .A2(_10143_),
    .A1(_10034_));
 sg13g2_buf_2 _17040_ (.A(_10148_),
    .X(_10149_));
 sg13g2_nand2_1 _17041_ (.Y(_10150_),
    .A(_10133_),
    .B(_10149_));
 sg13g2_nand2_1 _17042_ (.Y(_10151_),
    .A(net1098),
    .B(_10136_));
 sg13g2_buf_1 _17043_ (.A(_10151_),
    .X(_10152_));
 sg13g2_buf_2 _17044_ (.A(\cpu.ex.r_mult[16] ),
    .X(_10153_));
 sg13g2_nor2b_1 _17045_ (.A(net1099),
    .B_N(net1100),
    .Y(_10154_));
 sg13g2_buf_2 _17046_ (.A(_10154_),
    .X(_10155_));
 sg13g2_buf_8 _17047_ (.A(net1100),
    .X(_10156_));
 sg13g2_nor2b_1 _17048_ (.A(net1008),
    .B_N(_10139_),
    .Y(_10157_));
 sg13g2_buf_8 _17049_ (.A(_10157_),
    .X(_10158_));
 sg13g2_a22oi_1 _17050_ (.Y(_10159_),
    .B1(net746),
    .B2(\cpu.ex.r_11[0] ),
    .A2(_10155_),
    .A1(_10153_));
 sg13g2_or2_1 _17051_ (.X(_10160_),
    .B(_10159_),
    .A(_10152_));
 sg13g2_nor2b_1 _17052_ (.A(net1009),
    .B_N(net1099),
    .Y(_10161_));
 sg13g2_buf_2 _17053_ (.A(_10161_),
    .X(_10162_));
 sg13g2_buf_1 _17054_ (.A(_10162_),
    .X(_10163_));
 sg13g2_inv_1 _17055_ (.Y(_10164_),
    .A(\cpu.ex.r_8[0] ));
 sg13g2_buf_1 _17056_ (.A(net1098),
    .X(_10165_));
 sg13g2_or2_1 _17057_ (.X(_10166_),
    .B(net1008),
    .A(net1007));
 sg13g2_buf_1 _17058_ (.A(_10166_),
    .X(_10167_));
 sg13g2_buf_1 _17059_ (.A(net1007),
    .X(_10168_));
 sg13g2_buf_8 _17060_ (.A(net1008),
    .X(_10169_));
 sg13g2_nand3_1 _17061_ (.B(net869),
    .C(net868),
    .A(\cpu.ex.r_13[0] ),
    .Y(_10170_));
 sg13g2_o21ai_1 _17062_ (.B1(_10170_),
    .Y(_10171_),
    .A1(_10164_),
    .A2(_10167_));
 sg13g2_nand2_1 _17063_ (.Y(_10172_),
    .A(net663),
    .B(_10171_));
 sg13g2_buf_1 _17064_ (.A(_10144_),
    .X(_10173_));
 sg13g2_nand3b_1 _17065_ (.B(net867),
    .C(\cpu.ex.r_10[0] ),
    .Y(_10174_),
    .A_N(net868));
 sg13g2_nand3b_1 _17066_ (.B(net868),
    .C(\cpu.ex.r_12[0] ),
    .Y(_10175_),
    .A_N(_10173_));
 sg13g2_buf_8 _17067_ (.A(_10165_),
    .X(_10176_));
 sg13g2_buf_8 _17068_ (.A(net1010),
    .X(_10177_));
 sg13g2_buf_8 _17069_ (.A(net865),
    .X(_10178_));
 sg13g2_nand2b_1 _17070_ (.Y(_10179_),
    .B(net745),
    .A_N(net866));
 sg13g2_a21oi_1 _17071_ (.A1(_10174_),
    .A2(_10175_),
    .Y(_10180_),
    .B1(_10179_));
 sg13g2_buf_1 _17072_ (.A(\cpu.ex.genblk3.r_prev_supmode ),
    .X(_10181_));
 sg13g2_nand3b_1 _17073_ (.B(net867),
    .C(_10181_),
    .Y(_10182_),
    .A_N(net745));
 sg13g2_nand3b_1 _17074_ (.B(_10178_),
    .C(\cpu.ex.r_9[0] ),
    .Y(_10183_),
    .A_N(net867));
 sg13g2_nand2b_1 _17075_ (.Y(_10184_),
    .B(net869),
    .A_N(_10169_));
 sg13g2_a21oi_1 _17076_ (.A1(_10182_),
    .A2(_10183_),
    .Y(_10185_),
    .B1(_10184_));
 sg13g2_nor2_1 _17077_ (.A(_10180_),
    .B(_10185_),
    .Y(_10186_));
 sg13g2_buf_8 _17078_ (.A(net1009),
    .X(_10187_));
 sg13g2_mux2_1 _17079_ (.A0(_08966_),
    .A1(\cpu.ex.r_stmp[0] ),
    .S(net864),
    .X(_10188_));
 sg13g2_nor2_2 _17080_ (.A(net1098),
    .B(net1010),
    .Y(_10189_));
 sg13g2_mux2_1 _17081_ (.A0(\cpu.ex.r_14[0] ),
    .A1(\cpu.ex.r_15[0] ),
    .S(net866),
    .X(_10190_));
 sg13g2_and2_1 _17082_ (.A(_10136_),
    .B(net1099),
    .X(_10191_));
 sg13g2_buf_1 _17083_ (.A(_10191_),
    .X(_10192_));
 sg13g2_a22oi_1 _17084_ (.Y(_10193_),
    .B1(_10190_),
    .B2(_10192_),
    .A2(_10189_),
    .A1(_10188_));
 sg13g2_buf_8 _17085_ (.A(net868),
    .X(_10194_));
 sg13g2_nand2b_1 _17086_ (.Y(_10195_),
    .B(net744),
    .A_N(_10193_));
 sg13g2_and4_1 _17087_ (.A(_10160_),
    .B(_10172_),
    .C(_10186_),
    .D(_10195_),
    .X(_10196_));
 sg13g2_inv_1 _17088_ (.Y(_10197_),
    .A(net1101));
 sg13g2_nand2_1 _17089_ (.Y(_10198_),
    .A(_10197_),
    .B(_10130_));
 sg13g2_buf_1 _17090_ (.A(_10198_),
    .X(_10199_));
 sg13g2_nand2b_1 _17091_ (.Y(_10200_),
    .B(_10017_),
    .A_N(_10033_));
 sg13g2_buf_8 _17092_ (.A(_10200_),
    .X(_10201_));
 sg13g2_nand4_1 _17093_ (.B(_10137_),
    .C(_10140_),
    .A(_10135_),
    .Y(_10202_),
    .D(_10142_));
 sg13g2_buf_2 _17094_ (.A(_10202_),
    .X(_10203_));
 sg13g2_nor3_2 _17095_ (.A(_10199_),
    .B(_10201_),
    .C(_10203_),
    .Y(_10204_));
 sg13g2_buf_1 _17096_ (.A(\cpu.dec.imm[0] ),
    .X(_10205_));
 sg13g2_nor2_1 _17097_ (.A(net1101),
    .B(_10130_),
    .Y(_10206_));
 sg13g2_buf_2 _17098_ (.A(_10206_),
    .X(_10207_));
 sg13g2_and2_1 _17099_ (.A(_10205_),
    .B(_10207_),
    .X(_10208_));
 sg13g2_a21oi_1 _17100_ (.A1(net1118),
    .A2(_10204_),
    .Y(_10209_),
    .B1(_10208_));
 sg13g2_o21ai_1 _17101_ (.B1(_10209_),
    .Y(_10210_),
    .A1(_10150_),
    .A2(_10196_));
 sg13g2_buf_1 _17102_ (.A(_10210_),
    .X(_10211_));
 sg13g2_and2_1 _17103_ (.A(_10034_),
    .B(_10045_),
    .X(_10212_));
 sg13g2_buf_8 _17104_ (.A(_10212_),
    .X(_10213_));
 sg13g2_buf_1 _17105_ (.A(net871),
    .X(_10214_));
 sg13g2_nor2_1 _17106_ (.A(_10050_),
    .B(net742),
    .Y(_10215_));
 sg13g2_mux2_1 _17107_ (.A0(\cpu.ex.r_epc[1] ),
    .A1(\cpu.ex.r_11[1] ),
    .S(net742),
    .X(_10216_));
 sg13g2_a22oi_1 _17108_ (.Y(_10217_),
    .B1(_10216_),
    .B2(_10051_),
    .A2(_10215_),
    .A1(\cpu.ex.r_lr[1] ));
 sg13g2_nor2b_1 _17109_ (.A(net1011),
    .B_N(_10038_),
    .Y(_10218_));
 sg13g2_buf_2 _17110_ (.A(_10218_),
    .X(_10219_));
 sg13g2_nand2b_1 _17111_ (.Y(_10220_),
    .B(_10219_),
    .A_N(_10217_));
 sg13g2_and2_1 _17112_ (.A(net871),
    .B(net872),
    .X(_10221_));
 sg13g2_buf_2 _17113_ (.A(_10221_),
    .X(_10222_));
 sg13g2_buf_1 _17114_ (.A(\cpu.ex.r_sp[1] ),
    .X(_10223_));
 sg13g2_buf_1 _17115_ (.A(_10060_),
    .X(_10224_));
 sg13g2_mux2_1 _17116_ (.A0(_10223_),
    .A1(\cpu.ex.r_stmp[1] ),
    .S(net863),
    .X(_10225_));
 sg13g2_a22oi_1 _17117_ (.Y(_10226_),
    .B1(_10225_),
    .B2(net748),
    .A2(_10222_),
    .A1(\cpu.ex.r_14[1] ));
 sg13g2_nor2b_1 _17118_ (.A(_10038_),
    .B_N(net1013),
    .Y(_10227_));
 sg13g2_buf_1 _17119_ (.A(_10227_),
    .X(_10228_));
 sg13g2_buf_1 _17120_ (.A(_10228_),
    .X(_10229_));
 sg13g2_nand2b_1 _17121_ (.Y(_10230_),
    .B(_10229_),
    .A_N(_10226_));
 sg13g2_nor2b_2 _17122_ (.A(net752),
    .B_N(net863),
    .Y(_10231_));
 sg13g2_inv_1 _17123_ (.Y(_10232_),
    .A(\cpu.ex.mmu_read[1] ));
 sg13g2_nand2b_1 _17124_ (.Y(_10233_),
    .B(net1012),
    .A_N(net1014));
 sg13g2_buf_1 _17125_ (.A(_10233_),
    .X(_10234_));
 sg13g2_buf_1 _17126_ (.A(net1012),
    .X(_10235_));
 sg13g2_nand3b_1 _17127_ (.B(net742),
    .C(\cpu.ex.r_12[1] ),
    .Y(_10236_),
    .A_N(_10235_));
 sg13g2_o21ai_1 _17128_ (.B1(_10236_),
    .Y(_10237_),
    .A1(_10232_),
    .A2(_10234_));
 sg13g2_buf_1 _17129_ (.A(\cpu.ex.r_prev_ie ),
    .X(_10238_));
 sg13g2_nor2_1 _17130_ (.A(net874),
    .B(net873),
    .Y(_10239_));
 sg13g2_buf_1 _17131_ (.A(\cpu.ex.r_mult[17] ),
    .X(_10240_));
 sg13g2_and3_1 _17132_ (.X(_10241_),
    .A(net752),
    .B(net862),
    .C(_10240_));
 sg13g2_a21o_1 _17133_ (.A2(_10239_),
    .A1(_10238_),
    .B1(_10241_),
    .X(_10242_));
 sg13g2_a22oi_1 _17134_ (.Y(_10243_),
    .B1(_10242_),
    .B2(_10059_),
    .A2(_10237_),
    .A1(_10231_));
 sg13g2_nor2b_1 _17135_ (.A(net874),
    .B_N(net1012),
    .Y(_10244_));
 sg13g2_buf_1 _17136_ (.A(_10244_),
    .X(_10245_));
 sg13g2_nand3_1 _17137_ (.B(net668),
    .C(_10245_),
    .A(\cpu.ex.r_9[1] ),
    .Y(_10246_));
 sg13g2_and4_1 _17138_ (.A(_10220_),
    .B(_10230_),
    .C(_10243_),
    .D(_10246_),
    .X(_10247_));
 sg13g2_buf_1 _17139_ (.A(_10078_),
    .X(_10248_));
 sg13g2_nor2_2 _17140_ (.A(_10235_),
    .B(net863),
    .Y(_10249_));
 sg13g2_and2_1 _17141_ (.A(_10054_),
    .B(net872),
    .X(_10250_));
 sg13g2_buf_1 _17142_ (.A(_10250_),
    .X(_10251_));
 sg13g2_a22oi_1 _17143_ (.Y(_10252_),
    .B1(_10251_),
    .B2(\cpu.ex.r_13[1] ),
    .A2(_10249_),
    .A1(\cpu.ex.r_8[1] ));
 sg13g2_inv_1 _17144_ (.Y(_10253_),
    .A(_00237_));
 sg13g2_a221oi_1 _17145_ (.B2(_10253_),
    .C1(_10083_),
    .B1(_10251_),
    .A1(\cpu.ex.r_10[1] ),
    .Y(_10254_),
    .A2(_10249_));
 sg13g2_a21oi_1 _17146_ (.A1(_10084_),
    .A2(_10252_),
    .Y(_10255_),
    .B1(_10254_));
 sg13g2_a21oi_1 _17147_ (.A1(_10248_),
    .A2(_10255_),
    .Y(_10256_),
    .B1(_10213_));
 sg13g2_a22oi_1 _17148_ (.Y(_10257_),
    .B1(_10247_),
    .B2(_10256_),
    .A2(net594),
    .A1(_09872_));
 sg13g2_buf_2 _17149_ (.A(_10257_),
    .X(_10258_));
 sg13g2_nor2_2 _17150_ (.A(_08132_),
    .B(_10121_),
    .Y(_10259_));
 sg13g2_inv_1 _17151_ (.Y(_10260_),
    .A(_09013_));
 sg13g2_o21ai_1 _17152_ (.B1(_08966_),
    .Y(_10261_),
    .A1(_08979_),
    .A2(_09010_));
 sg13g2_and3_1 _17153_ (.X(_10262_),
    .A(_10260_),
    .B(_08220_),
    .C(_10261_));
 sg13g2_o21ai_1 _17154_ (.B1(_10262_),
    .Y(_10263_),
    .A1(_08131_),
    .A2(net460));
 sg13g2_buf_8 _17155_ (.A(_10263_),
    .X(_10264_));
 sg13g2_nand4_1 _17156_ (.B(_10258_),
    .C(_10259_),
    .A(net374),
    .Y(_10265_),
    .D(net373));
 sg13g2_buf_1 _17157_ (.A(_10224_),
    .X(_10266_));
 sg13g2_nor2_1 _17158_ (.A(net862),
    .B(_10214_),
    .Y(_10267_));
 sg13g2_a22oi_1 _17159_ (.Y(_10268_),
    .B1(_10071_),
    .B2(\cpu.ex.r_13[0] ),
    .A2(_10267_),
    .A1(_08966_));
 sg13g2_mux2_1 _17160_ (.A0(\cpu.ex.r_stmp[0] ),
    .A1(_10153_),
    .S(net862),
    .X(_10269_));
 sg13g2_nand2_1 _17161_ (.Y(_10270_),
    .A(net667),
    .B(_10269_));
 sg13g2_o21ai_1 _17162_ (.B1(_10270_),
    .Y(_10271_),
    .A1(_10051_),
    .A2(_10268_));
 sg13g2_buf_1 _17163_ (.A(net862),
    .X(_10272_));
 sg13g2_and2_1 _17164_ (.A(_10050_),
    .B(\cpu.ex.r_10[0] ),
    .X(_10273_));
 sg13g2_a21oi_1 _17165_ (.A1(_10083_),
    .A2(\cpu.ex.r_8[0] ),
    .Y(_10274_),
    .B1(_10273_));
 sg13g2_nand3_1 _17166_ (.B(net740),
    .C(\cpu.ex.r_9[0] ),
    .A(net666),
    .Y(_10275_));
 sg13g2_o21ai_1 _17167_ (.B1(_10275_),
    .Y(_10276_),
    .A1(net740),
    .A2(_10274_));
 sg13g2_and2_1 _17168_ (.A(net874),
    .B(net873),
    .X(_10277_));
 sg13g2_buf_2 _17169_ (.A(_10277_),
    .X(_10278_));
 sg13g2_a22oi_1 _17170_ (.Y(_10279_),
    .B1(_10278_),
    .B2(\cpu.ex.r_15[0] ),
    .A2(_10239_),
    .A1(\cpu.ex.r_12[0] ));
 sg13g2_nor2b_1 _17171_ (.A(_10279_),
    .B_N(_10222_),
    .Y(_10280_));
 sg13g2_a221oi_1 _17172_ (.B2(_10063_),
    .C1(_10280_),
    .B1(_10276_),
    .A1(net741),
    .Y(_10281_),
    .A2(_10271_));
 sg13g2_nand2b_1 _17173_ (.Y(_10282_),
    .B(net1012),
    .A_N(net1011));
 sg13g2_and2_1 _17174_ (.A(net749),
    .B(\cpu.ex.r_11[0] ),
    .X(_10283_));
 sg13g2_a21oi_1 _17175_ (.A1(_10181_),
    .A2(_10088_),
    .Y(_10284_),
    .B1(_10283_));
 sg13g2_nor2b_1 _17176_ (.A(_10053_),
    .B_N(net871),
    .Y(_10285_));
 sg13g2_buf_2 _17177_ (.A(_10285_),
    .X(_10286_));
 sg13g2_nand3_1 _17178_ (.B(\cpu.ex.r_14[0] ),
    .C(_10286_),
    .A(net741),
    .Y(_10287_));
 sg13g2_o21ai_1 _17179_ (.B1(_10287_),
    .Y(_10288_),
    .A1(_10282_),
    .A2(_10284_));
 sg13g2_a21oi_1 _17180_ (.A1(_10052_),
    .A2(_10288_),
    .Y(_10289_),
    .B1(net594));
 sg13g2_a22oi_1 _17181_ (.Y(_10290_),
    .B1(_10281_),
    .B2(_10289_),
    .A2(net594),
    .A1(_08190_));
 sg13g2_buf_1 _17182_ (.A(_10290_),
    .X(_10291_));
 sg13g2_and2_1 _17183_ (.A(net1099),
    .B(_10134_),
    .X(_10292_));
 sg13g2_buf_1 _17184_ (.A(_10292_),
    .X(_10293_));
 sg13g2_mux2_1 _17185_ (.A0(\cpu.ex.r_epc[1] ),
    .A1(_10240_),
    .S(net1008),
    .X(_10294_));
 sg13g2_inv_1 _17186_ (.Y(_10295_),
    .A(net1010));
 sg13g2_inv_2 _17187_ (.Y(_10296_),
    .A(net1098));
 sg13g2_a221oi_1 _17188_ (.B2(_10295_),
    .C1(_10296_),
    .B1(_10294_),
    .A1(_10253_),
    .Y(_10297_),
    .A2(_10293_));
 sg13g2_a21oi_1 _17189_ (.A1(\cpu.ex.r_10[1] ),
    .A2(_10157_),
    .Y(_10298_),
    .B1(_10165_));
 sg13g2_o21ai_1 _17190_ (.B1(_10187_),
    .Y(_10299_),
    .A1(_10297_),
    .A2(_10298_));
 sg13g2_inv_2 _17191_ (.Y(_10300_),
    .A(net1008));
 sg13g2_buf_1 _17192_ (.A(_10300_),
    .X(_10301_));
 sg13g2_nor2b_1 _17193_ (.A(_10141_),
    .B_N(net1010),
    .Y(_10302_));
 sg13g2_mux2_1 _17194_ (.A0(\cpu.ex.mmu_read[1] ),
    .A1(\cpu.ex.r_13[1] ),
    .S(_10139_),
    .X(_10303_));
 sg13g2_a22oi_1 _17195_ (.Y(_10304_),
    .B1(_10303_),
    .B2(net1007),
    .A2(_10302_),
    .A1(\cpu.ex.r_12[1] ));
 sg13g2_inv_1 _17196_ (.Y(_10305_),
    .A(net1009));
 sg13g2_buf_1 _17197_ (.A(_10305_),
    .X(_10306_));
 sg13g2_o21ai_1 _17198_ (.B1(_10306_),
    .Y(_10307_),
    .A1(net739),
    .A2(_10304_));
 sg13g2_nor2b_1 _17199_ (.A(_10138_),
    .B_N(_10136_),
    .Y(_10308_));
 sg13g2_buf_2 _17200_ (.A(_10308_),
    .X(_10309_));
 sg13g2_a22oi_1 _17201_ (.Y(_10310_),
    .B1(_10309_),
    .B2(_10223_),
    .A2(_10162_),
    .A1(\cpu.ex.r_8[1] ));
 sg13g2_nor2_1 _17202_ (.A(_10136_),
    .B(net1099),
    .Y(_10311_));
 sg13g2_buf_2 _17203_ (.A(_10311_),
    .X(_10312_));
 sg13g2_a221oi_1 _17204_ (.B2(_10238_),
    .C1(_10300_),
    .B1(_10312_),
    .A1(\cpu.ex.r_14[1] ),
    .Y(_10313_),
    .A2(_10192_));
 sg13g2_a21oi_1 _17205_ (.A1(net739),
    .A2(_10310_),
    .Y(_10314_),
    .B1(_10313_));
 sg13g2_nor2_1 _17206_ (.A(_10144_),
    .B(_10156_),
    .Y(_10315_));
 sg13g2_buf_2 _17207_ (.A(_10315_),
    .X(_10316_));
 sg13g2_and2_1 _17208_ (.A(\cpu.ex.r_lr[1] ),
    .B(net1007),
    .X(_10317_));
 sg13g2_nor2b_1 _17209_ (.A(net1007),
    .B_N(\cpu.ex.r_stmp[1] ),
    .Y(_10318_));
 sg13g2_and2_1 _17210_ (.A(_10136_),
    .B(net1100),
    .X(_10319_));
 sg13g2_buf_2 _17211_ (.A(_10319_),
    .X(_10320_));
 sg13g2_a22oi_1 _17212_ (.Y(_10321_),
    .B1(_10318_),
    .B2(_10320_),
    .A2(_10317_),
    .A1(_10316_));
 sg13g2_mux2_1 _17213_ (.A0(\cpu.ex.r_9[1] ),
    .A1(\cpu.ex.r_11[1] ),
    .S(net1009),
    .X(_10322_));
 sg13g2_nand3_1 _17214_ (.B(_10158_),
    .C(_10322_),
    .A(_10176_),
    .Y(_10323_));
 sg13g2_o21ai_1 _17215_ (.B1(_10323_),
    .Y(_10324_),
    .A1(_10177_),
    .A2(_10321_));
 sg13g2_a221oi_1 _17216_ (.B2(_10296_),
    .C1(_10324_),
    .B1(_10314_),
    .A1(_10299_),
    .Y(_10325_),
    .A2(_10307_));
 sg13g2_buf_2 _17217_ (.A(_00184_),
    .X(_10326_));
 sg13g2_buf_1 _17218_ (.A(\cpu.dec.imm[1] ),
    .X(_10327_));
 sg13g2_nor2_1 _17219_ (.A(_10327_),
    .B(net1101),
    .Y(_10328_));
 sg13g2_a22oi_1 _17220_ (.Y(_10329_),
    .B1(_10328_),
    .B2(_10131_),
    .A2(_10326_),
    .A1(net1101));
 sg13g2_nand2_1 _17221_ (.Y(_10330_),
    .A(_10149_),
    .B(_10329_));
 sg13g2_nor3_1 _17222_ (.A(_09872_),
    .B(_10201_),
    .C(_10203_),
    .Y(_10331_));
 sg13g2_o21ai_1 _17223_ (.B1(_10329_),
    .Y(_10332_),
    .A1(_10199_),
    .A2(_10331_));
 sg13g2_o21ai_1 _17224_ (.B1(_10332_),
    .Y(_10333_),
    .A1(_10325_),
    .A2(_10330_));
 sg13g2_buf_8 _17225_ (.A(_10333_),
    .X(_10334_));
 sg13g2_a22oi_1 _17226_ (.Y(_10335_),
    .B1(_10334_),
    .B2(_10258_),
    .A2(_10291_),
    .A1(net374));
 sg13g2_nor2_1 _17227_ (.A(_10258_),
    .B(_10334_),
    .Y(_10336_));
 sg13g2_or2_1 _17228_ (.X(_10337_),
    .B(_10336_),
    .A(_10335_));
 sg13g2_a21oi_1 _17229_ (.A1(_10117_),
    .A2(net460),
    .Y(_10338_),
    .B1(_10123_));
 sg13g2_buf_1 _17230_ (.A(_10338_),
    .X(_10339_));
 sg13g2_a21oi_1 _17231_ (.A1(_10265_),
    .A2(_10337_),
    .Y(_10340_),
    .B1(net303));
 sg13g2_and2_1 _17232_ (.A(_10259_),
    .B(net373),
    .X(_10341_));
 sg13g2_nand2_1 _17233_ (.Y(_10342_),
    .A(_10145_),
    .B(net747));
 sg13g2_o21ai_1 _17234_ (.B1(_10342_),
    .Y(_10343_),
    .A1(_10201_),
    .A2(_10203_));
 sg13g2_buf_2 _17235_ (.A(_10343_),
    .X(_10344_));
 sg13g2_nor2_1 _17236_ (.A(net743),
    .B(_10344_),
    .Y(_10345_));
 sg13g2_nand4_1 _17237_ (.B(_10172_),
    .C(_10186_),
    .A(_10160_),
    .Y(_10346_),
    .D(_10195_));
 sg13g2_a221oi_1 _17238_ (.B2(net1118),
    .C1(_10208_),
    .B1(_10204_),
    .A1(_10345_),
    .Y(_10347_),
    .A2(_10346_));
 sg13g2_buf_2 _17239_ (.A(_10347_),
    .X(_10348_));
 sg13g2_inv_1 _17240_ (.Y(_10349_),
    .A(_10334_));
 sg13g2_nor2_1 _17241_ (.A(_10348_),
    .B(_10349_),
    .Y(_10350_));
 sg13g2_and2_1 _17242_ (.A(_10341_),
    .B(_10350_),
    .X(_10351_));
 sg13g2_nor2_1 _17243_ (.A(_10326_),
    .B(net251),
    .Y(_10352_));
 sg13g2_and2_1 _17244_ (.A(_10211_),
    .B(_10259_),
    .X(_10353_));
 sg13g2_a21o_1 _17245_ (.A2(_10353_),
    .A1(net373),
    .B1(_10334_),
    .X(_10354_));
 sg13g2_and2_1 _17246_ (.A(_10352_),
    .B(_10354_),
    .X(_10355_));
 sg13g2_or4_1 _17247_ (.A(_10128_),
    .B(_10340_),
    .C(_10351_),
    .D(_10355_),
    .X(_10356_));
 sg13g2_buf_1 _17248_ (.A(net596),
    .X(_10357_));
 sg13g2_nor2_1 _17249_ (.A(_09103_),
    .B(net527),
    .Y(_10358_));
 sg13g2_buf_1 _17250_ (.A(\cpu.ex.r_sp[3] ),
    .X(_10359_));
 sg13g2_nor2_1 _17251_ (.A(net871),
    .B(_10065_),
    .Y(_10360_));
 sg13g2_buf_2 _17252_ (.A(_10360_),
    .X(_10361_));
 sg13g2_mux2_1 _17253_ (.A0(\cpu.ex.r_10[3] ),
    .A1(\cpu.ex.r_14[3] ),
    .S(net750),
    .X(_10362_));
 sg13g2_a22oi_1 _17254_ (.Y(_10363_),
    .B1(_10362_),
    .B2(net660),
    .A2(_10361_),
    .A1(_10359_));
 sg13g2_nand2b_1 _17255_ (.Y(_10364_),
    .B(net662),
    .A_N(_10363_));
 sg13g2_buf_1 _17256_ (.A(\cpu.ex.r_mult[19] ),
    .X(_10365_));
 sg13g2_a22oi_1 _17257_ (.Y(_10366_),
    .B1(net668),
    .B2(\cpu.ex.r_11[3] ),
    .A2(net669),
    .A1(_10365_));
 sg13g2_nand2b_1 _17258_ (.Y(_10367_),
    .B(_10278_),
    .A_N(_10366_));
 sg13g2_nand2_1 _17259_ (.Y(_10368_),
    .A(net740),
    .B(\cpu.ex.r_13[3] ));
 sg13g2_nand2b_1 _17260_ (.Y(_10369_),
    .B(\cpu.ex.r_12[3] ),
    .A_N(net751));
 sg13g2_a21oi_1 _17261_ (.A1(_10368_),
    .A2(_10369_),
    .Y(_10370_),
    .B1(net671));
 sg13g2_nand2_2 _17262_ (.Y(_10371_),
    .A(net752),
    .B(net751));
 sg13g2_nor2_1 _17263_ (.A(_00239_),
    .B(_10371_),
    .Y(_10372_));
 sg13g2_o21ai_1 _17264_ (.B1(_10222_),
    .Y(_10373_),
    .A1(_10370_),
    .A2(_10372_));
 sg13g2_nor2b_1 _17265_ (.A(_10054_),
    .B_N(_10065_),
    .Y(_10374_));
 sg13g2_buf_2 _17266_ (.A(_10374_),
    .X(_10375_));
 sg13g2_a22oi_1 _17267_ (.Y(_10376_),
    .B1(_10375_),
    .B2(\cpu.ex.r_stmp[3] ),
    .A2(_10219_),
    .A1(\cpu.ex.r_epc[3] ));
 sg13g2_nand2b_1 _17268_ (.Y(_10377_),
    .B(_10077_),
    .A_N(_10376_));
 sg13g2_nand4_1 _17269_ (.B(_10367_),
    .C(_10373_),
    .A(_10364_),
    .Y(_10378_),
    .D(_10377_));
 sg13g2_nor2b_1 _17270_ (.A(net660),
    .B_N(_10272_),
    .Y(_10379_));
 sg13g2_a22oi_1 _17271_ (.Y(_10380_),
    .B1(_10286_),
    .B2(\cpu.ex.r_8[3] ),
    .A2(_10379_),
    .A1(\cpu.ex.r_lr[3] ));
 sg13g2_nor2_1 _17272_ (.A(_10266_),
    .B(_10380_),
    .Y(_10381_));
 sg13g2_buf_1 _17273_ (.A(\cpu.ex.mmu_read[3] ),
    .X(_10382_));
 sg13g2_a22oi_1 _17274_ (.Y(_10383_),
    .B1(net668),
    .B2(\cpu.ex.r_9[3] ),
    .A2(_10059_),
    .A1(_10382_));
 sg13g2_a21oi_1 _17275_ (.A1(net1056),
    .A2(net669),
    .Y(_10384_),
    .B1(net670));
 sg13g2_a21oi_1 _17276_ (.A1(net670),
    .A2(_10383_),
    .Y(_10385_),
    .B1(_10384_));
 sg13g2_o21ai_1 _17277_ (.B1(net666),
    .Y(_10386_),
    .A1(_10381_),
    .A2(_10385_));
 sg13g2_nand3b_1 _17278_ (.B(_10386_),
    .C(net527),
    .Y(_10387_),
    .A_N(_10378_));
 sg13g2_nand2b_1 _17279_ (.Y(_10388_),
    .B(_10387_),
    .A_N(_10358_));
 sg13g2_mux2_1 _17280_ (.A0(_00175_),
    .A1(_10388_),
    .S(_10126_),
    .X(_10389_));
 sg13g2_buf_2 _17281_ (.A(_10389_),
    .X(_10390_));
 sg13g2_buf_1 _17282_ (.A(_10295_),
    .X(_10391_));
 sg13g2_nor2b_1 _17283_ (.A(net1100),
    .B_N(_10136_),
    .Y(_10392_));
 sg13g2_buf_2 _17284_ (.A(_10392_),
    .X(_10393_));
 sg13g2_mux2_1 _17285_ (.A0(\cpu.ex.r_lr[3] ),
    .A1(_10382_),
    .S(net1100),
    .X(_10394_));
 sg13g2_a22oi_1 _17286_ (.Y(_10395_),
    .B1(_10394_),
    .B2(_10305_),
    .A2(_10393_),
    .A1(\cpu.ex.r_epc[3] ));
 sg13g2_nand3_1 _17287_ (.B(_10296_),
    .C(_10320_),
    .A(\cpu.ex.r_stmp[3] ),
    .Y(_10396_));
 sg13g2_o21ai_1 _17288_ (.B1(_10396_),
    .Y(_10397_),
    .A1(_10296_),
    .A2(_10395_));
 sg13g2_and2_1 _17289_ (.A(net737),
    .B(_10397_),
    .X(_10398_));
 sg13g2_nor2b_1 _17290_ (.A(net1098),
    .B_N(net1009),
    .Y(_10399_));
 sg13g2_buf_2 _17291_ (.A(_10399_),
    .X(_10400_));
 sg13g2_nand2_2 _17292_ (.Y(_10401_),
    .A(net865),
    .B(_10400_));
 sg13g2_and2_1 _17293_ (.A(\cpu.ex.r_14[3] ),
    .B(_10156_),
    .X(_10402_));
 sg13g2_a21oi_1 _17294_ (.A1(\cpu.ex.r_10[3] ),
    .A2(net739),
    .Y(_10403_),
    .B1(_10402_));
 sg13g2_nor2_1 _17295_ (.A(_10401_),
    .B(_10403_),
    .Y(_10404_));
 sg13g2_nand2_1 _17296_ (.Y(_10405_),
    .A(_10187_),
    .B(net739));
 sg13g2_and2_1 _17297_ (.A(net1098),
    .B(net1099),
    .X(_10406_));
 sg13g2_buf_1 _17298_ (.A(_10406_),
    .X(_10407_));
 sg13g2_a22oi_1 _17299_ (.Y(_10408_),
    .B1(_10407_),
    .B2(\cpu.ex.r_11[3] ),
    .A2(_10189_),
    .A1(_10359_));
 sg13g2_nor2b_1 _17300_ (.A(_10152_),
    .B_N(_10155_),
    .Y(_10409_));
 sg13g2_mux2_1 _17301_ (.A0(\cpu.ex.r_8[3] ),
    .A1(\cpu.ex.r_9[3] ),
    .S(net1007),
    .X(_10410_));
 sg13g2_nand2b_1 _17302_ (.Y(_10411_),
    .B(net1099),
    .A_N(net1100));
 sg13g2_buf_1 _17303_ (.A(_10411_),
    .X(_10412_));
 sg13g2_nor2_2 _17304_ (.A(net1009),
    .B(_10412_),
    .Y(_10413_));
 sg13g2_a22oi_1 _17305_ (.Y(_10414_),
    .B1(_10410_),
    .B2(_10413_),
    .A2(_10409_),
    .A1(_10365_));
 sg13g2_o21ai_1 _17306_ (.B1(_10414_),
    .Y(_10415_),
    .A1(_10405_),
    .A2(_10408_));
 sg13g2_and2_1 _17307_ (.A(\cpu.ex.r_12[3] ),
    .B(_10145_),
    .X(_10416_));
 sg13g2_nor2_1 _17308_ (.A(_00239_),
    .B(_10152_),
    .Y(_10417_));
 sg13g2_o21ai_1 _17309_ (.B1(_10177_),
    .Y(_10418_),
    .A1(_10416_),
    .A2(_10417_));
 sg13g2_a22oi_1 _17310_ (.Y(_10419_),
    .B1(_10407_),
    .B2(\cpu.ex.r_13[3] ),
    .A2(_10189_),
    .A1(net1056));
 sg13g2_or2_1 _17311_ (.X(_10420_),
    .B(_10419_),
    .A(net1009));
 sg13g2_a21oi_1 _17312_ (.A1(_10418_),
    .A2(_10420_),
    .Y(_10421_),
    .B1(net739));
 sg13g2_or4_1 _17313_ (.A(_10398_),
    .B(_10404_),
    .C(_10415_),
    .D(_10421_),
    .X(_10422_));
 sg13g2_buf_1 _17314_ (.A(_10422_),
    .X(_10423_));
 sg13g2_buf_1 _17315_ (.A(_10130_),
    .X(_10424_));
 sg13g2_nor2_1 _17316_ (.A(_10201_),
    .B(_10203_),
    .Y(_10425_));
 sg13g2_nand3_1 _17317_ (.B(net1006),
    .C(_10425_),
    .A(_09050_),
    .Y(_10426_));
 sg13g2_buf_1 _17318_ (.A(\cpu.dec.imm[3] ),
    .X(_10427_));
 sg13g2_a21oi_1 _17319_ (.A1(_10427_),
    .A2(_10131_),
    .Y(_10428_),
    .B1(net1101));
 sg13g2_a22oi_1 _17320_ (.Y(_10429_),
    .B1(_10426_),
    .B2(_10428_),
    .A2(_00175_),
    .A1(net1101));
 sg13g2_a21oi_1 _17321_ (.A1(_10345_),
    .A2(_10423_),
    .Y(_10430_),
    .B1(_10429_));
 sg13g2_buf_1 _17322_ (.A(_10430_),
    .X(_10431_));
 sg13g2_a21o_1 _17323_ (.A2(_10337_),
    .A1(_10265_),
    .B1(net303),
    .X(_10432_));
 sg13g2_buf_8 _17324_ (.A(_10293_),
    .X(_10433_));
 sg13g2_nor2b_1 _17325_ (.A(_00238_),
    .B_N(net1007),
    .Y(_10434_));
 sg13g2_nor2b_1 _17326_ (.A(net1007),
    .B_N(_10093_),
    .Y(_10435_));
 sg13g2_a22oi_1 _17327_ (.Y(_10436_),
    .B1(_10435_),
    .B2(net747),
    .A2(_10434_),
    .A1(net736));
 sg13g2_nand4_1 _17328_ (.B(_10296_),
    .C(_10300_),
    .A(\cpu.ex.r_8[2] ),
    .Y(_10437_),
    .D(_10162_));
 sg13g2_o21ai_1 _17329_ (.B1(_10437_),
    .Y(_10438_),
    .A1(net738),
    .A2(_10436_));
 sg13g2_mux2_1 _17330_ (.A0(\cpu.ex.r_epc[2] ),
    .A1(\cpu.ex.r_11[2] ),
    .S(net1010),
    .X(_10439_));
 sg13g2_a22oi_1 _17331_ (.Y(_10440_),
    .B1(_10439_),
    .B2(_10173_),
    .A2(_10162_),
    .A1(\cpu.ex.r_9[2] ));
 sg13g2_nor2_1 _17332_ (.A(_10296_),
    .B(_10440_),
    .Y(_10441_));
 sg13g2_inv_1 _17333_ (.Y(_10442_),
    .A(\cpu.ex.r_10[2] ));
 sg13g2_nand3_1 _17334_ (.B(_10176_),
    .C(_10312_),
    .A(\cpu.ex.r_lr[2] ),
    .Y(_10443_));
 sg13g2_o21ai_1 _17335_ (.B1(_10443_),
    .Y(_10444_),
    .A1(_10442_),
    .A2(_10401_));
 sg13g2_nor4_2 _17336_ (.A(net744),
    .B(_10438_),
    .C(_10441_),
    .Y(_10445_),
    .D(_10444_));
 sg13g2_nand3_1 _17337_ (.B(net866),
    .C(_10312_),
    .A(_10079_),
    .Y(_10446_));
 sg13g2_mux2_1 _17338_ (.A0(\cpu.ex.r_stmp[2] ),
    .A1(\cpu.ex.r_14[2] ),
    .S(net865),
    .X(_10447_));
 sg13g2_nand2_1 _17339_ (.Y(_10448_),
    .A(_10400_),
    .B(_10447_));
 sg13g2_mux2_1 _17340_ (.A0(_08222_),
    .A1(\cpu.ex.r_12[2] ),
    .S(net1010),
    .X(_10449_));
 sg13g2_a21oi_1 _17341_ (.A1(_10145_),
    .A2(_10449_),
    .Y(_10450_),
    .B1(net739));
 sg13g2_nand3_1 _17342_ (.B(_10448_),
    .C(_10450_),
    .A(_10446_),
    .Y(_10451_));
 sg13g2_buf_1 _17343_ (.A(_10296_),
    .X(_10452_));
 sg13g2_a22oi_1 _17344_ (.Y(_10453_),
    .B1(_10309_),
    .B2(_10075_),
    .A2(_10162_),
    .A1(\cpu.ex.r_13[2] ));
 sg13g2_nor2_1 _17345_ (.A(_10452_),
    .B(_10453_),
    .Y(_10454_));
 sg13g2_nor3_1 _17346_ (.A(_10438_),
    .B(_10451_),
    .C(_10454_),
    .Y(_10455_));
 sg13g2_or3_1 _17347_ (.A(_10150_),
    .B(_10445_),
    .C(_10455_),
    .X(_10456_));
 sg13g2_nor3_1 _17348_ (.A(_09216_),
    .B(_10201_),
    .C(_10203_),
    .Y(_10457_));
 sg13g2_buf_1 _17349_ (.A(\cpu.dec.imm[2] ),
    .X(_10458_));
 sg13g2_nand3_1 _17350_ (.B(_10197_),
    .C(_10131_),
    .A(_10458_),
    .Y(_10459_));
 sg13g2_o21ai_1 _17351_ (.B1(_10459_),
    .Y(_10460_),
    .A1(_10197_),
    .A2(_00269_));
 sg13g2_a21oi_1 _17352_ (.A1(_10133_),
    .A2(_10457_),
    .Y(_10461_),
    .B1(_10460_));
 sg13g2_nand2_1 _17353_ (.Y(_10462_),
    .A(_10456_),
    .B(_10461_));
 sg13g2_buf_1 _17354_ (.A(_10462_),
    .X(_10463_));
 sg13g2_a221oi_1 _17355_ (.B2(_10352_),
    .C1(net371),
    .B1(_10354_),
    .A1(_10341_),
    .Y(_10464_),
    .A2(_10350_));
 sg13g2_nor2_1 _17356_ (.A(_10128_),
    .B(net371),
    .Y(_10465_));
 sg13g2_a221oi_1 _17357_ (.B2(_10464_),
    .C1(_10465_),
    .B1(_10432_),
    .A1(_10390_),
    .Y(_10466_),
    .A2(net372));
 sg13g2_nor2_1 _17358_ (.A(_10390_),
    .B(net372),
    .Y(_10467_));
 sg13g2_a21oi_2 _17359_ (.B1(_10467_),
    .Y(_10468_),
    .A2(_10466_),
    .A1(_10356_));
 sg13g2_buf_1 _17360_ (.A(_00276_),
    .X(_10469_));
 sg13g2_nand2b_1 _17361_ (.Y(_10470_),
    .B(_10120_),
    .A_N(_10469_));
 sg13g2_or3_1 _17362_ (.A(_08131_),
    .B(net460),
    .C(_10470_),
    .X(_10471_));
 sg13g2_buf_1 _17363_ (.A(_10471_),
    .X(_10472_));
 sg13g2_inv_2 _17364_ (.Y(_10473_),
    .A(_09781_));
 sg13g2_nand2_1 _17365_ (.Y(_10474_),
    .A(_10473_),
    .B(net594));
 sg13g2_nor2_1 _17366_ (.A(net1013),
    .B(_10060_),
    .Y(_10475_));
 sg13g2_and2_1 _17367_ (.A(net1013),
    .B(_10040_),
    .X(_10476_));
 sg13g2_buf_2 _17368_ (.A(_10476_),
    .X(_10477_));
 sg13g2_buf_1 _17369_ (.A(\cpu.ex.r_mult[21] ),
    .X(_10478_));
 sg13g2_a22oi_1 _17370_ (.Y(_10479_),
    .B1(_10477_),
    .B2(_10478_),
    .A2(_10475_),
    .A1(\cpu.ex.r_lr[5] ));
 sg13g2_nand3b_1 _17371_ (.B(net1014),
    .C(\cpu.ex.r_9[5] ),
    .Y(_10480_),
    .A_N(net1013));
 sg13g2_nand3b_1 _17372_ (.B(\cpu.ex.r_epc[5] ),
    .C(net1013),
    .Y(_10481_),
    .A_N(net1014));
 sg13g2_a21o_1 _17373_ (.A2(_10481_),
    .A1(_10480_),
    .B1(_10282_),
    .X(_10482_));
 sg13g2_o21ai_1 _17374_ (.B1(_10482_),
    .Y(_10483_),
    .A1(_10234_),
    .A2(_10479_));
 sg13g2_nand2_2 _17375_ (.Y(_10484_),
    .A(net874),
    .B(_10100_));
 sg13g2_buf_1 _17376_ (.A(\cpu.ex.r_sp[5] ),
    .X(_10485_));
 sg13g2_mux2_1 _17377_ (.A0(_10485_),
    .A1(\cpu.ex.r_10[5] ),
    .S(_10036_),
    .X(_10486_));
 sg13g2_a22oi_1 _17378_ (.Y(_10487_),
    .B1(_10486_),
    .B2(_10098_),
    .A2(_10058_),
    .A1(\cpu.ex.r_stmp[5] ));
 sg13g2_mux2_1 _17379_ (.A0(\cpu.ex.r_8[5] ),
    .A1(\cpu.ex.r_12[5] ),
    .S(net1011),
    .X(_10488_));
 sg13g2_nand3_1 _17380_ (.B(_10095_),
    .C(_10488_),
    .A(net870),
    .Y(_10489_));
 sg13g2_o21ai_1 _17381_ (.B1(_10489_),
    .Y(_10490_),
    .A1(_10484_),
    .A2(_10487_));
 sg13g2_nor2b_1 _17382_ (.A(_00241_),
    .B_N(net1012),
    .Y(_10491_));
 sg13g2_nor2b_1 _17383_ (.A(net1012),
    .B_N(\cpu.ex.r_14[5] ),
    .Y(_10492_));
 sg13g2_o21ai_1 _17384_ (.B1(_10477_),
    .Y(_10493_),
    .A1(_10491_),
    .A2(_10492_));
 sg13g2_and2_1 _17385_ (.A(net1011),
    .B(\cpu.ex.r_13[5] ),
    .X(_10494_));
 sg13g2_and2_1 _17386_ (.A(net874),
    .B(\cpu.ex.r_11[5] ),
    .X(_10495_));
 sg13g2_a22oi_1 _17387_ (.Y(_10496_),
    .B1(_10495_),
    .B2(_10219_),
    .A2(_10494_),
    .A1(_10244_));
 sg13g2_a21oi_1 _17388_ (.A1(_10493_),
    .A2(_10496_),
    .Y(_10497_),
    .B1(net748));
 sg13g2_or4_1 _17389_ (.A(net594),
    .B(_10483_),
    .C(_10490_),
    .D(_10497_),
    .X(_10498_));
 sg13g2_and2_1 _17390_ (.A(_10474_),
    .B(_10498_),
    .X(_10499_));
 sg13g2_and4_1 _17391_ (.A(_08220_),
    .B(_10115_),
    .C(_10474_),
    .D(_10498_),
    .X(_10500_));
 sg13g2_a21oi_1 _17392_ (.A1(_08220_),
    .A2(_10115_),
    .Y(_10501_),
    .B1(_10470_));
 sg13g2_a221oi_1 _17393_ (.B2(net460),
    .C1(_10501_),
    .B1(_10500_),
    .A1(_10123_),
    .Y(_10502_),
    .A2(_10499_));
 sg13g2_buf_2 _17394_ (.A(_10502_),
    .X(_10503_));
 sg13g2_nand2_1 _17395_ (.Y(_10504_),
    .A(_10472_),
    .B(_10503_));
 sg13g2_buf_1 _17396_ (.A(_10504_),
    .X(_10505_));
 sg13g2_buf_8 _17397_ (.A(_10178_),
    .X(_10506_));
 sg13g2_buf_1 _17398_ (.A(_10506_),
    .X(_10507_));
 sg13g2_buf_8 _17399_ (.A(net864),
    .X(_10508_));
 sg13g2_nand3_1 _17400_ (.B(_10508_),
    .C(net744),
    .A(net869),
    .Y(_10509_));
 sg13g2_mux2_1 _17401_ (.A0(\cpu.ex.r_8[5] ),
    .A1(\cpu.ex.r_12[5] ),
    .S(net868),
    .X(_10510_));
 sg13g2_buf_8 _17402_ (.A(net866),
    .X(_10511_));
 sg13g2_and2_1 _17403_ (.A(\cpu.ex.r_11[5] ),
    .B(net734),
    .X(_10512_));
 sg13g2_a22oi_1 _17404_ (.Y(_10513_),
    .B1(_10512_),
    .B2(_10393_),
    .A2(_10510_),
    .A1(_10145_));
 sg13g2_o21ai_1 _17405_ (.B1(_10513_),
    .Y(_10514_),
    .A1(_00241_),
    .A2(_10509_));
 sg13g2_inv_1 _17406_ (.Y(_10515_),
    .A(\cpu.ex.r_10[5] ));
 sg13g2_buf_8 _17407_ (.A(net734),
    .X(_10516_));
 sg13g2_nand3_1 _17408_ (.B(net658),
    .C(_10312_),
    .A(\cpu.ex.r_lr[5] ),
    .Y(_10517_));
 sg13g2_o21ai_1 _17409_ (.B1(_10517_),
    .Y(_10518_),
    .A1(_10515_),
    .A2(_10401_));
 sg13g2_buf_1 _17410_ (.A(_10301_),
    .X(_10519_));
 sg13g2_nand3b_1 _17411_ (.B(net869),
    .C(\cpu.ex.r_epc[5] ),
    .Y(_10520_),
    .A_N(_10169_));
 sg13g2_nand3b_1 _17412_ (.B(net744),
    .C(\cpu.ex.r_stmp[5] ),
    .Y(_10521_),
    .A_N(net869));
 sg13g2_nand2b_1 _17413_ (.Y(_10522_),
    .B(_10508_),
    .A_N(net745));
 sg13g2_a21oi_1 _17414_ (.A1(_10520_),
    .A2(_10521_),
    .Y(_10523_),
    .B1(_10522_));
 sg13g2_mux2_1 _17415_ (.A0(\cpu.ex.r_9[5] ),
    .A1(\cpu.ex.r_13[5] ),
    .S(net868),
    .X(_10524_));
 sg13g2_and3_1 _17416_ (.X(_10525_),
    .A(net734),
    .B(_10162_),
    .C(_10524_));
 sg13g2_and4_1 _17417_ (.A(_10485_),
    .B(net861),
    .C(net739),
    .D(_10309_),
    .X(_10526_));
 sg13g2_nand3b_1 _17418_ (.B(net734),
    .C(_10478_),
    .Y(_10527_),
    .A_N(net745));
 sg13g2_nand3b_1 _17419_ (.B(net745),
    .C(\cpu.ex.r_14[5] ),
    .Y(_10528_),
    .A_N(net869));
 sg13g2_nand2_1 _17420_ (.Y(_10529_),
    .A(net735),
    .B(net744));
 sg13g2_a21oi_1 _17421_ (.A1(_10527_),
    .A2(_10528_),
    .Y(_10530_),
    .B1(_10529_));
 sg13g2_or4_1 _17422_ (.A(_10523_),
    .B(_10525_),
    .C(_10526_),
    .D(_10530_),
    .X(_10531_));
 sg13g2_a221oi_1 _17423_ (.B2(net657),
    .C1(_10531_),
    .B1(_10518_),
    .A1(net593),
    .Y(_10532_),
    .A2(_10514_));
 sg13g2_buf_8 _17424_ (.A(_10425_),
    .X(_10533_));
 sg13g2_nand2_1 _17425_ (.Y(_10534_),
    .A(_09781_),
    .B(net526));
 sg13g2_o21ai_1 _17426_ (.B1(_10534_),
    .Y(_10535_),
    .A1(_10344_),
    .A2(_10532_));
 sg13g2_buf_2 _17427_ (.A(_10535_),
    .X(_10536_));
 sg13g2_nand2_1 _17428_ (.Y(_10537_),
    .A(\cpu.dec.imm[5] ),
    .B(_10207_));
 sg13g2_o21ai_1 _17429_ (.B1(_10537_),
    .Y(_10538_),
    .A1(_10197_),
    .A2(_10469_));
 sg13g2_a21o_1 _17430_ (.A2(_10536_),
    .A1(_10133_),
    .B1(_10538_),
    .X(_10539_));
 sg13g2_buf_1 _17431_ (.A(_10539_),
    .X(_10540_));
 sg13g2_buf_1 _17432_ (.A(_10540_),
    .X(_10541_));
 sg13g2_nand2_1 _17433_ (.Y(_10542_),
    .A(\cpu.ex.r_stmp[4] ),
    .B(_10189_));
 sg13g2_nor2b_1 _17434_ (.A(_00240_),
    .B_N(net865),
    .Y(_10543_));
 sg13g2_buf_1 _17435_ (.A(\cpu.ex.r_mult[20] ),
    .X(_10544_));
 sg13g2_nor2b_1 _17436_ (.A(net865),
    .B_N(_10544_),
    .Y(_10545_));
 sg13g2_o21ai_1 _17437_ (.B1(_10168_),
    .Y(_10546_),
    .A1(_10543_),
    .A2(_10545_));
 sg13g2_a21oi_1 _17438_ (.A1(_10542_),
    .A2(_10546_),
    .Y(_10547_),
    .B1(net738));
 sg13g2_and3_1 _17439_ (.X(_10548_),
    .A(\cpu.ex.r_12[4] ),
    .B(net738),
    .C(_10302_));
 sg13g2_buf_1 _17440_ (.A(_10194_),
    .X(_10549_));
 sg13g2_o21ai_1 _17441_ (.B1(_10549_),
    .Y(_10550_),
    .A1(_10547_),
    .A2(_10548_));
 sg13g2_nand3_1 _17442_ (.B(net861),
    .C(net736),
    .A(\cpu.ex.r_14[4] ),
    .Y(_10551_));
 sg13g2_nand3_1 _17443_ (.B(_10511_),
    .C(net747),
    .A(\cpu.ex.r_epc[4] ),
    .Y(_10552_));
 sg13g2_a21oi_1 _17444_ (.A1(_10551_),
    .A2(_10552_),
    .Y(_10553_),
    .B1(net738));
 sg13g2_nand3b_1 _17445_ (.B(net864),
    .C(\cpu.ex.r_11[4] ),
    .Y(_10554_),
    .A_N(net1008));
 sg13g2_nand3b_1 _17446_ (.B(net1008),
    .C(\cpu.ex.r_13[4] ),
    .Y(_10555_),
    .A_N(net864));
 sg13g2_nand2_1 _17447_ (.Y(_10556_),
    .A(net869),
    .B(net745));
 sg13g2_a21oi_1 _17448_ (.A1(_10554_),
    .A2(_10555_),
    .Y(_10557_),
    .B1(_10556_));
 sg13g2_buf_1 _17449_ (.A(\cpu.ex.r_sp[4] ),
    .X(_10558_));
 sg13g2_nand3b_1 _17450_ (.B(net864),
    .C(_10558_),
    .Y(_10559_),
    .A_N(net865));
 sg13g2_nand3b_1 _17451_ (.B(net865),
    .C(\cpu.ex.r_8[4] ),
    .Y(_10560_),
    .A_N(net864));
 sg13g2_a21oi_1 _17452_ (.A1(_10559_),
    .A2(_10560_),
    .Y(_10561_),
    .B1(_10167_));
 sg13g2_nand3b_1 _17453_ (.B(net868),
    .C(_08134_),
    .Y(_10562_),
    .A_N(net866));
 sg13g2_nand3b_1 _17454_ (.B(net866),
    .C(\cpu.ex.r_lr[4] ),
    .Y(_10563_),
    .A_N(net1008));
 sg13g2_or2_1 _17455_ (.X(_10564_),
    .B(net865),
    .A(net864));
 sg13g2_a21oi_1 _17456_ (.A1(_10562_),
    .A2(_10563_),
    .Y(_10565_),
    .B1(_10564_));
 sg13g2_nand3b_1 _17457_ (.B(net866),
    .C(\cpu.ex.r_9[4] ),
    .Y(_10566_),
    .A_N(net864));
 sg13g2_nand3b_1 _17458_ (.B(net867),
    .C(\cpu.ex.r_10[4] ),
    .Y(_10567_),
    .A_N(net866));
 sg13g2_a21oi_1 _17459_ (.A1(_10566_),
    .A2(_10567_),
    .Y(_10568_),
    .B1(_10412_));
 sg13g2_nor4_1 _17460_ (.A(_10557_),
    .B(_10561_),
    .C(_10565_),
    .D(_10568_),
    .Y(_10569_));
 sg13g2_nor2b_1 _17461_ (.A(_10553_),
    .B_N(_10569_),
    .Y(_10570_));
 sg13g2_a21oi_2 _17462_ (.B1(_10150_),
    .Y(_10571_),
    .A2(_10570_),
    .A1(_10550_));
 sg13g2_nand2_1 _17463_ (.Y(_10572_),
    .A(_09381_),
    .B(_10204_));
 sg13g2_a22oi_1 _17464_ (.Y(_10573_),
    .B1(\cpu.dec.imm[4] ),
    .B2(_10207_),
    .A2(_10129_),
    .A1(net1050));
 sg13g2_nand2_1 _17465_ (.Y(_10574_),
    .A(_10572_),
    .B(_10573_));
 sg13g2_or2_1 _17466_ (.X(_10575_),
    .B(_10574_),
    .A(_10571_));
 sg13g2_buf_2 _17467_ (.A(_10575_),
    .X(_10576_));
 sg13g2_nand2_1 _17468_ (.Y(_10577_),
    .A(net1050),
    .B(_10120_));
 sg13g2_or3_1 _17469_ (.A(_08131_),
    .B(net460),
    .C(_10577_),
    .X(_10578_));
 sg13g2_buf_1 _17470_ (.A(_10578_),
    .X(_10579_));
 sg13g2_nand2_1 _17471_ (.Y(_10580_),
    .A(_09173_),
    .B(net594));
 sg13g2_nand3_1 _17472_ (.B(net662),
    .C(_10062_),
    .A(\cpu.ex.r_10[4] ),
    .Y(_10581_));
 sg13g2_mux4_1 _17473_ (.S0(_10038_),
    .A0(_10558_),
    .A1(\cpu.ex.r_epc[4] ),
    .A2(\cpu.ex.r_stmp[4] ),
    .A3(_10544_),
    .S1(net1011),
    .X(_10582_));
 sg13g2_and2_1 _17474_ (.A(_10076_),
    .B(_10582_),
    .X(_10583_));
 sg13g2_nand3b_1 _17475_ (.B(\cpu.ex.r_lr[4] ),
    .C(net873),
    .Y(_10584_),
    .A_N(net872));
 sg13g2_nand3b_1 _17476_ (.B(net872),
    .C(_08134_),
    .Y(_10585_),
    .A_N(net1012));
 sg13g2_or2_1 _17477_ (.X(_10586_),
    .B(net871),
    .A(net874));
 sg13g2_a21oi_1 _17478_ (.A1(_10584_),
    .A2(_10585_),
    .Y(_10587_),
    .B1(_10586_));
 sg13g2_nand2_1 _17479_ (.Y(_10588_),
    .A(net873),
    .B(\cpu.ex.r_13[4] ));
 sg13g2_nand2b_1 _17480_ (.Y(_10589_),
    .B(\cpu.ex.r_12[4] ),
    .A_N(net873));
 sg13g2_nand3b_1 _17481_ (.B(net1014),
    .C(net1011),
    .Y(_10590_),
    .A_N(net1013));
 sg13g2_buf_1 _17482_ (.A(_10590_),
    .X(_10591_));
 sg13g2_a21oi_1 _17483_ (.A1(_10588_),
    .A2(_10589_),
    .Y(_10592_),
    .B1(_10591_));
 sg13g2_nand2b_1 _17484_ (.Y(_10593_),
    .B(net872),
    .A_N(_00240_));
 sg13g2_nand2b_1 _17485_ (.Y(_10594_),
    .B(\cpu.ex.r_11[4] ),
    .A_N(net872));
 sg13g2_nand3_1 _17486_ (.B(net873),
    .C(net871),
    .A(net874),
    .Y(_10595_));
 sg13g2_a21oi_1 _17487_ (.A1(_10593_),
    .A2(_10594_),
    .Y(_10596_),
    .B1(_10595_));
 sg13g2_nor4_1 _17488_ (.A(_10583_),
    .B(_10587_),
    .C(_10592_),
    .D(_10596_),
    .Y(_10597_));
 sg13g2_and3_1 _17489_ (.X(_10598_),
    .A(net863),
    .B(\cpu.ex.r_14[4] ),
    .C(_10228_));
 sg13g2_mux2_1 _17490_ (.A0(\cpu.ex.r_8[4] ),
    .A1(\cpu.ex.r_9[4] ),
    .S(_10053_),
    .X(_10599_));
 sg13g2_and3_1 _17491_ (.X(_10600_),
    .A(_10083_),
    .B(_10098_),
    .C(_10599_));
 sg13g2_buf_8 _17492_ (.A(_10214_),
    .X(_10601_));
 sg13g2_o21ai_1 _17493_ (.B1(net655),
    .Y(_10602_),
    .A1(_10598_),
    .A2(_10600_));
 sg13g2_nand4_1 _17494_ (.B(_10581_),
    .C(_10597_),
    .A(_10046_),
    .Y(_10603_),
    .D(_10602_));
 sg13g2_and2_1 _17495_ (.A(_10580_),
    .B(_10603_),
    .X(_10604_));
 sg13g2_buf_1 _17496_ (.A(_10604_),
    .X(_10605_));
 sg13g2_and4_1 _17497_ (.A(_08220_),
    .B(_10115_),
    .C(_10580_),
    .D(_10603_),
    .X(_10606_));
 sg13g2_a21oi_1 _17498_ (.A1(_08220_),
    .A2(_10115_),
    .Y(_10607_),
    .B1(_10577_));
 sg13g2_a221oi_1 _17499_ (.B2(net460),
    .C1(_10607_),
    .B1(_10606_),
    .A1(_10123_),
    .Y(_10608_),
    .A2(_10605_));
 sg13g2_buf_1 _17500_ (.A(_10608_),
    .X(_10609_));
 sg13g2_nand2_1 _17501_ (.Y(_10610_),
    .A(_10579_),
    .B(_10609_));
 sg13g2_buf_1 _17502_ (.A(_10610_),
    .X(_10611_));
 sg13g2_a22oi_1 _17503_ (.Y(_10612_),
    .B1(_10576_),
    .B2(net229),
    .A2(net230),
    .A1(_10505_));
 sg13g2_buf_1 _17504_ (.A(_10612_),
    .X(_10613_));
 sg13g2_nand2b_1 _17505_ (.Y(_10614_),
    .B(net735),
    .A_N(_00244_));
 sg13g2_nand2b_1 _17506_ (.Y(_10615_),
    .B(\cpu.ex.r_13[8] ),
    .A_N(net735));
 sg13g2_nand2_1 _17507_ (.Y(_10616_),
    .A(net659),
    .B(_10194_));
 sg13g2_a21oi_1 _17508_ (.A1(_10614_),
    .A2(_10615_),
    .Y(_10617_),
    .B1(_10616_));
 sg13g2_mux2_1 _17509_ (.A0(\cpu.ex.r_lr[8] ),
    .A1(\cpu.ex.r_epc[8] ),
    .S(net735),
    .X(_10618_));
 sg13g2_and2_1 _17510_ (.A(net747),
    .B(_10618_),
    .X(_10619_));
 sg13g2_buf_1 _17511_ (.A(net734),
    .X(_10620_));
 sg13g2_o21ai_1 _17512_ (.B1(_10620_),
    .Y(_10621_),
    .A1(_10617_),
    .A2(_10619_));
 sg13g2_and3_1 _17513_ (.X(_10622_),
    .A(\cpu.ex.r_stmp[8] ),
    .B(net861),
    .C(_10155_));
 sg13g2_and3_1 _17514_ (.X(_10623_),
    .A(\cpu.ex.r_11[8] ),
    .B(net658),
    .C(net746));
 sg13g2_buf_1 _17515_ (.A(net735),
    .X(_10624_));
 sg13g2_buf_1 _17516_ (.A(net653),
    .X(_10625_));
 sg13g2_o21ai_1 _17517_ (.B1(net592),
    .Y(_10626_),
    .A1(_10622_),
    .A2(_10623_));
 sg13g2_buf_1 _17518_ (.A(\cpu.ex.r_mult[24] ),
    .X(_10627_));
 sg13g2_mux2_1 _17519_ (.A0(\cpu.ex.r_12[8] ),
    .A1(\cpu.ex.r_14[8] ),
    .S(net653),
    .X(_10628_));
 sg13g2_nor2_2 _17520_ (.A(net658),
    .B(_10616_),
    .Y(_10629_));
 sg13g2_a22oi_1 _17521_ (.Y(_10630_),
    .B1(_10628_),
    .B2(_10629_),
    .A2(_10409_),
    .A1(_10627_));
 sg13g2_buf_1 _17522_ (.A(\cpu.ex.r_sp[8] ),
    .X(_10631_));
 sg13g2_nand3b_1 _17523_ (.B(net653),
    .C(_10631_),
    .Y(_10632_),
    .A_N(net659));
 sg13g2_nand3b_1 _17524_ (.B(net659),
    .C(\cpu.ex.r_8[8] ),
    .Y(_10633_),
    .A_N(net735));
 sg13g2_a21oi_1 _17525_ (.A1(_10632_),
    .A2(_10633_),
    .Y(_10634_),
    .B1(_10167_));
 sg13g2_nand3b_1 _17526_ (.B(net658),
    .C(\cpu.ex.r_9[8] ),
    .Y(_10635_),
    .A_N(net735));
 sg13g2_nand3b_1 _17527_ (.B(net653),
    .C(\cpu.ex.r_10[8] ),
    .Y(_10636_),
    .A_N(net734));
 sg13g2_a21oi_1 _17528_ (.A1(_10635_),
    .A2(_10636_),
    .Y(_10637_),
    .B1(_10412_));
 sg13g2_nor2_1 _17529_ (.A(_10634_),
    .B(_10637_),
    .Y(_10638_));
 sg13g2_nand4_1 _17530_ (.B(_10626_),
    .C(_10630_),
    .A(_10621_),
    .Y(_10639_),
    .D(_10638_));
 sg13g2_a221oi_1 _17531_ (.B2(_10639_),
    .C1(_10131_),
    .B1(_10149_),
    .A1(_09024_),
    .Y(_10640_),
    .A2(net526));
 sg13g2_o21ai_1 _17532_ (.B1(_10197_),
    .Y(_10641_),
    .A1(net1006),
    .A2(\cpu.dec.imm[8] ));
 sg13g2_buf_1 _17533_ (.A(net1101),
    .X(_10642_));
 sg13g2_inv_2 _17534_ (.Y(_10643_),
    .A(_00268_));
 sg13g2_nand2_1 _17535_ (.Y(_10644_),
    .A(net1005),
    .B(_10643_));
 sg13g2_o21ai_1 _17536_ (.B1(_10644_),
    .Y(_10645_),
    .A1(_10640_),
    .A2(_10641_));
 sg13g2_buf_2 _17537_ (.A(_10645_),
    .X(_10646_));
 sg13g2_nand2b_1 _17538_ (.Y(_10647_),
    .B(net862),
    .A_N(_00244_));
 sg13g2_nand2b_1 _17539_ (.Y(_10648_),
    .B(\cpu.ex.r_14[8] ),
    .A_N(net862));
 sg13g2_nand3_1 _17540_ (.B(net742),
    .C(net863),
    .A(net752),
    .Y(_10649_));
 sg13g2_a21o_1 _17541_ (.A2(_10648_),
    .A1(_10647_),
    .B1(_10649_),
    .X(_10650_));
 sg13g2_nand3_1 _17542_ (.B(net668),
    .C(net661),
    .A(\cpu.ex.r_9[8] ),
    .Y(_10651_));
 sg13g2_mux2_1 _17543_ (.A0(\cpu.ex.r_8[8] ),
    .A1(\cpu.ex.r_12[8] ),
    .S(net863),
    .X(_10652_));
 sg13g2_nand3_1 _17544_ (.B(_10095_),
    .C(_10652_),
    .A(net870),
    .Y(_10653_));
 sg13g2_nand3_1 _17545_ (.B(_10651_),
    .C(_10653_),
    .A(_10650_),
    .Y(_10654_));
 sg13g2_nand2_1 _17546_ (.Y(_10655_),
    .A(_10272_),
    .B(_10266_));
 sg13g2_a22oi_1 _17547_ (.Y(_10656_),
    .B1(net665),
    .B2(\cpu.ex.r_13[8] ),
    .A2(net667),
    .A1(\cpu.ex.r_mult[24] ));
 sg13g2_nor2_1 _17548_ (.A(_10655_),
    .B(_10656_),
    .Y(_10657_));
 sg13g2_mux2_1 _17549_ (.A0(\cpu.ex.r_epc[8] ),
    .A1(\cpu.ex.r_11[8] ),
    .S(net742),
    .X(_10658_));
 sg13g2_a22oi_1 _17550_ (.Y(_10659_),
    .B1(_10658_),
    .B2(net671),
    .A2(_10215_),
    .A1(\cpu.ex.r_lr[8] ));
 sg13g2_nor2_1 _17551_ (.A(_10282_),
    .B(_10659_),
    .Y(_10660_));
 sg13g2_mux2_1 _17552_ (.A0(_10631_),
    .A1(\cpu.ex.r_stmp[8] ),
    .S(net750),
    .X(_10661_));
 sg13g2_a22oi_1 _17553_ (.Y(_10662_),
    .B1(_10661_),
    .B2(net748),
    .A2(net668),
    .A1(\cpu.ex.r_10[8] ));
 sg13g2_nor2_1 _17554_ (.A(_10484_),
    .B(_10662_),
    .Y(_10663_));
 sg13g2_nor4_1 _17555_ (.A(_10654_),
    .B(_10657_),
    .C(_10660_),
    .D(_10663_),
    .Y(_10664_));
 sg13g2_nor2_1 _17556_ (.A(_09024_),
    .B(net596),
    .Y(_10665_));
 sg13g2_a21o_1 _17557_ (.A2(_10664_),
    .A1(net596),
    .B1(_10665_),
    .X(_10666_));
 sg13g2_buf_1 _17558_ (.A(_10666_),
    .X(_10667_));
 sg13g2_mux2_1 _17559_ (.A0(_00268_),
    .A1(_10667_),
    .S(net251),
    .X(_10668_));
 sg13g2_buf_1 _17560_ (.A(_10668_),
    .X(_10669_));
 sg13g2_nand2_1 _17561_ (.Y(_10670_),
    .A(_10646_),
    .B(_10669_));
 sg13g2_buf_2 _17562_ (.A(_10670_),
    .X(_10671_));
 sg13g2_nor2_1 _17563_ (.A(_10640_),
    .B(_10641_),
    .Y(_10672_));
 sg13g2_a21oi_1 _17564_ (.A1(_10642_),
    .A2(_10643_),
    .Y(_10673_),
    .B1(_10672_));
 sg13g2_buf_2 _17565_ (.A(_10673_),
    .X(_10674_));
 sg13g2_inv_1 _17566_ (.Y(_10675_),
    .A(_10667_));
 sg13g2_buf_8 _17567_ (.A(_10125_),
    .X(_10676_));
 sg13g2_mux2_1 _17568_ (.A0(_10643_),
    .A1(_10675_),
    .S(_10676_),
    .X(_10677_));
 sg13g2_buf_2 _17569_ (.A(_10677_),
    .X(_10678_));
 sg13g2_nand2_1 _17570_ (.Y(_10679_),
    .A(_10674_),
    .B(_10678_));
 sg13g2_nand2_1 _17571_ (.Y(_10680_),
    .A(_10671_),
    .B(_10679_));
 sg13g2_nand2_1 _17572_ (.Y(_10681_),
    .A(_09023_),
    .B(_10533_));
 sg13g2_and2_1 _17573_ (.A(net746),
    .B(_10400_),
    .X(_10682_));
 sg13g2_inv_1 _17574_ (.Y(_10683_),
    .A(\cpu.ex.r_9[6] ));
 sg13g2_nand2_1 _17575_ (.Y(_10684_),
    .A(\cpu.ex.r_13[6] ),
    .B(net744));
 sg13g2_o21ai_1 _17576_ (.B1(_10684_),
    .Y(_10685_),
    .A1(_10683_),
    .A2(net744));
 sg13g2_and2_1 _17577_ (.A(_10511_),
    .B(net663),
    .X(_10686_));
 sg13g2_a22oi_1 _17578_ (.Y(_10687_),
    .B1(_10685_),
    .B2(_10686_),
    .A2(_10682_),
    .A1(\cpu.ex.r_10[6] ));
 sg13g2_nor2_1 _17579_ (.A(net861),
    .B(net659),
    .Y(_10688_));
 sg13g2_and3_1 _17580_ (.X(_10689_),
    .A(\cpu.ex.r_mult[22] ),
    .B(net867),
    .C(net868));
 sg13g2_a21o_1 _17581_ (.A2(_10316_),
    .A1(\cpu.ex.r_lr[6] ),
    .B1(_10689_),
    .X(_10690_));
 sg13g2_inv_1 _17582_ (.Y(_10691_),
    .A(\cpu.ex.r_12[6] ));
 sg13g2_or2_1 _17583_ (.X(_10692_),
    .B(net867),
    .A(_10168_));
 sg13g2_nand3b_1 _17584_ (.B(net869),
    .C(net867),
    .Y(_10693_),
    .A_N(_00242_));
 sg13g2_o21ai_1 _17585_ (.B1(_10693_),
    .Y(_10694_),
    .A1(_10691_),
    .A2(_10692_));
 sg13g2_buf_1 _17586_ (.A(\cpu.ex.r_sp[6] ),
    .X(_10695_));
 sg13g2_nand3b_1 _17587_ (.B(net735),
    .C(_10695_),
    .Y(_10696_),
    .A_N(net745));
 sg13g2_nand3b_1 _17588_ (.B(net745),
    .C(\cpu.ex.r_8[6] ),
    .Y(_10697_),
    .A_N(net867));
 sg13g2_a21oi_1 _17589_ (.A1(_10696_),
    .A2(_10697_),
    .Y(_10698_),
    .B1(_10167_));
 sg13g2_a221oi_1 _17590_ (.B2(net736),
    .C1(_10698_),
    .B1(_10694_),
    .A1(_10688_),
    .Y(_10699_),
    .A2(_10690_));
 sg13g2_a21o_1 _17591_ (.A2(_10699_),
    .A1(_10687_),
    .B1(_10344_),
    .X(_10700_));
 sg13g2_nand3_1 _17592_ (.B(net734),
    .C(net746),
    .A(\cpu.ex.r_11[6] ),
    .Y(_10701_));
 sg13g2_nand3_1 _17593_ (.B(net861),
    .C(_10155_),
    .A(\cpu.ex.r_stmp[6] ),
    .Y(_10702_));
 sg13g2_nand3_1 _17594_ (.B(net861),
    .C(net736),
    .A(\cpu.ex.r_14[6] ),
    .Y(_10703_));
 sg13g2_nand3_1 _17595_ (.B(net734),
    .C(net747),
    .A(\cpu.ex.r_epc[6] ),
    .Y(_10704_));
 sg13g2_nand4_1 _17596_ (.B(_10702_),
    .C(_10703_),
    .A(_10701_),
    .Y(_10705_),
    .D(_10704_));
 sg13g2_nand3_1 _17597_ (.B(_10149_),
    .C(_10705_),
    .A(net592),
    .Y(_10706_));
 sg13g2_nand3_1 _17598_ (.B(_10700_),
    .C(_10706_),
    .A(_10681_),
    .Y(_10707_));
 sg13g2_buf_2 _17599_ (.A(_10707_),
    .X(_10708_));
 sg13g2_nor2_1 _17600_ (.A(net743),
    .B(_10708_),
    .Y(_10709_));
 sg13g2_buf_2 _17601_ (.A(_00275_),
    .X(_10710_));
 sg13g2_nor3_1 _17602_ (.A(_10129_),
    .B(net1006),
    .C(\cpu.dec.imm[6] ),
    .Y(_10711_));
 sg13g2_a21oi_1 _17603_ (.A1(net1005),
    .A2(_10710_),
    .Y(_10712_),
    .B1(_10711_));
 sg13g2_nor2b_1 _17604_ (.A(_10709_),
    .B_N(_10712_),
    .Y(_10713_));
 sg13g2_buf_1 _17605_ (.A(_10713_),
    .X(_10714_));
 sg13g2_inv_1 _17606_ (.Y(_10715_),
    .A(_00242_));
 sg13g2_a22oi_1 _17607_ (.Y(_10716_),
    .B1(_10477_),
    .B2(_10715_),
    .A2(_10475_),
    .A1(\cpu.ex.r_9[6] ));
 sg13g2_nand2b_1 _17608_ (.Y(_10717_),
    .B(_10071_),
    .A_N(_10716_));
 sg13g2_mux2_1 _17609_ (.A0(\cpu.ex.r_8[6] ),
    .A1(\cpu.ex.r_12[6] ),
    .S(net863),
    .X(_10718_));
 sg13g2_nand3_1 _17610_ (.B(net665),
    .C(_10718_),
    .A(net870),
    .Y(_10719_));
 sg13g2_nand3_1 _17611_ (.B(net662),
    .C(_10058_),
    .A(\cpu.ex.r_stmp[6] ),
    .Y(_10720_));
 sg13g2_and4_1 _17612_ (.A(_10046_),
    .B(_10717_),
    .C(_10719_),
    .D(_10720_),
    .X(_10721_));
 sg13g2_nand2_1 _17613_ (.Y(_10722_),
    .A(net748),
    .B(_10098_));
 sg13g2_a22oi_1 _17614_ (.Y(_10723_),
    .B1(net661),
    .B2(\cpu.ex.r_lr[6] ),
    .A2(net662),
    .A1(_10695_));
 sg13g2_nor2_1 _17615_ (.A(_10722_),
    .B(_10723_),
    .Y(_10724_));
 sg13g2_buf_1 _17616_ (.A(\cpu.ex.r_mult[22] ),
    .X(_10725_));
 sg13g2_a22oi_1 _17617_ (.Y(_10726_),
    .B1(_10062_),
    .B2(\cpu.ex.r_11[6] ),
    .A2(_10058_),
    .A1(_10725_));
 sg13g2_nor2_1 _17618_ (.A(_10371_),
    .B(_10726_),
    .Y(_10727_));
 sg13g2_mux2_1 _17619_ (.A0(\cpu.ex.r_10[6] ),
    .A1(\cpu.ex.r_14[6] ),
    .S(net863),
    .X(_10728_));
 sg13g2_nand3_1 _17620_ (.B(net662),
    .C(_10728_),
    .A(net655),
    .Y(_10729_));
 sg13g2_nand3_1 _17621_ (.B(net661),
    .C(_10222_),
    .A(\cpu.ex.r_13[6] ),
    .Y(_10730_));
 sg13g2_nand3_1 _17622_ (.B(_10361_),
    .C(_10278_),
    .A(\cpu.ex.r_epc[6] ),
    .Y(_10731_));
 sg13g2_nand3_1 _17623_ (.B(_10730_),
    .C(_10731_),
    .A(_10729_),
    .Y(_10732_));
 sg13g2_nor3_1 _17624_ (.A(_10724_),
    .B(_10727_),
    .C(_10732_),
    .Y(_10733_));
 sg13g2_nor2_1 _17625_ (.A(_09023_),
    .B(_10046_),
    .Y(_10734_));
 sg13g2_a21o_1 _17626_ (.A2(_10733_),
    .A1(_10721_),
    .B1(_10734_),
    .X(_10735_));
 sg13g2_buf_1 _17627_ (.A(_10735_),
    .X(_10736_));
 sg13g2_mux2_1 _17628_ (.A0(_10710_),
    .A1(_10736_),
    .S(net251),
    .X(_10737_));
 sg13g2_buf_1 _17629_ (.A(_10737_),
    .X(_10738_));
 sg13g2_xnor2_1 _17630_ (.Y(_10739_),
    .A(_10714_),
    .B(_10738_));
 sg13g2_buf_2 _17631_ (.A(_00274_),
    .X(_10740_));
 sg13g2_inv_1 _17632_ (.Y(_10741_),
    .A(_10740_));
 sg13g2_nand3_1 _17633_ (.B(\cpu.ex.r_9[7] ),
    .C(_10095_),
    .A(net664),
    .Y(_10742_));
 sg13g2_buf_1 _17634_ (.A(\cpu.ex.r_mult[23] ),
    .X(_10743_));
 sg13g2_nand3_1 _17635_ (.B(_10743_),
    .C(_10058_),
    .A(net752),
    .Y(_10744_));
 sg13g2_a21oi_1 _17636_ (.A1(_10742_),
    .A2(_10744_),
    .Y(_10745_),
    .B1(net870));
 sg13g2_nand2_1 _17637_ (.Y(_10746_),
    .A(net671),
    .B(net655));
 sg13g2_inv_1 _17638_ (.Y(_10747_),
    .A(_00243_));
 sg13g2_a22oi_1 _17639_ (.Y(_10748_),
    .B1(_10251_),
    .B2(_10747_),
    .A2(_10249_),
    .A1(\cpu.ex.r_10[7] ));
 sg13g2_nor2_1 _17640_ (.A(_10746_),
    .B(_10748_),
    .Y(_10749_));
 sg13g2_a22oi_1 _17641_ (.Y(_10750_),
    .B1(_10095_),
    .B2(\cpu.ex.r_12[7] ),
    .A2(net667),
    .A1(\cpu.ex.r_stmp[7] ));
 sg13g2_nor2b_1 _17642_ (.A(_10750_),
    .B_N(_10375_),
    .Y(_10751_));
 sg13g2_nor3_1 _17643_ (.A(_10745_),
    .B(_10749_),
    .C(_10751_),
    .Y(_10752_));
 sg13g2_buf_1 _17644_ (.A(\cpu.dec.user_io ),
    .X(_10753_));
 sg13g2_and3_1 _17645_ (.X(_10754_),
    .A(net666),
    .B(_10753_),
    .C(_10375_));
 sg13g2_buf_1 _17646_ (.A(\cpu.ex.r_sp[7] ),
    .X(_10755_));
 sg13g2_a22oi_1 _17647_ (.Y(_10756_),
    .B1(net661),
    .B2(\cpu.ex.r_lr[7] ),
    .A2(_10228_),
    .A1(_10755_));
 sg13g2_nand2_1 _17648_ (.Y(_10757_),
    .A(\cpu.ex.r_epc[7] ),
    .B(_10278_));
 sg13g2_a21oi_1 _17649_ (.A1(_10756_),
    .A2(_10757_),
    .Y(_10758_),
    .B1(net741));
 sg13g2_o21ai_1 _17650_ (.B1(net748),
    .Y(_10759_),
    .A1(_10754_),
    .A2(_10758_));
 sg13g2_nor2b_1 _17651_ (.A(_10224_),
    .B_N(_10049_),
    .Y(_10760_));
 sg13g2_a22oi_1 _17652_ (.Y(_10761_),
    .B1(_10760_),
    .B2(\cpu.ex.r_11[7] ),
    .A2(_10231_),
    .A1(\cpu.ex.r_13[7] ));
 sg13g2_a221oi_1 _17653_ (.B2(\cpu.ex.r_14[7] ),
    .C1(net751),
    .B1(_10477_),
    .A1(\cpu.ex.r_8[7] ),
    .Y(_10762_),
    .A2(_10475_));
 sg13g2_a21oi_1 _17654_ (.A1(net740),
    .A2(_10761_),
    .Y(_10763_),
    .B1(_10762_));
 sg13g2_nand2_1 _17655_ (.Y(_10764_),
    .A(net660),
    .B(_10763_));
 sg13g2_nand3_1 _17656_ (.B(_10759_),
    .C(_10764_),
    .A(_10752_),
    .Y(_10765_));
 sg13g2_mux2_1 _17657_ (.A0(_09026_),
    .A1(_10765_),
    .S(net596),
    .X(_10766_));
 sg13g2_buf_1 _17658_ (.A(_10766_),
    .X(_10767_));
 sg13g2_mux2_1 _17659_ (.A0(_10741_),
    .A1(_10767_),
    .S(net251),
    .X(_10768_));
 sg13g2_buf_1 _17660_ (.A(_10768_),
    .X(_10769_));
 sg13g2_inv_1 _17661_ (.Y(_10770_),
    .A(net207));
 sg13g2_buf_1 _17662_ (.A(_10452_),
    .X(_10771_));
 sg13g2_mux2_1 _17663_ (.A0(_10755_),
    .A1(\cpu.ex.r_stmp[7] ),
    .S(net656),
    .X(_10772_));
 sg13g2_a22oi_1 _17664_ (.Y(_10773_),
    .B1(_10772_),
    .B2(net737),
    .A2(net746),
    .A1(\cpu.ex.r_10[7] ));
 sg13g2_nand3_1 _17665_ (.B(net738),
    .C(net736),
    .A(\cpu.ex.r_12[7] ),
    .Y(_10774_));
 sg13g2_o21ai_1 _17666_ (.B1(_10774_),
    .Y(_10775_),
    .A1(net738),
    .A2(_10773_));
 sg13g2_and2_1 _17667_ (.A(net733),
    .B(_10775_),
    .X(_10776_));
 sg13g2_a22oi_1 _17668_ (.Y(_10777_),
    .B1(net736),
    .B2(_10747_),
    .A2(net747),
    .A1(\cpu.ex.r_epc[7] ));
 sg13g2_or2_1 _17669_ (.X(_10778_),
    .B(_10777_),
    .A(_10152_));
 sg13g2_mux2_1 _17670_ (.A0(\cpu.ex.r_8[7] ),
    .A1(\cpu.ex.r_9[7] ),
    .S(_10516_),
    .X(_10779_));
 sg13g2_and2_1 _17671_ (.A(\cpu.ex.r_11[7] ),
    .B(net654),
    .X(_10780_));
 sg13g2_and2_1 _17672_ (.A(net657),
    .B(_10192_),
    .X(_10781_));
 sg13g2_and4_1 _17673_ (.A(\cpu.ex.r_13[7] ),
    .B(net654),
    .C(net656),
    .D(net663),
    .X(_10782_));
 sg13g2_a221oi_1 _17674_ (.B2(_10781_),
    .C1(_10782_),
    .B1(_10780_),
    .A1(_10413_),
    .Y(_10783_),
    .A2(_10779_));
 sg13g2_inv_1 _17675_ (.Y(_10784_),
    .A(\cpu.ex.r_14[7] ));
 sg13g2_nand3b_1 _17676_ (.B(_10620_),
    .C(_10743_),
    .Y(_10785_),
    .A_N(_10506_));
 sg13g2_o21ai_1 _17677_ (.B1(_10785_),
    .Y(_10786_),
    .A1(_10784_),
    .A2(_10179_));
 sg13g2_inv_1 _17678_ (.Y(_10787_),
    .A(\cpu.ex.r_lr[7] ));
 sg13g2_nand3b_1 _17679_ (.B(net656),
    .C(_10753_),
    .Y(_10788_),
    .A_N(net658));
 sg13g2_o21ai_1 _17680_ (.B1(_10788_),
    .Y(_10789_),
    .A1(_10787_),
    .A2(_10184_));
 sg13g2_a22oi_1 _17681_ (.Y(_10790_),
    .B1(_10789_),
    .B2(_10312_),
    .A2(_10786_),
    .A1(_10320_));
 sg13g2_nand3_1 _17682_ (.B(_10783_),
    .C(_10790_),
    .A(_10778_),
    .Y(_10791_));
 sg13g2_buf_1 _17683_ (.A(_10149_),
    .X(_10792_));
 sg13g2_o21ai_1 _17684_ (.B1(net525),
    .Y(_10793_),
    .A1(_10776_),
    .A2(_10791_));
 sg13g2_a21oi_1 _17685_ (.A1(_09026_),
    .A2(net526),
    .Y(_10794_),
    .B1(net743));
 sg13g2_buf_1 _17686_ (.A(_10197_),
    .X(_10795_));
 sg13g2_nand2b_1 _17687_ (.Y(_10796_),
    .B(_10207_),
    .A_N(\cpu.dec.imm[7] ));
 sg13g2_o21ai_1 _17688_ (.B1(_10796_),
    .Y(_10797_),
    .A1(_10795_),
    .A2(_10741_));
 sg13g2_a21o_1 _17689_ (.A2(_10794_),
    .A1(_10793_),
    .B1(_10797_),
    .X(_10798_));
 sg13g2_buf_1 _17690_ (.A(_10798_),
    .X(_10799_));
 sg13g2_buf_1 _17691_ (.A(_10799_),
    .X(_10800_));
 sg13g2_nand2_1 _17692_ (.Y(_10801_),
    .A(_10770_),
    .B(net228));
 sg13g2_nand2_1 _17693_ (.Y(_10802_),
    .A(_10505_),
    .B(net230));
 sg13g2_nor2_1 _17694_ (.A(_10576_),
    .B(_10610_),
    .Y(_10803_));
 sg13g2_nor2_1 _17695_ (.A(_10505_),
    .B(net230),
    .Y(_10804_));
 sg13g2_a21oi_1 _17696_ (.A1(_10802_),
    .A2(_10803_),
    .Y(_10805_),
    .B1(_10804_));
 sg13g2_nand4_1 _17697_ (.B(_10739_),
    .C(_10801_),
    .A(_10680_),
    .Y(_10806_),
    .D(_10805_));
 sg13g2_a21oi_1 _17698_ (.A1(_10468_),
    .A2(_10613_),
    .Y(_10807_),
    .B1(_10806_));
 sg13g2_o21ai_1 _17699_ (.B1(_10712_),
    .Y(_10808_),
    .A1(net743),
    .A2(_10708_));
 sg13g2_buf_2 _17700_ (.A(_10808_),
    .X(_10809_));
 sg13g2_nor4_1 _17701_ (.A(_10674_),
    .B(_10809_),
    .C(_10799_),
    .D(_10738_),
    .Y(_10810_));
 sg13g2_a21oi_1 _17702_ (.A1(_10793_),
    .A2(_10794_),
    .Y(_10811_),
    .B1(_10797_));
 sg13g2_buf_1 _17703_ (.A(_10811_),
    .X(_10812_));
 sg13g2_and3_1 _17704_ (.X(_10813_),
    .A(net207),
    .B(_10646_),
    .C(net249));
 sg13g2_inv_1 _17705_ (.Y(_10814_),
    .A(_10710_));
 sg13g2_inv_1 _17706_ (.Y(_10815_),
    .A(_10736_));
 sg13g2_mux2_1 _17707_ (.A0(_10814_),
    .A1(_10815_),
    .S(net251),
    .X(_10816_));
 sg13g2_buf_1 _17708_ (.A(_10816_),
    .X(_10817_));
 sg13g2_and4_1 _17709_ (.A(net207),
    .B(_10646_),
    .C(_10714_),
    .D(net206),
    .X(_10818_));
 sg13g2_or4_1 _17710_ (.A(_10678_),
    .B(_10810_),
    .C(_10813_),
    .D(_10818_),
    .X(_10819_));
 sg13g2_buf_1 _17711_ (.A(_10674_),
    .X(_10820_));
 sg13g2_nor3_1 _17712_ (.A(_10740_),
    .B(_10710_),
    .C(_10809_),
    .Y(_10821_));
 sg13g2_nor2_1 _17713_ (.A(_10710_),
    .B(_10711_),
    .Y(_10822_));
 sg13g2_o21ai_1 _17714_ (.B1(_10822_),
    .Y(_10823_),
    .A1(net743),
    .A2(_10708_));
 sg13g2_a21oi_1 _17715_ (.A1(_10740_),
    .A2(_10823_),
    .Y(_10824_),
    .B1(_10799_));
 sg13g2_o21ai_1 _17716_ (.B1(net303),
    .Y(_10825_),
    .A1(_10821_),
    .A2(_10824_));
 sg13g2_buf_1 _17717_ (.A(net250),
    .X(_10826_));
 sg13g2_nand3_1 _17718_ (.B(_10767_),
    .C(net249),
    .A(net227),
    .Y(_10827_));
 sg13g2_nor3_1 _17719_ (.A(net303),
    .B(_10736_),
    .C(_10809_),
    .Y(_10828_));
 sg13g2_o21ai_1 _17720_ (.B1(_10828_),
    .Y(_10829_),
    .A1(_10767_),
    .A2(net249));
 sg13g2_nand4_1 _17721_ (.B(_10825_),
    .C(_10827_),
    .A(net205),
    .Y(_10830_),
    .D(_10829_));
 sg13g2_buf_2 _17722_ (.A(\cpu.addr[9] ),
    .X(_10831_));
 sg13g2_nand2b_1 _17723_ (.Y(_10832_),
    .B(_10213_),
    .A_N(_10831_));
 sg13g2_nand2_1 _17724_ (.Y(_10833_),
    .A(\cpu.ex.r_epc[9] ),
    .B(_10361_));
 sg13g2_nor2b_1 _17725_ (.A(_00245_),
    .B_N(net742),
    .Y(_10834_));
 sg13g2_buf_2 _17726_ (.A(\cpu.ex.r_mult[25] ),
    .X(_10835_));
 sg13g2_nor2b_1 _17727_ (.A(net742),
    .B_N(_10835_),
    .Y(_10836_));
 sg13g2_o21ai_1 _17728_ (.B1(net741),
    .Y(_10837_),
    .A1(_10834_),
    .A2(_10836_));
 sg13g2_a21oi_1 _17729_ (.A1(_10833_),
    .A2(_10837_),
    .Y(_10838_),
    .B1(net870));
 sg13g2_buf_1 _17730_ (.A(\cpu.ex.r_sp[9] ),
    .X(_10839_));
 sg13g2_and3_1 _17731_ (.X(_10840_),
    .A(net748),
    .B(_10839_),
    .C(_10249_));
 sg13g2_o21ai_1 _17732_ (.B1(net595),
    .Y(_10841_),
    .A1(_10838_),
    .A2(_10840_));
 sg13g2_a22oi_1 _17733_ (.Y(_10842_),
    .B1(_10062_),
    .B2(\cpu.ex.r_10[9] ),
    .A2(_10058_),
    .A1(\cpu.ex.r_stmp[9] ));
 sg13g2_nor2_1 _17734_ (.A(_10484_),
    .B(_10842_),
    .Y(_10843_));
 sg13g2_nand2_1 _17735_ (.Y(_10844_),
    .A(net751),
    .B(\cpu.ex.r_13[9] ));
 sg13g2_nand2_1 _17736_ (.Y(_10845_),
    .A(net870),
    .B(\cpu.ex.r_12[9] ));
 sg13g2_a21oi_1 _17737_ (.A1(_10844_),
    .A2(_10845_),
    .Y(_10846_),
    .B1(_10591_));
 sg13g2_a22oi_1 _17738_ (.Y(_10847_),
    .B1(_10375_),
    .B2(\cpu.ex.r_14[9] ),
    .A2(_10219_),
    .A1(\cpu.ex.r_11[9] ));
 sg13g2_nor2_1 _17739_ (.A(_10746_),
    .B(_10847_),
    .Y(_10848_));
 sg13g2_mux2_1 _17740_ (.A0(\cpu.ex.r_lr[9] ),
    .A1(\cpu.ex.r_9[9] ),
    .S(net742),
    .X(_10849_));
 sg13g2_a22oi_1 _17741_ (.Y(_10850_),
    .B1(_10849_),
    .B2(net740),
    .A2(_10286_),
    .A1(\cpu.ex.r_8[9] ));
 sg13g2_nor2b_1 _17742_ (.A(_10850_),
    .B_N(_10475_),
    .Y(_10851_));
 sg13g2_nor4_1 _17743_ (.A(_10843_),
    .B(_10846_),
    .C(_10848_),
    .D(_10851_),
    .Y(_10852_));
 sg13g2_nand3_1 _17744_ (.B(_10841_),
    .C(_10852_),
    .A(net596),
    .Y(_10853_));
 sg13g2_nand2_1 _17745_ (.Y(_10854_),
    .A(_10832_),
    .B(_10853_));
 sg13g2_mux2_1 _17746_ (.A0(_00273_),
    .A1(_10854_),
    .S(net250),
    .X(_10855_));
 sg13g2_buf_2 _17747_ (.A(_10855_),
    .X(_10856_));
 sg13g2_or2_1 _17748_ (.X(_10857_),
    .B(_10509_),
    .A(_00245_));
 sg13g2_nand3_1 _17749_ (.B(net861),
    .C(_10316_),
    .A(\cpu.ex.r_8[9] ),
    .Y(_10858_));
 sg13g2_a21oi_1 _17750_ (.A1(_10857_),
    .A2(_10858_),
    .Y(_10859_),
    .B1(net737));
 sg13g2_nand3_1 _17751_ (.B(net861),
    .C(_10309_),
    .A(\cpu.ex.r_stmp[9] ),
    .Y(_10860_));
 sg13g2_nand3_1 _17752_ (.B(net658),
    .C(net663),
    .A(\cpu.ex.r_13[9] ),
    .Y(_10861_));
 sg13g2_a21oi_1 _17753_ (.A1(_10860_),
    .A2(_10861_),
    .Y(_10862_),
    .B1(net657));
 sg13g2_nand3_1 _17754_ (.B(net733),
    .C(net736),
    .A(\cpu.ex.r_12[9] ),
    .Y(_10863_));
 sg13g2_mux2_1 _17755_ (.A0(\cpu.ex.r_lr[9] ),
    .A1(\cpu.ex.r_9[9] ),
    .S(net659),
    .X(_10864_));
 sg13g2_nand2b_1 _17756_ (.Y(_10865_),
    .B(_10864_),
    .A_N(_10184_));
 sg13g2_a21oi_1 _17757_ (.A1(_10863_),
    .A2(_10865_),
    .Y(_10866_),
    .B1(net653));
 sg13g2_mux2_1 _17758_ (.A0(\cpu.ex.r_epc[9] ),
    .A1(_10835_),
    .S(net744),
    .X(_10867_));
 sg13g2_a221oi_1 _17759_ (.B2(net737),
    .C1(net733),
    .B1(_10867_),
    .A1(\cpu.ex.r_11[9] ),
    .Y(_10868_),
    .A2(net746));
 sg13g2_mux2_1 _17760_ (.A0(_10839_),
    .A1(\cpu.ex.r_10[9] ),
    .S(net659),
    .X(_10869_));
 sg13g2_a221oi_1 _17761_ (.B2(net739),
    .C1(net658),
    .B1(_10869_),
    .A1(\cpu.ex.r_14[9] ),
    .Y(_10870_),
    .A2(net736));
 sg13g2_nor3_1 _17762_ (.A(net738),
    .B(_10868_),
    .C(_10870_),
    .Y(_10871_));
 sg13g2_or4_1 _17763_ (.A(_10859_),
    .B(_10862_),
    .C(_10866_),
    .D(_10871_),
    .X(_10872_));
 sg13g2_a22oi_1 _17764_ (.Y(_10873_),
    .B1(_10149_),
    .B2(_10872_),
    .A2(net526),
    .A1(_10831_));
 sg13g2_inv_2 _17765_ (.Y(_10874_),
    .A(_00273_));
 sg13g2_a22oi_1 _17766_ (.Y(_10875_),
    .B1(\cpu.dec.imm[9] ),
    .B2(_10207_),
    .A2(_10874_),
    .A1(net1005));
 sg13g2_o21ai_1 _17767_ (.B1(_10875_),
    .Y(_10876_),
    .A1(net743),
    .A2(_10873_));
 sg13g2_buf_1 _17768_ (.A(_10876_),
    .X(_10877_));
 sg13g2_inv_2 _17769_ (.Y(_10878_),
    .A(_10877_));
 sg13g2_nor2_1 _17770_ (.A(_10856_),
    .B(_10878_),
    .Y(_10879_));
 sg13g2_a21o_1 _17771_ (.A2(_10830_),
    .A1(_10819_),
    .B1(_10879_),
    .X(_10880_));
 sg13g2_buf_1 _17772_ (.A(_10880_),
    .X(_10881_));
 sg13g2_inv_1 _17773_ (.Y(_10882_),
    .A(_00271_));
 sg13g2_nand2_1 _17774_ (.Y(_10883_),
    .A(net1005),
    .B(_10882_));
 sg13g2_buf_2 _17775_ (.A(_10883_),
    .X(_10884_));
 sg13g2_or2_1 _17776_ (.X(_10885_),
    .B(\cpu.dec.imm[11] ),
    .A(net1006));
 sg13g2_nor2_1 _17777_ (.A(net733),
    .B(_10522_),
    .Y(_10886_));
 sg13g2_and2_1 _17778_ (.A(\cpu.ex.r_8[11] ),
    .B(net663),
    .X(_10887_));
 sg13g2_a22oi_1 _17779_ (.Y(_10888_),
    .B1(_10887_),
    .B2(net733),
    .A2(_10886_),
    .A1(\cpu.ex.r_epc[11] ));
 sg13g2_nor2_1 _17780_ (.A(_10516_),
    .B(_10522_),
    .Y(_10889_));
 sg13g2_a221oi_1 _17781_ (.B2(\cpu.ex.r_13[11] ),
    .C1(net657),
    .B1(_10686_),
    .A1(\cpu.ex.r_stmp[11] ),
    .Y(_10890_),
    .A2(_10889_));
 sg13g2_nor2_1 _17782_ (.A(_00247_),
    .B(_10152_),
    .Y(_10891_));
 sg13g2_nand2_1 _17783_ (.Y(_10892_),
    .A(\cpu.ex.r_14[11] ),
    .B(_10624_));
 sg13g2_nand2b_1 _17784_ (.Y(_10893_),
    .B(\cpu.ex.r_12[11] ),
    .A_N(_10624_));
 sg13g2_a21oi_1 _17785_ (.A1(_10892_),
    .A2(_10893_),
    .Y(_10894_),
    .B1(net654));
 sg13g2_o21ai_1 _17786_ (.B1(net593),
    .Y(_10895_),
    .A1(_10891_),
    .A2(_10894_));
 sg13g2_a22oi_1 _17787_ (.Y(_10896_),
    .B1(_10890_),
    .B2(_10895_),
    .A2(_10888_),
    .A1(net657));
 sg13g2_buf_1 _17788_ (.A(_10549_),
    .X(_10897_));
 sg13g2_buf_1 _17789_ (.A(\cpu.ex.r_sp[11] ),
    .X(_10898_));
 sg13g2_nor2_1 _17790_ (.A(net733),
    .B(net653),
    .Y(_10899_));
 sg13g2_mux2_1 _17791_ (.A0(\cpu.ex.r_lr[11] ),
    .A1(\cpu.ex.r_9[11] ),
    .S(net659),
    .X(_10900_));
 sg13g2_a22oi_1 _17792_ (.Y(_10901_),
    .B1(_10899_),
    .B2(_10900_),
    .A2(_10889_),
    .A1(_10898_));
 sg13g2_buf_1 _17793_ (.A(\cpu.ex.r_mult[27] ),
    .X(_10902_));
 sg13g2_mux2_1 _17794_ (.A0(\cpu.ex.r_10[11] ),
    .A1(\cpu.ex.r_11[11] ),
    .S(net654),
    .X(_10903_));
 sg13g2_a22oi_1 _17795_ (.Y(_10904_),
    .B1(_10781_),
    .B2(_10903_),
    .A2(_10409_),
    .A1(_10902_));
 sg13g2_o21ai_1 _17796_ (.B1(_10904_),
    .Y(_10905_),
    .A1(net591),
    .A2(_10901_));
 sg13g2_o21ai_1 _17797_ (.B1(net525),
    .Y(_10906_),
    .A1(_10896_),
    .A2(_10905_));
 sg13g2_buf_2 _17798_ (.A(\cpu.addr[11] ),
    .X(_10907_));
 sg13g2_nand2_1 _17799_ (.Y(_10908_),
    .A(_10907_),
    .B(net526));
 sg13g2_nand3_1 _17800_ (.B(_10906_),
    .C(_10908_),
    .A(net1006),
    .Y(_10909_));
 sg13g2_nand3_1 _17801_ (.B(_10885_),
    .C(_10909_),
    .A(net860),
    .Y(_10910_));
 sg13g2_buf_2 _17802_ (.A(_10910_),
    .X(_10911_));
 sg13g2_nand2_1 _17803_ (.Y(_10912_),
    .A(_10884_),
    .B(_10911_));
 sg13g2_buf_1 _17804_ (.A(_10912_),
    .X(_10913_));
 sg13g2_and2_1 _17805_ (.A(_10098_),
    .B(_10286_),
    .X(_10914_));
 sg13g2_mux2_1 _17806_ (.A0(\cpu.ex.r_8[11] ),
    .A1(\cpu.ex.r_10[11] ),
    .S(net595),
    .X(_10915_));
 sg13g2_nand2_1 _17807_ (.Y(_10916_),
    .A(_10914_),
    .B(_10915_));
 sg13g2_inv_1 _17808_ (.Y(_10917_),
    .A(_00247_));
 sg13g2_and3_1 _17809_ (.X(_10918_),
    .A(_10055_),
    .B(net749),
    .C(net750));
 sg13g2_nor3_1 _17810_ (.A(net862),
    .B(net749),
    .C(net750),
    .Y(_10919_));
 sg13g2_a22oi_1 _17811_ (.Y(_10920_),
    .B1(_10919_),
    .B2(_10898_),
    .A2(_10918_),
    .A1(_10917_));
 sg13g2_inv_1 _17812_ (.Y(_10921_),
    .A(_10920_));
 sg13g2_inv_1 _17813_ (.Y(_10922_),
    .A(\cpu.ex.r_13[11] ));
 sg13g2_nand3_1 _17814_ (.B(\cpu.ex.r_epc[11] ),
    .C(_10361_),
    .A(net671),
    .Y(_10923_));
 sg13g2_o21ai_1 _17815_ (.B1(_10923_),
    .Y(_10924_),
    .A1(_10922_),
    .A2(_10591_));
 sg13g2_a22oi_1 _17816_ (.Y(_10925_),
    .B1(_10924_),
    .B2(net670),
    .A2(_10921_),
    .A1(net595));
 sg13g2_a22oi_1 _17817_ (.Y(_10926_),
    .B1(_10375_),
    .B2(\cpu.ex.r_12[11] ),
    .A2(_10219_),
    .A1(\cpu.ex.r_9[11] ));
 sg13g2_a221oi_1 _17818_ (.B2(\cpu.ex.r_14[11] ),
    .C1(net666),
    .B1(_10375_),
    .A1(\cpu.ex.r_11[11] ),
    .Y(_10927_),
    .A2(_10219_));
 sg13g2_a21oi_1 _17819_ (.A1(net666),
    .A2(_10926_),
    .Y(_10928_),
    .B1(_10927_));
 sg13g2_nand2_1 _17820_ (.Y(_10929_),
    .A(net660),
    .B(_10928_));
 sg13g2_nand3_1 _17821_ (.B(\cpu.ex.r_lr[11] ),
    .C(net661),
    .A(net664),
    .Y(_10930_));
 sg13g2_mux2_1 _17822_ (.A0(\cpu.ex.r_stmp[11] ),
    .A1(_10902_),
    .S(net751),
    .X(_10931_));
 sg13g2_nand2_1 _17823_ (.Y(_10932_),
    .A(_10477_),
    .B(_10931_));
 sg13g2_a21o_1 _17824_ (.A2(_10932_),
    .A1(_10930_),
    .B1(net660),
    .X(_10933_));
 sg13g2_nand4_1 _17825_ (.B(_10925_),
    .C(_10929_),
    .A(_10916_),
    .Y(_10934_),
    .D(_10933_));
 sg13g2_mux2_1 _17826_ (.A0(_10907_),
    .A1(_10934_),
    .S(_10357_),
    .X(_10935_));
 sg13g2_buf_1 _17827_ (.A(_10935_),
    .X(_10936_));
 sg13g2_nor2_1 _17828_ (.A(_00271_),
    .B(net250),
    .Y(_10937_));
 sg13g2_a21o_1 _17829_ (.A2(_10936_),
    .A1(net227),
    .B1(_10937_),
    .X(_10938_));
 sg13g2_buf_1 _17830_ (.A(_10938_),
    .X(_10939_));
 sg13g2_nor2_1 _17831_ (.A(net183),
    .B(_10939_),
    .Y(_10940_));
 sg13g2_inv_1 _17832_ (.Y(_10941_),
    .A(_00272_));
 sg13g2_nand3_1 _17833_ (.B(_10063_),
    .C(_10278_),
    .A(\cpu.ex.r_11[10] ),
    .Y(_10942_));
 sg13g2_mux2_1 _17834_ (.A0(\cpu.ex.r_8[10] ),
    .A1(\cpu.ex.r_12[10] ),
    .S(_10066_),
    .X(_10943_));
 sg13g2_nand3_1 _17835_ (.B(_10096_),
    .C(_10943_),
    .A(net870),
    .Y(_10944_));
 sg13g2_nand2_1 _17836_ (.Y(_10945_),
    .A(_10942_),
    .B(_10944_));
 sg13g2_and2_1 _17837_ (.A(net751),
    .B(_10058_),
    .X(_10946_));
 sg13g2_buf_2 _17838_ (.A(\cpu.ex.r_mult[26] ),
    .X(_10947_));
 sg13g2_a22oi_1 _17839_ (.Y(_10948_),
    .B1(_10946_),
    .B2(_10947_),
    .A2(_10914_),
    .A1(\cpu.ex.r_10[10] ));
 sg13g2_inv_1 _17840_ (.Y(_10949_),
    .A(\cpu.ex.r_13[10] ));
 sg13g2_nor2_1 _17841_ (.A(_10949_),
    .B(_10591_),
    .Y(_10950_));
 sg13g2_and3_1 _17842_ (.X(_10951_),
    .A(net752),
    .B(\cpu.ex.r_epc[10] ),
    .C(_10361_));
 sg13g2_o21ai_1 _17843_ (.B1(net670),
    .Y(_10952_),
    .A1(_10950_),
    .A2(_10951_));
 sg13g2_o21ai_1 _17844_ (.B1(_10952_),
    .Y(_10953_),
    .A1(net666),
    .A2(_10948_));
 sg13g2_inv_1 _17845_ (.Y(_10954_),
    .A(_00246_));
 sg13g2_a22oi_1 _17846_ (.Y(_10955_),
    .B1(_10071_),
    .B2(_10954_),
    .A2(_10267_),
    .A1(\cpu.ex.r_stmp[10] ));
 sg13g2_nor2b_1 _17847_ (.A(_10955_),
    .B_N(_10477_),
    .Y(_10956_));
 sg13g2_buf_1 _17848_ (.A(\cpu.ex.r_sp[10] ),
    .X(_10957_));
 sg13g2_a22oi_1 _17849_ (.Y(_10958_),
    .B1(_10222_),
    .B2(\cpu.ex.r_14[10] ),
    .A2(_10361_),
    .A1(_10957_));
 sg13g2_mux2_1 _17850_ (.A0(\cpu.ex.r_lr[10] ),
    .A1(\cpu.ex.r_9[10] ),
    .S(net655),
    .X(_10959_));
 sg13g2_nand3_1 _17851_ (.B(net661),
    .C(_10959_),
    .A(net664),
    .Y(_10960_));
 sg13g2_o21ai_1 _17852_ (.B1(_10960_),
    .Y(_10961_),
    .A1(_10484_),
    .A2(_10958_));
 sg13g2_nor4_1 _17853_ (.A(_10945_),
    .B(_10953_),
    .C(_10956_),
    .D(_10961_),
    .Y(_10962_));
 sg13g2_buf_1 _17854_ (.A(\cpu.addr[10] ),
    .X(_10963_));
 sg13g2_nor2_1 _17855_ (.A(net1095),
    .B(net596),
    .Y(_10964_));
 sg13g2_a21oi_1 _17856_ (.A1(net527),
    .A2(_10962_),
    .Y(_10965_),
    .B1(_10964_));
 sg13g2_mux2_1 _17857_ (.A0(_10941_),
    .A1(_10965_),
    .S(net251),
    .X(_10966_));
 sg13g2_buf_8 _17858_ (.A(_10966_),
    .X(_10967_));
 sg13g2_nand2_1 _17859_ (.Y(_10968_),
    .A(net1005),
    .B(_10941_));
 sg13g2_buf_2 _17860_ (.A(_10968_),
    .X(_10969_));
 sg13g2_nor2_1 _17861_ (.A(net1006),
    .B(\cpu.dec.imm[10] ),
    .Y(_10970_));
 sg13g2_and2_1 _17862_ (.A(net658),
    .B(net747),
    .X(_10971_));
 sg13g2_buf_1 _17863_ (.A(_10971_),
    .X(_10972_));
 sg13g2_buf_1 _17864_ (.A(net654),
    .X(_10973_));
 sg13g2_mux2_1 _17865_ (.A0(_10957_),
    .A1(\cpu.ex.r_stmp[10] ),
    .S(net656),
    .X(_10974_));
 sg13g2_a22oi_1 _17866_ (.Y(_10975_),
    .B1(_10974_),
    .B2(net737),
    .A2(_10433_),
    .A1(\cpu.ex.r_14[10] ));
 sg13g2_nor2_1 _17867_ (.A(net590),
    .B(_10975_),
    .Y(_10976_));
 sg13g2_a21oi_1 _17868_ (.A1(\cpu.ex.r_epc[10] ),
    .A2(_10972_),
    .Y(_10977_),
    .B1(_10976_));
 sg13g2_nand2_1 _17869_ (.Y(_10978_),
    .A(\cpu.ex.r_lr[10] ),
    .B(_10312_));
 sg13g2_nand3_1 _17870_ (.B(net656),
    .C(_10192_),
    .A(_10954_),
    .Y(_10979_));
 sg13g2_o21ai_1 _17871_ (.B1(_10979_),
    .Y(_10980_),
    .A1(net591),
    .A2(_10978_));
 sg13g2_and2_1 _17872_ (.A(\cpu.ex.r_12[10] ),
    .B(net656),
    .X(_10981_));
 sg13g2_a21oi_1 _17873_ (.A1(\cpu.ex.r_8[10] ),
    .A2(_10301_),
    .Y(_10982_),
    .B1(_10981_));
 sg13g2_nand3_1 _17874_ (.B(net654),
    .C(net656),
    .A(\cpu.ex.r_13[10] ),
    .Y(_10983_));
 sg13g2_o21ai_1 _17875_ (.B1(_10983_),
    .Y(_10984_),
    .A1(net590),
    .A2(_10982_));
 sg13g2_mux2_1 _17876_ (.A0(\cpu.ex.r_9[10] ),
    .A1(\cpu.ex.r_11[10] ),
    .S(net653),
    .X(_10985_));
 sg13g2_nand3_1 _17877_ (.B(_10158_),
    .C(_10985_),
    .A(net654),
    .Y(_10986_));
 sg13g2_nand4_1 _17878_ (.B(net654),
    .C(net591),
    .A(_10947_),
    .Y(_10987_),
    .D(_10309_));
 sg13g2_nand3_1 _17879_ (.B(net746),
    .C(_10400_),
    .A(\cpu.ex.r_10[10] ),
    .Y(_10988_));
 sg13g2_nand3_1 _17880_ (.B(_10987_),
    .C(_10988_),
    .A(_10986_),
    .Y(_10989_));
 sg13g2_a221oi_1 _17881_ (.B2(net663),
    .C1(_10989_),
    .B1(_10984_),
    .A1(net590),
    .Y(_10990_),
    .A2(_10980_));
 sg13g2_o21ai_1 _17882_ (.B1(_10990_),
    .Y(_10991_),
    .A1(_10306_),
    .A2(_10977_));
 sg13g2_a221oi_1 _17883_ (.B2(_10991_),
    .C1(_10131_),
    .B1(net525),
    .A1(net1095),
    .Y(_10992_),
    .A2(_10533_));
 sg13g2_or3_1 _17884_ (.A(net1005),
    .B(_10970_),
    .C(_10992_),
    .X(_10993_));
 sg13g2_buf_2 _17885_ (.A(_10993_),
    .X(_10994_));
 sg13g2_nand2_1 _17886_ (.Y(_10995_),
    .A(_10969_),
    .B(_10994_));
 sg13g2_buf_1 _17887_ (.A(_10995_),
    .X(_10996_));
 sg13g2_nand2_1 _17888_ (.Y(_10997_),
    .A(net204),
    .B(net182));
 sg13g2_nand2_1 _17889_ (.Y(_10998_),
    .A(net183),
    .B(_10939_));
 sg13g2_o21ai_1 _17890_ (.B1(_10998_),
    .Y(_10999_),
    .A1(_10940_),
    .A2(_10997_));
 sg13g2_or3_1 _17891_ (.A(_10807_),
    .B(_10881_),
    .C(_10999_),
    .X(_11000_));
 sg13g2_buf_1 _17892_ (.A(_11000_),
    .X(_11001_));
 sg13g2_inv_1 _17893_ (.Y(_11002_),
    .A(_00270_));
 sg13g2_inv_1 _17894_ (.Y(_11003_),
    .A(_00248_));
 sg13g2_a22oi_1 _17895_ (.Y(_11004_),
    .B1(_10222_),
    .B2(_11003_),
    .A2(_10361_),
    .A1(\cpu.ex.r_epc[12] ));
 sg13g2_nand3b_1 _17896_ (.B(net741),
    .C(\cpu.ex.r_14[12] ),
    .Y(_11005_),
    .A_N(net751));
 sg13g2_nand3b_1 _17897_ (.B(\cpu.ex.r_11[12] ),
    .C(net740),
    .Y(_11006_),
    .A_N(net750));
 sg13g2_a21o_1 _17898_ (.A2(_11006_),
    .A1(_11005_),
    .B1(_10746_),
    .X(_11007_));
 sg13g2_o21ai_1 _17899_ (.B1(_11007_),
    .Y(_11008_),
    .A1(_10371_),
    .A2(_11004_));
 sg13g2_nand3_1 _17900_ (.B(\cpu.ex.r_8[12] ),
    .C(_10286_),
    .A(net664),
    .Y(_11009_));
 sg13g2_buf_2 _17901_ (.A(\cpu.ex.mmu_read[12] ),
    .X(_11010_));
 sg13g2_nand3_1 _17902_ (.B(_11010_),
    .C(net669),
    .A(net670),
    .Y(_11011_));
 sg13g2_a21oi_1 _17903_ (.A1(_11009_),
    .A2(_11011_),
    .Y(_11012_),
    .B1(net595));
 sg13g2_a221oi_1 _17904_ (.B2(\cpu.ex.r_12[12] ),
    .C1(_10056_),
    .B1(net665),
    .A1(\cpu.ex.r_stmp[12] ),
    .Y(_11013_),
    .A2(net667));
 sg13g2_buf_2 _17905_ (.A(\cpu.ex.r_mult[28] ),
    .X(_11014_));
 sg13g2_a221oi_1 _17906_ (.B2(\cpu.ex.r_13[12] ),
    .C1(_10101_),
    .B1(net665),
    .A1(_11014_),
    .Y(_11015_),
    .A2(_10077_));
 sg13g2_nor3_1 _17907_ (.A(net664),
    .B(_11013_),
    .C(_11015_),
    .Y(_11016_));
 sg13g2_mux2_1 _17908_ (.A0(\cpu.ex.r_lr[12] ),
    .A1(\cpu.ex.r_9[12] ),
    .S(_10601_),
    .X(_11017_));
 sg13g2_buf_1 _17909_ (.A(\cpu.ex.r_sp[12] ),
    .X(_11018_));
 sg13g2_mux2_1 _17910_ (.A0(_11018_),
    .A1(\cpu.ex.r_10[12] ),
    .S(_10601_),
    .X(_11019_));
 sg13g2_a22oi_1 _17911_ (.Y(_11020_),
    .B1(_11019_),
    .B2(net662),
    .A2(_11017_),
    .A1(_10245_));
 sg13g2_nor2_1 _17912_ (.A(net741),
    .B(_11020_),
    .Y(_11021_));
 sg13g2_nor4_2 _17913_ (.A(_11008_),
    .B(_11012_),
    .C(_11016_),
    .Y(_11022_),
    .D(_11021_));
 sg13g2_buf_1 _17914_ (.A(net679),
    .X(_11023_));
 sg13g2_nor2_1 _17915_ (.A(net589),
    .B(net527),
    .Y(_11024_));
 sg13g2_a21oi_1 _17916_ (.A1(net527),
    .A2(_11022_),
    .Y(_11025_),
    .B1(_11024_));
 sg13g2_and2_1 _17917_ (.A(net227),
    .B(_11025_),
    .X(_11026_));
 sg13g2_a21oi_1 _17918_ (.A1(_11002_),
    .A2(net303),
    .Y(_11027_),
    .B1(_11026_));
 sg13g2_buf_1 _17919_ (.A(_11027_),
    .X(_11028_));
 sg13g2_inv_1 _17920_ (.Y(_11029_),
    .A(_10884_));
 sg13g2_and3_1 _17921_ (.X(_11030_),
    .A(net860),
    .B(_10885_),
    .C(_10909_));
 sg13g2_buf_1 _17922_ (.A(_11030_),
    .X(_11031_));
 sg13g2_nor2_1 _17923_ (.A(_11029_),
    .B(_11031_),
    .Y(_11032_));
 sg13g2_buf_1 _17924_ (.A(_11032_),
    .X(_11033_));
 sg13g2_a21oi_2 _17925_ (.B1(_10937_),
    .Y(_11034_),
    .A2(_10936_),
    .A1(net227));
 sg13g2_nor2_1 _17926_ (.A(_11033_),
    .B(_11034_),
    .Y(_11035_));
 sg13g2_nand2_1 _17927_ (.Y(_11036_),
    .A(_10856_),
    .B(_10878_));
 sg13g2_nand2_1 _17928_ (.Y(_11037_),
    .A(net182),
    .B(_11036_));
 sg13g2_o21ai_1 _17929_ (.B1(net204),
    .Y(_11038_),
    .A1(net182),
    .A2(_11036_));
 sg13g2_a21oi_1 _17930_ (.A1(_11037_),
    .A2(_11038_),
    .Y(_11039_),
    .B1(_10940_));
 sg13g2_nor2_1 _17931_ (.A(_11035_),
    .B(_11039_),
    .Y(_11040_));
 sg13g2_nor2_1 _17932_ (.A(_11028_),
    .B(_11040_),
    .Y(_11041_));
 sg13g2_buf_1 _17933_ (.A(net886),
    .X(_11042_));
 sg13g2_buf_1 _17934_ (.A(net526),
    .X(_11043_));
 sg13g2_mux2_1 _17935_ (.A0(\cpu.ex.r_epc[14] ),
    .A1(\cpu.ex.r_11[14] ),
    .S(net593),
    .X(_11044_));
 sg13g2_nand2_1 _17936_ (.Y(_11045_),
    .A(net657),
    .B(_11044_));
 sg13g2_o21ai_1 _17937_ (.B1(_11045_),
    .Y(_11046_),
    .A1(_00250_),
    .A2(_10616_));
 sg13g2_buf_2 _17938_ (.A(\cpu.ex.r_mult[30] ),
    .X(_11047_));
 sg13g2_a22oi_1 _17939_ (.Y(_11048_),
    .B1(_10320_),
    .B2(_11047_),
    .A2(_10316_),
    .A1(\cpu.ex.r_lr[14] ));
 sg13g2_buf_1 _17940_ (.A(_10973_),
    .X(_11049_));
 sg13g2_o21ai_1 _17941_ (.B1(net524),
    .Y(_11050_),
    .A1(net593),
    .A2(_11048_));
 sg13g2_a221oi_1 _17942_ (.B2(net592),
    .C1(_11050_),
    .B1(_11046_),
    .A1(\cpu.ex.r_9[14] ),
    .Y(_11051_),
    .A2(_10413_));
 sg13g2_buf_1 _17943_ (.A(\cpu.ex.r_sp[14] ),
    .X(_11052_));
 sg13g2_a22oi_1 _17944_ (.Y(_11053_),
    .B1(_10309_),
    .B2(_11052_),
    .A2(net663),
    .A1(\cpu.ex.r_8[14] ));
 sg13g2_a221oi_1 _17945_ (.B2(\cpu.ex.r_stmp[14] ),
    .C1(net657),
    .B1(_10309_),
    .A1(\cpu.ex.r_12[14] ),
    .Y(_11054_),
    .A2(net663));
 sg13g2_a21oi_1 _17946_ (.A1(net657),
    .A2(_11053_),
    .Y(_11055_),
    .B1(_11054_));
 sg13g2_nor2_1 _17947_ (.A(_11049_),
    .B(_11055_),
    .Y(_11056_));
 sg13g2_nand3_1 _17948_ (.B(net733),
    .C(_10393_),
    .A(\cpu.ex.r_10[14] ),
    .Y(_11057_));
 sg13g2_nor2b_1 _17949_ (.A(net653),
    .B_N(net656),
    .Y(_11058_));
 sg13g2_nand3_1 _17950_ (.B(net524),
    .C(_11058_),
    .A(\cpu.ex.r_13[14] ),
    .Y(_11059_));
 sg13g2_nand2_1 _17951_ (.Y(_11060_),
    .A(_11057_),
    .B(_11059_));
 sg13g2_inv_1 _17952_ (.Y(_11061_),
    .A(\cpu.ex.r_14[14] ));
 sg13g2_buf_2 _17953_ (.A(\cpu.ex.mmu_read[14] ),
    .X(_11062_));
 sg13g2_nand3_1 _17954_ (.B(net524),
    .C(_10312_),
    .A(_11062_),
    .Y(_11063_));
 sg13g2_o21ai_1 _17955_ (.B1(_11063_),
    .Y(_11064_),
    .A1(_11061_),
    .A2(_10401_));
 sg13g2_a22oi_1 _17956_ (.Y(_11065_),
    .B1(_11064_),
    .B2(net591),
    .A2(_11060_),
    .A1(net593));
 sg13g2_o21ai_1 _17957_ (.B1(_11065_),
    .Y(_11066_),
    .A1(_11051_),
    .A2(_11056_));
 sg13g2_a22oi_1 _17958_ (.Y(_11067_),
    .B1(_10792_),
    .B2(_11066_),
    .A2(net459),
    .A1(net732));
 sg13g2_inv_1 _17959_ (.Y(_11068_),
    .A(_00179_));
 sg13g2_a22oi_1 _17960_ (.Y(_11069_),
    .B1(\cpu.dec.imm[14] ),
    .B2(_10207_),
    .A2(_11068_),
    .A1(net1005));
 sg13g2_o21ai_1 _17961_ (.B1(_11069_),
    .Y(_11070_),
    .A1(net743),
    .A2(_11067_));
 sg13g2_buf_2 _17962_ (.A(_11070_),
    .X(_11071_));
 sg13g2_inv_1 _17963_ (.Y(_11072_),
    .A(_11071_));
 sg13g2_buf_1 _17964_ (.A(_11072_),
    .X(_11073_));
 sg13g2_inv_1 _17965_ (.Y(_11074_),
    .A(\cpu.ex.r_epc[14] ));
 sg13g2_nand3b_1 _17966_ (.B(net655),
    .C(\cpu.ex.r_10[14] ),
    .Y(_11075_),
    .A_N(net740));
 sg13g2_o21ai_1 _17967_ (.B1(_11075_),
    .Y(_11076_),
    .A1(_11074_),
    .A2(_10234_));
 sg13g2_inv_1 _17968_ (.Y(_11077_),
    .A(\cpu.ex.r_lr[14] ));
 sg13g2_nand3_1 _17969_ (.B(net660),
    .C(\cpu.ex.r_11[14] ),
    .A(net671),
    .Y(_11078_));
 sg13g2_o21ai_1 _17970_ (.B1(_11078_),
    .Y(_11079_),
    .A1(_11077_),
    .A2(_10586_));
 sg13g2_a22oi_1 _17971_ (.Y(_11080_),
    .B1(_11079_),
    .B2(_10219_),
    .A2(_11076_),
    .A1(_10760_));
 sg13g2_and2_1 _17972_ (.A(net669),
    .B(_10278_),
    .X(_11081_));
 sg13g2_mux2_1 _17973_ (.A0(\cpu.ex.r_9[14] ),
    .A1(\cpu.ex.r_13[14] ),
    .S(net741),
    .X(_11082_));
 sg13g2_and2_1 _17974_ (.A(net660),
    .B(net661),
    .X(_11083_));
 sg13g2_nand2b_1 _17975_ (.Y(_11084_),
    .B(net740),
    .A_N(_00250_));
 sg13g2_nand2b_1 _17976_ (.Y(_11085_),
    .B(\cpu.ex.r_14[14] ),
    .A_N(net751));
 sg13g2_a21oi_1 _17977_ (.A1(_11084_),
    .A2(_11085_),
    .Y(_11086_),
    .B1(_10649_));
 sg13g2_a221oi_1 _17978_ (.B2(_11083_),
    .C1(_11086_),
    .B1(_11082_),
    .A1(_11047_),
    .Y(_11087_),
    .A2(_11081_));
 sg13g2_nand3_1 _17979_ (.B(\cpu.ex.r_8[14] ),
    .C(_10286_),
    .A(net664),
    .Y(_11088_));
 sg13g2_nand3_1 _17980_ (.B(_11062_),
    .C(net669),
    .A(_10056_),
    .Y(_11089_));
 sg13g2_a21o_1 _17981_ (.A2(_11089_),
    .A1(_11088_),
    .B1(net595),
    .X(_11090_));
 sg13g2_nand3_1 _17982_ (.B(\cpu.ex.r_12[14] ),
    .C(net665),
    .A(net741),
    .Y(_11091_));
 sg13g2_mux2_1 _17983_ (.A0(_11052_),
    .A1(\cpu.ex.r_stmp[14] ),
    .S(_10066_),
    .X(_11092_));
 sg13g2_nand2_1 _17984_ (.Y(_11093_),
    .A(net667),
    .B(_11092_));
 sg13g2_a21o_1 _17985_ (.A2(_11093_),
    .A1(_11091_),
    .B1(net670),
    .X(_11094_));
 sg13g2_nand4_1 _17986_ (.B(_11087_),
    .C(_11090_),
    .A(_11080_),
    .Y(_11095_),
    .D(_11094_));
 sg13g2_mux2_1 _17987_ (.A0(net732),
    .A1(_11095_),
    .S(net596),
    .X(_11096_));
 sg13g2_mux2_1 _17988_ (.A0(_11068_),
    .A1(_11096_),
    .S(_10826_),
    .X(_11097_));
 sg13g2_buf_2 _17989_ (.A(_11097_),
    .X(_11098_));
 sg13g2_inv_1 _17990_ (.Y(_11099_),
    .A(_11098_));
 sg13g2_buf_1 _17991_ (.A(_11099_),
    .X(_11100_));
 sg13g2_mux2_1 _17992_ (.A0(\cpu.ex.r_stmp[13] ),
    .A1(\cpu.ex.r_14[13] ),
    .S(net660),
    .X(_11101_));
 sg13g2_a22oi_1 _17993_ (.Y(_11102_),
    .B1(_11101_),
    .B2(net595),
    .A2(net665),
    .A1(\cpu.ex.r_12[13] ));
 sg13g2_nand2b_1 _17994_ (.Y(_11103_),
    .B(_10375_),
    .A_N(_11102_));
 sg13g2_inv_1 _17995_ (.Y(_11104_),
    .A(_00249_));
 sg13g2_buf_1 _17996_ (.A(\cpu.ex.r_sp[13] ),
    .X(_11105_));
 sg13g2_a22oi_1 _17997_ (.Y(_11106_),
    .B1(_10919_),
    .B2(_11105_),
    .A2(_10918_),
    .A1(_11104_));
 sg13g2_nand2b_1 _17998_ (.Y(_11107_),
    .B(net595),
    .A_N(_11106_));
 sg13g2_nand3_1 _17999_ (.B(net662),
    .C(net668),
    .A(\cpu.ex.r_10[13] ),
    .Y(_11108_));
 sg13g2_mux2_1 _18000_ (.A0(\cpu.ex.r_lr[13] ),
    .A1(\cpu.ex.r_9[13] ),
    .S(_10078_),
    .X(_11109_));
 sg13g2_nand3_1 _18001_ (.B(net661),
    .C(_11109_),
    .A(net664),
    .Y(_11110_));
 sg13g2_nand2_1 _18002_ (.Y(_11111_),
    .A(_11108_),
    .B(_11110_));
 sg13g2_buf_2 _18003_ (.A(\cpu.ex.r_mult[29] ),
    .X(_11112_));
 sg13g2_a22oi_1 _18004_ (.Y(_11113_),
    .B1(net668),
    .B2(\cpu.ex.r_11[13] ),
    .A2(net669),
    .A1(_11112_));
 sg13g2_nor2_1 _18005_ (.A(_10371_),
    .B(_11113_),
    .Y(_11114_));
 sg13g2_buf_1 _18006_ (.A(\cpu.ex.mmu_read[13] ),
    .X(_11115_));
 sg13g2_a22oi_1 _18007_ (.Y(_11116_),
    .B1(_10760_),
    .B2(\cpu.ex.r_epc[13] ),
    .A2(_10231_),
    .A1(_11115_));
 sg13g2_nor2_1 _18008_ (.A(_10234_),
    .B(_11116_),
    .Y(_11117_));
 sg13g2_a22oi_1 _18009_ (.Y(_11118_),
    .B1(_10251_),
    .B2(\cpu.ex.r_13[13] ),
    .A2(_10249_),
    .A1(\cpu.ex.r_8[13] ));
 sg13g2_nor2b_1 _18010_ (.A(_11118_),
    .B_N(_10096_),
    .Y(_11119_));
 sg13g2_nor4_1 _18011_ (.A(_11111_),
    .B(_11114_),
    .C(_11117_),
    .D(_11119_),
    .Y(_11120_));
 sg13g2_nand4_1 _18012_ (.B(_11103_),
    .C(_11107_),
    .A(net527),
    .Y(_11121_),
    .D(_11120_));
 sg13g2_nand2b_1 _18013_ (.Y(_11122_),
    .B(net594),
    .A_N(net678));
 sg13g2_and2_1 _18014_ (.A(_11121_),
    .B(_11122_),
    .X(_11123_));
 sg13g2_buf_1 _18015_ (.A(_11123_),
    .X(_11124_));
 sg13g2_buf_1 _18016_ (.A(_00180_),
    .X(_11125_));
 sg13g2_nor2_1 _18017_ (.A(_11125_),
    .B(net227),
    .Y(_11126_));
 sg13g2_a21oi_1 _18018_ (.A1(net227),
    .A2(_11124_),
    .Y(_11127_),
    .B1(_11126_));
 sg13g2_o21ai_1 _18019_ (.B1(_11127_),
    .Y(_11128_),
    .A1(net147),
    .A2(net119));
 sg13g2_nor2_1 _18020_ (.A(net860),
    .B(_11125_),
    .Y(_11129_));
 sg13g2_or2_1 _18021_ (.X(_11130_),
    .B(\cpu.dec.imm[13] ),
    .A(_10424_));
 sg13g2_a22oi_1 _18022_ (.Y(_11131_),
    .B1(_10629_),
    .B2(\cpu.ex.r_14[13] ),
    .A2(_10972_),
    .A1(\cpu.ex.r_epc[13] ));
 sg13g2_and2_1 _18023_ (.A(_11115_),
    .B(_10155_),
    .X(_11132_));
 sg13g2_nor2_1 _18024_ (.A(net590),
    .B(_10412_),
    .Y(_11133_));
 sg13g2_a221oi_1 _18025_ (.B2(\cpu.ex.r_8[13] ),
    .C1(_10625_),
    .B1(_11133_),
    .A1(net590),
    .Y(_11134_),
    .A2(_11132_));
 sg13g2_a21o_1 _18026_ (.A2(_11131_),
    .A1(net592),
    .B1(_11134_),
    .X(_11135_));
 sg13g2_a221oi_1 _18027_ (.B2(_11112_),
    .C1(net593),
    .B1(_10320_),
    .A1(\cpu.ex.r_lr[13] ),
    .Y(_11136_),
    .A2(_10316_));
 sg13g2_a221oi_1 _18028_ (.B2(_11104_),
    .C1(net737),
    .B1(_10320_),
    .A1(\cpu.ex.r_9[13] ),
    .Y(_11137_),
    .A2(_10316_));
 sg13g2_nor3_1 _18029_ (.A(net733),
    .B(_11136_),
    .C(_11137_),
    .Y(_11138_));
 sg13g2_a22oi_1 _18030_ (.Y(_11139_),
    .B1(_10407_),
    .B2(\cpu.ex.r_11[13] ),
    .A2(_10189_),
    .A1(_11105_));
 sg13g2_nor2_1 _18031_ (.A(_10405_),
    .B(_11139_),
    .Y(_11140_));
 sg13g2_a22oi_1 _18032_ (.Y(_11141_),
    .B1(_10309_),
    .B2(\cpu.ex.r_stmp[13] ),
    .A2(_10163_),
    .A1(\cpu.ex.r_12[13] ));
 sg13g2_nor3_1 _18033_ (.A(net590),
    .B(_10519_),
    .C(_11141_),
    .Y(_11142_));
 sg13g2_nand3_1 _18034_ (.B(_10771_),
    .C(_10393_),
    .A(\cpu.ex.r_10[13] ),
    .Y(_11143_));
 sg13g2_nand3_1 _18035_ (.B(net590),
    .C(_11058_),
    .A(\cpu.ex.r_13[13] ),
    .Y(_11144_));
 sg13g2_a21oi_1 _18036_ (.A1(_11143_),
    .A2(_11144_),
    .Y(_11145_),
    .B1(net737));
 sg13g2_nor4_1 _18037_ (.A(_11138_),
    .B(_11140_),
    .C(_11142_),
    .D(_11145_),
    .Y(_11146_));
 sg13g2_a21oi_1 _18038_ (.A1(_11135_),
    .A2(_11146_),
    .Y(_11147_),
    .B1(_10344_));
 sg13g2_nand2_1 _18039_ (.Y(_11148_),
    .A(net601),
    .B(net526));
 sg13g2_nand3b_1 _18040_ (.B(_11148_),
    .C(net1006),
    .Y(_11149_),
    .A_N(_11147_));
 sg13g2_and3_1 _18041_ (.X(_11150_),
    .A(net860),
    .B(_11130_),
    .C(_11149_));
 sg13g2_buf_1 _18042_ (.A(_11150_),
    .X(_11151_));
 sg13g2_nor2_1 _18043_ (.A(_11129_),
    .B(_11151_),
    .Y(_11152_));
 sg13g2_buf_1 _18044_ (.A(_11152_),
    .X(_11153_));
 sg13g2_o21ai_1 _18045_ (.B1(_11153_),
    .Y(_11154_),
    .A1(net147),
    .A2(net119));
 sg13g2_a21o_1 _18046_ (.A2(_10613_),
    .A1(_10468_),
    .B1(_10806_),
    .X(_11155_));
 sg13g2_a21o_1 _18047_ (.A2(net303),
    .A1(_11002_),
    .B1(_11026_),
    .X(_11156_));
 sg13g2_buf_2 _18048_ (.A(_11156_),
    .X(_11157_));
 sg13g2_nor3_1 _18049_ (.A(_11157_),
    .B(_10881_),
    .C(_10999_),
    .Y(_11158_));
 sg13g2_mux2_1 _18050_ (.A0(\cpu.ex.r_8[12] ),
    .A1(\cpu.ex.r_12[12] ),
    .S(_10897_),
    .X(_11159_));
 sg13g2_a22oi_1 _18051_ (.Y(_11160_),
    .B1(_11159_),
    .B2(net738),
    .A2(_10393_),
    .A1(\cpu.ex.r_10[12] ));
 sg13g2_nand2b_1 _18052_ (.Y(_11161_),
    .B(_11003_),
    .A_N(_10509_));
 sg13g2_o21ai_1 _18053_ (.B1(_11161_),
    .Y(_11162_),
    .A1(net524),
    .A2(_11160_));
 sg13g2_mux2_1 _18054_ (.A0(\cpu.ex.r_stmp[12] ),
    .A1(\cpu.ex.r_14[12] ),
    .S(_10507_),
    .X(_11163_));
 sg13g2_a22oi_1 _18055_ (.Y(_11164_),
    .B1(_11163_),
    .B2(net591),
    .A2(net747),
    .A1(_11018_));
 sg13g2_nand3_1 _18056_ (.B(net524),
    .C(net746),
    .A(\cpu.ex.r_11[12] ),
    .Y(_11165_));
 sg13g2_o21ai_1 _18057_ (.B1(_11165_),
    .Y(_11166_),
    .A1(net524),
    .A2(_11164_));
 sg13g2_mux4_1 _18058_ (.S0(_10625_),
    .A0(\cpu.ex.r_lr[12] ),
    .A1(\cpu.ex.r_epc[12] ),
    .A2(_11010_),
    .A3(_11014_),
    .S1(net591),
    .X(_11167_));
 sg13g2_mux2_1 _18059_ (.A0(\cpu.ex.r_9[12] ),
    .A1(\cpu.ex.r_13[12] ),
    .S(net591),
    .X(_11168_));
 sg13g2_a22oi_1 _18060_ (.Y(_11169_),
    .B1(_11168_),
    .B2(_10163_),
    .A2(_11167_),
    .A1(_10391_));
 sg13g2_nor2_1 _18061_ (.A(_10771_),
    .B(_11169_),
    .Y(_11170_));
 sg13g2_a221oi_1 _18062_ (.B2(net592),
    .C1(_11170_),
    .B1(_11166_),
    .A1(net593),
    .Y(_11171_),
    .A2(_11162_));
 sg13g2_nand2_1 _18063_ (.Y(_11172_),
    .A(net589),
    .B(net459));
 sg13g2_o21ai_1 _18064_ (.B1(_11172_),
    .Y(_11173_),
    .A1(_10344_),
    .A2(_11171_));
 sg13g2_nor2_1 _18065_ (.A(net860),
    .B(_00270_),
    .Y(_11174_));
 sg13g2_a221oi_1 _18066_ (.B2(_10133_),
    .C1(_11174_),
    .B1(_11173_),
    .A1(\cpu.dec.imm[12] ),
    .Y(_11175_),
    .A2(_10207_));
 sg13g2_buf_2 _18067_ (.A(_11175_),
    .X(_11176_));
 sg13g2_buf_1 _18068_ (.A(_11176_),
    .X(_11177_));
 sg13g2_a221oi_1 _18069_ (.B2(_11158_),
    .C1(net203),
    .B1(_11155_),
    .A1(_11028_),
    .Y(_11178_),
    .A2(_11040_));
 sg13g2_a221oi_1 _18070_ (.B2(_11154_),
    .C1(_11178_),
    .B1(_11128_),
    .A1(_11001_),
    .Y(_11179_),
    .A2(_11041_));
 sg13g2_buf_1 _18071_ (.A(_11179_),
    .X(_11180_));
 sg13g2_nor2_1 _18072_ (.A(_11072_),
    .B(net119),
    .Y(_11181_));
 sg13g2_nand2_1 _18073_ (.Y(_11182_),
    .A(_11153_),
    .B(_11127_));
 sg13g2_nor2_1 _18074_ (.A(_11181_),
    .B(_11182_),
    .Y(_11183_));
 sg13g2_a21oi_1 _18075_ (.A1(_11073_),
    .A2(net119),
    .Y(_11184_),
    .B1(_11183_));
 sg13g2_nand2b_1 _18076_ (.Y(_11185_),
    .B(_11184_),
    .A_N(_11180_));
 sg13g2_buf_1 _18077_ (.A(_09385_),
    .X(_11186_));
 sg13g2_inv_1 _18078_ (.Y(_11187_),
    .A(\cpu.ex.r_14[15] ));
 sg13g2_buf_2 _18079_ (.A(\cpu.ex.mmu_read[15] ),
    .X(_11188_));
 sg13g2_nand3_1 _18080_ (.B(_10973_),
    .C(_10312_),
    .A(_11188_),
    .Y(_11189_));
 sg13g2_o21ai_1 _18081_ (.B1(_11189_),
    .Y(_11190_),
    .A1(_11187_),
    .A2(_10401_));
 sg13g2_buf_1 _18082_ (.A(\cpu.ex.r_sp[15] ),
    .X(_11191_));
 sg13g2_and2_1 _18083_ (.A(\cpu.ex.r_10[15] ),
    .B(net659),
    .X(_11192_));
 sg13g2_a21oi_1 _18084_ (.A1(_11191_),
    .A2(_10391_),
    .Y(_11193_),
    .B1(_11192_));
 sg13g2_nor3_1 _18085_ (.A(net590),
    .B(_10405_),
    .C(_11193_),
    .Y(_11194_));
 sg13g2_a21o_1 _18086_ (.A2(_11190_),
    .A1(net591),
    .B1(_11194_),
    .X(_11195_));
 sg13g2_and2_1 _18087_ (.A(net592),
    .B(_10155_),
    .X(_11196_));
 sg13g2_and3_1 _18088_ (.X(_11197_),
    .A(\cpu.ex.r_13[15] ),
    .B(net593),
    .C(_11058_));
 sg13g2_a221oi_1 _18089_ (.B2(\cpu.ex.r_9[15] ),
    .C1(_11197_),
    .B1(_10413_),
    .A1(\cpu.ex.r_mult[31] ),
    .Y(_11198_),
    .A2(_11196_));
 sg13g2_a221oi_1 _18090_ (.B2(\cpu.ex.r_8[15] ),
    .C1(net524),
    .B1(_10413_),
    .A1(\cpu.ex.r_stmp[15] ),
    .Y(_11199_),
    .A2(_11196_));
 sg13g2_a21oi_1 _18091_ (.A1(net524),
    .A2(_11198_),
    .Y(_11200_),
    .B1(_11199_));
 sg13g2_a22oi_1 _18092_ (.Y(_11201_),
    .B1(_10629_),
    .B2(\cpu.ex.r_12[15] ),
    .A2(_10972_),
    .A1(\cpu.ex.r_lr[15] ));
 sg13g2_nor2_1 _18093_ (.A(net592),
    .B(_11201_),
    .Y(_11202_));
 sg13g2_inv_1 _18094_ (.Y(_11203_),
    .A(_00251_));
 sg13g2_mux2_1 _18095_ (.A0(\cpu.ex.r_epc[15] ),
    .A1(\cpu.ex.r_11[15] ),
    .S(_10507_),
    .X(_11204_));
 sg13g2_a22oi_1 _18096_ (.Y(_11205_),
    .B1(_11204_),
    .B2(_10519_),
    .A2(_10433_),
    .A1(_11203_));
 sg13g2_nor2_1 _18097_ (.A(_10152_),
    .B(_11205_),
    .Y(_11206_));
 sg13g2_or4_1 _18098_ (.A(_11195_),
    .B(_11200_),
    .C(_11202_),
    .D(_11206_),
    .X(_11207_));
 sg13g2_a22oi_1 _18099_ (.Y(_11208_),
    .B1(_10792_),
    .B2(_11207_),
    .A2(net459),
    .A1(net731));
 sg13g2_nor2_1 _18100_ (.A(_10424_),
    .B(\cpu.dec.imm[15] ),
    .Y(_11209_));
 sg13g2_a21oi_1 _18101_ (.A1(net1006),
    .A2(_11208_),
    .Y(_11210_),
    .B1(_11209_));
 sg13g2_nor2_1 _18102_ (.A(net860),
    .B(_00178_),
    .Y(_11211_));
 sg13g2_a21o_1 _18103_ (.A2(_11210_),
    .A1(net860),
    .B1(_11211_),
    .X(_11212_));
 sg13g2_buf_1 _18104_ (.A(_11212_),
    .X(_11213_));
 sg13g2_inv_1 _18105_ (.Y(_11214_),
    .A(_00178_));
 sg13g2_mux4_1 _18106_ (.S0(net752),
    .A0(\cpu.ex.r_lr[15] ),
    .A1(\cpu.ex.r_epc[15] ),
    .A2(\cpu.ex.r_9[15] ),
    .A3(\cpu.ex.r_11[15] ),
    .S1(net655),
    .X(_11215_));
 sg13g2_and2_1 _18107_ (.A(_10219_),
    .B(_11215_),
    .X(_11216_));
 sg13g2_mux2_1 _18108_ (.A0(\cpu.ex.r_12[15] ),
    .A1(\cpu.ex.r_13[15] ),
    .S(net862),
    .X(_11217_));
 sg13g2_mux2_1 _18109_ (.A0(\cpu.ex.r_10[15] ),
    .A1(\cpu.ex.r_14[15] ),
    .S(net750),
    .X(_11218_));
 sg13g2_a22oi_1 _18110_ (.Y(_11219_),
    .B1(_11218_),
    .B2(net662),
    .A2(_11217_),
    .A1(_10231_));
 sg13g2_nand3_1 _18111_ (.B(_10361_),
    .C(_10229_),
    .A(_11191_),
    .Y(_11220_));
 sg13g2_o21ai_1 _18112_ (.B1(_11220_),
    .Y(_11221_),
    .A1(net748),
    .A2(_11219_));
 sg13g2_nand3_1 _18113_ (.B(\cpu.ex.r_8[15] ),
    .C(net665),
    .A(net664),
    .Y(_11222_));
 sg13g2_nand3_1 _18114_ (.B(\cpu.ex.r_stmp[15] ),
    .C(net669),
    .A(net671),
    .Y(_11223_));
 sg13g2_a21oi_1 _18115_ (.A1(_11222_),
    .A2(_11223_),
    .Y(_11224_),
    .B1(net670));
 sg13g2_nor2b_1 _18116_ (.A(_00251_),
    .B_N(net655),
    .Y(_11225_));
 sg13g2_nor2b_1 _18117_ (.A(net655),
    .B_N(\cpu.ex.r_mult[31] ),
    .Y(_11226_));
 sg13g2_o21ai_1 _18118_ (.B1(net671),
    .Y(_11227_),
    .A1(_11225_),
    .A2(_11226_));
 sg13g2_nand2_1 _18119_ (.Y(_11228_),
    .A(_11188_),
    .B(_10215_));
 sg13g2_a21oi_1 _18120_ (.A1(_11227_),
    .A2(_11228_),
    .Y(_11229_),
    .B1(_10655_));
 sg13g2_nor4_1 _18121_ (.A(_11216_),
    .B(_11221_),
    .C(_11224_),
    .D(_11229_),
    .Y(_11230_));
 sg13g2_nor2_1 _18122_ (.A(net731),
    .B(_10047_),
    .Y(_11231_));
 sg13g2_a21oi_2 _18123_ (.B1(_11231_),
    .Y(_11232_),
    .A2(_11230_),
    .A1(net527));
 sg13g2_mux2_1 _18124_ (.A0(_11214_),
    .A1(_11232_),
    .S(net227),
    .X(_11233_));
 sg13g2_buf_2 _18125_ (.A(_11233_),
    .X(_11234_));
 sg13g2_buf_1 _18126_ (.A(_11234_),
    .X(_11235_));
 sg13g2_buf_1 _18127_ (.A(net146),
    .X(_11236_));
 sg13g2_nor2_1 _18128_ (.A(net202),
    .B(net118),
    .Y(_11237_));
 sg13g2_nand2_1 _18129_ (.Y(_11238_),
    .A(net202),
    .B(net146));
 sg13g2_o21ai_1 _18130_ (.B1(_11238_),
    .Y(_11239_),
    .A1(_11185_),
    .A2(_11237_));
 sg13g2_o21ai_1 _18131_ (.B1(_10947_),
    .Y(_11240_),
    .A1(_11029_),
    .A2(_11031_));
 sg13g2_inv_2 _18132_ (.Y(_11241_),
    .A(_10947_));
 sg13g2_nand3_1 _18133_ (.B(_10884_),
    .C(_10911_),
    .A(_11241_),
    .Y(_11242_));
 sg13g2_buf_1 _18134_ (.A(_10743_),
    .X(_11243_));
 sg13g2_buf_1 _18135_ (.A(_10646_),
    .X(_11244_));
 sg13g2_nand2_1 _18136_ (.Y(_11245_),
    .A(net1004),
    .B(net226));
 sg13g2_a21oi_1 _18137_ (.A1(_11240_),
    .A2(_11242_),
    .Y(_11246_),
    .B1(_11245_));
 sg13g2_nor4_1 _18138_ (.A(net1004),
    .B(_11241_),
    .C(net181),
    .D(net226),
    .Y(_11247_));
 sg13g2_buf_1 _18139_ (.A(_09146_),
    .X(_11248_));
 sg13g2_buf_1 _18140_ (.A(net652),
    .X(_11249_));
 sg13g2_o21ai_1 _18141_ (.B1(net588),
    .Y(_11250_),
    .A1(_11246_),
    .A2(_11247_));
 sg13g2_o21ai_1 _18142_ (.B1(net652),
    .Y(_11251_),
    .A1(_11243_),
    .A2(_10947_));
 sg13g2_nand3_1 _18143_ (.B(net205),
    .C(_11251_),
    .A(net181),
    .Y(_11252_));
 sg13g2_inv_2 _18144_ (.Y(_11253_),
    .A(_10835_));
 sg13g2_and2_1 _18145_ (.A(_10969_),
    .B(_10994_),
    .X(_11254_));
 sg13g2_buf_2 _18146_ (.A(_11254_),
    .X(_11255_));
 sg13g2_buf_1 _18147_ (.A(net248),
    .X(_11256_));
 sg13g2_nor4_1 _18148_ (.A(net1097),
    .B(_11253_),
    .C(_11255_),
    .D(net225),
    .Y(_11257_));
 sg13g2_a21o_1 _18149_ (.A2(_10994_),
    .A1(_10969_),
    .B1(_11253_),
    .X(_11258_));
 sg13g2_nand3_1 _18150_ (.B(_10969_),
    .C(_10994_),
    .A(_11253_),
    .Y(_11259_));
 sg13g2_nand2_1 _18151_ (.Y(_11260_),
    .A(net1097),
    .B(net225));
 sg13g2_a21oi_1 _18152_ (.A1(_11258_),
    .A2(_11259_),
    .Y(_11261_),
    .B1(_11260_));
 sg13g2_o21ai_1 _18153_ (.B1(net588),
    .Y(_11262_),
    .A1(_11257_),
    .A2(_11261_));
 sg13g2_buf_1 _18154_ (.A(_11255_),
    .X(_11263_));
 sg13g2_o21ai_1 _18155_ (.B1(net588),
    .Y(_11264_),
    .A1(_10627_),
    .A2(_10835_));
 sg13g2_nand3_1 _18156_ (.B(_10878_),
    .C(_11264_),
    .A(net145),
    .Y(_11265_));
 sg13g2_a22oi_1 _18157_ (.Y(_11266_),
    .B1(_11262_),
    .B2(_11265_),
    .A2(_11252_),
    .A1(_11250_));
 sg13g2_buf_1 _18158_ (.A(_09153_),
    .X(_11267_));
 sg13g2_nand2b_1 _18159_ (.Y(_11268_),
    .B(net249),
    .A_N(net1096));
 sg13g2_buf_1 _18160_ (.A(_10478_),
    .X(_11269_));
 sg13g2_buf_1 _18161_ (.A(_10544_),
    .X(_11270_));
 sg13g2_a21oi_1 _18162_ (.A1(_10133_),
    .A2(_10536_),
    .Y(_11271_),
    .B1(_10538_));
 sg13g2_nor2_1 _18163_ (.A(net1002),
    .B(_11271_),
    .Y(_11272_));
 sg13g2_nor2_1 _18164_ (.A(_10571_),
    .B(_10574_),
    .Y(_11273_));
 sg13g2_buf_1 _18165_ (.A(_11273_),
    .X(_11274_));
 sg13g2_buf_1 _18166_ (.A(_10365_),
    .X(_11275_));
 sg13g2_a22oi_1 _18167_ (.Y(_11276_),
    .B1(net302),
    .B2(_11275_),
    .A2(_11271_),
    .A1(_10544_));
 sg13g2_buf_1 _18168_ (.A(_10714_),
    .X(_11277_));
 sg13g2_o21ai_1 _18169_ (.B1(net201),
    .Y(_11278_),
    .A1(_11272_),
    .A2(_11276_));
 sg13g2_nor3_1 _18170_ (.A(net201),
    .B(_11272_),
    .C(_11276_),
    .Y(_11279_));
 sg13g2_a21o_1 _18171_ (.A2(_11278_),
    .A1(_11269_),
    .B1(_11279_),
    .X(_11280_));
 sg13g2_and2_1 _18172_ (.A(net1096),
    .B(net228),
    .X(_11281_));
 sg13g2_a21oi_1 _18173_ (.A1(_11268_),
    .A2(_11280_),
    .Y(_11282_),
    .B1(_11281_));
 sg13g2_xnor2_1 _18174_ (.Y(_11283_),
    .A(net1096),
    .B(net228));
 sg13g2_buf_8 _18175_ (.A(_10809_),
    .X(_11284_));
 sg13g2_nand2b_1 _18176_ (.Y(_11285_),
    .B(_10478_),
    .A_N(net224));
 sg13g2_inv_1 _18177_ (.Y(_11286_),
    .A(_10478_));
 sg13g2_nand4_1 _18178_ (.B(net1096),
    .C(net224),
    .A(_11286_),
    .Y(_11287_),
    .D(net249));
 sg13g2_o21ai_1 _18179_ (.B1(_11287_),
    .Y(_11288_),
    .A1(_11283_),
    .A2(_11285_));
 sg13g2_and2_1 _18180_ (.A(_10809_),
    .B(_10799_),
    .X(_11289_));
 sg13g2_buf_2 _18181_ (.A(_11289_),
    .X(_11290_));
 sg13g2_o21ai_1 _18182_ (.B1(net652),
    .Y(_11291_),
    .A1(_11269_),
    .A2(net1096));
 sg13g2_a22oi_1 _18183_ (.Y(_11292_),
    .B1(_11290_),
    .B2(_11291_),
    .A2(_11288_),
    .A1(_11248_));
 sg13g2_buf_1 _18184_ (.A(_10576_),
    .X(_11293_));
 sg13g2_nand2_1 _18185_ (.Y(_11294_),
    .A(net1001),
    .B(net247));
 sg13g2_buf_1 _18186_ (.A(_11271_),
    .X(_11295_));
 sg13g2_xnor2_1 _18187_ (.Y(_11296_),
    .A(net1002),
    .B(net246));
 sg13g2_inv_1 _18188_ (.Y(_11297_),
    .A(net1001));
 sg13g2_nand4_1 _18189_ (.B(net1002),
    .C(net230),
    .A(_11297_),
    .Y(_11298_),
    .D(net302));
 sg13g2_o21ai_1 _18190_ (.B1(_11298_),
    .Y(_11299_),
    .A1(_11294_),
    .A2(_11296_));
 sg13g2_nor2_1 _18191_ (.A(net230),
    .B(net247),
    .Y(_11300_));
 sg13g2_o21ai_1 _18192_ (.B1(net652),
    .Y(_11301_),
    .A1(net1001),
    .A2(net1002));
 sg13g2_a22oi_1 _18193_ (.Y(_11302_),
    .B1(_11300_),
    .B2(_11301_),
    .A2(_11299_),
    .A1(net652));
 sg13g2_or2_1 _18194_ (.X(_11303_),
    .B(_11302_),
    .A(_11292_));
 sg13g2_o21ai_1 _18195_ (.B1(_11303_),
    .Y(_11304_),
    .A1(_11267_),
    .A2(_11282_));
 sg13g2_a21oi_1 _18196_ (.A1(_11241_),
    .A2(net183),
    .Y(_11305_),
    .B1(_11253_));
 sg13g2_inv_1 _18197_ (.Y(_11306_),
    .A(net1097));
 sg13g2_nand2_1 _18198_ (.Y(_11307_),
    .A(_11306_),
    .B(net248));
 sg13g2_inv_1 _18199_ (.Y(_11308_),
    .A(_10743_));
 sg13g2_nor2_1 _18200_ (.A(_11308_),
    .B(_10646_),
    .Y(_11309_));
 sg13g2_nor2_1 _18201_ (.A(_11306_),
    .B(net248),
    .Y(_11310_));
 sg13g2_a21oi_1 _18202_ (.A1(_11307_),
    .A2(_11309_),
    .Y(_11311_),
    .B1(_11310_));
 sg13g2_o21ai_1 _18203_ (.B1(net182),
    .Y(_11312_),
    .A1(_09153_),
    .A2(_11311_));
 sg13g2_nor4_1 _18204_ (.A(_11241_),
    .B(_09153_),
    .C(net182),
    .D(_11311_),
    .Y(_11313_));
 sg13g2_a221oi_1 _18205_ (.B2(_11312_),
    .C1(_11313_),
    .B1(_11305_),
    .A1(_10947_),
    .Y(_11314_),
    .A2(net181));
 sg13g2_nor2_1 _18206_ (.A(_09153_),
    .B(_11311_),
    .Y(_11315_));
 sg13g2_nand3_1 _18207_ (.B(_11255_),
    .C(_11315_),
    .A(net181),
    .Y(_11316_));
 sg13g2_o21ai_1 _18208_ (.B1(_11316_),
    .Y(_11317_),
    .A1(net651),
    .A2(_11314_));
 sg13g2_buf_1 _18209_ (.A(_11317_),
    .X(_11318_));
 sg13g2_a21oi_1 _18210_ (.A1(_11266_),
    .A2(_11304_),
    .Y(_11319_),
    .B1(_11318_));
 sg13g2_nor2_1 _18211_ (.A(_11267_),
    .B(_11282_),
    .Y(_11320_));
 sg13g2_mux2_1 _18212_ (.A0(_11002_),
    .A1(_11068_),
    .S(net1109),
    .X(_11321_));
 sg13g2_nor3_1 _18213_ (.A(_09147_),
    .B(_09121_),
    .C(net1031),
    .Y(_11322_));
 sg13g2_buf_1 _18214_ (.A(_11322_),
    .X(_11323_));
 sg13g2_nor2_1 _18215_ (.A(_09153_),
    .B(net730),
    .Y(_11324_));
 sg13g2_buf_2 _18216_ (.A(_11324_),
    .X(_11325_));
 sg13g2_inv_1 _18217_ (.Y(_11326_),
    .A(_09140_));
 sg13g2_nor2_1 _18218_ (.A(_09141_),
    .B(\cpu.ex.r_mult_off[1] ),
    .Y(_11327_));
 sg13g2_nand2_1 _18219_ (.Y(_11328_),
    .A(_11326_),
    .B(_11327_));
 sg13g2_nand2_1 _18220_ (.Y(_11329_),
    .A(_11325_),
    .B(_11328_));
 sg13g2_nand2_1 _18221_ (.Y(_11330_),
    .A(_09146_),
    .B(_09149_));
 sg13g2_inv_1 _18222_ (.Y(_11331_),
    .A(_11125_));
 sg13g2_a21oi_1 _18223_ (.A1(net1109),
    .A2(_11331_),
    .Y(_11332_),
    .B1(_09141_));
 sg13g2_nor3_1 _18224_ (.A(_11326_),
    .B(_11330_),
    .C(_11332_),
    .Y(_11333_));
 sg13g2_a21o_1 _18225_ (.A2(_11329_),
    .A1(_11214_),
    .B1(_11333_),
    .X(_11334_));
 sg13g2_o21ai_1 _18226_ (.B1(_11334_),
    .Y(_11335_),
    .A1(\cpu.ex.c_mult_off[0] ),
    .A2(_11321_));
 sg13g2_nand2_1 _18227_ (.Y(_11336_),
    .A(net303),
    .B(_11335_));
 sg13g2_and4_1 _18228_ (.A(net1109),
    .B(_09140_),
    .C(_11325_),
    .D(_11122_),
    .X(_11337_));
 sg13g2_o21ai_1 _18229_ (.B1(_09140_),
    .Y(_11338_),
    .A1(_09141_),
    .A2(net1109));
 sg13g2_and3_1 _18230_ (.X(_11339_),
    .A(_11325_),
    .B(_11328_),
    .C(_11338_));
 sg13g2_buf_1 _18231_ (.A(_11339_),
    .X(_11340_));
 sg13g2_nor2_1 _18232_ (.A(\cpu.ex.c_mult_off[0] ),
    .B(_11340_),
    .Y(_11341_));
 sg13g2_a221oi_1 _18233_ (.B2(_11337_),
    .C1(_11341_),
    .B1(_11121_),
    .A1(_11329_),
    .Y(_11342_),
    .A2(_11232_));
 sg13g2_nand3_1 _18234_ (.B(net1109),
    .C(_11325_),
    .A(_09141_),
    .Y(_11343_));
 sg13g2_nor3_1 _18235_ (.A(_09139_),
    .B(\cpu.ex.c_mult_off[0] ),
    .C(net594),
    .Y(_11344_));
 sg13g2_nor4_1 _18236_ (.A(net679),
    .B(_09139_),
    .C(\cpu.ex.c_mult_off[0] ),
    .D(net527),
    .Y(_11345_));
 sg13g2_a21oi_1 _18237_ (.A1(_11022_),
    .A2(_11344_),
    .Y(_11346_),
    .B1(_11345_));
 sg13g2_o21ai_1 _18238_ (.B1(_11346_),
    .Y(_11347_),
    .A1(_11096_),
    .A2(_11343_));
 sg13g2_o21ai_1 _18239_ (.B1(net250),
    .Y(_11348_),
    .A1(_11342_),
    .A2(_11347_));
 sg13g2_and2_1 _18240_ (.A(_10832_),
    .B(_10853_),
    .X(_11349_));
 sg13g2_mux2_1 _18241_ (.A0(_10874_),
    .A1(_11349_),
    .S(_10125_),
    .X(_11350_));
 sg13g2_buf_2 _18242_ (.A(_11350_),
    .X(_11351_));
 sg13g2_xnor2_1 _18243_ (.Y(_11352_),
    .A(_09141_),
    .B(net1109));
 sg13g2_nor3_1 _18244_ (.A(_09141_),
    .B(_11330_),
    .C(_11352_),
    .Y(_11353_));
 sg13g2_and2_1 _18245_ (.A(_11340_),
    .B(_11353_),
    .X(_11354_));
 sg13g2_xor2_1 _18246_ (.B(_11328_),
    .A(\cpu.ex.r_mult_off[3] ),
    .X(_11355_));
 sg13g2_nand2_1 _18247_ (.Y(\cpu.ex.c_mult_off[3] ),
    .A(_11325_),
    .B(_11355_));
 sg13g2_inv_1 _18248_ (.Y(_11356_),
    .A(\cpu.ex.c_mult_off[3] ));
 sg13g2_a221oi_1 _18249_ (.B2(_11354_),
    .C1(_11356_),
    .B1(_11351_),
    .A1(_11336_),
    .Y(_11357_),
    .A2(_11348_));
 sg13g2_inv_1 _18250_ (.Y(_11358_),
    .A(_11343_));
 sg13g2_nand3_1 _18251_ (.B(_11358_),
    .C(net204),
    .A(_11340_),
    .Y(_11359_));
 sg13g2_nor2_1 _18252_ (.A(net1109),
    .B(\cpu.ex.c_mult_off[0] ),
    .Y(_11360_));
 sg13g2_nand2b_1 _18253_ (.Y(_11361_),
    .B(_11325_),
    .A_N(_11327_));
 sg13g2_a221oi_1 _18254_ (.B2(_10936_),
    .C1(_10338_),
    .B1(_11361_),
    .A1(_11360_),
    .Y(_11362_),
    .A2(_10675_));
 sg13g2_nand2_1 _18255_ (.Y(_11363_),
    .A(_10882_),
    .B(_11361_));
 sg13g2_nand2_1 _18256_ (.Y(_11364_),
    .A(_10643_),
    .B(_11360_));
 sg13g2_nand3_1 _18257_ (.B(_11363_),
    .C(_11364_),
    .A(net303),
    .Y(_11365_));
 sg13g2_nand3b_1 _18258_ (.B(_11365_),
    .C(_11340_),
    .Y(_11366_),
    .A_N(_11362_));
 sg13g2_and3_1 _18259_ (.X(_11367_),
    .A(_11357_),
    .B(_11359_),
    .C(_11366_));
 sg13g2_buf_1 _18260_ (.A(_11367_),
    .X(_11368_));
 sg13g2_buf_1 _18261_ (.A(_10334_),
    .X(_11369_));
 sg13g2_nand2_1 _18262_ (.Y(_11370_),
    .A(_10153_),
    .B(_09146_));
 sg13g2_o21ai_1 _18263_ (.B1(net374),
    .Y(_11371_),
    .A1(net370),
    .A2(_11370_));
 sg13g2_inv_1 _18264_ (.Y(_11372_),
    .A(_11371_));
 sg13g2_nor2_1 _18265_ (.A(_11330_),
    .B(_11352_),
    .Y(_11373_));
 sg13g2_inv_1 _18266_ (.Y(\cpu.ex.c_mult_off[1] ),
    .A(_11373_));
 sg13g2_mux4_1 _18267_ (.S0(\cpu.ex.c_mult_off[1] ),
    .A0(net1050),
    .A1(_10814_),
    .A2(_10605_),
    .A3(_10815_),
    .S1(net250),
    .X(_11374_));
 sg13g2_nand2b_1 _18268_ (.Y(_11375_),
    .B(\cpu.ex.c_mult_off[1] ),
    .A_N(net207));
 sg13g2_and2_1 _18269_ (.A(_10472_),
    .B(_10503_),
    .X(_11376_));
 sg13g2_buf_1 _18270_ (.A(_11376_),
    .X(_11377_));
 sg13g2_a221oi_1 _18271_ (.B2(_11377_),
    .C1(_11340_),
    .B1(_11373_),
    .A1(_09141_),
    .Y(_11378_),
    .A2(_11325_));
 sg13g2_a221oi_1 _18272_ (.B2(_11378_),
    .C1(_11371_),
    .B1(_11375_),
    .A1(_11341_),
    .Y(_11379_),
    .A2(_11374_));
 sg13g2_o21ai_1 _18273_ (.B1(_10117_),
    .Y(_11380_),
    .A1(_08131_),
    .A2(net460));
 sg13g2_nor2_1 _18274_ (.A(_10121_),
    .B(_10326_),
    .Y(_11381_));
 sg13g2_a22oi_1 _18275_ (.Y(_11382_),
    .B1(_10258_),
    .B2(_10676_),
    .A2(_11381_),
    .A1(_11380_));
 sg13g2_buf_1 _18276_ (.A(_11382_),
    .X(_11383_));
 sg13g2_a22oi_1 _18277_ (.Y(_11384_),
    .B1(_10291_),
    .B2(net251),
    .A2(_10264_),
    .A1(_10259_));
 sg13g2_buf_8 _18278_ (.A(_11384_),
    .X(_11385_));
 sg13g2_inv_1 _18279_ (.Y(\cpu.ex.c_mult_off[2] ),
    .A(_11340_));
 sg13g2_a221oi_1 _18280_ (.B2(_11360_),
    .C1(\cpu.ex.c_mult_off[2] ),
    .B1(_11385_),
    .A1(_11353_),
    .Y(_11386_),
    .A2(_11383_));
 sg13g2_or2_1 _18281_ (.X(_11387_),
    .B(_10103_),
    .A(_10048_));
 sg13g2_mux2_1 _18282_ (.A0(_00269_),
    .A1(_11387_),
    .S(_10126_),
    .X(_11388_));
 sg13g2_buf_2 _18283_ (.A(_11388_),
    .X(_11389_));
 sg13g2_a22oi_1 _18284_ (.Y(_11390_),
    .B1(_11389_),
    .B2(_11358_),
    .A2(_10390_),
    .A1(_11361_));
 sg13g2_a21oi_2 _18285_ (.B1(\cpu.ex.c_mult_off[3] ),
    .Y(_11391_),
    .A2(_11390_),
    .A1(_11386_));
 sg13g2_and2_1 _18286_ (.A(net370),
    .B(_11370_),
    .X(_11392_));
 sg13g2_a221oi_1 _18287_ (.B2(_11391_),
    .C1(_11392_),
    .B1(_11379_),
    .A1(_11368_),
    .Y(_11393_),
    .A2(_11372_));
 sg13g2_buf_2 _18288_ (.A(_11393_),
    .X(_11394_));
 sg13g2_buf_1 _18289_ (.A(_10240_),
    .X(_11395_));
 sg13g2_nand2_1 _18290_ (.Y(_11396_),
    .A(net1000),
    .B(net652));
 sg13g2_a21o_1 _18291_ (.A2(_10423_),
    .A1(_10345_),
    .B1(_10429_),
    .X(_11397_));
 sg13g2_buf_1 _18292_ (.A(_11397_),
    .X(_11398_));
 sg13g2_buf_1 _18293_ (.A(_11398_),
    .X(_11399_));
 sg13g2_buf_1 _18294_ (.A(net372),
    .X(_11400_));
 sg13g2_and2_1 _18295_ (.A(_10075_),
    .B(_09146_),
    .X(_11401_));
 sg13g2_buf_1 _18296_ (.A(_11401_),
    .X(_11402_));
 sg13g2_and2_1 _18297_ (.A(_10456_),
    .B(_10461_),
    .X(_11403_));
 sg13g2_buf_1 _18298_ (.A(_11403_),
    .X(_11404_));
 sg13g2_buf_1 _18299_ (.A(_11404_),
    .X(_11405_));
 sg13g2_o21ai_1 _18300_ (.B1(net299),
    .Y(_11406_),
    .A1(net300),
    .A2(_11402_));
 sg13g2_o21ai_1 _18301_ (.B1(_11406_),
    .Y(_11407_),
    .A1(_11396_),
    .A2(net301));
 sg13g2_and2_1 _18302_ (.A(_11394_),
    .B(_11407_),
    .X(_11408_));
 sg13g2_buf_1 _18303_ (.A(_10075_),
    .X(_11409_));
 sg13g2_and3_1 _18304_ (.X(_11410_),
    .A(net1000),
    .B(net999),
    .C(_09146_));
 sg13g2_buf_1 _18305_ (.A(_11410_),
    .X(_11411_));
 sg13g2_nor3_1 _18306_ (.A(_11396_),
    .B(net301),
    .C(net371),
    .Y(_11412_));
 sg13g2_a221oi_1 _18307_ (.B2(net372),
    .C1(_11412_),
    .B1(_11402_),
    .A1(_11411_),
    .Y(_11413_),
    .A2(net299));
 sg13g2_buf_1 _18308_ (.A(_11413_),
    .X(_11414_));
 sg13g2_inv_1 _18309_ (.Y(_11415_),
    .A(_11414_));
 sg13g2_a21o_1 _18310_ (.A2(_11411_),
    .A1(_11394_),
    .B1(_11415_),
    .X(_11416_));
 sg13g2_nor4_2 _18311_ (.A(_11318_),
    .B(_11320_),
    .C(_11408_),
    .Y(_11417_),
    .D(_11416_));
 sg13g2_buf_1 _18312_ (.A(net588),
    .X(_11418_));
 sg13g2_o21ai_1 _18313_ (.B1(_11014_),
    .Y(_11419_),
    .A1(_11129_),
    .A2(_11151_));
 sg13g2_inv_2 _18314_ (.Y(_11420_),
    .A(_11014_));
 sg13g2_nand2_1 _18315_ (.Y(_11421_),
    .A(net1005),
    .B(_11331_));
 sg13g2_nand3_1 _18316_ (.B(_11130_),
    .C(_11149_),
    .A(_10795_),
    .Y(_11422_));
 sg13g2_buf_1 _18317_ (.A(_11422_),
    .X(_11423_));
 sg13g2_nand3_1 _18318_ (.B(_11421_),
    .C(_11423_),
    .A(_11420_),
    .Y(_11424_));
 sg13g2_inv_1 _18319_ (.Y(_11425_),
    .A(_11173_));
 sg13g2_a21oi_1 _18320_ (.A1(\cpu.dec.imm[12] ),
    .A2(_10207_),
    .Y(_11426_),
    .B1(_11174_));
 sg13g2_o21ai_1 _18321_ (.B1(_11426_),
    .Y(_11427_),
    .A1(net743),
    .A2(_11425_));
 sg13g2_buf_2 _18322_ (.A(_11427_),
    .X(_11428_));
 sg13g2_nand2_1 _18323_ (.Y(_11429_),
    .A(_10902_),
    .B(_11428_));
 sg13g2_a21oi_1 _18324_ (.A1(_11419_),
    .A2(_11424_),
    .Y(_11430_),
    .B1(_11429_));
 sg13g2_buf_1 _18325_ (.A(_10902_),
    .X(_11431_));
 sg13g2_nor4_1 _18326_ (.A(net998),
    .B(_11420_),
    .C(_11153_),
    .D(_11428_),
    .Y(_11432_));
 sg13g2_o21ai_1 _18327_ (.B1(_11249_),
    .Y(_11433_),
    .A1(_11430_),
    .A2(_11432_));
 sg13g2_nand2_1 _18328_ (.Y(_11434_),
    .A(_11421_),
    .B(_11423_));
 sg13g2_buf_1 _18329_ (.A(_11434_),
    .X(_11435_));
 sg13g2_nor2_1 _18330_ (.A(net180),
    .B(_11428_),
    .Y(_11436_));
 sg13g2_o21ai_1 _18331_ (.B1(_11249_),
    .Y(_11437_),
    .A1(_11431_),
    .A2(_11014_));
 sg13g2_nand2_1 _18332_ (.Y(_11438_),
    .A(_11436_),
    .B(_11437_));
 sg13g2_nand2_1 _18333_ (.Y(_11439_),
    .A(_11112_),
    .B(net588));
 sg13g2_xnor2_1 _18334_ (.Y(_11440_),
    .A(_11071_),
    .B(_11439_));
 sg13g2_a21oi_1 _18335_ (.A1(_11433_),
    .A2(_11438_),
    .Y(_11441_),
    .B1(_11440_));
 sg13g2_nand3_1 _18336_ (.B(net523),
    .C(_11441_),
    .A(_11047_),
    .Y(_11442_));
 sg13g2_nor3_1 _18337_ (.A(_11319_),
    .B(_11417_),
    .C(_11442_),
    .Y(_11443_));
 sg13g2_a21oi_1 _18338_ (.A1(net860),
    .A2(_11210_),
    .Y(_11444_),
    .B1(_11211_));
 sg13g2_buf_1 _18339_ (.A(_11444_),
    .X(_11445_));
 sg13g2_a21o_1 _18340_ (.A2(_11304_),
    .A1(_11266_),
    .B1(_11318_),
    .X(_11446_));
 sg13g2_or4_1 _18341_ (.A(_11318_),
    .B(_11320_),
    .C(_11408_),
    .D(_11416_),
    .X(_11447_));
 sg13g2_and4_1 _18342_ (.A(net199),
    .B(_11446_),
    .C(_11447_),
    .D(_11441_),
    .X(_11448_));
 sg13g2_nand2_1 _18343_ (.Y(_11449_),
    .A(_11047_),
    .B(net523));
 sg13g2_nor2_1 _18344_ (.A(net202),
    .B(_11449_),
    .Y(_11450_));
 sg13g2_buf_1 _18345_ (.A(_11071_),
    .X(_11451_));
 sg13g2_nand2_1 _18346_ (.Y(_11452_),
    .A(_11420_),
    .B(net180));
 sg13g2_and2_1 _18347_ (.A(net998),
    .B(net203),
    .X(_11453_));
 sg13g2_nor2_1 _18348_ (.A(_11420_),
    .B(net180),
    .Y(_11454_));
 sg13g2_a21oi_1 _18349_ (.A1(_11452_),
    .A2(_11453_),
    .Y(_11455_),
    .B1(_11454_));
 sg13g2_inv_1 _18350_ (.Y(_11456_),
    .A(_11112_));
 sg13g2_a21oi_1 _18351_ (.A1(net179),
    .A2(_11455_),
    .Y(_11457_),
    .B1(_11456_));
 sg13g2_nor2_1 _18352_ (.A(net179),
    .B(_11455_),
    .Y(_11458_));
 sg13g2_o21ai_1 _18353_ (.B1(net523),
    .Y(_11459_),
    .A1(_11457_),
    .A2(_11458_));
 sg13g2_a21oi_1 _18354_ (.A1(net202),
    .A2(_11449_),
    .Y(_11460_),
    .B1(_11459_));
 sg13g2_nor4_1 _18355_ (.A(_11443_),
    .B(_11448_),
    .C(_11450_),
    .D(_11460_),
    .Y(_11461_));
 sg13g2_buf_2 _18356_ (.A(_11461_),
    .X(_11462_));
 sg13g2_nand2b_1 _18357_ (.Y(_11463_),
    .B(_10030_),
    .A_N(_10028_));
 sg13g2_buf_1 _18358_ (.A(_11463_),
    .X(_11464_));
 sg13g2_buf_1 _18359_ (.A(_11464_),
    .X(_11465_));
 sg13g2_buf_1 _18360_ (.A(net374),
    .X(_11466_));
 sg13g2_buf_1 _18361_ (.A(net298),
    .X(_11467_));
 sg13g2_a22oi_1 _18362_ (.Y(_11468_),
    .B1(_11375_),
    .B2(_11378_),
    .A2(_11374_),
    .A1(_11341_));
 sg13g2_a21oi_1 _18363_ (.A1(_11468_),
    .A2(_11391_),
    .Y(_11469_),
    .B1(_11368_));
 sg13g2_buf_8 _18364_ (.A(_11469_),
    .X(_11470_));
 sg13g2_buf_1 _18365_ (.A(_11470_),
    .X(_11471_));
 sg13g2_buf_1 _18366_ (.A(_09155_),
    .X(_11472_));
 sg13g2_buf_1 _18367_ (.A(net730),
    .X(_11473_));
 sg13g2_nor2_1 _18368_ (.A(net997),
    .B(net650),
    .Y(_11474_));
 sg13g2_buf_2 _18369_ (.A(_11474_),
    .X(_11475_));
 sg13g2_a21oi_1 _18370_ (.A1(net245),
    .A2(net80),
    .Y(_11476_),
    .B1(_11475_));
 sg13g2_nor2_1 _18371_ (.A(net458),
    .B(_11476_),
    .Y(_11477_));
 sg13g2_nand4_1 _18372_ (.B(_10911_),
    .C(_10969_),
    .A(_10884_),
    .Y(_11478_),
    .D(_10994_));
 sg13g2_nor2_1 _18373_ (.A(net301),
    .B(net371),
    .Y(_11479_));
 sg13g2_buf_2 _18374_ (.A(_11479_),
    .X(_11480_));
 sg13g2_nor2_2 _18375_ (.A(net374),
    .B(net370),
    .Y(_11481_));
 sg13g2_nand2_2 _18376_ (.Y(_11482_),
    .A(_11480_),
    .B(_11481_));
 sg13g2_nand3_1 _18377_ (.B(_11290_),
    .C(_11300_),
    .A(net205),
    .Y(_11483_));
 sg13g2_nor4_1 _18378_ (.A(net225),
    .B(_11478_),
    .C(_11482_),
    .D(_11483_),
    .Y(_11484_));
 sg13g2_buf_1 _18379_ (.A(_11428_),
    .X(_11485_));
 sg13g2_nor4_1 _18380_ (.A(net202),
    .B(_11071_),
    .C(net180),
    .D(net178),
    .Y(_11486_));
 sg13g2_nor2_1 _18381_ (.A(_09138_),
    .B(net651),
    .Y(_11487_));
 sg13g2_a21oi_1 _18382_ (.A1(_11484_),
    .A2(_11486_),
    .Y(_11488_),
    .B1(_11487_));
 sg13g2_nand2_1 _18383_ (.Y(_11489_),
    .A(_11477_),
    .B(_11488_));
 sg13g2_buf_2 _18384_ (.A(\cpu.ex.r_mult[0] ),
    .X(_11490_));
 sg13g2_a21o_1 _18385_ (.A2(_11487_),
    .A1(_11490_),
    .B1(_09158_),
    .X(_11491_));
 sg13g2_a22oi_1 _18386_ (.Y(_11492_),
    .B1(_11477_),
    .B2(_11491_),
    .A2(_10028_),
    .A1(_11490_));
 sg13g2_o21ai_1 _18387_ (.B1(_11492_),
    .Y(_11493_),
    .A1(_11462_),
    .A2(_11489_));
 sg13g2_a21oi_2 _18388_ (.B1(_11493_),
    .Y(_11494_),
    .A2(_11239_),
    .A1(_10031_));
 sg13g2_inv_1 _18389_ (.Y(\cpu.ex.c_mult[0] ),
    .A(_11494_));
 sg13g2_buf_1 _18390_ (.A(\cpu.dec.load ),
    .X(_11495_));
 sg13g2_inv_2 _18391_ (.Y(_11496_),
    .A(net387));
 sg13g2_nand2_1 _18392_ (.Y(_11497_),
    .A(_09164_),
    .B(_11496_));
 sg13g2_or2_1 _18393_ (.X(_11498_),
    .B(net997),
    .A(_09138_));
 sg13g2_o21ai_1 _18394_ (.B1(_11498_),
    .Y(_11499_),
    .A1(_09121_),
    .A2(_09151_));
 sg13g2_buf_2 _18395_ (.A(_11499_),
    .X(_11500_));
 sg13g2_nor2_1 _18396_ (.A(_09121_),
    .B(_09144_),
    .Y(_11501_));
 sg13g2_nor2_1 _18397_ (.A(\cpu.ex.c_div_running ),
    .B(\cpu.ex.c_mult_running ),
    .Y(_11502_));
 sg13g2_buf_1 _18398_ (.A(_00236_),
    .X(_11503_));
 sg13g2_nand2_1 _18399_ (.Y(_11504_),
    .A(_10120_),
    .B(\cpu.cond[2] ));
 sg13g2_inv_2 _18400_ (.Y(_11505_),
    .A(net1038));
 sg13g2_a21o_1 _18401_ (.A2(_11504_),
    .A1(_11503_),
    .B1(_11505_),
    .X(_11506_));
 sg13g2_buf_1 _18402_ (.A(_11506_),
    .X(_11507_));
 sg13g2_buf_1 _18403_ (.A(\cpu.dec.jmp ),
    .X(_11508_));
 sg13g2_or2_1 _18404_ (.X(_11509_),
    .B(_11508_),
    .A(_10120_));
 sg13g2_a22oi_1 _18405_ (.Y(_11510_),
    .B1(net649),
    .B2(_11509_),
    .A2(\cpu.dec.r_swapsp ),
    .A1(_10181_));
 sg13g2_nand4_1 _18406_ (.B(_11501_),
    .C(_11502_),
    .A(net1119),
    .Y(_11511_),
    .D(_11510_));
 sg13g2_nand3_1 _18407_ (.B(_11500_),
    .C(_11511_),
    .A(_11497_),
    .Y(_11512_));
 sg13g2_buf_1 _18408_ (.A(_11512_),
    .X(_11513_));
 sg13g2_and2_1 _18409_ (.A(net1039),
    .B(_11513_),
    .X(_11514_));
 sg13g2_buf_2 _18410_ (.A(_11514_),
    .X(_11515_));
 sg13g2_nand2_1 _18411_ (.Y(_11516_),
    .A(_00277_),
    .B(_11515_));
 sg13g2_nand2_1 _18412_ (.Y(_11517_),
    .A(_08962_),
    .B(_11513_));
 sg13g2_buf_1 _18413_ (.A(_11517_),
    .X(_11518_));
 sg13g2_nand3_1 _18414_ (.B(_09581_),
    .C(_09593_),
    .A(_09570_),
    .Y(_11519_));
 sg13g2_nor4_1 _18415_ (.A(_09234_),
    .B(_09373_),
    .C(_09511_),
    .D(_11519_),
    .Y(_11520_));
 sg13g2_nor4_1 _18416_ (.A(_09278_),
    .B(_09312_),
    .C(_09400_),
    .D(_09430_),
    .Y(_11521_));
 sg13g2_nor4_1 _18417_ (.A(_09347_),
    .B(_09456_),
    .C(_09624_),
    .D(_09646_),
    .Y(_11522_));
 sg13g2_nand4_1 _18418_ (.B(_11520_),
    .C(_11521_),
    .A(_09175_),
    .Y(_11523_),
    .D(_11522_));
 sg13g2_buf_1 _18419_ (.A(_11523_),
    .X(_11524_));
 sg13g2_and2_1 _18420_ (.A(_09182_),
    .B(_09180_),
    .X(_11525_));
 sg13g2_o21ai_1 _18421_ (.B1(_09168_),
    .Y(_11526_),
    .A1(_11524_),
    .A2(_11525_));
 sg13g2_and2_1 _18422_ (.A(_09022_),
    .B(_11526_),
    .X(_11527_));
 sg13g2_buf_1 _18423_ (.A(_11527_),
    .X(_11528_));
 sg13g2_nand2_1 _18424_ (.Y(_11529_),
    .A(net144),
    .B(_11528_));
 sg13g2_a21o_1 _18425_ (.A2(_11529_),
    .A1(_11516_),
    .B1(_09018_),
    .X(_11530_));
 sg13g2_o21ai_1 _18426_ (.B1(_11530_),
    .Y(_00054_),
    .A1(_11495_),
    .A2(_11516_));
 sg13g2_inv_1 _18427_ (.Y(_11531_),
    .A(_11184_));
 sg13g2_nor3_1 _18428_ (.A(net199),
    .B(_11180_),
    .C(_11531_),
    .Y(_11532_));
 sg13g2_inv_1 _18429_ (.Y(_11533_),
    .A(net1123));
 sg13g2_nor3_2 _18430_ (.A(_11533_),
    .B(_10028_),
    .C(_10030_),
    .Y(_11534_));
 sg13g2_and2_1 _18431_ (.A(net118),
    .B(_11534_),
    .X(_11535_));
 sg13g2_o21ai_1 _18432_ (.B1(_11445_),
    .Y(_11536_),
    .A1(_11180_),
    .A2(_11531_));
 sg13g2_a22oi_1 _18433_ (.Y(_11537_),
    .B1(_11535_),
    .B2(_11536_),
    .A2(_11534_),
    .A1(_11532_));
 sg13g2_buf_8 _18434_ (.A(_11537_),
    .X(_11538_));
 sg13g2_buf_1 _18435_ (.A(_11538_),
    .X(_11539_));
 sg13g2_nor2b_1 _18436_ (.A(_10028_),
    .B_N(_10030_),
    .Y(_11540_));
 sg13g2_buf_1 _18437_ (.A(_11540_),
    .X(_11541_));
 sg13g2_buf_1 _18438_ (.A(net370),
    .X(_11542_));
 sg13g2_buf_1 _18439_ (.A(net297),
    .X(_11543_));
 sg13g2_nand2_1 _18440_ (.Y(_11544_),
    .A(net80),
    .B(net244));
 sg13g2_buf_1 _18441_ (.A(_09157_),
    .X(_11545_));
 sg13g2_buf_1 _18442_ (.A(net587),
    .X(_11546_));
 sg13g2_nand3_1 _18443_ (.B(net521),
    .C(_11544_),
    .A(_11490_),
    .Y(_11547_));
 sg13g2_o21ai_1 _18444_ (.B1(_11547_),
    .Y(_11548_),
    .A1(_11490_),
    .A2(_11544_));
 sg13g2_and2_1 _18445_ (.A(_11475_),
    .B(_11488_),
    .X(_11549_));
 sg13g2_buf_1 _18446_ (.A(_11549_),
    .X(_11550_));
 sg13g2_nand2_1 _18447_ (.Y(_11551_),
    .A(_11490_),
    .B(_11550_));
 sg13g2_o21ai_1 _18448_ (.B1(_11551_),
    .Y(_11552_),
    .A1(net521),
    .A2(_11544_));
 sg13g2_a21o_1 _18449_ (.A2(_11548_),
    .A1(net997),
    .B1(_11552_),
    .X(_11553_));
 sg13g2_nor2_1 _18450_ (.A(_09138_),
    .B(net997),
    .Y(_11554_));
 sg13g2_nand2_1 _18451_ (.Y(_11555_),
    .A(_11325_),
    .B(_11554_));
 sg13g2_buf_2 _18452_ (.A(_11555_),
    .X(_11556_));
 sg13g2_nor2_1 _18453_ (.A(_11464_),
    .B(_11556_),
    .Y(_11557_));
 sg13g2_or2_1 _18454_ (.X(_11558_),
    .B(_11557_),
    .A(_10028_));
 sg13g2_buf_1 _18455_ (.A(_11558_),
    .X(_11559_));
 sg13g2_buf_1 _18456_ (.A(_11559_),
    .X(_11560_));
 sg13g2_buf_2 _18457_ (.A(\cpu.ex.r_mult[1] ),
    .X(_11561_));
 sg13g2_a22oi_1 _18458_ (.Y(_11562_),
    .B1(net243),
    .B2(_11561_),
    .A2(_11553_),
    .A1(net522));
 sg13g2_nand2_1 _18459_ (.Y(\cpu.ex.c_mult[1] ),
    .A(net27),
    .B(_11562_));
 sg13g2_buf_1 _18460_ (.A(_11550_),
    .X(_11563_));
 sg13g2_buf_1 _18461_ (.A(net80),
    .X(_11564_));
 sg13g2_buf_1 _18462_ (.A(net371),
    .X(_11565_));
 sg13g2_nand2_1 _18463_ (.Y(_11566_),
    .A(_11490_),
    .B(net297));
 sg13g2_xnor2_1 _18464_ (.Y(_11567_),
    .A(net296),
    .B(_11566_));
 sg13g2_buf_1 _18465_ (.A(net650),
    .X(_11568_));
 sg13g2_a21oi_1 _18466_ (.A1(_11564_),
    .A2(_11567_),
    .Y(_11569_),
    .B1(_11568_));
 sg13g2_nor3_1 _18467_ (.A(net650),
    .B(net296),
    .C(_11566_),
    .Y(_11570_));
 sg13g2_a21oi_1 _18468_ (.A1(net296),
    .A2(_11566_),
    .Y(_11571_),
    .B1(_11570_));
 sg13g2_nand2_1 _18469_ (.Y(_11572_),
    .A(net586),
    .B(net296));
 sg13g2_o21ai_1 _18470_ (.B1(_11572_),
    .Y(_11573_),
    .A1(_11561_),
    .A2(_11571_));
 sg13g2_a22oi_1 _18471_ (.Y(_11574_),
    .B1(_11573_),
    .B2(_11564_),
    .A2(_11569_),
    .A1(_11561_));
 sg13g2_inv_1 _18472_ (.Y(_11575_),
    .A(_11574_));
 sg13g2_a22oi_1 _18473_ (.Y(_11576_),
    .B1(_11575_),
    .B2(_09158_),
    .A2(_11563_),
    .A1(_11561_));
 sg13g2_buf_1 _18474_ (.A(\cpu.ex.r_mult[2] ),
    .X(_11577_));
 sg13g2_nand2_1 _18475_ (.Y(_11578_),
    .A(_11577_),
    .B(net243));
 sg13g2_o21ai_1 _18476_ (.B1(_11578_),
    .Y(_11579_),
    .A1(net458),
    .A2(_11576_));
 sg13g2_nand2b_1 _18477_ (.Y(\cpu.ex.c_mult[2] ),
    .B(net27),
    .A_N(_11579_));
 sg13g2_a21o_1 _18478_ (.A2(_11391_),
    .A1(_11468_),
    .B1(_11368_),
    .X(_11580_));
 sg13g2_buf_1 _18479_ (.A(_11580_),
    .X(_11581_));
 sg13g2_buf_8 _18480_ (.A(_11581_),
    .X(_11582_));
 sg13g2_buf_1 _18481_ (.A(net78),
    .X(_11583_));
 sg13g2_buf_1 _18482_ (.A(net301),
    .X(_11584_));
 sg13g2_inv_1 _18483_ (.Y(_11585_),
    .A(_11561_));
 sg13g2_buf_1 _18484_ (.A(net299),
    .X(_11586_));
 sg13g2_nor2_1 _18485_ (.A(_10445_),
    .B(_10455_),
    .Y(_11587_));
 sg13g2_nand2_1 _18486_ (.Y(_11588_),
    .A(_11561_),
    .B(_10133_));
 sg13g2_nor2_1 _18487_ (.A(_10344_),
    .B(_11588_),
    .Y(_11589_));
 sg13g2_nand2_1 _18488_ (.Y(_11590_),
    .A(_09035_),
    .B(net526));
 sg13g2_nand2_1 _18489_ (.Y(_11591_),
    .A(_11561_),
    .B(_10460_));
 sg13g2_o21ai_1 _18490_ (.B1(_11591_),
    .Y(_11592_),
    .A1(_11590_),
    .A2(_11588_));
 sg13g2_a221oi_1 _18491_ (.B2(_11589_),
    .C1(_11592_),
    .B1(_11587_),
    .A1(_11490_),
    .Y(_11593_),
    .A2(_10334_));
 sg13g2_a21oi_2 _18492_ (.B1(_11593_),
    .Y(_11594_),
    .A2(net241),
    .A1(_11585_));
 sg13g2_nand3_1 _18493_ (.B(net300),
    .C(_11594_),
    .A(net587),
    .Y(_11595_));
 sg13g2_o21ai_1 _18494_ (.B1(_11595_),
    .Y(_11596_),
    .A1(net300),
    .A2(_11594_));
 sg13g2_inv_1 _18495_ (.Y(_11597_),
    .A(_11577_));
 sg13g2_a22oi_1 _18496_ (.Y(_11598_),
    .B1(_11596_),
    .B2(_11597_),
    .A2(net242),
    .A1(_11568_));
 sg13g2_xnor2_1 _18497_ (.Y(_11599_),
    .A(net300),
    .B(_11594_));
 sg13g2_nand2_1 _18498_ (.Y(_11600_),
    .A(net73),
    .B(_11599_));
 sg13g2_nand3_1 _18499_ (.B(net521),
    .C(_11600_),
    .A(_11577_),
    .Y(_11601_));
 sg13g2_o21ai_1 _18500_ (.B1(_11601_),
    .Y(_11602_),
    .A1(net72),
    .A2(_11598_));
 sg13g2_a22oi_1 _18501_ (.Y(_11603_),
    .B1(_11602_),
    .B2(_09158_),
    .A2(_11563_),
    .A1(_11577_));
 sg13g2_buf_2 _18502_ (.A(\cpu.ex.r_mult[3] ),
    .X(_11604_));
 sg13g2_nand2_1 _18503_ (.Y(_11605_),
    .A(_11604_),
    .B(net243));
 sg13g2_o21ai_1 _18504_ (.B1(_11605_),
    .Y(_11606_),
    .A1(net458),
    .A2(_11603_));
 sg13g2_nand2b_1 _18505_ (.Y(\cpu.ex.c_mult[3] ),
    .B(net27),
    .A_N(_11606_));
 sg13g2_buf_2 _18506_ (.A(\cpu.ex.r_mult[4] ),
    .X(_11607_));
 sg13g2_a221oi_1 _18507_ (.B2(_11585_),
    .C1(_11593_),
    .B1(_11404_),
    .A1(_11597_),
    .Y(_11608_),
    .A2(net372));
 sg13g2_buf_1 _18508_ (.A(_11608_),
    .X(_11609_));
 sg13g2_nor2_1 _18509_ (.A(_11597_),
    .B(net372),
    .Y(_11610_));
 sg13g2_nor2_1 _18510_ (.A(_11609_),
    .B(_11610_),
    .Y(_11611_));
 sg13g2_nor3_1 _18511_ (.A(_11473_),
    .B(net247),
    .C(_11611_),
    .Y(_11612_));
 sg13g2_a21oi_1 _18512_ (.A1(net247),
    .A2(_11611_),
    .Y(_11613_),
    .B1(_11612_));
 sg13g2_nand2_1 _18513_ (.Y(_11614_),
    .A(net586),
    .B(_11293_));
 sg13g2_o21ai_1 _18514_ (.B1(_11614_),
    .Y(_11615_),
    .A1(_11604_),
    .A2(_11613_));
 sg13g2_xnor2_1 _18515_ (.Y(_11616_),
    .A(_11293_),
    .B(_11611_));
 sg13g2_nand2_1 _18516_ (.Y(_11617_),
    .A(_11604_),
    .B(net587));
 sg13g2_a21oi_1 _18517_ (.A1(net73),
    .A2(_11616_),
    .Y(_11618_),
    .B1(_11617_));
 sg13g2_a21oi_1 _18518_ (.A1(net73),
    .A2(_11615_),
    .Y(_11619_),
    .B1(_11618_));
 sg13g2_nor2_1 _18519_ (.A(_11330_),
    .B(_11498_),
    .Y(_11620_));
 sg13g2_buf_2 _18520_ (.A(_11620_),
    .X(_11621_));
 sg13g2_a22oi_1 _18521_ (.Y(_11622_),
    .B1(_11621_),
    .B2(_11607_),
    .A2(_11550_),
    .A1(_11604_));
 sg13g2_o21ai_1 _18522_ (.B1(_11622_),
    .Y(_11623_),
    .A1(_11475_),
    .A2(_11619_));
 sg13g2_a22oi_1 _18523_ (.Y(_11624_),
    .B1(net522),
    .B2(_11623_),
    .A2(_10029_),
    .A1(_11607_));
 sg13g2_nand2_1 _18524_ (.Y(\cpu.ex.c_mult[4] ),
    .A(_11538_),
    .B(_11624_));
 sg13g2_nand2b_1 _18525_ (.Y(_11625_),
    .B(net302),
    .A_N(_11604_));
 sg13g2_and2_1 _18526_ (.A(_11604_),
    .B(_10576_),
    .X(_11626_));
 sg13g2_or3_1 _18527_ (.A(_11609_),
    .B(_11610_),
    .C(_11626_),
    .X(_11627_));
 sg13g2_buf_1 _18528_ (.A(_11627_),
    .X(_11628_));
 sg13g2_nand3_1 _18529_ (.B(_11625_),
    .C(_11628_),
    .A(net587),
    .Y(_11629_));
 sg13g2_xnor2_1 _18530_ (.Y(_11630_),
    .A(net246),
    .B(_11629_));
 sg13g2_nor2_1 _18531_ (.A(net72),
    .B(_11630_),
    .Y(_11631_));
 sg13g2_o21ai_1 _18532_ (.B1(net521),
    .Y(_11632_),
    .A1(_09156_),
    .A2(_11607_));
 sg13g2_nand2_2 _18533_ (.Y(_11633_),
    .A(net997),
    .B(net587));
 sg13g2_nand2_1 _18534_ (.Y(_11634_),
    .A(_11475_),
    .B(_11488_));
 sg13g2_o21ai_1 _18535_ (.B1(_11634_),
    .Y(_11635_),
    .A1(_11631_),
    .A2(_11633_));
 sg13g2_a22oi_1 _18536_ (.Y(_11636_),
    .B1(_11635_),
    .B2(_11607_),
    .A2(_11632_),
    .A1(_11631_));
 sg13g2_buf_2 _18537_ (.A(\cpu.ex.r_mult[5] ),
    .X(_11637_));
 sg13g2_nand2_1 _18538_ (.Y(_11638_),
    .A(_11637_),
    .B(net243));
 sg13g2_o21ai_1 _18539_ (.B1(_11638_),
    .Y(_11639_),
    .A1(_11465_),
    .A2(_11636_));
 sg13g2_nand2b_1 _18540_ (.Y(\cpu.ex.c_mult[5] ),
    .B(_11538_),
    .A_N(_11639_));
 sg13g2_nor2_1 _18541_ (.A(_11475_),
    .B(_11464_),
    .Y(_11640_));
 sg13g2_buf_1 _18542_ (.A(_11640_),
    .X(_11641_));
 sg13g2_nand2_1 _18543_ (.Y(_11642_),
    .A(_11637_),
    .B(net521));
 sg13g2_nand2_1 _18544_ (.Y(_11643_),
    .A(_11607_),
    .B(_10541_));
 sg13g2_nor2_1 _18545_ (.A(_11607_),
    .B(_10540_),
    .Y(_11644_));
 sg13g2_inv_1 _18546_ (.Y(_11645_),
    .A(_11644_));
 sg13g2_nand3_1 _18547_ (.B(_11628_),
    .C(_11645_),
    .A(_11625_),
    .Y(_11646_));
 sg13g2_buf_1 _18548_ (.A(_11646_),
    .X(_11647_));
 sg13g2_or2_1 _18549_ (.X(_11648_),
    .B(_10809_),
    .A(net730));
 sg13g2_buf_1 _18550_ (.A(_11648_),
    .X(_11649_));
 sg13g2_a21oi_1 _18551_ (.A1(_11643_),
    .A2(_11647_),
    .Y(_11650_),
    .B1(_11649_));
 sg13g2_nor2_1 _18552_ (.A(net586),
    .B(_11647_),
    .Y(_11651_));
 sg13g2_buf_1 _18553_ (.A(_11284_),
    .X(_11652_));
 sg13g2_o21ai_1 _18554_ (.B1(net198),
    .Y(_11653_),
    .A1(net586),
    .A2(_11643_));
 sg13g2_nor2_1 _18555_ (.A(_11651_),
    .B(_11653_),
    .Y(_11654_));
 sg13g2_nor3_1 _18556_ (.A(net72),
    .B(_11650_),
    .C(_11654_),
    .Y(_11655_));
 sg13g2_xnor2_1 _18557_ (.Y(_11656_),
    .A(_11642_),
    .B(_11655_));
 sg13g2_nand2_1 _18558_ (.Y(_11657_),
    .A(net422),
    .B(_11656_));
 sg13g2_buf_1 _18559_ (.A(\cpu.ex.r_mult[6] ),
    .X(_11658_));
 sg13g2_nor2_1 _18560_ (.A(_11464_),
    .B(_11634_),
    .Y(_11659_));
 sg13g2_buf_2 _18561_ (.A(_11659_),
    .X(_11660_));
 sg13g2_buf_1 _18562_ (.A(_11660_),
    .X(_11661_));
 sg13g2_a22oi_1 _18563_ (.Y(_11662_),
    .B1(net71),
    .B2(_11637_),
    .A2(net243),
    .A1(_11658_));
 sg13g2_nand2_1 _18564_ (.Y(_11663_),
    .A(_11657_),
    .B(_11662_));
 sg13g2_nand2b_1 _18565_ (.Y(\cpu.ex.c_mult[6] ),
    .B(_11538_),
    .A_N(_11663_));
 sg13g2_nand2_1 _18566_ (.Y(_11664_),
    .A(_11658_),
    .B(_09149_));
 sg13g2_buf_1 _18567_ (.A(_10812_),
    .X(_11665_));
 sg13g2_inv_1 _18568_ (.Y(_11666_),
    .A(_11637_));
 sg13g2_inv_1 _18569_ (.Y(_11667_),
    .A(_11607_));
 sg13g2_nor3_1 _18570_ (.A(_11604_),
    .B(_10571_),
    .C(_10574_),
    .Y(_11668_));
 sg13g2_a221oi_1 _18571_ (.B2(_11667_),
    .C1(_11668_),
    .B1(net246),
    .A1(_11666_),
    .Y(_11669_),
    .A2(net224));
 sg13g2_o21ai_1 _18572_ (.B1(_11669_),
    .Y(_11670_),
    .A1(_11609_),
    .A2(_11610_));
 sg13g2_a21oi_1 _18573_ (.A1(_11666_),
    .A2(net224),
    .Y(_11671_),
    .B1(_11295_));
 sg13g2_o21ai_1 _18574_ (.B1(_11604_),
    .Y(_11672_),
    .A1(_10571_),
    .A2(_10574_));
 sg13g2_a221oi_1 _18575_ (.B2(_11672_),
    .C1(_11667_),
    .B1(_11295_),
    .A1(_11666_),
    .Y(_11673_),
    .A2(_10809_));
 sg13g2_a221oi_1 _18576_ (.B2(_11671_),
    .C1(_11673_),
    .B1(_11626_),
    .A1(_11637_),
    .Y(_11674_),
    .A2(net201));
 sg13g2_buf_1 _18577_ (.A(_11674_),
    .X(_11675_));
 sg13g2_a21oi_1 _18578_ (.A1(_11670_),
    .A2(_11675_),
    .Y(_11676_),
    .B1(net650));
 sg13g2_xnor2_1 _18579_ (.Y(_11677_),
    .A(net223),
    .B(_11676_));
 sg13g2_nor2_1 _18580_ (.A(net72),
    .B(_11677_),
    .Y(_11678_));
 sg13g2_xnor2_1 _18581_ (.Y(_11679_),
    .A(_11664_),
    .B(_11678_));
 sg13g2_buf_1 _18582_ (.A(\cpu.ex.r_mult[7] ),
    .X(_11680_));
 sg13g2_and2_1 _18583_ (.A(net1094),
    .B(_11559_),
    .X(_11681_));
 sg13g2_a221oi_1 _18584_ (.B2(net422),
    .C1(_11681_),
    .B1(_11679_),
    .A1(_11658_),
    .Y(_11682_),
    .A2(_11660_));
 sg13g2_nand2_1 _18585_ (.Y(\cpu.ex.c_mult[7] ),
    .A(net27),
    .B(_11682_));
 sg13g2_nand2_1 _18586_ (.Y(_11683_),
    .A(net1094),
    .B(net683));
 sg13g2_and2_1 _18587_ (.A(_10809_),
    .B(_11643_),
    .X(_11684_));
 sg13g2_nand2_1 _18588_ (.Y(_11685_),
    .A(_11647_),
    .B(_11684_));
 sg13g2_o21ai_1 _18589_ (.B1(_11637_),
    .Y(_11686_),
    .A1(_11658_),
    .A2(net249));
 sg13g2_nor2_1 _18590_ (.A(_11473_),
    .B(_11686_),
    .Y(_11687_));
 sg13g2_nor2_1 _18591_ (.A(_11644_),
    .B(_11649_),
    .Y(_11688_));
 sg13g2_nand3_1 _18592_ (.B(_11628_),
    .C(_11688_),
    .A(_11625_),
    .Y(_11689_));
 sg13g2_nor2_1 _18593_ (.A(_11643_),
    .B(_11649_),
    .Y(_11690_));
 sg13g2_nor2_1 _18594_ (.A(net249),
    .B(_11690_),
    .Y(_11691_));
 sg13g2_a21oi_1 _18595_ (.A1(_11689_),
    .A2(_11691_),
    .Y(_11692_),
    .B1(_11664_));
 sg13g2_a221oi_1 _18596_ (.B2(_11687_),
    .C1(_11692_),
    .B1(_11685_),
    .A1(net223),
    .Y(_11693_),
    .A2(_11650_));
 sg13g2_xnor2_1 _18597_ (.Y(_11694_),
    .A(net226),
    .B(_11693_));
 sg13g2_nand2_1 _18598_ (.Y(_11695_),
    .A(net80),
    .B(_11694_));
 sg13g2_mux2_1 _18599_ (.A0(net1094),
    .A1(_11683_),
    .S(_11695_),
    .X(_11696_));
 sg13g2_nand3_1 _18600_ (.B(net73),
    .C(_11694_),
    .A(net586),
    .Y(_11697_));
 sg13g2_buf_1 _18601_ (.A(\cpu.ex.r_mult[8] ),
    .X(_11698_));
 sg13g2_a22oi_1 _18602_ (.Y(_11699_),
    .B1(_11621_),
    .B2(net1093),
    .A2(_11550_),
    .A1(net1094));
 sg13g2_and2_1 _18603_ (.A(_11697_),
    .B(_11699_),
    .X(_11700_));
 sg13g2_o21ai_1 _18604_ (.B1(_11700_),
    .Y(_11701_),
    .A1(_09156_),
    .A2(_11696_));
 sg13g2_and2_1 _18605_ (.A(net1093),
    .B(_10028_),
    .X(_11702_));
 sg13g2_a221oi_1 _18606_ (.B2(net522),
    .C1(_11702_),
    .B1(_11701_),
    .A1(_11239_),
    .Y(_11703_),
    .A2(_11534_));
 sg13g2_inv_1 _18607_ (.Y(\cpu.ex.c_mult[8] ),
    .A(_11703_));
 sg13g2_nand3_1 _18608_ (.B(net73),
    .C(net225),
    .A(net586),
    .Y(_11704_));
 sg13g2_o21ai_1 _18609_ (.B1(_11658_),
    .Y(_11705_),
    .A1(net1094),
    .A2(net226));
 sg13g2_nand2b_1 _18610_ (.Y(_11706_),
    .B(net683),
    .A_N(_11705_));
 sg13g2_nand3_1 _18611_ (.B(net226),
    .C(net223),
    .A(net683),
    .Y(_11707_));
 sg13g2_a22oi_1 _18612_ (.Y(_11708_),
    .B1(_11706_),
    .B2(_11707_),
    .A2(_11675_),
    .A1(_11670_));
 sg13g2_or2_1 _18613_ (.X(_11709_),
    .B(_11683_),
    .A(net228));
 sg13g2_a21oi_1 _18614_ (.A1(_11670_),
    .A2(_11675_),
    .Y(_11710_),
    .B1(_11709_));
 sg13g2_nor3_1 _18615_ (.A(net730),
    .B(_10800_),
    .C(_11705_),
    .Y(_11711_));
 sg13g2_nor2_1 _18616_ (.A(net205),
    .B(_11683_),
    .Y(_11712_));
 sg13g2_nor4_2 _18617_ (.A(_11708_),
    .B(_11710_),
    .C(_11711_),
    .Y(_11713_),
    .D(_11712_));
 sg13g2_xnor2_1 _18618_ (.Y(_11714_),
    .A(net225),
    .B(_11713_));
 sg13g2_nand2_1 _18619_ (.Y(_11715_),
    .A(net80),
    .B(_11714_));
 sg13g2_nand4_1 _18620_ (.B(_11698_),
    .C(_11546_),
    .A(_11472_),
    .Y(_11716_),
    .D(_11715_));
 sg13g2_inv_1 _18621_ (.Y(_11717_),
    .A(net1093));
 sg13g2_nand4_1 _18622_ (.B(_11717_),
    .C(net73),
    .A(_11472_),
    .Y(_11718_),
    .D(_11714_));
 sg13g2_nand3_1 _18623_ (.B(_11716_),
    .C(_11718_),
    .A(_11704_),
    .Y(_11719_));
 sg13g2_buf_1 _18624_ (.A(\cpu.ex.r_mult[9] ),
    .X(_11720_));
 sg13g2_and2_1 _18625_ (.A(_11720_),
    .B(_11559_),
    .X(_11721_));
 sg13g2_a221oi_1 _18626_ (.B2(net522),
    .C1(_11721_),
    .B1(_11719_),
    .A1(net1093),
    .Y(_11722_),
    .A2(_11660_));
 sg13g2_nand2_1 _18627_ (.Y(\cpu.ex.c_mult[9] ),
    .A(_11539_),
    .B(_11722_));
 sg13g2_nand2_1 _18628_ (.Y(_11723_),
    .A(_11720_),
    .B(net683));
 sg13g2_a221oi_1 _18629_ (.B2(_11684_),
    .C1(_11686_),
    .B1(_11647_),
    .A1(\cpu.dec.mult ),
    .Y(_11724_),
    .A2(_11501_));
 sg13g2_nand2_1 _18630_ (.Y(_11725_),
    .A(net1093),
    .B(net248));
 sg13g2_nand2b_1 _18631_ (.Y(_11726_),
    .B(_11717_),
    .A_N(net248));
 sg13g2_and4_1 _18632_ (.A(net1094),
    .B(_10674_),
    .C(_11725_),
    .D(_11726_),
    .X(_11727_));
 sg13g2_nor4_1 _18633_ (.A(net1094),
    .B(_11717_),
    .C(net248),
    .D(_10674_),
    .Y(_11728_));
 sg13g2_o21ai_1 _18634_ (.B1(_09149_),
    .Y(_11729_),
    .A1(_11727_),
    .A2(_11728_));
 sg13g2_o21ai_1 _18635_ (.B1(_09149_),
    .Y(_11730_),
    .A1(_11680_),
    .A2(net1093));
 sg13g2_nand3_1 _18636_ (.B(_10646_),
    .C(_11730_),
    .A(net248),
    .Y(_11731_));
 sg13g2_nand2_1 _18637_ (.Y(_11732_),
    .A(_11729_),
    .B(_11731_));
 sg13g2_o21ai_1 _18638_ (.B1(_11732_),
    .Y(_11733_),
    .A1(_11724_),
    .A2(_11692_));
 sg13g2_buf_1 _18639_ (.A(_11733_),
    .X(_11734_));
 sg13g2_nand2_1 _18640_ (.Y(_11735_),
    .A(net1094),
    .B(_10646_));
 sg13g2_nor2_1 _18641_ (.A(net1093),
    .B(net248),
    .Y(_11736_));
 sg13g2_o21ai_1 _18642_ (.B1(_11725_),
    .Y(_11737_),
    .A1(_11735_),
    .A2(_11736_));
 sg13g2_a21oi_1 _18643_ (.A1(_11729_),
    .A2(_11731_),
    .Y(_11738_),
    .B1(_10800_));
 sg13g2_a22oi_1 _18644_ (.Y(_11739_),
    .B1(_11738_),
    .B2(_11650_),
    .A2(_11737_),
    .A1(net683));
 sg13g2_buf_1 _18645_ (.A(_11739_),
    .X(_11740_));
 sg13g2_a21o_1 _18646_ (.A2(_11740_),
    .A1(_11734_),
    .B1(net182),
    .X(_11741_));
 sg13g2_nand3_1 _18647_ (.B(_11734_),
    .C(_11740_),
    .A(net182),
    .Y(_11742_));
 sg13g2_a21oi_1 _18648_ (.A1(_11741_),
    .A2(_11742_),
    .Y(_11743_),
    .B1(net72));
 sg13g2_xnor2_1 _18649_ (.Y(_11744_),
    .A(_11723_),
    .B(_11743_));
 sg13g2_buf_1 _18650_ (.A(\cpu.ex.r_mult[10] ),
    .X(_11745_));
 sg13g2_and2_1 _18651_ (.A(_11745_),
    .B(net243),
    .X(_11746_));
 sg13g2_a221oi_1 _18652_ (.B2(net422),
    .C1(_11746_),
    .B1(_11744_),
    .A1(_11720_),
    .Y(_11747_),
    .A2(_11661_));
 sg13g2_nand2_1 _18653_ (.Y(\cpu.ex.c_mult[10] ),
    .A(net27),
    .B(_11747_));
 sg13g2_inv_1 _18654_ (.Y(_11748_),
    .A(_11720_));
 sg13g2_a21oi_1 _18655_ (.A1(_11748_),
    .A2(net145),
    .Y(_11749_),
    .B1(_11725_));
 sg13g2_a21oi_2 _18656_ (.B1(_11748_),
    .Y(_11750_),
    .A2(_10994_),
    .A1(_10969_));
 sg13g2_o21ai_1 _18657_ (.B1(net587),
    .Y(_11751_),
    .A1(_11749_),
    .A2(_11750_));
 sg13g2_nand2_1 _18658_ (.Y(_11752_),
    .A(_11713_),
    .B(_11751_));
 sg13g2_o21ai_1 _18659_ (.B1(_11545_),
    .Y(_11753_),
    .A1(net1093),
    .A2(_11750_));
 sg13g2_a221oi_1 _18660_ (.B2(_10878_),
    .C1(net78),
    .B1(_11753_),
    .A1(net145),
    .Y(_11754_),
    .A2(_11723_));
 sg13g2_nand2_1 _18661_ (.Y(_11755_),
    .A(_11752_),
    .B(_11754_));
 sg13g2_nand2_1 _18662_ (.Y(_11756_),
    .A(_11745_),
    .B(_09149_));
 sg13g2_nor2_1 _18663_ (.A(net78),
    .B(net181),
    .Y(_11757_));
 sg13g2_xnor2_1 _18664_ (.Y(_11758_),
    .A(_11756_),
    .B(_11757_));
 sg13g2_xnor2_1 _18665_ (.Y(_11759_),
    .A(_11755_),
    .B(_11758_));
 sg13g2_nand2_1 _18666_ (.Y(_11760_),
    .A(net422),
    .B(_11759_));
 sg13g2_buf_2 _18667_ (.A(\cpu.ex.r_mult[11] ),
    .X(_11761_));
 sg13g2_a22oi_1 _18668_ (.Y(_11762_),
    .B1(_11660_),
    .B2(_11745_),
    .A2(_11560_),
    .A1(_11761_));
 sg13g2_nand3_1 _18669_ (.B(_11760_),
    .C(_11762_),
    .A(_11538_),
    .Y(\cpu.ex.c_mult[11] ));
 sg13g2_buf_1 _18670_ (.A(\cpu.ex.r_mult[12] ),
    .X(_11763_));
 sg13g2_inv_1 _18671_ (.Y(_11764_),
    .A(_11745_));
 sg13g2_o21ai_1 _18672_ (.B1(_11764_),
    .Y(_11765_),
    .A1(_11029_),
    .A2(_11031_));
 sg13g2_o21ai_1 _18673_ (.B1(_11765_),
    .Y(_11766_),
    .A1(net183),
    .A2(_11756_));
 sg13g2_a221oi_1 _18674_ (.B2(_11748_),
    .C1(_11255_),
    .B1(_11766_),
    .A1(net730),
    .Y(_11767_),
    .A2(net183));
 sg13g2_xnor2_1 _18675_ (.Y(_11768_),
    .A(_11764_),
    .B(_11032_));
 sg13g2_o21ai_1 _18676_ (.B1(_11255_),
    .Y(_11769_),
    .A1(_11723_),
    .A2(_11768_));
 sg13g2_nand3b_1 _18677_ (.B(_11769_),
    .C(_11470_),
    .Y(_11770_),
    .A_N(_11767_));
 sg13g2_a21oi_1 _18678_ (.A1(_11734_),
    .A2(_11740_),
    .Y(_11771_),
    .B1(_11770_));
 sg13g2_nand2_1 _18679_ (.Y(_11772_),
    .A(net80),
    .B(net178));
 sg13g2_nand3_1 _18680_ (.B(_10884_),
    .C(_10911_),
    .A(_11764_),
    .Y(_11773_));
 sg13g2_a21oi_1 _18681_ (.A1(_10884_),
    .A2(_10911_),
    .Y(_11774_),
    .B1(_11764_));
 sg13g2_a21oi_1 _18682_ (.A1(_11750_),
    .A2(_11773_),
    .Y(_11775_),
    .B1(_11774_));
 sg13g2_nand2_1 _18683_ (.Y(_11776_),
    .A(_11176_),
    .B(_11775_));
 sg13g2_nand2_1 _18684_ (.Y(_11777_),
    .A(net80),
    .B(_11776_));
 sg13g2_inv_1 _18685_ (.Y(_11778_),
    .A(_11761_));
 sg13g2_a21o_1 _18686_ (.A2(_11773_),
    .A1(_11750_),
    .B1(_11774_),
    .X(_11779_));
 sg13g2_nand2_1 _18687_ (.Y(_11780_),
    .A(_11761_),
    .B(net683));
 sg13g2_nor4_1 _18688_ (.A(_11582_),
    .B(_11177_),
    .C(_11779_),
    .D(_11780_),
    .Y(_11781_));
 sg13g2_a221oi_1 _18689_ (.B2(_11778_),
    .C1(_11781_),
    .B1(_11777_),
    .A1(net586),
    .Y(_11782_),
    .A2(_11772_));
 sg13g2_nor2_1 _18690_ (.A(_11771_),
    .B(_11782_),
    .Y(_11783_));
 sg13g2_nor2_1 _18691_ (.A(_11778_),
    .B(net730),
    .Y(_11784_));
 sg13g2_xnor2_1 _18692_ (.Y(_11785_),
    .A(_11772_),
    .B(_11784_));
 sg13g2_nand2_1 _18693_ (.Y(_11786_),
    .A(_11778_),
    .B(net203));
 sg13g2_nand2_1 _18694_ (.Y(_11787_),
    .A(_11761_),
    .B(net178));
 sg13g2_nand4_1 _18695_ (.B(_11779_),
    .C(_11786_),
    .A(net80),
    .Y(_11788_),
    .D(_11787_));
 sg13g2_a21oi_1 _18696_ (.A1(net997),
    .A2(_11788_),
    .Y(_11789_),
    .B1(net586));
 sg13g2_a21o_1 _18697_ (.A2(_11785_),
    .A1(_11771_),
    .B1(_11789_),
    .X(_11790_));
 sg13g2_nand2_1 _18698_ (.Y(_11791_),
    .A(_11761_),
    .B(net79));
 sg13g2_o21ai_1 _18699_ (.B1(_11791_),
    .Y(_11792_),
    .A1(_11783_),
    .A2(_11790_));
 sg13g2_a22oi_1 _18700_ (.Y(_11793_),
    .B1(_11792_),
    .B2(_11541_),
    .A2(net243),
    .A1(net1092));
 sg13g2_nand2_1 _18701_ (.Y(\cpu.ex.c_mult[12] ),
    .A(_11539_),
    .B(_11793_));
 sg13g2_buf_2 _18702_ (.A(\cpu.ex.r_mult[13] ),
    .X(_11794_));
 sg13g2_buf_1 _18703_ (.A(_11153_),
    .X(_11795_));
 sg13g2_nand2_1 _18704_ (.Y(_11796_),
    .A(_11774_),
    .B(_11786_));
 sg13g2_a21oi_2 _18705_ (.B1(net650),
    .Y(_11797_),
    .A2(_11796_),
    .A1(_11787_));
 sg13g2_nand3_1 _18706_ (.B(_11795_),
    .C(_11797_),
    .A(_11471_),
    .Y(_11798_));
 sg13g2_nor2_1 _18707_ (.A(_11761_),
    .B(_11176_),
    .Y(_11799_));
 sg13g2_a21oi_1 _18708_ (.A1(_11176_),
    .A2(_11784_),
    .Y(_11800_),
    .B1(_11799_));
 sg13g2_nand2_1 _18709_ (.Y(_11801_),
    .A(net730),
    .B(_11428_));
 sg13g2_o21ai_1 _18710_ (.B1(_11801_),
    .Y(_11802_),
    .A1(_11745_),
    .A2(_11800_));
 sg13g2_nor3_1 _18711_ (.A(_11761_),
    .B(net183),
    .C(_11756_),
    .Y(_11803_));
 sg13g2_a22oi_1 _18712_ (.Y(_11804_),
    .B1(_11803_),
    .B2(net178),
    .A2(_11802_),
    .A1(_10913_));
 sg13g2_nand2b_1 _18713_ (.Y(_11805_),
    .B(_11470_),
    .A_N(_11804_));
 sg13g2_nor2_1 _18714_ (.A(net178),
    .B(_10913_),
    .Y(_11806_));
 sg13g2_nor2_1 _18715_ (.A(_11764_),
    .B(_11780_),
    .Y(_11807_));
 sg13g2_o21ai_1 _18716_ (.B1(_11807_),
    .Y(_11808_),
    .A1(_11582_),
    .A2(_11806_));
 sg13g2_nand2_1 _18717_ (.Y(_11809_),
    .A(_11805_),
    .B(_11808_));
 sg13g2_nand4_1 _18718_ (.B(_11752_),
    .C(_11754_),
    .A(_11795_),
    .Y(_11810_),
    .D(_11809_));
 sg13g2_nor3_1 _18719_ (.A(net78),
    .B(_11153_),
    .C(_11797_),
    .Y(_11811_));
 sg13g2_nand2_1 _18720_ (.Y(_11812_),
    .A(_11755_),
    .B(_11811_));
 sg13g2_nand3_1 _18721_ (.B(_11808_),
    .C(_11811_),
    .A(_11805_),
    .Y(_11813_));
 sg13g2_nand4_1 _18722_ (.B(_11810_),
    .C(_11812_),
    .A(_11798_),
    .Y(_11814_),
    .D(_11813_));
 sg13g2_nor2_2 _18723_ (.A(_09156_),
    .B(net650),
    .Y(_11815_));
 sg13g2_nand2_1 _18724_ (.Y(_11816_),
    .A(net522),
    .B(_11815_));
 sg13g2_buf_2 _18725_ (.A(_11816_),
    .X(_11817_));
 sg13g2_nand2_1 _18726_ (.Y(_11818_),
    .A(net522),
    .B(net79));
 sg13g2_o21ai_1 _18727_ (.B1(_11818_),
    .Y(_11819_),
    .A1(_11814_),
    .A2(_11817_));
 sg13g2_nand2_1 _18728_ (.Y(_11820_),
    .A(\cpu.ex.r_mult[12] ),
    .B(_09149_));
 sg13g2_and3_1 _18729_ (.X(_11821_),
    .A(_11641_),
    .B(_11814_),
    .C(_11820_));
 sg13g2_a221oi_1 _18730_ (.B2(_11763_),
    .C1(_11821_),
    .B1(_11819_),
    .A1(_11794_),
    .Y(_11822_),
    .A2(_11560_));
 sg13g2_buf_1 _18731_ (.A(_11822_),
    .X(_11823_));
 sg13g2_nand2_1 _18732_ (.Y(\cpu.ex.c_mult[13] ),
    .A(net27),
    .B(_11823_));
 sg13g2_and2_1 _18733_ (.A(net1092),
    .B(_11784_),
    .X(_11824_));
 sg13g2_o21ai_1 _18734_ (.B1(_11824_),
    .Y(_11825_),
    .A1(_11581_),
    .A2(_11436_));
 sg13g2_nor3_1 _18735_ (.A(_11129_),
    .B(_11151_),
    .C(_11820_),
    .Y(_11826_));
 sg13g2_a21oi_1 _18736_ (.A1(_11421_),
    .A2(_11423_),
    .Y(_11827_),
    .B1(net1092));
 sg13g2_o21ai_1 _18737_ (.B1(_11778_),
    .Y(_11828_),
    .A1(_11826_),
    .A2(_11827_));
 sg13g2_nand2_1 _18738_ (.Y(_11829_),
    .A(net730),
    .B(net180));
 sg13g2_a21oi_1 _18739_ (.A1(_11828_),
    .A2(_11829_),
    .Y(_11830_),
    .B1(_11176_));
 sg13g2_nor4_1 _18740_ (.A(net1092),
    .B(_11153_),
    .C(_11428_),
    .D(_11780_),
    .Y(_11831_));
 sg13g2_o21ai_1 _18741_ (.B1(_11470_),
    .Y(_11832_),
    .A1(_11830_),
    .A2(_11831_));
 sg13g2_a221oi_1 _18742_ (.B2(_11832_),
    .C1(_11770_),
    .B1(_11825_),
    .A1(_11734_),
    .Y(_11833_),
    .A2(_11740_));
 sg13g2_buf_1 _18743_ (.A(_11833_),
    .X(_11834_));
 sg13g2_o21ai_1 _18744_ (.B1(_11778_),
    .Y(_11835_),
    .A1(_11176_),
    .A2(_11775_));
 sg13g2_a22oi_1 _18745_ (.Y(_11836_),
    .B1(_11776_),
    .B2(_11835_),
    .A2(net180),
    .A1(net1092));
 sg13g2_o21ai_1 _18746_ (.B1(_11545_),
    .Y(_11837_),
    .A1(_11763_),
    .A2(net180));
 sg13g2_nor3_1 _18747_ (.A(net72),
    .B(_11836_),
    .C(_11837_),
    .Y(_11838_));
 sg13g2_nor2_1 _18748_ (.A(_11834_),
    .B(_11838_),
    .Y(_11839_));
 sg13g2_nand2_2 _18749_ (.Y(_11840_),
    .A(_11794_),
    .B(_09157_));
 sg13g2_nor2_1 _18750_ (.A(_11583_),
    .B(net147),
    .Y(_11841_));
 sg13g2_xnor2_1 _18751_ (.Y(_11842_),
    .A(_11840_),
    .B(_11841_));
 sg13g2_xnor2_1 _18752_ (.Y(_11843_),
    .A(_11839_),
    .B(_11842_));
 sg13g2_and2_1 _18753_ (.A(\cpu.ex.r_mult[14] ),
    .B(net243),
    .X(_11844_));
 sg13g2_a221oi_1 _18754_ (.B2(net422),
    .C1(_11844_),
    .B1(_11843_),
    .A1(_11794_),
    .Y(_11845_),
    .A2(net71));
 sg13g2_nand2_1 _18755_ (.Y(\cpu.ex.c_mult[14] ),
    .A(net27),
    .B(_11845_));
 sg13g2_buf_1 _18756_ (.A(net180),
    .X(_11846_));
 sg13g2_inv_1 _18757_ (.Y(_11847_),
    .A(_11794_));
 sg13g2_nor2_1 _18758_ (.A(_11071_),
    .B(_11840_),
    .Y(_11848_));
 sg13g2_a21oi_1 _18759_ (.A1(_11847_),
    .A2(net179),
    .Y(_11849_),
    .B1(_11848_));
 sg13g2_nand2_1 _18760_ (.Y(_11850_),
    .A(net650),
    .B(net179));
 sg13g2_o21ai_1 _18761_ (.B1(_11850_),
    .Y(_11851_),
    .A1(net1092),
    .A2(_11849_));
 sg13g2_nor3_1 _18762_ (.A(_11794_),
    .B(_11435_),
    .C(_11820_),
    .Y(_11852_));
 sg13g2_a22oi_1 _18763_ (.Y(_11853_),
    .B1(_11852_),
    .B2(net179),
    .A2(_11851_),
    .A1(net142));
 sg13g2_nor2_1 _18764_ (.A(net78),
    .B(_11853_),
    .Y(_11854_));
 sg13g2_inv_1 _18765_ (.Y(_11855_),
    .A(_11840_));
 sg13g2_o21ai_1 _18766_ (.B1(_11471_),
    .Y(_11856_),
    .A1(_11451_),
    .A2(net142));
 sg13g2_and3_1 _18767_ (.X(_11857_),
    .A(net1092),
    .B(_11855_),
    .C(_11856_));
 sg13g2_o21ai_1 _18768_ (.B1(_11809_),
    .Y(_11858_),
    .A1(_11854_),
    .A2(_11857_));
 sg13g2_or2_1 _18769_ (.X(_11859_),
    .B(_11858_),
    .A(_11755_));
 sg13g2_buf_2 _18770_ (.A(_00149_),
    .X(_11860_));
 sg13g2_nor2_1 _18771_ (.A(_11860_),
    .B(_11323_),
    .Y(_11861_));
 sg13g2_buf_1 _18772_ (.A(_11861_),
    .X(_11862_));
 sg13g2_xnor2_1 _18773_ (.Y(_11863_),
    .A(net199),
    .B(_11862_));
 sg13g2_nand2_1 _18774_ (.Y(_11864_),
    .A(_11583_),
    .B(_11862_));
 sg13g2_o21ai_1 _18775_ (.B1(_11864_),
    .Y(_11865_),
    .A1(_11859_),
    .A2(_11863_));
 sg13g2_nand2_1 _18776_ (.Y(_11866_),
    .A(net142),
    .B(_11797_));
 sg13g2_a21oi_1 _18777_ (.A1(net147),
    .A2(_11866_),
    .Y(_11867_),
    .B1(_11840_));
 sg13g2_o21ai_1 _18778_ (.B1(net1092),
    .Y(_11868_),
    .A1(_11794_),
    .A2(_11451_));
 sg13g2_nor2_1 _18779_ (.A(net650),
    .B(_11868_),
    .Y(_11869_));
 sg13g2_o21ai_1 _18780_ (.B1(_11869_),
    .Y(_11870_),
    .A1(net142),
    .A2(_11797_));
 sg13g2_o21ai_1 _18781_ (.B1(_11870_),
    .Y(_11871_),
    .A1(net147),
    .A2(_11866_));
 sg13g2_nor2_1 _18782_ (.A(_11867_),
    .B(_11871_),
    .Y(_11872_));
 sg13g2_nor2_1 _18783_ (.A(net78),
    .B(_11862_),
    .Y(_11873_));
 sg13g2_mux2_1 _18784_ (.A0(_11862_),
    .A1(_11873_),
    .S(net202),
    .X(_11874_));
 sg13g2_and3_1 _18785_ (.X(_11875_),
    .A(net422),
    .B(_11872_),
    .C(_11874_));
 sg13g2_mux2_1 _18786_ (.A0(_11862_),
    .A1(_11873_),
    .S(net199),
    .X(_11876_));
 sg13g2_nand2_1 _18787_ (.Y(_11877_),
    .A(net422),
    .B(_11876_));
 sg13g2_inv_1 _18788_ (.Y(_11878_),
    .A(_11860_));
 sg13g2_a22oi_1 _18789_ (.Y(_11879_),
    .B1(_11660_),
    .B2(_11878_),
    .A2(_11559_),
    .A1(\cpu.ex.r_mult[15] ));
 sg13g2_o21ai_1 _18790_ (.B1(_11879_),
    .Y(_11880_),
    .A1(_11872_),
    .A2(_11877_));
 sg13g2_a221oi_1 _18791_ (.B2(_11859_),
    .C1(_11880_),
    .B1(_11875_),
    .A1(net422),
    .Y(_11881_),
    .A2(_11865_));
 sg13g2_nand2_1 _18792_ (.Y(\cpu.ex.c_mult[15] ),
    .A(net27),
    .B(_11881_));
 sg13g2_inv_1 _18793_ (.Y(_00000_),
    .A(net2));
 sg13g2_inv_1 _18794_ (.Y(_11882_),
    .A(_09677_));
 sg13g2_and3_1 _18795_ (.X(_00008_),
    .A(_09678_),
    .B(net779),
    .C(_11882_));
 sg13g2_and3_1 _18796_ (.X(_00005_),
    .A(net1107),
    .B(net779),
    .C(_09669_));
 sg13g2_buf_1 _18797_ (.A(\cpu.qspi.r_state[11] ),
    .X(_11883_));
 sg13g2_buf_1 _18798_ (.A(net783),
    .X(_11884_));
 sg13g2_and2_1 _18799_ (.A(_11883_),
    .B(net648),
    .X(_00004_));
 sg13g2_buf_2 _18800_ (.A(\cpu.qspi.r_state[10] ),
    .X(_11885_));
 sg13g2_and2_1 _18801_ (.A(_11885_),
    .B(_11884_),
    .X(_00003_));
 sg13g2_buf_2 _18802_ (.A(\cpu.qspi.r_state[15] ),
    .X(_11886_));
 sg13g2_and2_1 _18803_ (.A(_11886_),
    .B(net779),
    .X(_00002_));
 sg13g2_inv_1 _18804_ (.Y(_11887_),
    .A(_09673_));
 sg13g2_nor3_1 _18805_ (.A(_11887_),
    .B(net684),
    .C(net600),
    .Y(_00001_));
 sg13g2_nor2_1 _18806_ (.A(_09700_),
    .B(_09702_),
    .Y(_00007_));
 sg13g2_inv_1 _18807_ (.Y(_11888_),
    .A(\cpu.cond[1] ));
 sg13g2_a21o_1 _18808_ (.A2(_10962_),
    .A1(_10357_),
    .B1(_10964_),
    .X(_11889_));
 sg13g2_nand4_1 _18809_ (.B(_10667_),
    .C(_11889_),
    .A(_10854_),
    .Y(_11890_),
    .D(_11387_));
 sg13g2_nor3_1 _18810_ (.A(_11124_),
    .B(_11096_),
    .C(_11890_),
    .Y(_11891_));
 sg13g2_nor4_1 _18811_ (.A(_11025_),
    .B(_10936_),
    .C(_10605_),
    .D(_10291_),
    .Y(_11892_));
 sg13g2_nor2b_1 _18812_ (.A(_10358_),
    .B_N(_10387_),
    .Y(_11893_));
 sg13g2_nor4_1 _18813_ (.A(_10767_),
    .B(_10499_),
    .C(_10258_),
    .D(_11893_),
    .Y(_11894_));
 sg13g2_nand4_1 _18814_ (.B(_11891_),
    .C(_11892_),
    .A(_10736_),
    .Y(_11895_),
    .D(_11894_));
 sg13g2_a21oi_1 _18815_ (.A1(_11888_),
    .A2(_11895_),
    .Y(_11896_),
    .B1(_11232_));
 sg13g2_xnor2_1 _18816_ (.Y(_11897_),
    .A(_09021_),
    .B(_11896_));
 sg13g2_a21oi_2 _18817_ (.B1(_10121_),
    .Y(_11898_),
    .A2(_11897_),
    .A1(_10107_));
 sg13g2_nor2_1 _18818_ (.A(_11508_),
    .B(_11898_),
    .Y(_11899_));
 sg13g2_buf_1 _18819_ (.A(_11501_),
    .X(_11900_));
 sg13g2_nor2b_1 _18820_ (.A(_11899_),
    .B_N(net729),
    .Y(_00053_));
 sg13g2_buf_2 _18821_ (.A(\cpu.qspi.r_state[13] ),
    .X(_11901_));
 sg13g2_and2_1 _18822_ (.A(_11901_),
    .B(net779),
    .X(_00006_));
 sg13g2_buf_2 _18823_ (.A(\cpu.qspi.r_state[3] ),
    .X(_11902_));
 sg13g2_and2_1 _18824_ (.A(_11902_),
    .B(net779),
    .X(_00009_));
 sg13g2_buf_1 _18825_ (.A(\cpu.qspi.r_state[6] ),
    .X(_11903_));
 sg13g2_and2_1 _18826_ (.A(_11903_),
    .B(net779),
    .X(_00010_));
 sg13g2_buf_1 _18827_ (.A(net778),
    .X(_11904_));
 sg13g2_nor3_1 _18828_ (.A(_08260_),
    .B(_08923_),
    .C(_11904_),
    .Y(_00052_));
 sg13g2_or2_1 _18829_ (.X(_11905_),
    .B(_09117_),
    .A(_09057_));
 sg13g2_buf_1 _18830_ (.A(_11905_),
    .X(_11906_));
 sg13g2_nor3_1 _18831_ (.A(_09111_),
    .B(_09132_),
    .C(_11906_),
    .Y(_11907_));
 sg13g2_a21oi_1 _18832_ (.A1(net378),
    .A2(_11906_),
    .Y(_11908_),
    .B1(_11907_));
 sg13g2_nand2_1 _18833_ (.Y(_11909_),
    .A(_09162_),
    .B(_11908_));
 sg13g2_buf_1 _18834_ (.A(_00205_),
    .X(_11910_));
 sg13g2_nor2_1 _18835_ (.A(_09117_),
    .B(net1110),
    .Y(_11911_));
 sg13g2_buf_1 _18836_ (.A(\cpu.spi.r_sel[1] ),
    .X(_11912_));
 sg13g2_buf_1 _18837_ (.A(_11912_),
    .X(_11913_));
 sg13g2_buf_1 _18838_ (.A(_11913_),
    .X(_11914_));
 sg13g2_buf_1 _18839_ (.A(\cpu.spi.r_src[2] ),
    .X(_11915_));
 sg13g2_inv_1 _18840_ (.Y(_11916_),
    .A(_00261_));
 sg13g2_buf_1 _18841_ (.A(\cpu.spi.r_sel[0] ),
    .X(_11917_));
 sg13g2_buf_1 _18842_ (.A(_11917_),
    .X(_11918_));
 sg13g2_mux2_1 _18843_ (.A0(_11915_),
    .A1(_11916_),
    .S(_11918_),
    .X(_11919_));
 sg13g2_nand2_1 _18844_ (.Y(_11920_),
    .A(net995),
    .B(_00262_));
 sg13g2_o21ai_1 _18845_ (.B1(_11920_),
    .Y(_11921_),
    .A1(net995),
    .A2(_11916_));
 sg13g2_nor2_1 _18846_ (.A(_11913_),
    .B(_11921_),
    .Y(_11922_));
 sg13g2_a21oi_2 _18847_ (.B1(_11922_),
    .Y(_11923_),
    .A2(_11919_),
    .A1(_11914_));
 sg13g2_a21oi_1 _18848_ (.A1(_11910_),
    .A2(_11911_),
    .Y(_11924_),
    .B1(_11923_));
 sg13g2_nor2_1 _18849_ (.A(_09058_),
    .B(net1110),
    .Y(_11925_));
 sg13g2_inv_2 _18850_ (.Y(_11926_),
    .A(_11912_));
 sg13g2_buf_1 _18851_ (.A(\cpu.spi.r_mode[0][1] ),
    .X(_11927_));
 sg13g2_buf_1 _18852_ (.A(\cpu.spi.r_mode[1][1] ),
    .X(_11928_));
 sg13g2_buf_1 _18853_ (.A(net995),
    .X(_11929_));
 sg13g2_buf_1 _18854_ (.A(net858),
    .X(_11930_));
 sg13g2_mux2_1 _18855_ (.A0(_11927_),
    .A1(_11928_),
    .S(net728),
    .X(_11931_));
 sg13g2_nor2_1 _18856_ (.A(_11926_),
    .B(_11917_),
    .Y(_11932_));
 sg13g2_buf_1 _18857_ (.A(\cpu.spi.r_mode[2][1] ),
    .X(_11933_));
 sg13g2_a22oi_1 _18858_ (.Y(_11934_),
    .B1(_11932_),
    .B2(_11933_),
    .A2(_11931_),
    .A1(_11926_));
 sg13g2_xnor2_1 _18859_ (.Y(_11935_),
    .A(_11925_),
    .B(_11934_));
 sg13g2_nand2_1 _18860_ (.Y(_11936_),
    .A(_11910_),
    .B(_11911_));
 sg13g2_buf_1 _18861_ (.A(_09781_),
    .X(_11937_));
 sg13g2_buf_1 _18862_ (.A(net994),
    .X(_11938_));
 sg13g2_buf_1 _18863_ (.A(net763),
    .X(_11939_));
 sg13g2_nand2_1 _18864_ (.Y(_11940_),
    .A(net646),
    .B(_00262_));
 sg13g2_o21ai_1 _18865_ (.B1(_11940_),
    .Y(_11941_),
    .A1(net646),
    .A2(_11916_));
 sg13g2_buf_1 _18866_ (.A(_09174_),
    .X(_11942_));
 sg13g2_nand3_1 _18867_ (.B(net645),
    .C(_11915_),
    .A(_11938_),
    .Y(_11943_));
 sg13g2_o21ai_1 _18868_ (.B1(_11943_),
    .Y(_11944_),
    .A1(net857),
    .A2(_11941_));
 sg13g2_nor2b_1 _18869_ (.A(_11936_),
    .B_N(_11944_),
    .Y(_11945_));
 sg13g2_buf_1 _18870_ (.A(net857),
    .X(_11946_));
 sg13g2_buf_1 _18871_ (.A(net646),
    .X(_11947_));
 sg13g2_buf_1 _18872_ (.A(net585),
    .X(_11948_));
 sg13g2_nand2b_1 _18873_ (.Y(_11949_),
    .B(net585),
    .A_N(_11927_));
 sg13g2_o21ai_1 _18874_ (.B1(_11949_),
    .Y(_11950_),
    .A1(_11948_),
    .A2(_11933_));
 sg13g2_mux2_1 _18875_ (.A0(_11927_),
    .A1(_11928_),
    .S(net585),
    .X(_11951_));
 sg13g2_nor2_1 _18876_ (.A(net727),
    .B(_11951_),
    .Y(_11952_));
 sg13g2_a21oi_1 _18877_ (.A1(net727),
    .A2(_11950_),
    .Y(_11953_),
    .B1(_11952_));
 sg13g2_a22oi_1 _18878_ (.Y(_11954_),
    .B1(_11945_),
    .B2(_11953_),
    .A2(_11935_),
    .A1(_11924_));
 sg13g2_nor2_1 _18879_ (.A(_11924_),
    .B(_11945_),
    .Y(_11955_));
 sg13g2_buf_1 _18880_ (.A(\cpu.gpio.genblk1[3].srcs_o[5] ),
    .X(_11956_));
 sg13g2_o21ai_1 _18881_ (.B1(net1091),
    .Y(_11957_),
    .A1(_11909_),
    .A2(_11955_));
 sg13g2_o21ai_1 _18882_ (.B1(_11957_),
    .Y(_00295_),
    .A1(_11909_),
    .A2(_11954_));
 sg13g2_nor2b_1 _18883_ (.A(_11909_),
    .B_N(_11955_),
    .Y(_11958_));
 sg13g2_buf_1 _18884_ (.A(_11936_),
    .X(_11959_));
 sg13g2_nor2b_1 _18885_ (.A(net726),
    .B_N(_11953_),
    .Y(_11960_));
 sg13g2_a21oi_1 _18886_ (.A1(net726),
    .A2(_11935_),
    .Y(_11961_),
    .B1(_11960_));
 sg13g2_buf_1 _18887_ (.A(\cpu.gpio.genblk1[3].srcs_o[4] ),
    .X(_11962_));
 sg13g2_nor2_1 _18888_ (.A(net1090),
    .B(_11958_),
    .Y(_11963_));
 sg13g2_a21oi_1 _18889_ (.A1(_11958_),
    .A2(_11961_),
    .Y(_00296_),
    .B1(_11963_));
 sg13g2_buf_1 _18890_ (.A(\cpu.gpio.genblk1[3].srcs_o[3] ),
    .X(_11964_));
 sg13g2_buf_1 _18891_ (.A(net1033),
    .X(_11965_));
 sg13g2_mux2_1 _18892_ (.A0(\cpu.spi.r_out[7] ),
    .A1(net1104),
    .S(_11965_),
    .X(_11966_));
 sg13g2_inv_1 _18893_ (.Y(_11967_),
    .A(_00203_));
 sg13g2_mux2_1 _18894_ (.A0(_11967_),
    .A1(\cpu.spi.r_mode[1][0] ),
    .S(_11917_),
    .X(_11968_));
 sg13g2_a22oi_1 _18895_ (.Y(_11969_),
    .B1(_11968_),
    .B2(_11926_),
    .A2(_11932_),
    .A1(\cpu.spi.r_mode[2][0] ));
 sg13g2_buf_1 _18896_ (.A(_11969_),
    .X(_11970_));
 sg13g2_nand3_1 _18897_ (.B(_09108_),
    .C(_11970_),
    .A(net1033),
    .Y(_11971_));
 sg13g2_o21ai_1 _18898_ (.B1(_09125_),
    .Y(_11972_),
    .A1(net1110),
    .A2(_11906_));
 sg13g2_nand2_1 _18899_ (.Y(_11973_),
    .A(net379),
    .B(_11970_));
 sg13g2_a21o_1 _18900_ (.A2(_09061_),
    .A1(_00199_),
    .B1(_09117_),
    .X(_11974_));
 sg13g2_o21ai_1 _18901_ (.B1(_09117_),
    .Y(_11975_),
    .A1(net378),
    .A2(_11970_));
 sg13g2_nand2_1 _18902_ (.Y(_11976_),
    .A(_09114_),
    .B(_11975_));
 sg13g2_o21ai_1 _18903_ (.B1(_11976_),
    .Y(_11977_),
    .A1(_11973_),
    .A2(_11974_));
 sg13g2_nand2_1 _18904_ (.Y(_11978_),
    .A(net901),
    .B(_11977_));
 sg13g2_a21oi_1 _18905_ (.A1(_11971_),
    .A2(_11972_),
    .Y(_11979_),
    .B1(_11978_));
 sg13g2_nor2b_1 _18906_ (.A(_11923_),
    .B_N(_11979_),
    .Y(_11980_));
 sg13g2_mux2_1 _18907_ (.A0(net1089),
    .A1(_11966_),
    .S(_11980_),
    .X(_00297_));
 sg13g2_buf_1 _18908_ (.A(\cpu.gpio.genblk1[3].srcs_o[2] ),
    .X(_11981_));
 sg13g2_nand2_1 _18909_ (.Y(_11982_),
    .A(_11923_),
    .B(_11979_));
 sg13g2_mux2_1 _18910_ (.A0(_11966_),
    .A1(net1088),
    .S(_11982_),
    .X(_00298_));
 sg13g2_nand2_1 _18911_ (.Y(_11983_),
    .A(_08125_),
    .B(_09166_));
 sg13g2_buf_2 _18912_ (.A(_00254_),
    .X(_11984_));
 sg13g2_buf_2 _18913_ (.A(_11984_),
    .X(_11985_));
 sg13g2_o21ai_1 _18914_ (.B1(net993),
    .Y(_11986_),
    .A1(_08127_),
    .A2(_11983_));
 sg13g2_buf_2 _18915_ (.A(_11986_),
    .X(_11987_));
 sg13g2_buf_2 _18916_ (.A(net768),
    .X(_11988_));
 sg13g2_nand2_1 _18917_ (.Y(_11989_),
    .A(net644),
    .B(_09210_));
 sg13g2_buf_2 _18918_ (.A(\cpu.dcache.r_offset[2] ),
    .X(_11990_));
 sg13g2_buf_1 _18919_ (.A(\cpu.dcache.r_offset[1] ),
    .X(_11991_));
 sg13g2_and2_1 _18920_ (.A(_11991_),
    .B(\cpu.dcache.r_offset[0] ),
    .X(_11992_));
 sg13g2_buf_1 _18921_ (.A(_11992_),
    .X(_11993_));
 sg13g2_nand3_1 _18922_ (.B(\cpu.d_wstrobe_d ),
    .C(_11993_),
    .A(_11990_),
    .Y(_11994_));
 sg13g2_buf_1 _18923_ (.A(_11994_),
    .X(_11995_));
 sg13g2_nor2_1 _18924_ (.A(_09182_),
    .B(_08180_),
    .Y(_11996_));
 sg13g2_nand2_1 _18925_ (.Y(_11997_),
    .A(_09168_),
    .B(_11996_));
 sg13g2_a21o_1 _18926_ (.A2(net643),
    .A1(_11524_),
    .B1(_11997_),
    .X(_11998_));
 sg13g2_buf_1 _18927_ (.A(_11998_),
    .X(_11999_));
 sg13g2_or2_1 _18928_ (.X(_12000_),
    .B(_11999_),
    .A(_11989_));
 sg13g2_buf_1 _18929_ (.A(_12000_),
    .X(_12001_));
 sg13g2_nor2_1 _18930_ (.A(_11987_),
    .B(_12001_),
    .Y(_12002_));
 sg13g2_buf_2 _18931_ (.A(_12002_),
    .X(_12003_));
 sg13g2_buf_1 _18932_ (.A(_12003_),
    .X(_12004_));
 sg13g2_buf_1 _18933_ (.A(uio_in[0]),
    .X(_12005_));
 sg13g2_buf_1 _18934_ (.A(_12005_),
    .X(_12006_));
 sg13g2_buf_2 _18935_ (.A(net1087),
    .X(_12007_));
 sg13g2_buf_1 _18936_ (.A(_11989_),
    .X(_12008_));
 sg13g2_buf_1 _18937_ (.A(\cpu.d_wstrobe_d ),
    .X(_12009_));
 sg13g2_buf_1 _18938_ (.A(_00255_),
    .X(_12010_));
 sg13g2_buf_1 _18939_ (.A(_12010_),
    .X(_12011_));
 sg13g2_buf_1 _18940_ (.A(\cpu.dcache.r_offset[0] ),
    .X(_12012_));
 sg13g2_inv_2 _18941_ (.Y(_12013_),
    .A(net1085));
 sg13g2_nor2_1 _18942_ (.A(_11991_),
    .B(_12013_),
    .Y(_12014_));
 sg13g2_nand3_1 _18943_ (.B(net991),
    .C(_12014_),
    .A(net1086),
    .Y(_12015_));
 sg13g2_buf_2 _18944_ (.A(_12015_),
    .X(_12016_));
 sg13g2_nor2_1 _18945_ (.A(net519),
    .B(_12016_),
    .Y(_12017_));
 sg13g2_buf_2 _18946_ (.A(_12017_),
    .X(_12018_));
 sg13g2_nor2b_1 _18947_ (.A(_12018_),
    .B_N(\cpu.dcache.r_data[0][0] ),
    .Y(_12019_));
 sg13g2_a21oi_1 _18948_ (.A1(net992),
    .A2(_12018_),
    .Y(_12020_),
    .B1(_12019_));
 sg13g2_nand2_1 _18949_ (.Y(_12021_),
    .A(_09927_),
    .B(net62));
 sg13g2_o21ai_1 _18950_ (.B1(_12021_),
    .Y(_00299_),
    .A1(_12004_),
    .A2(_12020_));
 sg13g2_nor2_1 _18951_ (.A(_08126_),
    .B(_08181_),
    .Y(_12022_));
 sg13g2_mux2_1 _18952_ (.A0(_09873_),
    .A1(_11984_),
    .S(_08128_),
    .X(_12023_));
 sg13g2_nand2_1 _18953_ (.Y(_12024_),
    .A(_12022_),
    .B(_12023_));
 sg13g2_buf_2 _18954_ (.A(_12024_),
    .X(_12025_));
 sg13g2_nor2_1 _18955_ (.A(_12001_),
    .B(_12025_),
    .Y(_12026_));
 sg13g2_buf_2 _18956_ (.A(_12026_),
    .X(_12027_));
 sg13g2_buf_1 _18957_ (.A(_12027_),
    .X(_12028_));
 sg13g2_buf_1 _18958_ (.A(uio_in[2]),
    .X(_12029_));
 sg13g2_buf_1 _18959_ (.A(_12029_),
    .X(_12030_));
 sg13g2_buf_2 _18960_ (.A(net1084),
    .X(_12031_));
 sg13g2_nand3_1 _18961_ (.B(net991),
    .C(_11993_),
    .A(net1086),
    .Y(_12032_));
 sg13g2_buf_2 _18962_ (.A(_12032_),
    .X(_12033_));
 sg13g2_nor2_1 _18963_ (.A(net519),
    .B(_12033_),
    .Y(_12034_));
 sg13g2_buf_2 _18964_ (.A(_12034_),
    .X(_12035_));
 sg13g2_nor2b_1 _18965_ (.A(_12035_),
    .B_N(\cpu.dcache.r_data[0][10] ),
    .Y(_12036_));
 sg13g2_a21oi_1 _18966_ (.A1(net990),
    .A2(_12035_),
    .Y(_12037_),
    .B1(_12036_));
 sg13g2_nand2_1 _18967_ (.Y(_12038_),
    .A(_08127_),
    .B(_12022_));
 sg13g2_buf_1 _18968_ (.A(_12038_),
    .X(_12039_));
 sg13g2_buf_1 _18969_ (.A(_12039_),
    .X(_12040_));
 sg13g2_mux2_1 _18970_ (.A0(_09986_),
    .A1(_09881_),
    .S(_12040_),
    .X(_12041_));
 sg13g2_buf_2 _18971_ (.A(_12041_),
    .X(_12042_));
 sg13g2_buf_1 _18972_ (.A(_12042_),
    .X(_12043_));
 sg13g2_nand2_1 _18973_ (.Y(_12044_),
    .A(net421),
    .B(_12027_));
 sg13g2_o21ai_1 _18974_ (.B1(_12044_),
    .Y(_00300_),
    .A1(_12028_),
    .A2(_12037_));
 sg13g2_buf_1 _18975_ (.A(uio_in[3]),
    .X(_12045_));
 sg13g2_buf_1 _18976_ (.A(_12045_),
    .X(_12046_));
 sg13g2_buf_2 _18977_ (.A(net1083),
    .X(_12047_));
 sg13g2_nor2b_1 _18978_ (.A(_12035_),
    .B_N(\cpu.dcache.r_data[0][11] ),
    .Y(_12048_));
 sg13g2_a21oi_1 _18979_ (.A1(net989),
    .A2(_12035_),
    .Y(_12049_),
    .B1(_12048_));
 sg13g2_mux2_1 _18980_ (.A0(_09991_),
    .A1(_09890_),
    .S(net584),
    .X(_12050_));
 sg13g2_buf_2 _18981_ (.A(_12050_),
    .X(_12051_));
 sg13g2_nand2_1 _18982_ (.Y(_12052_),
    .A(_12028_),
    .B(_12051_));
 sg13g2_o21ai_1 _18983_ (.B1(_12052_),
    .Y(_00301_),
    .A1(net61),
    .A2(_12049_));
 sg13g2_nor2b_1 _18984_ (.A(net1085),
    .B_N(_11991_),
    .Y(_12053_));
 sg13g2_nand3_1 _18985_ (.B(_12011_),
    .C(_12053_),
    .A(net1086),
    .Y(_12054_));
 sg13g2_buf_2 _18986_ (.A(_12054_),
    .X(_12055_));
 sg13g2_nor2_1 _18987_ (.A(net519),
    .B(_12055_),
    .Y(_12056_));
 sg13g2_buf_2 _18988_ (.A(_12056_),
    .X(_12057_));
 sg13g2_nor2b_1 _18989_ (.A(_12057_),
    .B_N(\cpu.dcache.r_data[0][12] ),
    .Y(_12058_));
 sg13g2_a21oi_1 _18990_ (.A1(net992),
    .A2(_12057_),
    .Y(_12059_),
    .B1(_12058_));
 sg13g2_inv_2 _18991_ (.Y(_12060_),
    .A(\cpu.dcache.wdata[12] ));
 sg13g2_nand2_1 _18992_ (.Y(_12061_),
    .A(net1105),
    .B(net584));
 sg13g2_o21ai_1 _18993_ (.B1(_12061_),
    .Y(_12062_),
    .A1(_12060_),
    .A2(net584));
 sg13g2_buf_2 _18994_ (.A(_12062_),
    .X(_12063_));
 sg13g2_nand2_1 _18995_ (.Y(_12064_),
    .A(net61),
    .B(_12063_));
 sg13g2_o21ai_1 _18996_ (.B1(_12064_),
    .Y(_00302_),
    .A1(net61),
    .A2(_12059_));
 sg13g2_buf_1 _18997_ (.A(uio_in[1]),
    .X(_12065_));
 sg13g2_buf_1 _18998_ (.A(_12065_),
    .X(_12066_));
 sg13g2_buf_2 _18999_ (.A(net1082),
    .X(_12067_));
 sg13g2_nor2b_1 _19000_ (.A(_12057_),
    .B_N(\cpu.dcache.r_data[0][13] ),
    .Y(_12068_));
 sg13g2_a21oi_1 _19001_ (.A1(net988),
    .A2(_12057_),
    .Y(_12069_),
    .B1(_12068_));
 sg13g2_inv_2 _19002_ (.Y(_12070_),
    .A(\cpu.dcache.wdata[13] ));
 sg13g2_nand2_1 _19003_ (.Y(_12071_),
    .A(_09901_),
    .B(_12039_));
 sg13g2_o21ai_1 _19004_ (.B1(_12071_),
    .Y(_12072_),
    .A1(_12070_),
    .A2(net584));
 sg13g2_buf_2 _19005_ (.A(_12072_),
    .X(_12073_));
 sg13g2_nand2_1 _19006_ (.Y(_12074_),
    .A(_12027_),
    .B(_12073_));
 sg13g2_o21ai_1 _19007_ (.B1(_12074_),
    .Y(_00303_),
    .A1(net61),
    .A2(_12069_));
 sg13g2_nor2b_1 _19008_ (.A(_12057_),
    .B_N(\cpu.dcache.r_data[0][14] ),
    .Y(_12075_));
 sg13g2_a21oi_1 _19009_ (.A1(net990),
    .A2(_12057_),
    .Y(_12076_),
    .B1(_12075_));
 sg13g2_inv_2 _19010_ (.Y(_12077_),
    .A(\cpu.dcache.wdata[14] ));
 sg13g2_nand2_1 _19011_ (.Y(_12078_),
    .A(_09907_),
    .B(_12039_));
 sg13g2_o21ai_1 _19012_ (.B1(_12078_),
    .Y(_12079_),
    .A1(_12077_),
    .A2(net584));
 sg13g2_buf_2 _19013_ (.A(_12079_),
    .X(_12080_));
 sg13g2_nand2_1 _19014_ (.Y(_12081_),
    .A(_12027_),
    .B(_12080_));
 sg13g2_o21ai_1 _19015_ (.B1(_12081_),
    .Y(_00304_),
    .A1(net61),
    .A2(_12076_));
 sg13g2_nor2b_1 _19016_ (.A(_12057_),
    .B_N(\cpu.dcache.r_data[0][15] ),
    .Y(_12082_));
 sg13g2_a21oi_1 _19017_ (.A1(net989),
    .A2(_12057_),
    .Y(_12083_),
    .B1(_12082_));
 sg13g2_inv_2 _19018_ (.Y(_12084_),
    .A(\cpu.dcache.wdata[15] ));
 sg13g2_nand2_1 _19019_ (.Y(_12085_),
    .A(net1104),
    .B(_12039_));
 sg13g2_o21ai_1 _19020_ (.B1(_12085_),
    .Y(_12086_),
    .A1(_12084_),
    .A2(_12040_));
 sg13g2_buf_2 _19021_ (.A(_12086_),
    .X(_12087_));
 sg13g2_nand2_1 _19022_ (.Y(_12088_),
    .A(_12027_),
    .B(_12087_));
 sg13g2_o21ai_1 _19023_ (.B1(_12088_),
    .Y(_00305_),
    .A1(net61),
    .A2(_12083_));
 sg13g2_o21ai_1 _19024_ (.B1(net755),
    .Y(_12089_),
    .A1(_08127_),
    .A2(_11983_));
 sg13g2_buf_2 _19025_ (.A(_12089_),
    .X(_12090_));
 sg13g2_nor2_1 _19026_ (.A(_12001_),
    .B(_12090_),
    .Y(_12091_));
 sg13g2_buf_1 _19027_ (.A(_12091_),
    .X(_12092_));
 sg13g2_buf_1 _19028_ (.A(_12092_),
    .X(_12093_));
 sg13g2_buf_1 _19029_ (.A(_11990_),
    .X(_12094_));
 sg13g2_nand3_1 _19030_ (.B(net1086),
    .C(_12014_),
    .A(net987),
    .Y(_12095_));
 sg13g2_buf_2 _19031_ (.A(_12095_),
    .X(_12096_));
 sg13g2_nor2_1 _19032_ (.A(net519),
    .B(_12096_),
    .Y(_12097_));
 sg13g2_buf_2 _19033_ (.A(_12097_),
    .X(_12098_));
 sg13g2_nor2b_1 _19034_ (.A(_12098_),
    .B_N(\cpu.dcache.r_data[0][16] ),
    .Y(_12099_));
 sg13g2_a21oi_1 _19035_ (.A1(net992),
    .A2(_12098_),
    .Y(_12100_),
    .B1(_12099_));
 sg13g2_nand2_1 _19036_ (.Y(_12101_),
    .A(_09927_),
    .B(net60));
 sg13g2_o21ai_1 _19037_ (.B1(_12101_),
    .Y(_00306_),
    .A1(net60),
    .A2(_12100_));
 sg13g2_nor2b_1 _19038_ (.A(_12098_),
    .B_N(\cpu.dcache.r_data[0][17] ),
    .Y(_12102_));
 sg13g2_a21oi_1 _19039_ (.A1(net988),
    .A2(_12098_),
    .Y(_12103_),
    .B1(_12102_));
 sg13g2_buf_1 _19040_ (.A(_09871_),
    .X(_12104_));
 sg13g2_nand2_1 _19041_ (.Y(_12105_),
    .A(net855),
    .B(net60));
 sg13g2_o21ai_1 _19042_ (.B1(_12105_),
    .Y(_00307_),
    .A1(net60),
    .A2(_12103_));
 sg13g2_buf_1 _19043_ (.A(_09883_),
    .X(_12106_));
 sg13g2_buf_2 _19044_ (.A(_12029_),
    .X(_12107_));
 sg13g2_mux2_1 _19045_ (.A0(\cpu.dcache.r_data[0][18] ),
    .A1(net1081),
    .S(_12098_),
    .X(_12108_));
 sg13g2_nor2_1 _19046_ (.A(_12092_),
    .B(_12108_),
    .Y(_12109_));
 sg13g2_a21oi_1 _19047_ (.A1(net725),
    .A2(net60),
    .Y(_00308_),
    .B1(_12109_));
 sg13g2_inv_1 _19048_ (.Y(_12110_),
    .A(net1106));
 sg13g2_buf_1 _19049_ (.A(_12110_),
    .X(_12111_));
 sg13g2_buf_1 _19050_ (.A(net854),
    .X(_12112_));
 sg13g2_buf_1 _19051_ (.A(_12045_),
    .X(_12113_));
 sg13g2_mux2_1 _19052_ (.A0(\cpu.dcache.r_data[0][19] ),
    .A1(net1080),
    .S(_12098_),
    .X(_12114_));
 sg13g2_nor2_1 _19053_ (.A(_12092_),
    .B(_12114_),
    .Y(_12115_));
 sg13g2_a21oi_1 _19054_ (.A1(net724),
    .A2(net60),
    .Y(_00309_),
    .B1(_12115_));
 sg13g2_nor2b_1 _19055_ (.A(_12018_),
    .B_N(\cpu.dcache.r_data[0][1] ),
    .Y(_12116_));
 sg13g2_a21oi_1 _19056_ (.A1(net988),
    .A2(_12018_),
    .Y(_12117_),
    .B1(_12116_));
 sg13g2_nand2_1 _19057_ (.Y(_12118_),
    .A(_12104_),
    .B(net62));
 sg13g2_o21ai_1 _19058_ (.B1(_12118_),
    .Y(_00310_),
    .A1(net62),
    .A2(_12117_));
 sg13g2_inv_1 _19059_ (.Y(_12119_),
    .A(net1105));
 sg13g2_buf_1 _19060_ (.A(_12119_),
    .X(_12120_));
 sg13g2_buf_1 _19061_ (.A(net853),
    .X(_12121_));
 sg13g2_buf_1 _19062_ (.A(_12005_),
    .X(_12122_));
 sg13g2_nor2_1 _19063_ (.A(_11991_),
    .B(net1085),
    .Y(_12123_));
 sg13g2_nand3_1 _19064_ (.B(net1086),
    .C(_12123_),
    .A(_11990_),
    .Y(_12124_));
 sg13g2_buf_2 _19065_ (.A(_12124_),
    .X(_12125_));
 sg13g2_nor2_1 _19066_ (.A(net519),
    .B(_12125_),
    .Y(_12126_));
 sg13g2_buf_2 _19067_ (.A(_12126_),
    .X(_12127_));
 sg13g2_mux2_1 _19068_ (.A0(\cpu.dcache.r_data[0][20] ),
    .A1(net1079),
    .S(_12127_),
    .X(_12128_));
 sg13g2_nor2_1 _19069_ (.A(_12092_),
    .B(_12128_),
    .Y(_12129_));
 sg13g2_a21oi_1 _19070_ (.A1(_12121_),
    .A2(net60),
    .Y(_00311_),
    .B1(_12129_));
 sg13g2_nor2b_1 _19071_ (.A(_12127_),
    .B_N(\cpu.dcache.r_data[0][21] ),
    .Y(_12130_));
 sg13g2_a21oi_1 _19072_ (.A1(net988),
    .A2(_12127_),
    .Y(_12131_),
    .B1(_12130_));
 sg13g2_buf_1 _19073_ (.A(_09901_),
    .X(_12132_));
 sg13g2_nand2_1 _19074_ (.Y(_12133_),
    .A(_12132_),
    .B(_12092_));
 sg13g2_o21ai_1 _19075_ (.B1(_12133_),
    .Y(_00312_),
    .A1(net60),
    .A2(_12131_));
 sg13g2_nor2b_1 _19076_ (.A(_12127_),
    .B_N(\cpu.dcache.r_data[0][22] ),
    .Y(_12134_));
 sg13g2_a21oi_1 _19077_ (.A1(net990),
    .A2(_12127_),
    .Y(_12135_),
    .B1(_12134_));
 sg13g2_buf_1 _19078_ (.A(_09907_),
    .X(_12136_));
 sg13g2_nand2_1 _19079_ (.Y(_12137_),
    .A(_12136_),
    .B(_12092_));
 sg13g2_o21ai_1 _19080_ (.B1(_12137_),
    .Y(_00313_),
    .A1(_12093_),
    .A2(_12135_));
 sg13g2_inv_1 _19081_ (.Y(_12138_),
    .A(net1104));
 sg13g2_buf_1 _19082_ (.A(_12138_),
    .X(_12139_));
 sg13g2_buf_1 _19083_ (.A(net852),
    .X(_12140_));
 sg13g2_mux2_1 _19084_ (.A0(\cpu.dcache.r_data[0][23] ),
    .A1(net1080),
    .S(_12127_),
    .X(_12141_));
 sg13g2_nor2_1 _19085_ (.A(_12092_),
    .B(_12141_),
    .Y(_12142_));
 sg13g2_a21oi_1 _19086_ (.A1(net722),
    .A2(_12093_),
    .Y(_00314_),
    .B1(_12142_));
 sg13g2_buf_2 _19087_ (.A(_12005_),
    .X(_12143_));
 sg13g2_or2_1 _19088_ (.X(_12144_),
    .B(net643),
    .A(_12008_));
 sg13g2_buf_2 _19089_ (.A(_12144_),
    .X(_12145_));
 sg13g2_mux2_1 _19090_ (.A0(_12143_),
    .A1(\cpu.dcache.r_data[0][24] ),
    .S(_12145_),
    .X(_12146_));
 sg13g2_mux2_1 _19091_ (.A0(_09975_),
    .A1(_09859_),
    .S(net584),
    .X(_12147_));
 sg13g2_buf_2 _19092_ (.A(_12147_),
    .X(_12148_));
 sg13g2_buf_1 _19093_ (.A(_12148_),
    .X(_12149_));
 sg13g2_nor2_1 _19094_ (.A(_08127_),
    .B(_09776_),
    .Y(_12150_));
 sg13g2_a21oi_1 _19095_ (.A1(_08127_),
    .A2(_11984_),
    .Y(_12151_),
    .B1(_12150_));
 sg13g2_nand2_1 _19096_ (.Y(_12152_),
    .A(_12022_),
    .B(_12151_));
 sg13g2_buf_2 _19097_ (.A(_12152_),
    .X(_12153_));
 sg13g2_nor2_1 _19098_ (.A(_12001_),
    .B(_12153_),
    .Y(_12154_));
 sg13g2_buf_2 _19099_ (.A(_12154_),
    .X(_12155_));
 sg13g2_mux2_1 _19100_ (.A0(_12146_),
    .A1(_12149_),
    .S(net70),
    .X(_00315_));
 sg13g2_mux2_1 _19101_ (.A0(net1082),
    .A1(\cpu.dcache.r_data[0][25] ),
    .S(_12145_),
    .X(_12156_));
 sg13g2_inv_2 _19102_ (.Y(_12157_),
    .A(\cpu.dcache.wdata[9] ));
 sg13g2_nand2_1 _19103_ (.Y(_12158_),
    .A(_09870_),
    .B(net584));
 sg13g2_o21ai_1 _19104_ (.B1(_12158_),
    .Y(_12159_),
    .A1(_12157_),
    .A2(net584));
 sg13g2_buf_2 _19105_ (.A(_12159_),
    .X(_12160_));
 sg13g2_buf_1 _19106_ (.A(_12160_),
    .X(_12161_));
 sg13g2_mux2_1 _19107_ (.A0(_12156_),
    .A1(net369),
    .S(_12155_),
    .X(_00316_));
 sg13g2_mux2_1 _19108_ (.A0(net1081),
    .A1(\cpu.dcache.r_data[0][26] ),
    .S(_12145_),
    .X(_12162_));
 sg13g2_mux2_1 _19109_ (.A0(_12162_),
    .A1(_12043_),
    .S(net70),
    .X(_00317_));
 sg13g2_mux2_1 _19110_ (.A0(net1080),
    .A1(\cpu.dcache.r_data[0][27] ),
    .S(_12145_),
    .X(_12163_));
 sg13g2_buf_1 _19111_ (.A(_12051_),
    .X(_12164_));
 sg13g2_mux2_1 _19112_ (.A0(_12163_),
    .A1(_12164_),
    .S(_12155_),
    .X(_00318_));
 sg13g2_nand3_1 _19113_ (.B(net1086),
    .C(_12053_),
    .A(_12094_),
    .Y(_12165_));
 sg13g2_buf_2 _19114_ (.A(_12165_),
    .X(_12166_));
 sg13g2_nor2_1 _19115_ (.A(net519),
    .B(_12166_),
    .Y(_12167_));
 sg13g2_buf_2 _19116_ (.A(_12167_),
    .X(_12168_));
 sg13g2_nor2b_1 _19117_ (.A(_12168_),
    .B_N(\cpu.dcache.r_data[0][28] ),
    .Y(_12169_));
 sg13g2_a21oi_1 _19118_ (.A1(net992),
    .A2(_12168_),
    .Y(_12170_),
    .B1(_12169_));
 sg13g2_buf_1 _19119_ (.A(_12063_),
    .X(_12171_));
 sg13g2_nand2_1 _19120_ (.Y(_12172_),
    .A(net368),
    .B(net70));
 sg13g2_o21ai_1 _19121_ (.B1(_12172_),
    .Y(_00319_),
    .A1(net70),
    .A2(_12170_));
 sg13g2_nor2b_1 _19122_ (.A(_12168_),
    .B_N(\cpu.dcache.r_data[0][29] ),
    .Y(_12173_));
 sg13g2_a21oi_1 _19123_ (.A1(net988),
    .A2(_12168_),
    .Y(_12174_),
    .B1(_12173_));
 sg13g2_buf_1 _19124_ (.A(_12073_),
    .X(_12175_));
 sg13g2_nand2_1 _19125_ (.Y(_12176_),
    .A(net418),
    .B(net70));
 sg13g2_o21ai_1 _19126_ (.B1(_12176_),
    .Y(_00320_),
    .A1(net70),
    .A2(_12174_));
 sg13g2_mux2_1 _19127_ (.A0(\cpu.dcache.r_data[0][2] ),
    .A1(net1081),
    .S(_12018_),
    .X(_12177_));
 sg13g2_nor2_1 _19128_ (.A(_12003_),
    .B(_12177_),
    .Y(_12178_));
 sg13g2_a21oi_1 _19129_ (.A1(_12106_),
    .A2(_12004_),
    .Y(_00321_),
    .B1(_12178_));
 sg13g2_nor2b_1 _19130_ (.A(_12168_),
    .B_N(\cpu.dcache.r_data[0][30] ),
    .Y(_12179_));
 sg13g2_a21oi_1 _19131_ (.A1(net990),
    .A2(_12168_),
    .Y(_12180_),
    .B1(_12179_));
 sg13g2_buf_1 _19132_ (.A(_12080_),
    .X(_12181_));
 sg13g2_nand2_1 _19133_ (.Y(_12182_),
    .A(net417),
    .B(_12154_));
 sg13g2_o21ai_1 _19134_ (.B1(_12182_),
    .Y(_00322_),
    .A1(net70),
    .A2(_12180_));
 sg13g2_nor2b_1 _19135_ (.A(_12168_),
    .B_N(\cpu.dcache.r_data[0][31] ),
    .Y(_12183_));
 sg13g2_a21oi_1 _19136_ (.A1(net989),
    .A2(_12168_),
    .Y(_12184_),
    .B1(_12183_));
 sg13g2_buf_1 _19137_ (.A(_12087_),
    .X(_12185_));
 sg13g2_nand2_1 _19138_ (.Y(_12186_),
    .A(_12185_),
    .B(_12154_));
 sg13g2_o21ai_1 _19139_ (.B1(_12186_),
    .Y(_00323_),
    .A1(net70),
    .A2(_12184_));
 sg13g2_mux2_1 _19140_ (.A0(\cpu.dcache.r_data[0][3] ),
    .A1(net1080),
    .S(_12018_),
    .X(_12187_));
 sg13g2_nor2_1 _19141_ (.A(_12003_),
    .B(_12187_),
    .Y(_12188_));
 sg13g2_a21oi_1 _19142_ (.A1(_12112_),
    .A2(net62),
    .Y(_00324_),
    .B1(_12188_));
 sg13g2_nand3_1 _19143_ (.B(net991),
    .C(_12123_),
    .A(net1086),
    .Y(_12189_));
 sg13g2_buf_2 _19144_ (.A(_12189_),
    .X(_12190_));
 sg13g2_nor2_1 _19145_ (.A(net519),
    .B(_12190_),
    .Y(_12191_));
 sg13g2_buf_2 _19146_ (.A(_12191_),
    .X(_12192_));
 sg13g2_mux2_1 _19147_ (.A0(\cpu.dcache.r_data[0][4] ),
    .A1(_12122_),
    .S(_12192_),
    .X(_12193_));
 sg13g2_nor2_1 _19148_ (.A(_12003_),
    .B(_12193_),
    .Y(_12194_));
 sg13g2_a21oi_1 _19149_ (.A1(net723),
    .A2(net62),
    .Y(_00325_),
    .B1(_12194_));
 sg13g2_nor2b_1 _19150_ (.A(_12192_),
    .B_N(\cpu.dcache.r_data[0][5] ),
    .Y(_12195_));
 sg13g2_a21oi_1 _19151_ (.A1(net988),
    .A2(_12192_),
    .Y(_12196_),
    .B1(_12195_));
 sg13g2_buf_1 _19152_ (.A(_09901_),
    .X(_12197_));
 sg13g2_nand2_1 _19153_ (.Y(_12198_),
    .A(_12197_),
    .B(_12003_));
 sg13g2_o21ai_1 _19154_ (.B1(_12198_),
    .Y(_00326_),
    .A1(net62),
    .A2(_12196_));
 sg13g2_nor2b_1 _19155_ (.A(_12192_),
    .B_N(\cpu.dcache.r_data[0][6] ),
    .Y(_12199_));
 sg13g2_a21oi_1 _19156_ (.A1(net990),
    .A2(_12192_),
    .Y(_12200_),
    .B1(_12199_));
 sg13g2_nand2_1 _19157_ (.Y(_12201_),
    .A(net985),
    .B(_12003_));
 sg13g2_o21ai_1 _19158_ (.B1(_12201_),
    .Y(_00327_),
    .A1(net62),
    .A2(_12200_));
 sg13g2_buf_1 _19159_ (.A(net1083),
    .X(_12202_));
 sg13g2_mux2_1 _19160_ (.A0(\cpu.dcache.r_data[0][7] ),
    .A1(_12202_),
    .S(_12192_),
    .X(_12203_));
 sg13g2_nor2_1 _19161_ (.A(_12003_),
    .B(_12203_),
    .Y(_12204_));
 sg13g2_a21oi_1 _19162_ (.A1(net722),
    .A2(net62),
    .Y(_00328_),
    .B1(_12204_));
 sg13g2_nor2b_1 _19163_ (.A(_12035_),
    .B_N(\cpu.dcache.r_data[0][8] ),
    .Y(_12205_));
 sg13g2_a21oi_1 _19164_ (.A1(net992),
    .A2(_12035_),
    .Y(_12206_),
    .B1(_12205_));
 sg13g2_nand2_1 _19165_ (.Y(_12207_),
    .A(_12027_),
    .B(_12148_));
 sg13g2_o21ai_1 _19166_ (.B1(_12207_),
    .Y(_00329_),
    .A1(net61),
    .A2(_12206_));
 sg13g2_buf_1 _19167_ (.A(_12066_),
    .X(_12208_));
 sg13g2_nor2b_1 _19168_ (.A(_12035_),
    .B_N(\cpu.dcache.r_data[0][9] ),
    .Y(_12209_));
 sg13g2_a21oi_1 _19169_ (.A1(net982),
    .A2(_12035_),
    .Y(_12210_),
    .B1(_12209_));
 sg13g2_nand2_1 _19170_ (.Y(_12211_),
    .A(_12027_),
    .B(_12160_));
 sg13g2_o21ai_1 _19171_ (.B1(_12211_),
    .Y(_00330_),
    .A1(net61),
    .A2(_12210_));
 sg13g2_buf_1 _19172_ (.A(net531),
    .X(_12212_));
 sg13g2_or2_1 _19173_ (.X(_12213_),
    .B(_11999_),
    .A(_12212_));
 sg13g2_buf_1 _19174_ (.A(_12213_),
    .X(_12214_));
 sg13g2_nor2_1 _19175_ (.A(_11987_),
    .B(_12214_),
    .Y(_12215_));
 sg13g2_buf_1 _19176_ (.A(_12215_),
    .X(_12216_));
 sg13g2_buf_1 _19177_ (.A(_12216_),
    .X(_12217_));
 sg13g2_nor2_1 _19178_ (.A(net457),
    .B(_12016_),
    .Y(_12218_));
 sg13g2_buf_2 _19179_ (.A(_12218_),
    .X(_12219_));
 sg13g2_nor2b_1 _19180_ (.A(_12219_),
    .B_N(\cpu.dcache.r_data[1][0] ),
    .Y(_12220_));
 sg13g2_a21oi_1 _19181_ (.A1(net992),
    .A2(_12219_),
    .Y(_12221_),
    .B1(_12220_));
 sg13g2_buf_1 _19182_ (.A(_09860_),
    .X(_12222_));
 sg13g2_nand2_1 _19183_ (.Y(_12223_),
    .A(net851),
    .B(net59));
 sg13g2_o21ai_1 _19184_ (.B1(_12223_),
    .Y(_00331_),
    .A1(net59),
    .A2(_12221_));
 sg13g2_nor2_1 _19185_ (.A(_12025_),
    .B(_12214_),
    .Y(_12224_));
 sg13g2_buf_2 _19186_ (.A(_12224_),
    .X(_12225_));
 sg13g2_buf_1 _19187_ (.A(_12225_),
    .X(_12226_));
 sg13g2_nor2_1 _19188_ (.A(net457),
    .B(_12033_),
    .Y(_12227_));
 sg13g2_buf_2 _19189_ (.A(_12227_),
    .X(_12228_));
 sg13g2_nor2b_1 _19190_ (.A(_12228_),
    .B_N(\cpu.dcache.r_data[1][10] ),
    .Y(_12229_));
 sg13g2_a21oi_1 _19191_ (.A1(net990),
    .A2(_12228_),
    .Y(_12230_),
    .B1(_12229_));
 sg13g2_nand2_1 _19192_ (.Y(_12231_),
    .A(net421),
    .B(net58));
 sg13g2_o21ai_1 _19193_ (.B1(_12231_),
    .Y(_00332_),
    .A1(net58),
    .A2(_12230_));
 sg13g2_nor2b_1 _19194_ (.A(_12228_),
    .B_N(\cpu.dcache.r_data[1][11] ),
    .Y(_12232_));
 sg13g2_a21oi_1 _19195_ (.A1(net989),
    .A2(_12228_),
    .Y(_12233_),
    .B1(_12232_));
 sg13g2_nand2_1 _19196_ (.Y(_12234_),
    .A(net419),
    .B(_12226_));
 sg13g2_o21ai_1 _19197_ (.B1(_12234_),
    .Y(_00333_),
    .A1(_12226_),
    .A2(_12233_));
 sg13g2_buf_1 _19198_ (.A(net1087),
    .X(_12235_));
 sg13g2_nor2_1 _19199_ (.A(net457),
    .B(_12055_),
    .Y(_12236_));
 sg13g2_buf_2 _19200_ (.A(_12236_),
    .X(_12237_));
 sg13g2_nor2b_1 _19201_ (.A(_12237_),
    .B_N(\cpu.dcache.r_data[1][12] ),
    .Y(_12238_));
 sg13g2_a21oi_1 _19202_ (.A1(net981),
    .A2(_12237_),
    .Y(_12239_),
    .B1(_12238_));
 sg13g2_nand2_1 _19203_ (.Y(_12240_),
    .A(net368),
    .B(_12225_));
 sg13g2_o21ai_1 _19204_ (.B1(_12240_),
    .Y(_00334_),
    .A1(net58),
    .A2(_12239_));
 sg13g2_nor2b_1 _19205_ (.A(_12237_),
    .B_N(\cpu.dcache.r_data[1][13] ),
    .Y(_12241_));
 sg13g2_a21oi_1 _19206_ (.A1(net982),
    .A2(_12237_),
    .Y(_12242_),
    .B1(_12241_));
 sg13g2_nand2_1 _19207_ (.Y(_12243_),
    .A(net418),
    .B(_12225_));
 sg13g2_o21ai_1 _19208_ (.B1(_12243_),
    .Y(_00335_),
    .A1(net58),
    .A2(_12242_));
 sg13g2_buf_1 _19209_ (.A(net1084),
    .X(_12244_));
 sg13g2_nor2b_1 _19210_ (.A(_12237_),
    .B_N(\cpu.dcache.r_data[1][14] ),
    .Y(_12245_));
 sg13g2_a21oi_1 _19211_ (.A1(net980),
    .A2(_12237_),
    .Y(_12246_),
    .B1(_12245_));
 sg13g2_nand2_1 _19212_ (.Y(_12247_),
    .A(net417),
    .B(_12225_));
 sg13g2_o21ai_1 _19213_ (.B1(_12247_),
    .Y(_00336_),
    .A1(net58),
    .A2(_12246_));
 sg13g2_nor2b_1 _19214_ (.A(_12237_),
    .B_N(\cpu.dcache.r_data[1][15] ),
    .Y(_12248_));
 sg13g2_a21oi_1 _19215_ (.A1(net989),
    .A2(_12237_),
    .Y(_12249_),
    .B1(_12248_));
 sg13g2_nand2_1 _19216_ (.Y(_12250_),
    .A(net416),
    .B(_12225_));
 sg13g2_o21ai_1 _19217_ (.B1(_12250_),
    .Y(_00337_),
    .A1(net58),
    .A2(_12249_));
 sg13g2_nor2_1 _19218_ (.A(_12090_),
    .B(_12214_),
    .Y(_12251_));
 sg13g2_buf_1 _19219_ (.A(_12251_),
    .X(_12252_));
 sg13g2_buf_1 _19220_ (.A(_12252_),
    .X(_12253_));
 sg13g2_nor2_1 _19221_ (.A(net457),
    .B(_12096_),
    .Y(_12254_));
 sg13g2_buf_2 _19222_ (.A(_12254_),
    .X(_12255_));
 sg13g2_nor2b_1 _19223_ (.A(_12255_),
    .B_N(\cpu.dcache.r_data[1][16] ),
    .Y(_12256_));
 sg13g2_a21oi_1 _19224_ (.A1(net981),
    .A2(_12255_),
    .Y(_12257_),
    .B1(_12256_));
 sg13g2_nand2_1 _19225_ (.Y(_12258_),
    .A(net851),
    .B(net57));
 sg13g2_o21ai_1 _19226_ (.B1(_12258_),
    .Y(_00338_),
    .A1(net57),
    .A2(_12257_));
 sg13g2_nor2b_1 _19227_ (.A(_12255_),
    .B_N(\cpu.dcache.r_data[1][17] ),
    .Y(_12259_));
 sg13g2_a21oi_1 _19228_ (.A1(net982),
    .A2(_12255_),
    .Y(_12260_),
    .B1(_12259_));
 sg13g2_nand2_1 _19229_ (.Y(_12261_),
    .A(net855),
    .B(net57));
 sg13g2_o21ai_1 _19230_ (.B1(_12261_),
    .Y(_00339_),
    .A1(net57),
    .A2(_12260_));
 sg13g2_buf_1 _19231_ (.A(_12029_),
    .X(_12262_));
 sg13g2_mux2_1 _19232_ (.A0(\cpu.dcache.r_data[1][18] ),
    .A1(net1078),
    .S(_12255_),
    .X(_12263_));
 sg13g2_nor2_1 _19233_ (.A(_12252_),
    .B(_12263_),
    .Y(_12264_));
 sg13g2_a21oi_1 _19234_ (.A1(net725),
    .A2(_12253_),
    .Y(_00340_),
    .B1(_12264_));
 sg13g2_mux2_1 _19235_ (.A0(\cpu.dcache.r_data[1][19] ),
    .A1(net983),
    .S(_12255_),
    .X(_12265_));
 sg13g2_nor2_1 _19236_ (.A(_12252_),
    .B(_12265_),
    .Y(_12266_));
 sg13g2_a21oi_1 _19237_ (.A1(net724),
    .A2(net57),
    .Y(_00341_),
    .B1(_12266_));
 sg13g2_nor2b_1 _19238_ (.A(_12219_),
    .B_N(\cpu.dcache.r_data[1][1] ),
    .Y(_12267_));
 sg13g2_a21oi_1 _19239_ (.A1(net982),
    .A2(_12219_),
    .Y(_12268_),
    .B1(_12267_));
 sg13g2_nand2_1 _19240_ (.Y(_12269_),
    .A(net855),
    .B(net59));
 sg13g2_o21ai_1 _19241_ (.B1(_12269_),
    .Y(_00342_),
    .A1(net59),
    .A2(_12268_));
 sg13g2_nor2_1 _19242_ (.A(net457),
    .B(_12125_),
    .Y(_12270_));
 sg13g2_buf_2 _19243_ (.A(_12270_),
    .X(_12271_));
 sg13g2_mux2_1 _19244_ (.A0(\cpu.dcache.r_data[1][20] ),
    .A1(net1079),
    .S(_12271_),
    .X(_12272_));
 sg13g2_nor2_1 _19245_ (.A(_12252_),
    .B(_12272_),
    .Y(_12273_));
 sg13g2_a21oi_1 _19246_ (.A1(net723),
    .A2(net57),
    .Y(_00343_),
    .B1(_12273_));
 sg13g2_nor2b_1 _19247_ (.A(_12271_),
    .B_N(\cpu.dcache.r_data[1][21] ),
    .Y(_12274_));
 sg13g2_a21oi_1 _19248_ (.A1(net982),
    .A2(_12271_),
    .Y(_12275_),
    .B1(_12274_));
 sg13g2_nand2_1 _19249_ (.Y(_12276_),
    .A(net984),
    .B(_12252_));
 sg13g2_o21ai_1 _19250_ (.B1(_12276_),
    .Y(_00344_),
    .A1(_12253_),
    .A2(_12275_));
 sg13g2_nor2b_1 _19251_ (.A(_12271_),
    .B_N(\cpu.dcache.r_data[1][22] ),
    .Y(_12277_));
 sg13g2_a21oi_1 _19252_ (.A1(net980),
    .A2(_12271_),
    .Y(_12278_),
    .B1(_12277_));
 sg13g2_nand2_1 _19253_ (.Y(_12279_),
    .A(net985),
    .B(_12252_));
 sg13g2_o21ai_1 _19254_ (.B1(_12279_),
    .Y(_00345_),
    .A1(net57),
    .A2(_12278_));
 sg13g2_mux2_1 _19255_ (.A0(\cpu.dcache.r_data[1][23] ),
    .A1(net983),
    .S(_12271_),
    .X(_12280_));
 sg13g2_nor2_1 _19256_ (.A(_12252_),
    .B(_12280_),
    .Y(_12281_));
 sg13g2_a21oi_1 _19257_ (.A1(net722),
    .A2(net57),
    .Y(_00346_),
    .B1(_12281_));
 sg13g2_nor2_1 _19258_ (.A(_12153_),
    .B(_12214_),
    .Y(_12282_));
 sg13g2_buf_2 _19259_ (.A(_12282_),
    .X(_12283_));
 sg13g2_buf_1 _19260_ (.A(_12283_),
    .X(_12284_));
 sg13g2_nor2_1 _19261_ (.A(net457),
    .B(net643),
    .Y(_12285_));
 sg13g2_buf_1 _19262_ (.A(_12285_),
    .X(_12286_));
 sg13g2_nor2b_1 _19263_ (.A(net367),
    .B_N(\cpu.dcache.r_data[1][24] ),
    .Y(_12287_));
 sg13g2_a21oi_1 _19264_ (.A1(net981),
    .A2(net367),
    .Y(_12288_),
    .B1(_12287_));
 sg13g2_nand2_1 _19265_ (.Y(_12289_),
    .A(net420),
    .B(net56));
 sg13g2_o21ai_1 _19266_ (.B1(_12289_),
    .Y(_00347_),
    .A1(net56),
    .A2(_12288_));
 sg13g2_nor2b_1 _19267_ (.A(net367),
    .B_N(\cpu.dcache.r_data[1][25] ),
    .Y(_12290_));
 sg13g2_a21oi_1 _19268_ (.A1(_12208_),
    .A2(net367),
    .Y(_12291_),
    .B1(_12290_));
 sg13g2_nand2_1 _19269_ (.Y(_12292_),
    .A(_12161_),
    .B(net56));
 sg13g2_o21ai_1 _19270_ (.B1(_12292_),
    .Y(_00348_),
    .A1(_12284_),
    .A2(_12291_));
 sg13g2_nor2b_1 _19271_ (.A(net367),
    .B_N(\cpu.dcache.r_data[1][26] ),
    .Y(_12293_));
 sg13g2_a21oi_1 _19272_ (.A1(net980),
    .A2(net367),
    .Y(_12294_),
    .B1(_12293_));
 sg13g2_nand2_1 _19273_ (.Y(_12295_),
    .A(net421),
    .B(_12283_));
 sg13g2_o21ai_1 _19274_ (.B1(_12295_),
    .Y(_00349_),
    .A1(net56),
    .A2(_12294_));
 sg13g2_nor2b_1 _19275_ (.A(net367),
    .B_N(\cpu.dcache.r_data[1][27] ),
    .Y(_12296_));
 sg13g2_a21oi_1 _19276_ (.A1(net989),
    .A2(net367),
    .Y(_12297_),
    .B1(_12296_));
 sg13g2_nand2_1 _19277_ (.Y(_12298_),
    .A(net419),
    .B(_12283_));
 sg13g2_o21ai_1 _19278_ (.B1(_12298_),
    .Y(_00350_),
    .A1(_12284_),
    .A2(_12297_));
 sg13g2_nor2_1 _19279_ (.A(net457),
    .B(_12166_),
    .Y(_12299_));
 sg13g2_buf_2 _19280_ (.A(_12299_),
    .X(_12300_));
 sg13g2_nor2b_1 _19281_ (.A(_12300_),
    .B_N(\cpu.dcache.r_data[1][28] ),
    .Y(_12301_));
 sg13g2_a21oi_1 _19282_ (.A1(net981),
    .A2(_12300_),
    .Y(_12302_),
    .B1(_12301_));
 sg13g2_nand2_1 _19283_ (.Y(_12303_),
    .A(net368),
    .B(_12283_));
 sg13g2_o21ai_1 _19284_ (.B1(_12303_),
    .Y(_00351_),
    .A1(net56),
    .A2(_12302_));
 sg13g2_nor2b_1 _19285_ (.A(_12300_),
    .B_N(\cpu.dcache.r_data[1][29] ),
    .Y(_12304_));
 sg13g2_a21oi_1 _19286_ (.A1(_12208_),
    .A2(_12300_),
    .Y(_12305_),
    .B1(_12304_));
 sg13g2_nand2_1 _19287_ (.Y(_12306_),
    .A(net418),
    .B(_12283_));
 sg13g2_o21ai_1 _19288_ (.B1(_12306_),
    .Y(_00352_),
    .A1(net56),
    .A2(_12305_));
 sg13g2_mux2_1 _19289_ (.A0(\cpu.dcache.r_data[1][2] ),
    .A1(net1078),
    .S(_12219_),
    .X(_12307_));
 sg13g2_nor2_1 _19290_ (.A(_12216_),
    .B(_12307_),
    .Y(_12308_));
 sg13g2_a21oi_1 _19291_ (.A1(net725),
    .A2(_12217_),
    .Y(_00353_),
    .B1(_12308_));
 sg13g2_nor2b_1 _19292_ (.A(_12300_),
    .B_N(\cpu.dcache.r_data[1][30] ),
    .Y(_12309_));
 sg13g2_a21oi_1 _19293_ (.A1(net980),
    .A2(_12300_),
    .Y(_12310_),
    .B1(_12309_));
 sg13g2_nand2_1 _19294_ (.Y(_12311_),
    .A(net417),
    .B(_12283_));
 sg13g2_o21ai_1 _19295_ (.B1(_12311_),
    .Y(_00354_),
    .A1(net56),
    .A2(_12310_));
 sg13g2_buf_1 _19296_ (.A(net1083),
    .X(_12312_));
 sg13g2_nor2b_1 _19297_ (.A(_12300_),
    .B_N(\cpu.dcache.r_data[1][31] ),
    .Y(_12313_));
 sg13g2_a21oi_1 _19298_ (.A1(net979),
    .A2(_12300_),
    .Y(_12314_),
    .B1(_12313_));
 sg13g2_nand2_1 _19299_ (.Y(_12315_),
    .A(net416),
    .B(_12283_));
 sg13g2_o21ai_1 _19300_ (.B1(_12315_),
    .Y(_00355_),
    .A1(net56),
    .A2(_12314_));
 sg13g2_mux2_1 _19301_ (.A0(\cpu.dcache.r_data[1][3] ),
    .A1(net983),
    .S(_12219_),
    .X(_12316_));
 sg13g2_nor2_1 _19302_ (.A(_12216_),
    .B(_12316_),
    .Y(_12317_));
 sg13g2_a21oi_1 _19303_ (.A1(net724),
    .A2(net59),
    .Y(_00356_),
    .B1(_12317_));
 sg13g2_nor2_1 _19304_ (.A(net457),
    .B(_12190_),
    .Y(_12318_));
 sg13g2_buf_2 _19305_ (.A(_12318_),
    .X(_12319_));
 sg13g2_mux2_1 _19306_ (.A0(\cpu.dcache.r_data[1][4] ),
    .A1(net1079),
    .S(_12319_),
    .X(_12320_));
 sg13g2_nor2_1 _19307_ (.A(_12216_),
    .B(_12320_),
    .Y(_12321_));
 sg13g2_a21oi_1 _19308_ (.A1(net723),
    .A2(net59),
    .Y(_00357_),
    .B1(_12321_));
 sg13g2_nor2b_1 _19309_ (.A(_12319_),
    .B_N(\cpu.dcache.r_data[1][5] ),
    .Y(_12322_));
 sg13g2_a21oi_1 _19310_ (.A1(net982),
    .A2(_12319_),
    .Y(_12323_),
    .B1(_12322_));
 sg13g2_nand2_1 _19311_ (.Y(_12324_),
    .A(net984),
    .B(_12216_));
 sg13g2_o21ai_1 _19312_ (.B1(_12324_),
    .Y(_00358_),
    .A1(_12217_),
    .A2(_12323_));
 sg13g2_nor2b_1 _19313_ (.A(_12319_),
    .B_N(\cpu.dcache.r_data[1][6] ),
    .Y(_12325_));
 sg13g2_a21oi_1 _19314_ (.A1(net980),
    .A2(_12319_),
    .Y(_12326_),
    .B1(_12325_));
 sg13g2_nand2_1 _19315_ (.Y(_12327_),
    .A(net985),
    .B(_12216_));
 sg13g2_o21ai_1 _19316_ (.B1(_12327_),
    .Y(_00359_),
    .A1(net59),
    .A2(_12326_));
 sg13g2_mux2_1 _19317_ (.A0(\cpu.dcache.r_data[1][7] ),
    .A1(net983),
    .S(_12319_),
    .X(_12328_));
 sg13g2_nor2_1 _19318_ (.A(_12216_),
    .B(_12328_),
    .Y(_12329_));
 sg13g2_a21oi_1 _19319_ (.A1(net722),
    .A2(net59),
    .Y(_00360_),
    .B1(_12329_));
 sg13g2_nor2b_1 _19320_ (.A(_12228_),
    .B_N(\cpu.dcache.r_data[1][8] ),
    .Y(_12330_));
 sg13g2_a21oi_1 _19321_ (.A1(net981),
    .A2(_12228_),
    .Y(_12331_),
    .B1(_12330_));
 sg13g2_nand2_1 _19322_ (.Y(_12332_),
    .A(net420),
    .B(_12225_));
 sg13g2_o21ai_1 _19323_ (.B1(_12332_),
    .Y(_00361_),
    .A1(net58),
    .A2(_12331_));
 sg13g2_nor2b_1 _19324_ (.A(_12228_),
    .B_N(\cpu.dcache.r_data[1][9] ),
    .Y(_12333_));
 sg13g2_a21oi_1 _19325_ (.A1(net982),
    .A2(_12228_),
    .Y(_12334_),
    .B1(_12333_));
 sg13g2_nand2_1 _19326_ (.Y(_12335_),
    .A(net369),
    .B(_12225_));
 sg13g2_o21ai_1 _19327_ (.B1(_12335_),
    .Y(_00362_),
    .A1(net58),
    .A2(_12334_));
 sg13g2_nand2_1 _19328_ (.Y(_12336_),
    .A(net644),
    .B(net890));
 sg13g2_buf_1 _19329_ (.A(_12336_),
    .X(_12337_));
 sg13g2_or2_1 _19330_ (.X(_12338_),
    .B(_11999_),
    .A(net518));
 sg13g2_buf_1 _19331_ (.A(_12338_),
    .X(_12339_));
 sg13g2_nor2_1 _19332_ (.A(_11987_),
    .B(_12339_),
    .Y(_12340_));
 sg13g2_buf_1 _19333_ (.A(_12340_),
    .X(_12341_));
 sg13g2_buf_1 _19334_ (.A(_12341_),
    .X(_12342_));
 sg13g2_nor2_1 _19335_ (.A(net518),
    .B(_12016_),
    .Y(_12343_));
 sg13g2_buf_2 _19336_ (.A(_12343_),
    .X(_12344_));
 sg13g2_nor2b_1 _19337_ (.A(_12344_),
    .B_N(\cpu.dcache.r_data[2][0] ),
    .Y(_12345_));
 sg13g2_a21oi_1 _19338_ (.A1(net981),
    .A2(_12344_),
    .Y(_12346_),
    .B1(_12345_));
 sg13g2_nand2_1 _19339_ (.Y(_12347_),
    .A(net851),
    .B(net55));
 sg13g2_o21ai_1 _19340_ (.B1(_12347_),
    .Y(_00363_),
    .A1(net55),
    .A2(_12346_));
 sg13g2_nor2_1 _19341_ (.A(_12025_),
    .B(_12339_),
    .Y(_12348_));
 sg13g2_buf_2 _19342_ (.A(_12348_),
    .X(_12349_));
 sg13g2_buf_1 _19343_ (.A(_12349_),
    .X(_12350_));
 sg13g2_nor2_1 _19344_ (.A(net518),
    .B(_12033_),
    .Y(_12351_));
 sg13g2_buf_2 _19345_ (.A(_12351_),
    .X(_12352_));
 sg13g2_nor2b_1 _19346_ (.A(_12352_),
    .B_N(\cpu.dcache.r_data[2][10] ),
    .Y(_12353_));
 sg13g2_a21oi_1 _19347_ (.A1(_12244_),
    .A2(_12352_),
    .Y(_12354_),
    .B1(_12353_));
 sg13g2_nand2_1 _19348_ (.Y(_12355_),
    .A(net421),
    .B(net54));
 sg13g2_o21ai_1 _19349_ (.B1(_12355_),
    .Y(_00364_),
    .A1(net54),
    .A2(_12354_));
 sg13g2_nor2b_1 _19350_ (.A(_12352_),
    .B_N(\cpu.dcache.r_data[2][11] ),
    .Y(_12356_));
 sg13g2_a21oi_1 _19351_ (.A1(net979),
    .A2(_12352_),
    .Y(_12357_),
    .B1(_12356_));
 sg13g2_nand2_1 _19352_ (.Y(_12358_),
    .A(net419),
    .B(_12350_));
 sg13g2_o21ai_1 _19353_ (.B1(_12358_),
    .Y(_00365_),
    .A1(net54),
    .A2(_12357_));
 sg13g2_nor2_1 _19354_ (.A(net518),
    .B(_12055_),
    .Y(_12359_));
 sg13g2_buf_2 _19355_ (.A(_12359_),
    .X(_12360_));
 sg13g2_nor2b_1 _19356_ (.A(_12360_),
    .B_N(\cpu.dcache.r_data[2][12] ),
    .Y(_12361_));
 sg13g2_a21oi_1 _19357_ (.A1(net981),
    .A2(_12360_),
    .Y(_12362_),
    .B1(_12361_));
 sg13g2_nand2_1 _19358_ (.Y(_12363_),
    .A(net368),
    .B(_12349_));
 sg13g2_o21ai_1 _19359_ (.B1(_12363_),
    .Y(_00366_),
    .A1(net54),
    .A2(_12362_));
 sg13g2_nor2b_1 _19360_ (.A(_12360_),
    .B_N(\cpu.dcache.r_data[2][13] ),
    .Y(_12364_));
 sg13g2_a21oi_1 _19361_ (.A1(net982),
    .A2(_12360_),
    .Y(_12365_),
    .B1(_12364_));
 sg13g2_nand2_1 _19362_ (.Y(_12366_),
    .A(net418),
    .B(_12349_));
 sg13g2_o21ai_1 _19363_ (.B1(_12366_),
    .Y(_00367_),
    .A1(net54),
    .A2(_12365_));
 sg13g2_nor2b_1 _19364_ (.A(_12360_),
    .B_N(\cpu.dcache.r_data[2][14] ),
    .Y(_12367_));
 sg13g2_a21oi_1 _19365_ (.A1(_12244_),
    .A2(_12360_),
    .Y(_12368_),
    .B1(_12367_));
 sg13g2_nand2_1 _19366_ (.Y(_12369_),
    .A(net417),
    .B(_12349_));
 sg13g2_o21ai_1 _19367_ (.B1(_12369_),
    .Y(_00368_),
    .A1(net54),
    .A2(_12368_));
 sg13g2_nor2b_1 _19368_ (.A(_12360_),
    .B_N(\cpu.dcache.r_data[2][15] ),
    .Y(_12370_));
 sg13g2_a21oi_1 _19369_ (.A1(net979),
    .A2(_12360_),
    .Y(_12371_),
    .B1(_12370_));
 sg13g2_nand2_1 _19370_ (.Y(_12372_),
    .A(net416),
    .B(_12349_));
 sg13g2_o21ai_1 _19371_ (.B1(_12372_),
    .Y(_00369_),
    .A1(net54),
    .A2(_12371_));
 sg13g2_nor2_1 _19372_ (.A(_12090_),
    .B(_12339_),
    .Y(_12373_));
 sg13g2_buf_1 _19373_ (.A(_12373_),
    .X(_12374_));
 sg13g2_buf_1 _19374_ (.A(_12374_),
    .X(_12375_));
 sg13g2_nor2_1 _19375_ (.A(net518),
    .B(_12096_),
    .Y(_12376_));
 sg13g2_buf_2 _19376_ (.A(_12376_),
    .X(_12377_));
 sg13g2_nor2b_1 _19377_ (.A(_12377_),
    .B_N(\cpu.dcache.r_data[2][16] ),
    .Y(_12378_));
 sg13g2_a21oi_1 _19378_ (.A1(net981),
    .A2(_12377_),
    .Y(_12379_),
    .B1(_12378_));
 sg13g2_nand2_1 _19379_ (.Y(_12380_),
    .A(net851),
    .B(net53));
 sg13g2_o21ai_1 _19380_ (.B1(_12380_),
    .Y(_00370_),
    .A1(net53),
    .A2(_12379_));
 sg13g2_buf_1 _19381_ (.A(_12066_),
    .X(_12381_));
 sg13g2_nor2b_1 _19382_ (.A(_12377_),
    .B_N(\cpu.dcache.r_data[2][17] ),
    .Y(_12382_));
 sg13g2_a21oi_1 _19383_ (.A1(net978),
    .A2(_12377_),
    .Y(_12383_),
    .B1(_12382_));
 sg13g2_nand2_1 _19384_ (.Y(_12384_),
    .A(net855),
    .B(net53));
 sg13g2_o21ai_1 _19385_ (.B1(_12384_),
    .Y(_00371_),
    .A1(net53),
    .A2(_12383_));
 sg13g2_mux2_1 _19386_ (.A0(\cpu.dcache.r_data[2][18] ),
    .A1(net1078),
    .S(_12377_),
    .X(_12385_));
 sg13g2_nor2_1 _19387_ (.A(_12374_),
    .B(_12385_),
    .Y(_12386_));
 sg13g2_a21oi_1 _19388_ (.A1(net725),
    .A2(_12375_),
    .Y(_00372_),
    .B1(_12386_));
 sg13g2_mux2_1 _19389_ (.A0(\cpu.dcache.r_data[2][19] ),
    .A1(net983),
    .S(_12377_),
    .X(_12387_));
 sg13g2_nor2_1 _19390_ (.A(_12374_),
    .B(_12387_),
    .Y(_12388_));
 sg13g2_a21oi_1 _19391_ (.A1(net724),
    .A2(_12375_),
    .Y(_00373_),
    .B1(_12388_));
 sg13g2_nor2b_1 _19392_ (.A(_12344_),
    .B_N(\cpu.dcache.r_data[2][1] ),
    .Y(_12389_));
 sg13g2_a21oi_1 _19393_ (.A1(net978),
    .A2(_12344_),
    .Y(_12390_),
    .B1(_12389_));
 sg13g2_buf_1 _19394_ (.A(_09871_),
    .X(_12391_));
 sg13g2_nand2_1 _19395_ (.Y(_12392_),
    .A(net850),
    .B(net55));
 sg13g2_o21ai_1 _19396_ (.B1(_12392_),
    .Y(_00374_),
    .A1(net55),
    .A2(_12390_));
 sg13g2_nor2_1 _19397_ (.A(net518),
    .B(_12125_),
    .Y(_12393_));
 sg13g2_buf_2 _19398_ (.A(_12393_),
    .X(_12394_));
 sg13g2_mux2_1 _19399_ (.A0(\cpu.dcache.r_data[2][20] ),
    .A1(net1079),
    .S(_12394_),
    .X(_12395_));
 sg13g2_nor2_1 _19400_ (.A(_12374_),
    .B(_12395_),
    .Y(_12396_));
 sg13g2_a21oi_1 _19401_ (.A1(net723),
    .A2(net53),
    .Y(_00375_),
    .B1(_12396_));
 sg13g2_nor2b_1 _19402_ (.A(_12394_),
    .B_N(\cpu.dcache.r_data[2][21] ),
    .Y(_12397_));
 sg13g2_a21oi_1 _19403_ (.A1(net978),
    .A2(_12394_),
    .Y(_12398_),
    .B1(_12397_));
 sg13g2_nand2_1 _19404_ (.Y(_12399_),
    .A(net984),
    .B(_12374_));
 sg13g2_o21ai_1 _19405_ (.B1(_12399_),
    .Y(_00376_),
    .A1(net53),
    .A2(_12398_));
 sg13g2_nor2b_1 _19406_ (.A(_12394_),
    .B_N(\cpu.dcache.r_data[2][22] ),
    .Y(_12400_));
 sg13g2_a21oi_1 _19407_ (.A1(net980),
    .A2(_12394_),
    .Y(_12401_),
    .B1(_12400_));
 sg13g2_nand2_1 _19408_ (.Y(_12402_),
    .A(net985),
    .B(_12374_));
 sg13g2_o21ai_1 _19409_ (.B1(_12402_),
    .Y(_00377_),
    .A1(net53),
    .A2(_12401_));
 sg13g2_mux2_1 _19410_ (.A0(\cpu.dcache.r_data[2][23] ),
    .A1(net983),
    .S(_12394_),
    .X(_12403_));
 sg13g2_nor2_1 _19411_ (.A(_12374_),
    .B(_12403_),
    .Y(_12404_));
 sg13g2_a21oi_1 _19412_ (.A1(net722),
    .A2(net53),
    .Y(_00378_),
    .B1(_12404_));
 sg13g2_nor2_1 _19413_ (.A(_12153_),
    .B(_12339_),
    .Y(_12405_));
 sg13g2_buf_2 _19414_ (.A(_12405_),
    .X(_12406_));
 sg13g2_buf_1 _19415_ (.A(_12406_),
    .X(_12407_));
 sg13g2_nor2_1 _19416_ (.A(net518),
    .B(net643),
    .Y(_12408_));
 sg13g2_buf_1 _19417_ (.A(_12408_),
    .X(_12409_));
 sg13g2_nor2b_1 _19418_ (.A(net415),
    .B_N(\cpu.dcache.r_data[2][24] ),
    .Y(_12410_));
 sg13g2_a21oi_1 _19419_ (.A1(_12235_),
    .A2(net415),
    .Y(_12411_),
    .B1(_12410_));
 sg13g2_nand2_1 _19420_ (.Y(_12412_),
    .A(net420),
    .B(net52));
 sg13g2_o21ai_1 _19421_ (.B1(_12412_),
    .Y(_00379_),
    .A1(net52),
    .A2(_12411_));
 sg13g2_nor2b_1 _19422_ (.A(net415),
    .B_N(\cpu.dcache.r_data[2][25] ),
    .Y(_12413_));
 sg13g2_a21oi_1 _19423_ (.A1(_12381_),
    .A2(net415),
    .Y(_12414_),
    .B1(_12413_));
 sg13g2_nand2_1 _19424_ (.Y(_12415_),
    .A(net369),
    .B(net52));
 sg13g2_o21ai_1 _19425_ (.B1(_12415_),
    .Y(_00380_),
    .A1(net52),
    .A2(_12414_));
 sg13g2_nor2b_1 _19426_ (.A(net415),
    .B_N(\cpu.dcache.r_data[2][26] ),
    .Y(_12416_));
 sg13g2_a21oi_1 _19427_ (.A1(net980),
    .A2(net415),
    .Y(_12417_),
    .B1(_12416_));
 sg13g2_nand2_1 _19428_ (.Y(_12418_),
    .A(net421),
    .B(_12406_));
 sg13g2_o21ai_1 _19429_ (.B1(_12418_),
    .Y(_00381_),
    .A1(_12407_),
    .A2(_12417_));
 sg13g2_nor2b_1 _19430_ (.A(net415),
    .B_N(\cpu.dcache.r_data[2][27] ),
    .Y(_12419_));
 sg13g2_a21oi_1 _19431_ (.A1(_12312_),
    .A2(net415),
    .Y(_12420_),
    .B1(_12419_));
 sg13g2_nand2_1 _19432_ (.Y(_12421_),
    .A(net419),
    .B(_12406_));
 sg13g2_o21ai_1 _19433_ (.B1(_12421_),
    .Y(_00382_),
    .A1(_12407_),
    .A2(_12420_));
 sg13g2_nor2_1 _19434_ (.A(_12337_),
    .B(_12166_),
    .Y(_12422_));
 sg13g2_buf_2 _19435_ (.A(_12422_),
    .X(_12423_));
 sg13g2_nor2b_1 _19436_ (.A(_12423_),
    .B_N(\cpu.dcache.r_data[2][28] ),
    .Y(_12424_));
 sg13g2_a21oi_1 _19437_ (.A1(_12235_),
    .A2(_12423_),
    .Y(_12425_),
    .B1(_12424_));
 sg13g2_nand2_1 _19438_ (.Y(_12426_),
    .A(net368),
    .B(_12406_));
 sg13g2_o21ai_1 _19439_ (.B1(_12426_),
    .Y(_00383_),
    .A1(net52),
    .A2(_12425_));
 sg13g2_nor2b_1 _19440_ (.A(_12423_),
    .B_N(\cpu.dcache.r_data[2][29] ),
    .Y(_12427_));
 sg13g2_a21oi_1 _19441_ (.A1(_12381_),
    .A2(_12423_),
    .Y(_12428_),
    .B1(_12427_));
 sg13g2_nand2_1 _19442_ (.Y(_12429_),
    .A(net418),
    .B(_12406_));
 sg13g2_o21ai_1 _19443_ (.B1(_12429_),
    .Y(_00384_),
    .A1(net52),
    .A2(_12428_));
 sg13g2_mux2_1 _19444_ (.A0(\cpu.dcache.r_data[2][2] ),
    .A1(net1078),
    .S(_12344_),
    .X(_12430_));
 sg13g2_nor2_1 _19445_ (.A(_12341_),
    .B(_12430_),
    .Y(_12431_));
 sg13g2_a21oi_1 _19446_ (.A1(net725),
    .A2(net55),
    .Y(_00385_),
    .B1(_12431_));
 sg13g2_nor2b_1 _19447_ (.A(_12423_),
    .B_N(\cpu.dcache.r_data[2][30] ),
    .Y(_12432_));
 sg13g2_a21oi_1 _19448_ (.A1(net980),
    .A2(_12423_),
    .Y(_12433_),
    .B1(_12432_));
 sg13g2_nand2_1 _19449_ (.Y(_12434_),
    .A(_12181_),
    .B(_12406_));
 sg13g2_o21ai_1 _19450_ (.B1(_12434_),
    .Y(_00386_),
    .A1(net52),
    .A2(_12433_));
 sg13g2_nor2b_1 _19451_ (.A(_12423_),
    .B_N(\cpu.dcache.r_data[2][31] ),
    .Y(_12435_));
 sg13g2_a21oi_1 _19452_ (.A1(_12312_),
    .A2(_12423_),
    .Y(_12436_),
    .B1(_12435_));
 sg13g2_nand2_1 _19453_ (.Y(_12437_),
    .A(net416),
    .B(_12406_));
 sg13g2_o21ai_1 _19454_ (.B1(_12437_),
    .Y(_00387_),
    .A1(net52),
    .A2(_12436_));
 sg13g2_mux2_1 _19455_ (.A0(\cpu.dcache.r_data[2][3] ),
    .A1(net983),
    .S(_12344_),
    .X(_12438_));
 sg13g2_nor2_1 _19456_ (.A(_12341_),
    .B(_12438_),
    .Y(_12439_));
 sg13g2_a21oi_1 _19457_ (.A1(net724),
    .A2(net55),
    .Y(_00388_),
    .B1(_12439_));
 sg13g2_nor2_1 _19458_ (.A(net518),
    .B(_12190_),
    .Y(_12440_));
 sg13g2_buf_2 _19459_ (.A(_12440_),
    .X(_12441_));
 sg13g2_mux2_1 _19460_ (.A0(\cpu.dcache.r_data[2][4] ),
    .A1(net1079),
    .S(_12441_),
    .X(_12442_));
 sg13g2_nor2_1 _19461_ (.A(_12341_),
    .B(_12442_),
    .Y(_12443_));
 sg13g2_a21oi_1 _19462_ (.A1(net723),
    .A2(_12342_),
    .Y(_00389_),
    .B1(_12443_));
 sg13g2_nor2b_1 _19463_ (.A(_12441_),
    .B_N(\cpu.dcache.r_data[2][5] ),
    .Y(_12444_));
 sg13g2_a21oi_1 _19464_ (.A1(net978),
    .A2(_12441_),
    .Y(_12445_),
    .B1(_12444_));
 sg13g2_nand2_1 _19465_ (.Y(_12446_),
    .A(net984),
    .B(_12341_));
 sg13g2_o21ai_1 _19466_ (.B1(_12446_),
    .Y(_00390_),
    .A1(_12342_),
    .A2(_12445_));
 sg13g2_buf_1 _19467_ (.A(net1084),
    .X(_12447_));
 sg13g2_nor2b_1 _19468_ (.A(_12441_),
    .B_N(\cpu.dcache.r_data[2][6] ),
    .Y(_12448_));
 sg13g2_a21oi_1 _19469_ (.A1(net977),
    .A2(_12441_),
    .Y(_12449_),
    .B1(_12448_));
 sg13g2_nand2_1 _19470_ (.Y(_12450_),
    .A(net985),
    .B(_12341_));
 sg13g2_o21ai_1 _19471_ (.B1(_12450_),
    .Y(_00391_),
    .A1(net55),
    .A2(_12449_));
 sg13g2_mux2_1 _19472_ (.A0(\cpu.dcache.r_data[2][7] ),
    .A1(net983),
    .S(_12441_),
    .X(_12451_));
 sg13g2_nor2_1 _19473_ (.A(_12341_),
    .B(_12451_),
    .Y(_12452_));
 sg13g2_a21oi_1 _19474_ (.A1(net722),
    .A2(net55),
    .Y(_00392_),
    .B1(_12452_));
 sg13g2_buf_1 _19475_ (.A(net1087),
    .X(_12453_));
 sg13g2_nor2b_1 _19476_ (.A(_12352_),
    .B_N(\cpu.dcache.r_data[2][8] ),
    .Y(_12454_));
 sg13g2_a21oi_1 _19477_ (.A1(net976),
    .A2(_12352_),
    .Y(_12455_),
    .B1(_12454_));
 sg13g2_nand2_1 _19478_ (.Y(_12456_),
    .A(net420),
    .B(_12349_));
 sg13g2_o21ai_1 _19479_ (.B1(_12456_),
    .Y(_00393_),
    .A1(_12350_),
    .A2(_12455_));
 sg13g2_nor2b_1 _19480_ (.A(_12352_),
    .B_N(\cpu.dcache.r_data[2][9] ),
    .Y(_12457_));
 sg13g2_a21oi_1 _19481_ (.A1(net978),
    .A2(_12352_),
    .Y(_12458_),
    .B1(_12457_));
 sg13g2_nand2_1 _19482_ (.Y(_12459_),
    .A(net369),
    .B(_12349_));
 sg13g2_o21ai_1 _19483_ (.B1(_12459_),
    .Y(_00394_),
    .A1(net54),
    .A2(_12458_));
 sg13g2_buf_1 _19484_ (.A(net609),
    .X(_12460_));
 sg13g2_buf_1 _19485_ (.A(net517),
    .X(_12461_));
 sg13g2_nand2_1 _19486_ (.Y(_12462_),
    .A(net456),
    .B(net890));
 sg13g2_buf_1 _19487_ (.A(_12462_),
    .X(_12463_));
 sg13g2_or2_1 _19488_ (.X(_12464_),
    .B(_11999_),
    .A(net366));
 sg13g2_buf_1 _19489_ (.A(_12464_),
    .X(_12465_));
 sg13g2_nor2_1 _19490_ (.A(_11987_),
    .B(_12465_),
    .Y(_12466_));
 sg13g2_buf_1 _19491_ (.A(_12466_),
    .X(_12467_));
 sg13g2_buf_1 _19492_ (.A(_12467_),
    .X(_12468_));
 sg13g2_nor2_1 _19493_ (.A(net366),
    .B(_12016_),
    .Y(_12469_));
 sg13g2_buf_2 _19494_ (.A(_12469_),
    .X(_12470_));
 sg13g2_nor2b_1 _19495_ (.A(_12470_),
    .B_N(\cpu.dcache.r_data[3][0] ),
    .Y(_12471_));
 sg13g2_a21oi_1 _19496_ (.A1(net976),
    .A2(_12470_),
    .Y(_12472_),
    .B1(_12471_));
 sg13g2_nand2_1 _19497_ (.Y(_12473_),
    .A(net851),
    .B(net51));
 sg13g2_o21ai_1 _19498_ (.B1(_12473_),
    .Y(_00395_),
    .A1(_12468_),
    .A2(_12472_));
 sg13g2_nor2_1 _19499_ (.A(_12025_),
    .B(_12465_),
    .Y(_12474_));
 sg13g2_buf_2 _19500_ (.A(_12474_),
    .X(_12475_));
 sg13g2_buf_1 _19501_ (.A(_12475_),
    .X(_12476_));
 sg13g2_nor2_1 _19502_ (.A(net366),
    .B(_12033_),
    .Y(_12477_));
 sg13g2_buf_2 _19503_ (.A(_12477_),
    .X(_12478_));
 sg13g2_nor2b_1 _19504_ (.A(_12478_),
    .B_N(\cpu.dcache.r_data[3][10] ),
    .Y(_12479_));
 sg13g2_a21oi_1 _19505_ (.A1(net977),
    .A2(_12478_),
    .Y(_12480_),
    .B1(_12479_));
 sg13g2_nand2_1 _19506_ (.Y(_12481_),
    .A(net421),
    .B(net50));
 sg13g2_o21ai_1 _19507_ (.B1(_12481_),
    .Y(_00396_),
    .A1(_12476_),
    .A2(_12480_));
 sg13g2_nor2b_1 _19508_ (.A(_12478_),
    .B_N(\cpu.dcache.r_data[3][11] ),
    .Y(_12482_));
 sg13g2_a21oi_1 _19509_ (.A1(net979),
    .A2(_12478_),
    .Y(_12483_),
    .B1(_12482_));
 sg13g2_nand2_1 _19510_ (.Y(_12484_),
    .A(net419),
    .B(net50));
 sg13g2_o21ai_1 _19511_ (.B1(_12484_),
    .Y(_00397_),
    .A1(net50),
    .A2(_12483_));
 sg13g2_nor2_1 _19512_ (.A(net366),
    .B(_12055_),
    .Y(_12485_));
 sg13g2_buf_2 _19513_ (.A(_12485_),
    .X(_12486_));
 sg13g2_nor2b_1 _19514_ (.A(_12486_),
    .B_N(\cpu.dcache.r_data[3][12] ),
    .Y(_12487_));
 sg13g2_a21oi_1 _19515_ (.A1(net976),
    .A2(_12486_),
    .Y(_12488_),
    .B1(_12487_));
 sg13g2_nand2_1 _19516_ (.Y(_12489_),
    .A(net368),
    .B(_12475_));
 sg13g2_o21ai_1 _19517_ (.B1(_12489_),
    .Y(_00398_),
    .A1(net50),
    .A2(_12488_));
 sg13g2_nor2b_1 _19518_ (.A(_12486_),
    .B_N(\cpu.dcache.r_data[3][13] ),
    .Y(_12490_));
 sg13g2_a21oi_1 _19519_ (.A1(net978),
    .A2(_12486_),
    .Y(_12491_),
    .B1(_12490_));
 sg13g2_nand2_1 _19520_ (.Y(_12492_),
    .A(net418),
    .B(_12475_));
 sg13g2_o21ai_1 _19521_ (.B1(_12492_),
    .Y(_00399_),
    .A1(net50),
    .A2(_12491_));
 sg13g2_nor2b_1 _19522_ (.A(_12486_),
    .B_N(\cpu.dcache.r_data[3][14] ),
    .Y(_12493_));
 sg13g2_a21oi_1 _19523_ (.A1(net977),
    .A2(_12486_),
    .Y(_12494_),
    .B1(_12493_));
 sg13g2_nand2_1 _19524_ (.Y(_12495_),
    .A(net417),
    .B(_12475_));
 sg13g2_o21ai_1 _19525_ (.B1(_12495_),
    .Y(_00400_),
    .A1(net50),
    .A2(_12494_));
 sg13g2_nor2b_1 _19526_ (.A(_12486_),
    .B_N(\cpu.dcache.r_data[3][15] ),
    .Y(_12496_));
 sg13g2_a21oi_1 _19527_ (.A1(net979),
    .A2(_12486_),
    .Y(_12497_),
    .B1(_12496_));
 sg13g2_nand2_1 _19528_ (.Y(_12498_),
    .A(net416),
    .B(_12475_));
 sg13g2_o21ai_1 _19529_ (.B1(_12498_),
    .Y(_00401_),
    .A1(net50),
    .A2(_12497_));
 sg13g2_nor2_1 _19530_ (.A(_12090_),
    .B(_12465_),
    .Y(_12499_));
 sg13g2_buf_1 _19531_ (.A(_12499_),
    .X(_12500_));
 sg13g2_buf_1 _19532_ (.A(_12500_),
    .X(_12501_));
 sg13g2_nor2_1 _19533_ (.A(net366),
    .B(_12096_),
    .Y(_12502_));
 sg13g2_buf_2 _19534_ (.A(_12502_),
    .X(_12503_));
 sg13g2_nor2b_1 _19535_ (.A(_12503_),
    .B_N(\cpu.dcache.r_data[3][16] ),
    .Y(_12504_));
 sg13g2_a21oi_1 _19536_ (.A1(net976),
    .A2(_12503_),
    .Y(_12505_),
    .B1(_12504_));
 sg13g2_nand2_1 _19537_ (.Y(_12506_),
    .A(net851),
    .B(net49));
 sg13g2_o21ai_1 _19538_ (.B1(_12506_),
    .Y(_00402_),
    .A1(net49),
    .A2(_12505_));
 sg13g2_nor2b_1 _19539_ (.A(_12503_),
    .B_N(\cpu.dcache.r_data[3][17] ),
    .Y(_12507_));
 sg13g2_a21oi_1 _19540_ (.A1(net978),
    .A2(_12503_),
    .Y(_12508_),
    .B1(_12507_));
 sg13g2_nand2_1 _19541_ (.Y(_12509_),
    .A(net850),
    .B(net49));
 sg13g2_o21ai_1 _19542_ (.B1(_12509_),
    .Y(_00403_),
    .A1(net49),
    .A2(_12508_));
 sg13g2_mux2_1 _19543_ (.A0(\cpu.dcache.r_data[3][18] ),
    .A1(net1078),
    .S(_12503_),
    .X(_12510_));
 sg13g2_nor2_1 _19544_ (.A(_12500_),
    .B(_12510_),
    .Y(_12511_));
 sg13g2_a21oi_1 _19545_ (.A1(net725),
    .A2(_12501_),
    .Y(_00404_),
    .B1(_12511_));
 sg13g2_mux2_1 _19546_ (.A0(\cpu.dcache.r_data[3][19] ),
    .A1(_12202_),
    .S(_12503_),
    .X(_12512_));
 sg13g2_nor2_1 _19547_ (.A(_12500_),
    .B(_12512_),
    .Y(_12513_));
 sg13g2_a21oi_1 _19548_ (.A1(net724),
    .A2(_12501_),
    .Y(_00405_),
    .B1(_12513_));
 sg13g2_nor2b_1 _19549_ (.A(_12470_),
    .B_N(\cpu.dcache.r_data[3][1] ),
    .Y(_12514_));
 sg13g2_a21oi_1 _19550_ (.A1(net978),
    .A2(_12470_),
    .Y(_12515_),
    .B1(_12514_));
 sg13g2_nand2_1 _19551_ (.Y(_12516_),
    .A(net850),
    .B(net51));
 sg13g2_o21ai_1 _19552_ (.B1(_12516_),
    .Y(_00406_),
    .A1(net51),
    .A2(_12515_));
 sg13g2_or2_1 _19553_ (.X(_12517_),
    .B(_12125_),
    .A(net366));
 sg13g2_buf_1 _19554_ (.A(_12517_),
    .X(_12518_));
 sg13g2_mux2_1 _19555_ (.A0(net1079),
    .A1(\cpu.dcache.r_data[3][20] ),
    .S(_12518_),
    .X(_12519_));
 sg13g2_nor2_1 _19556_ (.A(_12500_),
    .B(_12519_),
    .Y(_12520_));
 sg13g2_a21oi_1 _19557_ (.A1(net723),
    .A2(net49),
    .Y(_00407_),
    .B1(_12520_));
 sg13g2_mux2_1 _19558_ (.A0(net1082),
    .A1(\cpu.dcache.r_data[3][21] ),
    .S(_12518_),
    .X(_12521_));
 sg13g2_buf_1 _19559_ (.A(net1021),
    .X(_12522_));
 sg13g2_mux2_1 _19560_ (.A0(_12521_),
    .A1(net849),
    .S(net49),
    .X(_00408_));
 sg13g2_mux2_1 _19561_ (.A0(net1081),
    .A1(\cpu.dcache.r_data[3][22] ),
    .S(_12518_),
    .X(_12523_));
 sg13g2_mux2_1 _19562_ (.A0(_12523_),
    .A1(net875),
    .S(net49),
    .X(_00409_));
 sg13g2_mux2_1 _19563_ (.A0(net1080),
    .A1(\cpu.dcache.r_data[3][23] ),
    .S(_12518_),
    .X(_12524_));
 sg13g2_nor2_1 _19564_ (.A(_12500_),
    .B(_12524_),
    .Y(_12525_));
 sg13g2_a21oi_1 _19565_ (.A1(net722),
    .A2(net49),
    .Y(_00410_),
    .B1(_12525_));
 sg13g2_nor2_1 _19566_ (.A(_12153_),
    .B(_12465_),
    .Y(_12526_));
 sg13g2_buf_2 _19567_ (.A(_12526_),
    .X(_12527_));
 sg13g2_buf_1 _19568_ (.A(_12527_),
    .X(_12528_));
 sg13g2_nor2_1 _19569_ (.A(_12463_),
    .B(net643),
    .Y(_12529_));
 sg13g2_buf_1 _19570_ (.A(_12529_),
    .X(_12530_));
 sg13g2_nor2b_1 _19571_ (.A(net240),
    .B_N(\cpu.dcache.r_data[3][24] ),
    .Y(_12531_));
 sg13g2_a21oi_1 _19572_ (.A1(net976),
    .A2(net240),
    .Y(_12532_),
    .B1(_12531_));
 sg13g2_nand2_1 _19573_ (.Y(_12533_),
    .A(net420),
    .B(net48));
 sg13g2_o21ai_1 _19574_ (.B1(_12533_),
    .Y(_00411_),
    .A1(net48),
    .A2(_12532_));
 sg13g2_buf_1 _19575_ (.A(net1082),
    .X(_12534_));
 sg13g2_nor2b_1 _19576_ (.A(net240),
    .B_N(\cpu.dcache.r_data[3][25] ),
    .Y(_12535_));
 sg13g2_a21oi_1 _19577_ (.A1(net975),
    .A2(net240),
    .Y(_12536_),
    .B1(_12535_));
 sg13g2_nand2_1 _19578_ (.Y(_12537_),
    .A(net369),
    .B(net48));
 sg13g2_o21ai_1 _19579_ (.B1(_12537_),
    .Y(_00412_),
    .A1(net48),
    .A2(_12536_));
 sg13g2_nor2b_1 _19580_ (.A(net240),
    .B_N(\cpu.dcache.r_data[3][26] ),
    .Y(_12538_));
 sg13g2_a21oi_1 _19581_ (.A1(net977),
    .A2(net240),
    .Y(_12539_),
    .B1(_12538_));
 sg13g2_nand2_1 _19582_ (.Y(_12540_),
    .A(net421),
    .B(_12527_));
 sg13g2_o21ai_1 _19583_ (.B1(_12540_),
    .Y(_00413_),
    .A1(_12528_),
    .A2(_12539_));
 sg13g2_nor2b_1 _19584_ (.A(net240),
    .B_N(\cpu.dcache.r_data[3][27] ),
    .Y(_12541_));
 sg13g2_a21oi_1 _19585_ (.A1(net979),
    .A2(net240),
    .Y(_12542_),
    .B1(_12541_));
 sg13g2_nand2_1 _19586_ (.Y(_12543_),
    .A(net419),
    .B(_12527_));
 sg13g2_o21ai_1 _19587_ (.B1(_12543_),
    .Y(_00414_),
    .A1(_12528_),
    .A2(_12542_));
 sg13g2_nor2_1 _19588_ (.A(net366),
    .B(_12166_),
    .Y(_12544_));
 sg13g2_buf_2 _19589_ (.A(_12544_),
    .X(_12545_));
 sg13g2_nor2b_1 _19590_ (.A(_12545_),
    .B_N(\cpu.dcache.r_data[3][28] ),
    .Y(_12546_));
 sg13g2_a21oi_1 _19591_ (.A1(net976),
    .A2(_12545_),
    .Y(_12547_),
    .B1(_12546_));
 sg13g2_nand2_1 _19592_ (.Y(_12548_),
    .A(_12171_),
    .B(_12527_));
 sg13g2_o21ai_1 _19593_ (.B1(_12548_),
    .Y(_00415_),
    .A1(net48),
    .A2(_12547_));
 sg13g2_nor2b_1 _19594_ (.A(_12545_),
    .B_N(\cpu.dcache.r_data[3][29] ),
    .Y(_12549_));
 sg13g2_a21oi_1 _19595_ (.A1(net975),
    .A2(_12545_),
    .Y(_12550_),
    .B1(_12549_));
 sg13g2_nand2_1 _19596_ (.Y(_12551_),
    .A(_12175_),
    .B(_12527_));
 sg13g2_o21ai_1 _19597_ (.B1(_12551_),
    .Y(_00416_),
    .A1(net48),
    .A2(_12550_));
 sg13g2_mux2_1 _19598_ (.A0(\cpu.dcache.r_data[3][2] ),
    .A1(net1078),
    .S(_12470_),
    .X(_12552_));
 sg13g2_nor2_1 _19599_ (.A(_12467_),
    .B(_12552_),
    .Y(_12553_));
 sg13g2_a21oi_1 _19600_ (.A1(net725),
    .A2(_12468_),
    .Y(_00417_),
    .B1(_12553_));
 sg13g2_nor2b_1 _19601_ (.A(_12545_),
    .B_N(\cpu.dcache.r_data[3][30] ),
    .Y(_12554_));
 sg13g2_a21oi_1 _19602_ (.A1(_12447_),
    .A2(_12545_),
    .Y(_12555_),
    .B1(_12554_));
 sg13g2_nand2_1 _19603_ (.Y(_12556_),
    .A(_12181_),
    .B(_12527_));
 sg13g2_o21ai_1 _19604_ (.B1(_12556_),
    .Y(_00418_),
    .A1(net48),
    .A2(_12555_));
 sg13g2_nor2b_1 _19605_ (.A(_12545_),
    .B_N(\cpu.dcache.r_data[3][31] ),
    .Y(_12557_));
 sg13g2_a21oi_1 _19606_ (.A1(net979),
    .A2(_12545_),
    .Y(_12558_),
    .B1(_12557_));
 sg13g2_nand2_1 _19607_ (.Y(_12559_),
    .A(net416),
    .B(_12527_));
 sg13g2_o21ai_1 _19608_ (.B1(_12559_),
    .Y(_00419_),
    .A1(net48),
    .A2(_12558_));
 sg13g2_buf_1 _19609_ (.A(_12045_),
    .X(_12560_));
 sg13g2_mux2_1 _19610_ (.A0(\cpu.dcache.r_data[3][3] ),
    .A1(net1077),
    .S(_12470_),
    .X(_12561_));
 sg13g2_nor2_1 _19611_ (.A(_12467_),
    .B(_12561_),
    .Y(_12562_));
 sg13g2_a21oi_1 _19612_ (.A1(net724),
    .A2(net51),
    .Y(_00420_),
    .B1(_12562_));
 sg13g2_or2_1 _19613_ (.X(_12563_),
    .B(_12190_),
    .A(net366));
 sg13g2_buf_1 _19614_ (.A(_12563_),
    .X(_12564_));
 sg13g2_mux2_1 _19615_ (.A0(net1079),
    .A1(\cpu.dcache.r_data[3][4] ),
    .S(_12564_),
    .X(_12565_));
 sg13g2_nor2_1 _19616_ (.A(_12467_),
    .B(_12565_),
    .Y(_12566_));
 sg13g2_a21oi_1 _19617_ (.A1(net723),
    .A2(net51),
    .Y(_00421_),
    .B1(_12566_));
 sg13g2_mux2_1 _19618_ (.A0(net1082),
    .A1(\cpu.dcache.r_data[3][5] ),
    .S(_12564_),
    .X(_12567_));
 sg13g2_mux2_1 _19619_ (.A0(_12567_),
    .A1(net849),
    .S(net51),
    .X(_00422_));
 sg13g2_mux2_1 _19620_ (.A0(net1081),
    .A1(\cpu.dcache.r_data[3][6] ),
    .S(_12564_),
    .X(_12568_));
 sg13g2_buf_1 _19621_ (.A(_09907_),
    .X(_12569_));
 sg13g2_mux2_1 _19622_ (.A0(_12568_),
    .A1(net974),
    .S(net51),
    .X(_00423_));
 sg13g2_mux2_1 _19623_ (.A0(net1080),
    .A1(\cpu.dcache.r_data[3][7] ),
    .S(_12564_),
    .X(_12570_));
 sg13g2_nor2_1 _19624_ (.A(_12467_),
    .B(_12570_),
    .Y(_12571_));
 sg13g2_a21oi_1 _19625_ (.A1(net722),
    .A2(net51),
    .Y(_00424_),
    .B1(_12571_));
 sg13g2_nor2b_1 _19626_ (.A(_12478_),
    .B_N(\cpu.dcache.r_data[3][8] ),
    .Y(_12572_));
 sg13g2_a21oi_1 _19627_ (.A1(_12453_),
    .A2(_12478_),
    .Y(_12573_),
    .B1(_12572_));
 sg13g2_nand2_1 _19628_ (.Y(_12574_),
    .A(net420),
    .B(_12475_));
 sg13g2_o21ai_1 _19629_ (.B1(_12574_),
    .Y(_00425_),
    .A1(_12476_),
    .A2(_12573_));
 sg13g2_nor2b_1 _19630_ (.A(_12478_),
    .B_N(\cpu.dcache.r_data[3][9] ),
    .Y(_12575_));
 sg13g2_a21oi_1 _19631_ (.A1(net975),
    .A2(_12478_),
    .Y(_12576_),
    .B1(_12575_));
 sg13g2_nand2_1 _19632_ (.Y(_12577_),
    .A(net369),
    .B(_12475_));
 sg13g2_o21ai_1 _19633_ (.B1(_12577_),
    .Y(_00426_),
    .A1(net50),
    .A2(_12576_));
 sg13g2_buf_1 _19634_ (.A(_09920_),
    .X(_12578_));
 sg13g2_or2_1 _19635_ (.X(_12579_),
    .B(_11999_),
    .A(net583));
 sg13g2_buf_1 _19636_ (.A(_12579_),
    .X(_12580_));
 sg13g2_nor2_1 _19637_ (.A(_11987_),
    .B(_12580_),
    .Y(_12581_));
 sg13g2_buf_1 _19638_ (.A(_12581_),
    .X(_12582_));
 sg13g2_buf_1 _19639_ (.A(_12582_),
    .X(_12583_));
 sg13g2_nor2_1 _19640_ (.A(net583),
    .B(_12016_),
    .Y(_12584_));
 sg13g2_buf_2 _19641_ (.A(_12584_),
    .X(_12585_));
 sg13g2_nor2b_1 _19642_ (.A(_12585_),
    .B_N(\cpu.dcache.r_data[4][0] ),
    .Y(_12586_));
 sg13g2_a21oi_1 _19643_ (.A1(net976),
    .A2(_12585_),
    .Y(_12587_),
    .B1(_12586_));
 sg13g2_nand2_1 _19644_ (.Y(_12588_),
    .A(net851),
    .B(net47));
 sg13g2_o21ai_1 _19645_ (.B1(_12588_),
    .Y(_00427_),
    .A1(net47),
    .A2(_12587_));
 sg13g2_nor2_1 _19646_ (.A(_12025_),
    .B(_12580_),
    .Y(_12589_));
 sg13g2_buf_2 _19647_ (.A(_12589_),
    .X(_12590_));
 sg13g2_buf_1 _19648_ (.A(_12590_),
    .X(_12591_));
 sg13g2_nor2_1 _19649_ (.A(net583),
    .B(_12033_),
    .Y(_12592_));
 sg13g2_buf_2 _19650_ (.A(_12592_),
    .X(_12593_));
 sg13g2_nor2b_1 _19651_ (.A(_12593_),
    .B_N(\cpu.dcache.r_data[4][10] ),
    .Y(_12594_));
 sg13g2_a21oi_1 _19652_ (.A1(net977),
    .A2(_12593_),
    .Y(_12595_),
    .B1(_12594_));
 sg13g2_nand2_1 _19653_ (.Y(_12596_),
    .A(net421),
    .B(net46));
 sg13g2_o21ai_1 _19654_ (.B1(_12596_),
    .Y(_00428_),
    .A1(net46),
    .A2(_12595_));
 sg13g2_nor2b_1 _19655_ (.A(_12593_),
    .B_N(\cpu.dcache.r_data[4][11] ),
    .Y(_12597_));
 sg13g2_a21oi_1 _19656_ (.A1(net979),
    .A2(_12593_),
    .Y(_12598_),
    .B1(_12597_));
 sg13g2_nand2_1 _19657_ (.Y(_12599_),
    .A(net419),
    .B(_12591_));
 sg13g2_o21ai_1 _19658_ (.B1(_12599_),
    .Y(_00429_),
    .A1(net46),
    .A2(_12598_));
 sg13g2_nor2_1 _19659_ (.A(net583),
    .B(_12055_),
    .Y(_12600_));
 sg13g2_buf_2 _19660_ (.A(_12600_),
    .X(_12601_));
 sg13g2_nor2b_1 _19661_ (.A(_12601_),
    .B_N(\cpu.dcache.r_data[4][12] ),
    .Y(_12602_));
 sg13g2_a21oi_1 _19662_ (.A1(_12453_),
    .A2(_12601_),
    .Y(_12603_),
    .B1(_12602_));
 sg13g2_nand2_1 _19663_ (.Y(_12604_),
    .A(net368),
    .B(_12590_));
 sg13g2_o21ai_1 _19664_ (.B1(_12604_),
    .Y(_00430_),
    .A1(net46),
    .A2(_12603_));
 sg13g2_nor2b_1 _19665_ (.A(_12601_),
    .B_N(\cpu.dcache.r_data[4][13] ),
    .Y(_12605_));
 sg13g2_a21oi_1 _19666_ (.A1(_12534_),
    .A2(_12601_),
    .Y(_12606_),
    .B1(_12605_));
 sg13g2_nand2_1 _19667_ (.Y(_12607_),
    .A(net418),
    .B(_12590_));
 sg13g2_o21ai_1 _19668_ (.B1(_12607_),
    .Y(_00431_),
    .A1(net46),
    .A2(_12606_));
 sg13g2_nor2b_1 _19669_ (.A(_12601_),
    .B_N(\cpu.dcache.r_data[4][14] ),
    .Y(_12608_));
 sg13g2_a21oi_1 _19670_ (.A1(net977),
    .A2(_12601_),
    .Y(_12609_),
    .B1(_12608_));
 sg13g2_nand2_1 _19671_ (.Y(_12610_),
    .A(net417),
    .B(_12590_));
 sg13g2_o21ai_1 _19672_ (.B1(_12610_),
    .Y(_00432_),
    .A1(net46),
    .A2(_12609_));
 sg13g2_buf_1 _19673_ (.A(net1083),
    .X(_12611_));
 sg13g2_nor2b_1 _19674_ (.A(_12601_),
    .B_N(\cpu.dcache.r_data[4][15] ),
    .Y(_12612_));
 sg13g2_a21oi_1 _19675_ (.A1(net973),
    .A2(_12601_),
    .Y(_12613_),
    .B1(_12612_));
 sg13g2_nand2_1 _19676_ (.Y(_12614_),
    .A(net416),
    .B(_12590_));
 sg13g2_o21ai_1 _19677_ (.B1(_12614_),
    .Y(_00433_),
    .A1(net46),
    .A2(_12613_));
 sg13g2_nor2_1 _19678_ (.A(_12090_),
    .B(_12580_),
    .Y(_12615_));
 sg13g2_buf_1 _19679_ (.A(_12615_),
    .X(_12616_));
 sg13g2_buf_1 _19680_ (.A(_12616_),
    .X(_12617_));
 sg13g2_nor2_1 _19681_ (.A(net583),
    .B(_12096_),
    .Y(_12618_));
 sg13g2_buf_2 _19682_ (.A(_12618_),
    .X(_12619_));
 sg13g2_nor2b_1 _19683_ (.A(_12619_),
    .B_N(\cpu.dcache.r_data[4][16] ),
    .Y(_12620_));
 sg13g2_a21oi_1 _19684_ (.A1(net976),
    .A2(_12619_),
    .Y(_12621_),
    .B1(_12620_));
 sg13g2_nand2_1 _19685_ (.Y(_12622_),
    .A(net851),
    .B(net45));
 sg13g2_o21ai_1 _19686_ (.B1(_12622_),
    .Y(_00434_),
    .A1(net45),
    .A2(_12621_));
 sg13g2_nor2b_1 _19687_ (.A(_12619_),
    .B_N(\cpu.dcache.r_data[4][17] ),
    .Y(_12623_));
 sg13g2_a21oi_1 _19688_ (.A1(net975),
    .A2(_12619_),
    .Y(_12624_),
    .B1(_12623_));
 sg13g2_nand2_1 _19689_ (.Y(_12625_),
    .A(net850),
    .B(net45));
 sg13g2_o21ai_1 _19690_ (.B1(_12625_),
    .Y(_00435_),
    .A1(net45),
    .A2(_12624_));
 sg13g2_mux2_1 _19691_ (.A0(\cpu.dcache.r_data[4][18] ),
    .A1(net1078),
    .S(_12619_),
    .X(_12626_));
 sg13g2_nor2_1 _19692_ (.A(_12616_),
    .B(_12626_),
    .Y(_12627_));
 sg13g2_a21oi_1 _19693_ (.A1(net725),
    .A2(net45),
    .Y(_00436_),
    .B1(_12627_));
 sg13g2_mux2_1 _19694_ (.A0(\cpu.dcache.r_data[4][19] ),
    .A1(net1077),
    .S(_12619_),
    .X(_12628_));
 sg13g2_nor2_1 _19695_ (.A(_12616_),
    .B(_12628_),
    .Y(_12629_));
 sg13g2_a21oi_1 _19696_ (.A1(net724),
    .A2(net45),
    .Y(_00437_),
    .B1(_12629_));
 sg13g2_nor2b_1 _19697_ (.A(_12585_),
    .B_N(\cpu.dcache.r_data[4][1] ),
    .Y(_12630_));
 sg13g2_a21oi_1 _19698_ (.A1(net975),
    .A2(_12585_),
    .Y(_12631_),
    .B1(_12630_));
 sg13g2_nand2_1 _19699_ (.Y(_12632_),
    .A(net850),
    .B(net47));
 sg13g2_o21ai_1 _19700_ (.B1(_12632_),
    .Y(_00438_),
    .A1(net47),
    .A2(_12631_));
 sg13g2_nor2_1 _19701_ (.A(net583),
    .B(_12125_),
    .Y(_12633_));
 sg13g2_buf_2 _19702_ (.A(_12633_),
    .X(_12634_));
 sg13g2_mux2_1 _19703_ (.A0(\cpu.dcache.r_data[4][20] ),
    .A1(net1087),
    .S(_12634_),
    .X(_12635_));
 sg13g2_nor2_1 _19704_ (.A(_12616_),
    .B(_12635_),
    .Y(_12636_));
 sg13g2_a21oi_1 _19705_ (.A1(net723),
    .A2(net45),
    .Y(_00439_),
    .B1(_12636_));
 sg13g2_nor2b_1 _19706_ (.A(_12634_),
    .B_N(\cpu.dcache.r_data[4][21] ),
    .Y(_12637_));
 sg13g2_a21oi_1 _19707_ (.A1(net975),
    .A2(_12634_),
    .Y(_12638_),
    .B1(_12637_));
 sg13g2_nand2_1 _19708_ (.Y(_12639_),
    .A(net984),
    .B(_12616_));
 sg13g2_o21ai_1 _19709_ (.B1(_12639_),
    .Y(_00440_),
    .A1(_12617_),
    .A2(_12638_));
 sg13g2_nor2b_1 _19710_ (.A(_12634_),
    .B_N(\cpu.dcache.r_data[4][22] ),
    .Y(_12640_));
 sg13g2_a21oi_1 _19711_ (.A1(net977),
    .A2(_12634_),
    .Y(_12641_),
    .B1(_12640_));
 sg13g2_nand2_1 _19712_ (.Y(_12642_),
    .A(net985),
    .B(_12616_));
 sg13g2_o21ai_1 _19713_ (.B1(_12642_),
    .Y(_00441_),
    .A1(_12617_),
    .A2(_12641_));
 sg13g2_mux2_1 _19714_ (.A0(\cpu.dcache.r_data[4][23] ),
    .A1(net1077),
    .S(_12634_),
    .X(_12643_));
 sg13g2_nor2_1 _19715_ (.A(_12616_),
    .B(_12643_),
    .Y(_12644_));
 sg13g2_a21oi_1 _19716_ (.A1(_12140_),
    .A2(net45),
    .Y(_00442_),
    .B1(_12644_));
 sg13g2_or2_1 _19717_ (.X(_12645_),
    .B(net643),
    .A(_12578_));
 sg13g2_buf_2 _19718_ (.A(_12645_),
    .X(_12646_));
 sg13g2_mux2_1 _19719_ (.A0(_12143_),
    .A1(\cpu.dcache.r_data[4][24] ),
    .S(_12646_),
    .X(_12647_));
 sg13g2_nor2_1 _19720_ (.A(_12153_),
    .B(_12580_),
    .Y(_12648_));
 sg13g2_buf_2 _19721_ (.A(_12648_),
    .X(_12649_));
 sg13g2_mux2_1 _19722_ (.A0(_12647_),
    .A1(net420),
    .S(net69),
    .X(_00443_));
 sg13g2_mux2_1 _19723_ (.A0(net1082),
    .A1(\cpu.dcache.r_data[4][25] ),
    .S(_12646_),
    .X(_12650_));
 sg13g2_mux2_1 _19724_ (.A0(_12650_),
    .A1(net369),
    .S(net69),
    .X(_00444_));
 sg13g2_mux2_1 _19725_ (.A0(net1081),
    .A1(\cpu.dcache.r_data[4][26] ),
    .S(_12646_),
    .X(_12651_));
 sg13g2_mux2_1 _19726_ (.A0(_12651_),
    .A1(_12043_),
    .S(_12649_),
    .X(_00445_));
 sg13g2_mux2_1 _19727_ (.A0(_12113_),
    .A1(\cpu.dcache.r_data[4][27] ),
    .S(_12646_),
    .X(_02658_));
 sg13g2_mux2_1 _19728_ (.A0(_02658_),
    .A1(_12164_),
    .S(_12649_),
    .X(_00446_));
 sg13g2_buf_1 _19729_ (.A(net1087),
    .X(_02659_));
 sg13g2_nor2_1 _19730_ (.A(_12578_),
    .B(_12166_),
    .Y(_02660_));
 sg13g2_buf_2 _19731_ (.A(_02660_),
    .X(_02661_));
 sg13g2_nor2b_1 _19732_ (.A(_02661_),
    .B_N(\cpu.dcache.r_data[4][28] ),
    .Y(_02662_));
 sg13g2_a21oi_1 _19733_ (.A1(net972),
    .A2(_02661_),
    .Y(_02663_),
    .B1(_02662_));
 sg13g2_nand2_1 _19734_ (.Y(_02664_),
    .A(_12171_),
    .B(net69));
 sg13g2_o21ai_1 _19735_ (.B1(_02664_),
    .Y(_00447_),
    .A1(net69),
    .A2(_02663_));
 sg13g2_nor2b_1 _19736_ (.A(_02661_),
    .B_N(\cpu.dcache.r_data[4][29] ),
    .Y(_02665_));
 sg13g2_a21oi_1 _19737_ (.A1(_12534_),
    .A2(_02661_),
    .Y(_02666_),
    .B1(_02665_));
 sg13g2_nand2_1 _19738_ (.Y(_02667_),
    .A(_12175_),
    .B(net69));
 sg13g2_o21ai_1 _19739_ (.B1(_02667_),
    .Y(_00448_),
    .A1(net69),
    .A2(_02666_));
 sg13g2_mux2_1 _19740_ (.A0(\cpu.dcache.r_data[4][2] ),
    .A1(_12262_),
    .S(_12585_),
    .X(_02668_));
 sg13g2_nor2_1 _19741_ (.A(_12582_),
    .B(_02668_),
    .Y(_02669_));
 sg13g2_a21oi_1 _19742_ (.A1(_12106_),
    .A2(net47),
    .Y(_00449_),
    .B1(_02669_));
 sg13g2_nor2b_1 _19743_ (.A(_02661_),
    .B_N(\cpu.dcache.r_data[4][30] ),
    .Y(_02670_));
 sg13g2_a21oi_1 _19744_ (.A1(_12447_),
    .A2(_02661_),
    .Y(_02671_),
    .B1(_02670_));
 sg13g2_nand2_1 _19745_ (.Y(_02672_),
    .A(net417),
    .B(_12648_));
 sg13g2_o21ai_1 _19746_ (.B1(_02672_),
    .Y(_00450_),
    .A1(net69),
    .A2(_02671_));
 sg13g2_nor2b_1 _19747_ (.A(_02661_),
    .B_N(\cpu.dcache.r_data[4][31] ),
    .Y(_02673_));
 sg13g2_a21oi_1 _19748_ (.A1(net973),
    .A2(_02661_),
    .Y(_02674_),
    .B1(_02673_));
 sg13g2_nand2_1 _19749_ (.Y(_02675_),
    .A(_12185_),
    .B(_12648_));
 sg13g2_o21ai_1 _19750_ (.B1(_02675_),
    .Y(_00451_),
    .A1(net69),
    .A2(_02674_));
 sg13g2_mux2_1 _19751_ (.A0(\cpu.dcache.r_data[4][3] ),
    .A1(net1077),
    .S(_12585_),
    .X(_02676_));
 sg13g2_nor2_1 _19752_ (.A(_12582_),
    .B(_02676_),
    .Y(_02677_));
 sg13g2_a21oi_1 _19753_ (.A1(_12112_),
    .A2(net47),
    .Y(_00452_),
    .B1(_02677_));
 sg13g2_nor2_1 _19754_ (.A(net583),
    .B(_12190_),
    .Y(_02678_));
 sg13g2_buf_2 _19755_ (.A(_02678_),
    .X(_02679_));
 sg13g2_mux2_1 _19756_ (.A0(\cpu.dcache.r_data[4][4] ),
    .A1(net1087),
    .S(_02679_),
    .X(_02680_));
 sg13g2_nor2_1 _19757_ (.A(_12582_),
    .B(_02680_),
    .Y(_02681_));
 sg13g2_a21oi_1 _19758_ (.A1(_12121_),
    .A2(net47),
    .Y(_00453_),
    .B1(_02681_));
 sg13g2_nor2b_1 _19759_ (.A(_02679_),
    .B_N(\cpu.dcache.r_data[4][5] ),
    .Y(_02682_));
 sg13g2_a21oi_1 _19760_ (.A1(net975),
    .A2(_02679_),
    .Y(_02683_),
    .B1(_02682_));
 sg13g2_nand2_1 _19761_ (.Y(_02684_),
    .A(_12197_),
    .B(_12582_));
 sg13g2_o21ai_1 _19762_ (.B1(_02684_),
    .Y(_00454_),
    .A1(_12583_),
    .A2(_02683_));
 sg13g2_nor2b_1 _19763_ (.A(_02679_),
    .B_N(\cpu.dcache.r_data[4][6] ),
    .Y(_02685_));
 sg13g2_a21oi_1 _19764_ (.A1(net977),
    .A2(_02679_),
    .Y(_02686_),
    .B1(_02685_));
 sg13g2_nand2_1 _19765_ (.Y(_02687_),
    .A(net985),
    .B(_12582_));
 sg13g2_o21ai_1 _19766_ (.B1(_02687_),
    .Y(_00455_),
    .A1(_12583_),
    .A2(_02686_));
 sg13g2_mux2_1 _19767_ (.A0(\cpu.dcache.r_data[4][7] ),
    .A1(net1077),
    .S(_02679_),
    .X(_02688_));
 sg13g2_nor2_1 _19768_ (.A(_12582_),
    .B(_02688_),
    .Y(_02689_));
 sg13g2_a21oi_1 _19769_ (.A1(_12140_),
    .A2(net47),
    .Y(_00456_),
    .B1(_02689_));
 sg13g2_nor2b_1 _19770_ (.A(_12593_),
    .B_N(\cpu.dcache.r_data[4][8] ),
    .Y(_02690_));
 sg13g2_a21oi_1 _19771_ (.A1(net972),
    .A2(_12593_),
    .Y(_02691_),
    .B1(_02690_));
 sg13g2_nand2_1 _19772_ (.Y(_02692_),
    .A(net420),
    .B(_12590_));
 sg13g2_o21ai_1 _19773_ (.B1(_02692_),
    .Y(_00457_),
    .A1(_12591_),
    .A2(_02691_));
 sg13g2_nor2b_1 _19774_ (.A(_12593_),
    .B_N(\cpu.dcache.r_data[4][9] ),
    .Y(_02693_));
 sg13g2_a21oi_1 _19775_ (.A1(net975),
    .A2(_12593_),
    .Y(_02694_),
    .B1(_02693_));
 sg13g2_nand2_1 _19776_ (.Y(_02695_),
    .A(net369),
    .B(_12590_));
 sg13g2_o21ai_1 _19777_ (.B1(_02695_),
    .Y(_00458_),
    .A1(net46),
    .A2(_02694_));
 sg13g2_nand2_1 _19778_ (.Y(_02696_),
    .A(net781),
    .B(_09331_));
 sg13g2_buf_2 _19779_ (.A(_02696_),
    .X(_02697_));
 sg13g2_buf_1 _19780_ (.A(_02697_),
    .X(_02698_));
 sg13g2_or2_1 _19781_ (.X(_02699_),
    .B(_11999_),
    .A(net516));
 sg13g2_buf_1 _19782_ (.A(_02699_),
    .X(_02700_));
 sg13g2_nor2_1 _19783_ (.A(_11987_),
    .B(_02700_),
    .Y(_02701_));
 sg13g2_buf_1 _19784_ (.A(_02701_),
    .X(_02702_));
 sg13g2_buf_1 _19785_ (.A(_02702_),
    .X(_02703_));
 sg13g2_nor2_1 _19786_ (.A(net516),
    .B(_12016_),
    .Y(_02704_));
 sg13g2_buf_2 _19787_ (.A(_02704_),
    .X(_02705_));
 sg13g2_nor2b_1 _19788_ (.A(_02705_),
    .B_N(\cpu.dcache.r_data[5][0] ),
    .Y(_02706_));
 sg13g2_a21oi_1 _19789_ (.A1(_02659_),
    .A2(_02705_),
    .Y(_02707_),
    .B1(_02706_));
 sg13g2_nand2_1 _19790_ (.Y(_02708_),
    .A(_12222_),
    .B(net44));
 sg13g2_o21ai_1 _19791_ (.B1(_02708_),
    .Y(_00459_),
    .A1(net44),
    .A2(_02707_));
 sg13g2_nor2_1 _19792_ (.A(_12025_),
    .B(_02700_),
    .Y(_02709_));
 sg13g2_buf_2 _19793_ (.A(_02709_),
    .X(_02710_));
 sg13g2_buf_1 _19794_ (.A(_02710_),
    .X(_02711_));
 sg13g2_buf_1 _19795_ (.A(_12030_),
    .X(_02712_));
 sg13g2_nor2_1 _19796_ (.A(net516),
    .B(_12033_),
    .Y(_02713_));
 sg13g2_buf_2 _19797_ (.A(_02713_),
    .X(_02714_));
 sg13g2_nor2b_1 _19798_ (.A(_02714_),
    .B_N(\cpu.dcache.r_data[5][10] ),
    .Y(_02715_));
 sg13g2_a21oi_1 _19799_ (.A1(net971),
    .A2(_02714_),
    .Y(_02716_),
    .B1(_02715_));
 sg13g2_nand2_1 _19800_ (.Y(_02717_),
    .A(_12042_),
    .B(net43));
 sg13g2_o21ai_1 _19801_ (.B1(_02717_),
    .Y(_00460_),
    .A1(_02711_),
    .A2(_02716_));
 sg13g2_nor2b_1 _19802_ (.A(_02714_),
    .B_N(\cpu.dcache.r_data[5][11] ),
    .Y(_02718_));
 sg13g2_a21oi_1 _19803_ (.A1(net973),
    .A2(_02714_),
    .Y(_02719_),
    .B1(_02718_));
 sg13g2_nand2_1 _19804_ (.Y(_02720_),
    .A(net419),
    .B(net43));
 sg13g2_o21ai_1 _19805_ (.B1(_02720_),
    .Y(_00461_),
    .A1(net43),
    .A2(_02719_));
 sg13g2_nor2_1 _19806_ (.A(net516),
    .B(_12055_),
    .Y(_02721_));
 sg13g2_buf_2 _19807_ (.A(_02721_),
    .X(_02722_));
 sg13g2_nor2b_1 _19808_ (.A(_02722_),
    .B_N(\cpu.dcache.r_data[5][12] ),
    .Y(_02723_));
 sg13g2_a21oi_1 _19809_ (.A1(net972),
    .A2(_02722_),
    .Y(_02724_),
    .B1(_02723_));
 sg13g2_nand2_1 _19810_ (.Y(_02725_),
    .A(net368),
    .B(_02710_));
 sg13g2_o21ai_1 _19811_ (.B1(_02725_),
    .Y(_00462_),
    .A1(net43),
    .A2(_02724_));
 sg13g2_buf_1 _19812_ (.A(_12065_),
    .X(_02726_));
 sg13g2_nor2b_1 _19813_ (.A(_02722_),
    .B_N(\cpu.dcache.r_data[5][13] ),
    .Y(_02727_));
 sg13g2_a21oi_1 _19814_ (.A1(net1076),
    .A2(_02722_),
    .Y(_02728_),
    .B1(_02727_));
 sg13g2_nand2_1 _19815_ (.Y(_02729_),
    .A(net418),
    .B(_02710_));
 sg13g2_o21ai_1 _19816_ (.B1(_02729_),
    .Y(_00463_),
    .A1(net43),
    .A2(_02728_));
 sg13g2_nor2b_1 _19817_ (.A(_02722_),
    .B_N(\cpu.dcache.r_data[5][14] ),
    .Y(_02730_));
 sg13g2_a21oi_1 _19818_ (.A1(net971),
    .A2(_02722_),
    .Y(_02731_),
    .B1(_02730_));
 sg13g2_nand2_1 _19819_ (.Y(_02732_),
    .A(net417),
    .B(_02710_));
 sg13g2_o21ai_1 _19820_ (.B1(_02732_),
    .Y(_00464_),
    .A1(net43),
    .A2(_02731_));
 sg13g2_nor2b_1 _19821_ (.A(_02722_),
    .B_N(\cpu.dcache.r_data[5][15] ),
    .Y(_02733_));
 sg13g2_a21oi_1 _19822_ (.A1(net973),
    .A2(_02722_),
    .Y(_02734_),
    .B1(_02733_));
 sg13g2_nand2_1 _19823_ (.Y(_02735_),
    .A(net416),
    .B(_02710_));
 sg13g2_o21ai_1 _19824_ (.B1(_02735_),
    .Y(_00465_),
    .A1(net43),
    .A2(_02734_));
 sg13g2_nor2_1 _19825_ (.A(_12090_),
    .B(_02700_),
    .Y(_02736_));
 sg13g2_buf_1 _19826_ (.A(_02736_),
    .X(_02737_));
 sg13g2_buf_1 _19827_ (.A(_02737_),
    .X(_02738_));
 sg13g2_nor2_1 _19828_ (.A(net516),
    .B(_12096_),
    .Y(_02739_));
 sg13g2_buf_2 _19829_ (.A(_02739_),
    .X(_02740_));
 sg13g2_nor2b_1 _19830_ (.A(_02740_),
    .B_N(\cpu.dcache.r_data[5][16] ),
    .Y(_02741_));
 sg13g2_a21oi_1 _19831_ (.A1(net972),
    .A2(_02740_),
    .Y(_02742_),
    .B1(_02741_));
 sg13g2_nand2_1 _19832_ (.Y(_02743_),
    .A(_12222_),
    .B(net42));
 sg13g2_o21ai_1 _19833_ (.B1(_02743_),
    .Y(_00466_),
    .A1(net42),
    .A2(_02742_));
 sg13g2_nor2b_1 _19834_ (.A(_02740_),
    .B_N(\cpu.dcache.r_data[5][17] ),
    .Y(_02744_));
 sg13g2_a21oi_1 _19835_ (.A1(net1076),
    .A2(_02740_),
    .Y(_02745_),
    .B1(_02744_));
 sg13g2_nand2_1 _19836_ (.Y(_02746_),
    .A(net850),
    .B(net42));
 sg13g2_o21ai_1 _19837_ (.B1(_02746_),
    .Y(_00467_),
    .A1(net42),
    .A2(_02745_));
 sg13g2_mux2_1 _19838_ (.A0(\cpu.dcache.r_data[5][18] ),
    .A1(_12262_),
    .S(_02740_),
    .X(_02747_));
 sg13g2_nor2_1 _19839_ (.A(_02737_),
    .B(_02747_),
    .Y(_02748_));
 sg13g2_a21oi_1 _19840_ (.A1(net753),
    .A2(net42),
    .Y(_00468_),
    .B1(_02748_));
 sg13g2_buf_1 _19841_ (.A(net854),
    .X(_02749_));
 sg13g2_mux2_1 _19842_ (.A0(\cpu.dcache.r_data[5][19] ),
    .A1(net1077),
    .S(_02740_),
    .X(_02750_));
 sg13g2_nor2_1 _19843_ (.A(_02737_),
    .B(_02750_),
    .Y(_02751_));
 sg13g2_a21oi_1 _19844_ (.A1(net721),
    .A2(net42),
    .Y(_00469_),
    .B1(_02751_));
 sg13g2_nor2b_1 _19845_ (.A(_02705_),
    .B_N(\cpu.dcache.r_data[5][1] ),
    .Y(_02752_));
 sg13g2_a21oi_1 _19846_ (.A1(net1076),
    .A2(_02705_),
    .Y(_02753_),
    .B1(_02752_));
 sg13g2_nand2_1 _19847_ (.Y(_02754_),
    .A(net850),
    .B(net44));
 sg13g2_o21ai_1 _19848_ (.B1(_02754_),
    .Y(_00470_),
    .A1(net44),
    .A2(_02753_));
 sg13g2_buf_1 _19849_ (.A(net853),
    .X(_02755_));
 sg13g2_nor2_1 _19850_ (.A(net516),
    .B(_12125_),
    .Y(_02756_));
 sg13g2_buf_2 _19851_ (.A(_02756_),
    .X(_02757_));
 sg13g2_mux2_1 _19852_ (.A0(\cpu.dcache.r_data[5][20] ),
    .A1(net1087),
    .S(_02757_),
    .X(_02758_));
 sg13g2_nor2_1 _19853_ (.A(_02737_),
    .B(_02758_),
    .Y(_02759_));
 sg13g2_a21oi_1 _19854_ (.A1(net720),
    .A2(_02738_),
    .Y(_00471_),
    .B1(_02759_));
 sg13g2_nor2b_1 _19855_ (.A(_02757_),
    .B_N(\cpu.dcache.r_data[5][21] ),
    .Y(_02760_));
 sg13g2_a21oi_1 _19856_ (.A1(net1076),
    .A2(_02757_),
    .Y(_02761_),
    .B1(_02760_));
 sg13g2_nand2_1 _19857_ (.Y(_02762_),
    .A(net984),
    .B(_02737_));
 sg13g2_o21ai_1 _19858_ (.B1(_02762_),
    .Y(_00472_),
    .A1(net42),
    .A2(_02761_));
 sg13g2_nor2b_1 _19859_ (.A(_02757_),
    .B_N(\cpu.dcache.r_data[5][22] ),
    .Y(_02763_));
 sg13g2_a21oi_1 _19860_ (.A1(net971),
    .A2(_02757_),
    .Y(_02764_),
    .B1(_02763_));
 sg13g2_nand2_1 _19861_ (.Y(_02765_),
    .A(net985),
    .B(_02737_));
 sg13g2_o21ai_1 _19862_ (.B1(_02765_),
    .Y(_00473_),
    .A1(_02738_),
    .A2(_02764_));
 sg13g2_buf_1 _19863_ (.A(net852),
    .X(_02766_));
 sg13g2_mux2_1 _19864_ (.A0(\cpu.dcache.r_data[5][23] ),
    .A1(_12560_),
    .S(_02757_),
    .X(_02767_));
 sg13g2_nor2_1 _19865_ (.A(_02737_),
    .B(_02767_),
    .Y(_02768_));
 sg13g2_a21oi_1 _19866_ (.A1(net719),
    .A2(net42),
    .Y(_00474_),
    .B1(_02768_));
 sg13g2_nor2_1 _19867_ (.A(_12153_),
    .B(_02700_),
    .Y(_02769_));
 sg13g2_buf_2 _19868_ (.A(_02769_),
    .X(_02770_));
 sg13g2_buf_1 _19869_ (.A(_02770_),
    .X(_02771_));
 sg13g2_nor2_1 _19870_ (.A(net516),
    .B(net643),
    .Y(_02772_));
 sg13g2_buf_1 _19871_ (.A(_02772_),
    .X(_02773_));
 sg13g2_nor2b_1 _19872_ (.A(net414),
    .B_N(\cpu.dcache.r_data[5][24] ),
    .Y(_02774_));
 sg13g2_a21oi_1 _19873_ (.A1(net972),
    .A2(net414),
    .Y(_02775_),
    .B1(_02774_));
 sg13g2_nand2_1 _19874_ (.Y(_02776_),
    .A(_12149_),
    .B(net41));
 sg13g2_o21ai_1 _19875_ (.B1(_02776_),
    .Y(_00475_),
    .A1(net41),
    .A2(_02775_));
 sg13g2_nor2b_1 _19876_ (.A(net414),
    .B_N(\cpu.dcache.r_data[5][25] ),
    .Y(_02777_));
 sg13g2_a21oi_1 _19877_ (.A1(net1076),
    .A2(net414),
    .Y(_02778_),
    .B1(_02777_));
 sg13g2_nand2_1 _19878_ (.Y(_02779_),
    .A(_12161_),
    .B(net41));
 sg13g2_o21ai_1 _19879_ (.B1(_02779_),
    .Y(_00476_),
    .A1(net41),
    .A2(_02778_));
 sg13g2_nor2b_1 _19880_ (.A(net414),
    .B_N(\cpu.dcache.r_data[5][26] ),
    .Y(_02780_));
 sg13g2_a21oi_1 _19881_ (.A1(net971),
    .A2(net414),
    .Y(_02781_),
    .B1(_02780_));
 sg13g2_nand2_1 _19882_ (.Y(_02782_),
    .A(_12042_),
    .B(_02770_));
 sg13g2_o21ai_1 _19883_ (.B1(_02782_),
    .Y(_00477_),
    .A1(_02771_),
    .A2(_02781_));
 sg13g2_nor2b_1 _19884_ (.A(net414),
    .B_N(\cpu.dcache.r_data[5][27] ),
    .Y(_02783_));
 sg13g2_a21oi_1 _19885_ (.A1(net973),
    .A2(net414),
    .Y(_02784_),
    .B1(_02783_));
 sg13g2_nand2_1 _19886_ (.Y(_02785_),
    .A(_12051_),
    .B(_02770_));
 sg13g2_o21ai_1 _19887_ (.B1(_02785_),
    .Y(_00478_),
    .A1(_02771_),
    .A2(_02784_));
 sg13g2_nor2_1 _19888_ (.A(_02698_),
    .B(_12166_),
    .Y(_02786_));
 sg13g2_buf_2 _19889_ (.A(_02786_),
    .X(_02787_));
 sg13g2_nor2b_1 _19890_ (.A(_02787_),
    .B_N(\cpu.dcache.r_data[5][28] ),
    .Y(_02788_));
 sg13g2_a21oi_1 _19891_ (.A1(net972),
    .A2(_02787_),
    .Y(_02789_),
    .B1(_02788_));
 sg13g2_nand2_1 _19892_ (.Y(_02790_),
    .A(_12063_),
    .B(_02770_));
 sg13g2_o21ai_1 _19893_ (.B1(_02790_),
    .Y(_00479_),
    .A1(net41),
    .A2(_02789_));
 sg13g2_nor2b_1 _19894_ (.A(_02787_),
    .B_N(\cpu.dcache.r_data[5][29] ),
    .Y(_02791_));
 sg13g2_a21oi_1 _19895_ (.A1(net1076),
    .A2(_02787_),
    .Y(_02792_),
    .B1(_02791_));
 sg13g2_nand2_1 _19896_ (.Y(_02793_),
    .A(_12073_),
    .B(_02770_));
 sg13g2_o21ai_1 _19897_ (.B1(_02793_),
    .Y(_00480_),
    .A1(net41),
    .A2(_02792_));
 sg13g2_mux2_1 _19898_ (.A0(\cpu.dcache.r_data[5][2] ),
    .A1(net1078),
    .S(_02705_),
    .X(_02794_));
 sg13g2_nor2_1 _19899_ (.A(_02702_),
    .B(_02794_),
    .Y(_02795_));
 sg13g2_a21oi_1 _19900_ (.A1(net753),
    .A2(_02703_),
    .Y(_00481_),
    .B1(_02795_));
 sg13g2_nor2b_1 _19901_ (.A(_02787_),
    .B_N(\cpu.dcache.r_data[5][30] ),
    .Y(_02796_));
 sg13g2_a21oi_1 _19902_ (.A1(net971),
    .A2(_02787_),
    .Y(_02797_),
    .B1(_02796_));
 sg13g2_nand2_1 _19903_ (.Y(_02798_),
    .A(_12080_),
    .B(_02770_));
 sg13g2_o21ai_1 _19904_ (.B1(_02798_),
    .Y(_00482_),
    .A1(net41),
    .A2(_02797_));
 sg13g2_nor2b_1 _19905_ (.A(_02787_),
    .B_N(\cpu.dcache.r_data[5][31] ),
    .Y(_02799_));
 sg13g2_a21oi_1 _19906_ (.A1(net973),
    .A2(_02787_),
    .Y(_02800_),
    .B1(_02799_));
 sg13g2_nand2_1 _19907_ (.Y(_02801_),
    .A(_12087_),
    .B(_02770_));
 sg13g2_o21ai_1 _19908_ (.B1(_02801_),
    .Y(_00483_),
    .A1(net41),
    .A2(_02800_));
 sg13g2_mux2_1 _19909_ (.A0(\cpu.dcache.r_data[5][3] ),
    .A1(net1077),
    .S(_02705_),
    .X(_02802_));
 sg13g2_nor2_1 _19910_ (.A(_02702_),
    .B(_02802_),
    .Y(_02803_));
 sg13g2_a21oi_1 _19911_ (.A1(net721),
    .A2(_02703_),
    .Y(_00484_),
    .B1(_02803_));
 sg13g2_nor2_1 _19912_ (.A(net516),
    .B(_12190_),
    .Y(_02804_));
 sg13g2_buf_2 _19913_ (.A(_02804_),
    .X(_02805_));
 sg13g2_mux2_1 _19914_ (.A0(\cpu.dcache.r_data[5][4] ),
    .A1(_12006_),
    .S(_02805_),
    .X(_02806_));
 sg13g2_nor2_1 _19915_ (.A(_02702_),
    .B(_02806_),
    .Y(_02807_));
 sg13g2_a21oi_1 _19916_ (.A1(net720),
    .A2(net44),
    .Y(_00485_),
    .B1(_02807_));
 sg13g2_nor2b_1 _19917_ (.A(_02805_),
    .B_N(\cpu.dcache.r_data[5][5] ),
    .Y(_02808_));
 sg13g2_a21oi_1 _19918_ (.A1(net1076),
    .A2(_02805_),
    .Y(_02809_),
    .B1(_02808_));
 sg13g2_nand2_1 _19919_ (.Y(_02810_),
    .A(net984),
    .B(_02702_));
 sg13g2_o21ai_1 _19920_ (.B1(_02810_),
    .Y(_00486_),
    .A1(net44),
    .A2(_02809_));
 sg13g2_nor2b_1 _19921_ (.A(_02805_),
    .B_N(\cpu.dcache.r_data[5][6] ),
    .Y(_02811_));
 sg13g2_a21oi_1 _19922_ (.A1(net971),
    .A2(_02805_),
    .Y(_02812_),
    .B1(_02811_));
 sg13g2_nand2_1 _19923_ (.Y(_02813_),
    .A(net1020),
    .B(_02702_));
 sg13g2_o21ai_1 _19924_ (.B1(_02813_),
    .Y(_00487_),
    .A1(net44),
    .A2(_02812_));
 sg13g2_mux2_1 _19925_ (.A0(\cpu.dcache.r_data[5][7] ),
    .A1(_12560_),
    .S(_02805_),
    .X(_02814_));
 sg13g2_nor2_1 _19926_ (.A(_02702_),
    .B(_02814_),
    .Y(_02815_));
 sg13g2_a21oi_1 _19927_ (.A1(net719),
    .A2(net44),
    .Y(_00488_),
    .B1(_02815_));
 sg13g2_nor2b_1 _19928_ (.A(_02714_),
    .B_N(\cpu.dcache.r_data[5][8] ),
    .Y(_02816_));
 sg13g2_a21oi_1 _19929_ (.A1(net972),
    .A2(_02714_),
    .Y(_02817_),
    .B1(_02816_));
 sg13g2_nand2_1 _19930_ (.Y(_02818_),
    .A(_12148_),
    .B(_02710_));
 sg13g2_o21ai_1 _19931_ (.B1(_02818_),
    .Y(_00489_),
    .A1(_02711_),
    .A2(_02817_));
 sg13g2_nor2b_1 _19932_ (.A(_02714_),
    .B_N(\cpu.dcache.r_data[5][9] ),
    .Y(_02819_));
 sg13g2_a21oi_1 _19933_ (.A1(_02726_),
    .A2(_02714_),
    .Y(_02820_),
    .B1(_02819_));
 sg13g2_nand2_1 _19934_ (.Y(_02821_),
    .A(_12160_),
    .B(_02710_));
 sg13g2_o21ai_1 _19935_ (.B1(_02821_),
    .Y(_00490_),
    .A1(net43),
    .A2(_02820_));
 sg13g2_buf_1 _19936_ (.A(_09340_),
    .X(_02822_));
 sg13g2_or2_1 _19937_ (.X(_02823_),
    .B(_11999_),
    .A(net642));
 sg13g2_buf_1 _19938_ (.A(_02823_),
    .X(_02824_));
 sg13g2_nor2_1 _19939_ (.A(_11987_),
    .B(_02824_),
    .Y(_02825_));
 sg13g2_buf_2 _19940_ (.A(_02825_),
    .X(_02826_));
 sg13g2_buf_1 _19941_ (.A(_02826_),
    .X(_02827_));
 sg13g2_nor2_1 _19942_ (.A(net642),
    .B(_12016_),
    .Y(_02828_));
 sg13g2_buf_2 _19943_ (.A(_02828_),
    .X(_02829_));
 sg13g2_nor2b_1 _19944_ (.A(_02829_),
    .B_N(\cpu.dcache.r_data[6][0] ),
    .Y(_02830_));
 sg13g2_a21oi_1 _19945_ (.A1(_02659_),
    .A2(_02829_),
    .Y(_02831_),
    .B1(_02830_));
 sg13g2_buf_1 _19946_ (.A(_09859_),
    .X(_02832_));
 sg13g2_nand2_1 _19947_ (.Y(_02833_),
    .A(net970),
    .B(net40));
 sg13g2_o21ai_1 _19948_ (.B1(_02833_),
    .Y(_00491_),
    .A1(net40),
    .A2(_02831_));
 sg13g2_nor2_1 _19949_ (.A(_12025_),
    .B(_02824_),
    .Y(_02834_));
 sg13g2_buf_2 _19950_ (.A(_02834_),
    .X(_02835_));
 sg13g2_buf_1 _19951_ (.A(_02835_),
    .X(_02836_));
 sg13g2_nor2_1 _19952_ (.A(net642),
    .B(_12033_),
    .Y(_02837_));
 sg13g2_buf_2 _19953_ (.A(_02837_),
    .X(_02838_));
 sg13g2_nor2b_1 _19954_ (.A(_02838_),
    .B_N(\cpu.dcache.r_data[6][10] ),
    .Y(_02839_));
 sg13g2_a21oi_1 _19955_ (.A1(net971),
    .A2(_02838_),
    .Y(_02840_),
    .B1(_02839_));
 sg13g2_nand2_1 _19956_ (.Y(_02841_),
    .A(_12042_),
    .B(_02836_));
 sg13g2_o21ai_1 _19957_ (.B1(_02841_),
    .Y(_00492_),
    .A1(net39),
    .A2(_02840_));
 sg13g2_nor2b_1 _19958_ (.A(_02838_),
    .B_N(\cpu.dcache.r_data[6][11] ),
    .Y(_02842_));
 sg13g2_a21oi_1 _19959_ (.A1(net973),
    .A2(_02838_),
    .Y(_02843_),
    .B1(_02842_));
 sg13g2_nand2_1 _19960_ (.Y(_02844_),
    .A(_12051_),
    .B(_02836_));
 sg13g2_o21ai_1 _19961_ (.B1(_02844_),
    .Y(_00493_),
    .A1(net39),
    .A2(_02843_));
 sg13g2_nor2_1 _19962_ (.A(net642),
    .B(_12055_),
    .Y(_02845_));
 sg13g2_buf_2 _19963_ (.A(_02845_),
    .X(_02846_));
 sg13g2_nor2b_1 _19964_ (.A(_02846_),
    .B_N(\cpu.dcache.r_data[6][12] ),
    .Y(_02847_));
 sg13g2_a21oi_1 _19965_ (.A1(net972),
    .A2(_02846_),
    .Y(_02848_),
    .B1(_02847_));
 sg13g2_nand2_1 _19966_ (.Y(_02849_),
    .A(_12063_),
    .B(_02835_));
 sg13g2_o21ai_1 _19967_ (.B1(_02849_),
    .Y(_00494_),
    .A1(net39),
    .A2(_02848_));
 sg13g2_nor2b_1 _19968_ (.A(_02846_),
    .B_N(\cpu.dcache.r_data[6][13] ),
    .Y(_02850_));
 sg13g2_a21oi_1 _19969_ (.A1(_02726_),
    .A2(_02846_),
    .Y(_02851_),
    .B1(_02850_));
 sg13g2_nand2_1 _19970_ (.Y(_02852_),
    .A(_12073_),
    .B(_02835_));
 sg13g2_o21ai_1 _19971_ (.B1(_02852_),
    .Y(_00495_),
    .A1(net39),
    .A2(_02851_));
 sg13g2_nor2b_1 _19972_ (.A(_02846_),
    .B_N(\cpu.dcache.r_data[6][14] ),
    .Y(_02853_));
 sg13g2_a21oi_1 _19973_ (.A1(_02712_),
    .A2(_02846_),
    .Y(_02854_),
    .B1(_02853_));
 sg13g2_nand2_1 _19974_ (.Y(_02855_),
    .A(_12080_),
    .B(_02835_));
 sg13g2_o21ai_1 _19975_ (.B1(_02855_),
    .Y(_00496_),
    .A1(net39),
    .A2(_02854_));
 sg13g2_nor2b_1 _19976_ (.A(_02846_),
    .B_N(\cpu.dcache.r_data[6][15] ),
    .Y(_02856_));
 sg13g2_a21oi_1 _19977_ (.A1(net973),
    .A2(_02846_),
    .Y(_02857_),
    .B1(_02856_));
 sg13g2_nand2_1 _19978_ (.Y(_02858_),
    .A(_12087_),
    .B(_02835_));
 sg13g2_o21ai_1 _19979_ (.B1(_02858_),
    .Y(_00497_),
    .A1(net39),
    .A2(_02857_));
 sg13g2_nor2_1 _19980_ (.A(_12090_),
    .B(_02824_),
    .Y(_02859_));
 sg13g2_buf_1 _19981_ (.A(_02859_),
    .X(_02860_));
 sg13g2_buf_1 _19982_ (.A(_02860_),
    .X(_02861_));
 sg13g2_buf_1 _19983_ (.A(_12005_),
    .X(_02862_));
 sg13g2_nor2_1 _19984_ (.A(net642),
    .B(_12096_),
    .Y(_02863_));
 sg13g2_buf_2 _19985_ (.A(_02863_),
    .X(_02864_));
 sg13g2_nor2b_1 _19986_ (.A(_02864_),
    .B_N(\cpu.dcache.r_data[6][16] ),
    .Y(_02865_));
 sg13g2_a21oi_1 _19987_ (.A1(net1075),
    .A2(_02864_),
    .Y(_02866_),
    .B1(_02865_));
 sg13g2_nand2_1 _19988_ (.Y(_02867_),
    .A(net970),
    .B(net38));
 sg13g2_o21ai_1 _19989_ (.B1(_02867_),
    .Y(_00498_),
    .A1(net38),
    .A2(_02866_));
 sg13g2_nor2b_1 _19990_ (.A(_02864_),
    .B_N(\cpu.dcache.r_data[6][17] ),
    .Y(_02868_));
 sg13g2_a21oi_1 _19991_ (.A1(net1076),
    .A2(_02864_),
    .Y(_02869_),
    .B1(_02868_));
 sg13g2_nand2_1 _19992_ (.Y(_02870_),
    .A(_12391_),
    .B(net38));
 sg13g2_o21ai_1 _19993_ (.B1(_02870_),
    .Y(_00499_),
    .A1(net38),
    .A2(_02869_));
 sg13g2_mux2_1 _19994_ (.A0(\cpu.dcache.r_data[6][18] ),
    .A1(net1084),
    .S(_02864_),
    .X(_02871_));
 sg13g2_nor2_1 _19995_ (.A(_02860_),
    .B(_02871_),
    .Y(_02872_));
 sg13g2_a21oi_1 _19996_ (.A1(net753),
    .A2(net38),
    .Y(_00500_),
    .B1(_02872_));
 sg13g2_mux2_1 _19997_ (.A0(\cpu.dcache.r_data[6][19] ),
    .A1(net1077),
    .S(_02864_),
    .X(_02873_));
 sg13g2_nor2_1 _19998_ (.A(_02860_),
    .B(_02873_),
    .Y(_02874_));
 sg13g2_a21oi_1 _19999_ (.A1(net721),
    .A2(_02861_),
    .Y(_00501_),
    .B1(_02874_));
 sg13g2_buf_1 _20000_ (.A(_12065_),
    .X(_02875_));
 sg13g2_nor2b_1 _20001_ (.A(_02829_),
    .B_N(\cpu.dcache.r_data[6][1] ),
    .Y(_02876_));
 sg13g2_a21oi_1 _20002_ (.A1(net1074),
    .A2(_02829_),
    .Y(_02877_),
    .B1(_02876_));
 sg13g2_nand2_1 _20003_ (.Y(_02878_),
    .A(_12391_),
    .B(net40));
 sg13g2_o21ai_1 _20004_ (.B1(_02878_),
    .Y(_00502_),
    .A1(net40),
    .A2(_02877_));
 sg13g2_nor2_1 _20005_ (.A(net642),
    .B(_12125_),
    .Y(_02879_));
 sg13g2_buf_2 _20006_ (.A(_02879_),
    .X(_02880_));
 sg13g2_mux2_1 _20007_ (.A0(\cpu.dcache.r_data[6][20] ),
    .A1(net1087),
    .S(_02880_),
    .X(_02881_));
 sg13g2_nor2_1 _20008_ (.A(_02860_),
    .B(_02881_),
    .Y(_02882_));
 sg13g2_a21oi_1 _20009_ (.A1(_02755_),
    .A2(net38),
    .Y(_00503_),
    .B1(_02882_));
 sg13g2_nor2b_1 _20010_ (.A(_02880_),
    .B_N(\cpu.dcache.r_data[6][21] ),
    .Y(_02883_));
 sg13g2_a21oi_1 _20011_ (.A1(net1074),
    .A2(_02880_),
    .Y(_02884_),
    .B1(_02883_));
 sg13g2_nand2_1 _20012_ (.Y(_02885_),
    .A(net984),
    .B(_02860_));
 sg13g2_o21ai_1 _20013_ (.B1(_02885_),
    .Y(_00504_),
    .A1(_02861_),
    .A2(_02884_));
 sg13g2_nor2b_1 _20014_ (.A(_02880_),
    .B_N(\cpu.dcache.r_data[6][22] ),
    .Y(_02886_));
 sg13g2_a21oi_1 _20015_ (.A1(net971),
    .A2(_02880_),
    .Y(_02887_),
    .B1(_02886_));
 sg13g2_nand2_1 _20016_ (.Y(_02888_),
    .A(net1020),
    .B(_02860_));
 sg13g2_o21ai_1 _20017_ (.B1(_02888_),
    .Y(_00505_),
    .A1(net38),
    .A2(_02887_));
 sg13g2_mux2_1 _20018_ (.A0(\cpu.dcache.r_data[6][23] ),
    .A1(net1083),
    .S(_02880_),
    .X(_02889_));
 sg13g2_nor2_1 _20019_ (.A(_02860_),
    .B(_02889_),
    .Y(_02890_));
 sg13g2_a21oi_1 _20020_ (.A1(net719),
    .A2(net38),
    .Y(_00506_),
    .B1(_02890_));
 sg13g2_nor2_1 _20021_ (.A(_12153_),
    .B(_02824_),
    .Y(_02891_));
 sg13g2_buf_2 _20022_ (.A(_02891_),
    .X(_02892_));
 sg13g2_buf_1 _20023_ (.A(_02892_),
    .X(_02893_));
 sg13g2_nor2_1 _20024_ (.A(net642),
    .B(_11995_),
    .Y(_02894_));
 sg13g2_buf_1 _20025_ (.A(_02894_),
    .X(_02895_));
 sg13g2_nor2b_1 _20026_ (.A(net515),
    .B_N(\cpu.dcache.r_data[6][24] ),
    .Y(_02896_));
 sg13g2_a21oi_1 _20027_ (.A1(net1075),
    .A2(net515),
    .Y(_02897_),
    .B1(_02896_));
 sg13g2_nand2_1 _20028_ (.Y(_02898_),
    .A(_12148_),
    .B(net37));
 sg13g2_o21ai_1 _20029_ (.B1(_02898_),
    .Y(_00507_),
    .A1(net37),
    .A2(_02897_));
 sg13g2_nor2b_1 _20030_ (.A(net515),
    .B_N(\cpu.dcache.r_data[6][25] ),
    .Y(_02899_));
 sg13g2_a21oi_1 _20031_ (.A1(net1074),
    .A2(net515),
    .Y(_02900_),
    .B1(_02899_));
 sg13g2_nand2_1 _20032_ (.Y(_02901_),
    .A(_12160_),
    .B(net37));
 sg13g2_o21ai_1 _20033_ (.B1(_02901_),
    .Y(_00508_),
    .A1(net37),
    .A2(_02900_));
 sg13g2_nor2b_1 _20034_ (.A(net515),
    .B_N(\cpu.dcache.r_data[6][26] ),
    .Y(_02902_));
 sg13g2_a21oi_1 _20035_ (.A1(_02712_),
    .A2(net515),
    .Y(_02903_),
    .B1(_02902_));
 sg13g2_nand2_1 _20036_ (.Y(_02904_),
    .A(_12042_),
    .B(_02892_));
 sg13g2_o21ai_1 _20037_ (.B1(_02904_),
    .Y(_00509_),
    .A1(_02893_),
    .A2(_02903_));
 sg13g2_nor2b_1 _20038_ (.A(net515),
    .B_N(\cpu.dcache.r_data[6][27] ),
    .Y(_02905_));
 sg13g2_a21oi_1 _20039_ (.A1(_12611_),
    .A2(net515),
    .Y(_02906_),
    .B1(_02905_));
 sg13g2_nand2_1 _20040_ (.Y(_02907_),
    .A(_12051_),
    .B(_02892_));
 sg13g2_o21ai_1 _20041_ (.B1(_02907_),
    .Y(_00510_),
    .A1(_02893_),
    .A2(_02906_));
 sg13g2_nor2_1 _20042_ (.A(_02822_),
    .B(_12166_),
    .Y(_02908_));
 sg13g2_buf_2 _20043_ (.A(_02908_),
    .X(_02909_));
 sg13g2_nor2b_1 _20044_ (.A(_02909_),
    .B_N(\cpu.dcache.r_data[6][28] ),
    .Y(_02910_));
 sg13g2_a21oi_1 _20045_ (.A1(net1075),
    .A2(_02909_),
    .Y(_02911_),
    .B1(_02910_));
 sg13g2_nand2_1 _20046_ (.Y(_02912_),
    .A(_12063_),
    .B(_02892_));
 sg13g2_o21ai_1 _20047_ (.B1(_02912_),
    .Y(_00511_),
    .A1(net37),
    .A2(_02911_));
 sg13g2_nor2b_1 _20048_ (.A(_02909_),
    .B_N(\cpu.dcache.r_data[6][29] ),
    .Y(_02913_));
 sg13g2_a21oi_1 _20049_ (.A1(net1074),
    .A2(_02909_),
    .Y(_02914_),
    .B1(_02913_));
 sg13g2_nand2_1 _20050_ (.Y(_02915_),
    .A(_12073_),
    .B(_02892_));
 sg13g2_o21ai_1 _20051_ (.B1(_02915_),
    .Y(_00512_),
    .A1(net37),
    .A2(_02914_));
 sg13g2_mux2_1 _20052_ (.A0(\cpu.dcache.r_data[6][2] ),
    .A1(net1084),
    .S(_02829_),
    .X(_02916_));
 sg13g2_nor2_1 _20053_ (.A(_02826_),
    .B(_02916_),
    .Y(_02917_));
 sg13g2_a21oi_1 _20054_ (.A1(net753),
    .A2(net40),
    .Y(_00513_),
    .B1(_02917_));
 sg13g2_buf_2 _20055_ (.A(net1084),
    .X(_02918_));
 sg13g2_nor2b_1 _20056_ (.A(_02909_),
    .B_N(\cpu.dcache.r_data[6][30] ),
    .Y(_02919_));
 sg13g2_a21oi_1 _20057_ (.A1(net969),
    .A2(_02909_),
    .Y(_02920_),
    .B1(_02919_));
 sg13g2_nand2_1 _20058_ (.Y(_02921_),
    .A(_12080_),
    .B(_02892_));
 sg13g2_o21ai_1 _20059_ (.B1(_02921_),
    .Y(_00514_),
    .A1(net37),
    .A2(_02920_));
 sg13g2_nor2b_1 _20060_ (.A(_02909_),
    .B_N(\cpu.dcache.r_data[6][31] ),
    .Y(_02922_));
 sg13g2_a21oi_1 _20061_ (.A1(_12611_),
    .A2(_02909_),
    .Y(_02923_),
    .B1(_02922_));
 sg13g2_nand2_1 _20062_ (.Y(_02924_),
    .A(_12087_),
    .B(_02892_));
 sg13g2_o21ai_1 _20063_ (.B1(_02924_),
    .Y(_00515_),
    .A1(net37),
    .A2(_02923_));
 sg13g2_mux2_1 _20064_ (.A0(\cpu.dcache.r_data[6][3] ),
    .A1(net1083),
    .S(_02829_),
    .X(_02925_));
 sg13g2_nor2_1 _20065_ (.A(_02826_),
    .B(_02925_),
    .Y(_02926_));
 sg13g2_a21oi_1 _20066_ (.A1(net721),
    .A2(net40),
    .Y(_00516_),
    .B1(_02926_));
 sg13g2_nor2_1 _20067_ (.A(net642),
    .B(_12190_),
    .Y(_02927_));
 sg13g2_buf_2 _20068_ (.A(_02927_),
    .X(_02928_));
 sg13g2_mux2_1 _20069_ (.A0(\cpu.dcache.r_data[6][4] ),
    .A1(_12006_),
    .S(_02928_),
    .X(_02929_));
 sg13g2_nor2_1 _20070_ (.A(_02826_),
    .B(_02929_),
    .Y(_02930_));
 sg13g2_a21oi_1 _20071_ (.A1(net720),
    .A2(net40),
    .Y(_00517_),
    .B1(_02930_));
 sg13g2_nor2b_1 _20072_ (.A(_02928_),
    .B_N(\cpu.dcache.r_data[6][5] ),
    .Y(_02931_));
 sg13g2_a21oi_1 _20073_ (.A1(net1074),
    .A2(_02928_),
    .Y(_02932_),
    .B1(_02931_));
 sg13g2_nand2_1 _20074_ (.Y(_02933_),
    .A(net1021),
    .B(_02826_));
 sg13g2_o21ai_1 _20075_ (.B1(_02933_),
    .Y(_00518_),
    .A1(_02827_),
    .A2(_02932_));
 sg13g2_nor2b_1 _20076_ (.A(_02928_),
    .B_N(\cpu.dcache.r_data[6][6] ),
    .Y(_02934_));
 sg13g2_a21oi_1 _20077_ (.A1(net969),
    .A2(_02928_),
    .Y(_02935_),
    .B1(_02934_));
 sg13g2_nand2_1 _20078_ (.Y(_02936_),
    .A(net1020),
    .B(_02826_));
 sg13g2_o21ai_1 _20079_ (.B1(_02936_),
    .Y(_00519_),
    .A1(net40),
    .A2(_02935_));
 sg13g2_mux2_1 _20080_ (.A0(\cpu.dcache.r_data[6][7] ),
    .A1(net1083),
    .S(_02928_),
    .X(_02937_));
 sg13g2_nor2_1 _20081_ (.A(_02826_),
    .B(_02937_),
    .Y(_02938_));
 sg13g2_a21oi_1 _20082_ (.A1(net719),
    .A2(_02827_),
    .Y(_00520_),
    .B1(_02938_));
 sg13g2_nor2b_1 _20083_ (.A(_02838_),
    .B_N(\cpu.dcache.r_data[6][8] ),
    .Y(_02939_));
 sg13g2_a21oi_1 _20084_ (.A1(net1075),
    .A2(_02838_),
    .Y(_02940_),
    .B1(_02939_));
 sg13g2_nand2_1 _20085_ (.Y(_02941_),
    .A(_12148_),
    .B(_02835_));
 sg13g2_o21ai_1 _20086_ (.B1(_02941_),
    .Y(_00521_),
    .A1(net39),
    .A2(_02940_));
 sg13g2_nor2b_1 _20087_ (.A(_02838_),
    .B_N(\cpu.dcache.r_data[6][9] ),
    .Y(_02942_));
 sg13g2_a21oi_1 _20088_ (.A1(_02875_),
    .A2(_02838_),
    .Y(_02943_),
    .B1(_02942_));
 sg13g2_nand2_1 _20089_ (.Y(_02944_),
    .A(_12160_),
    .B(_02835_));
 sg13g2_o21ai_1 _20090_ (.B1(_02944_),
    .Y(_00522_),
    .A1(net39),
    .A2(_02943_));
 sg13g2_or2_1 _20091_ (.X(_02945_),
    .B(_11999_),
    .A(_09616_));
 sg13g2_buf_1 _20092_ (.A(_02945_),
    .X(_02946_));
 sg13g2_nor2_1 _20093_ (.A(_11987_),
    .B(_02946_),
    .Y(_02947_));
 sg13g2_buf_1 _20094_ (.A(_02947_),
    .X(_02948_));
 sg13g2_buf_1 _20095_ (.A(_02948_),
    .X(_02949_));
 sg13g2_nor2_1 _20096_ (.A(net672),
    .B(_12016_),
    .Y(_02950_));
 sg13g2_buf_2 _20097_ (.A(_02950_),
    .X(_02951_));
 sg13g2_nor2b_1 _20098_ (.A(_02951_),
    .B_N(\cpu.dcache.r_data[7][0] ),
    .Y(_02952_));
 sg13g2_a21oi_1 _20099_ (.A1(net1075),
    .A2(_02951_),
    .Y(_02953_),
    .B1(_02952_));
 sg13g2_nand2_1 _20100_ (.Y(_02954_),
    .A(_02832_),
    .B(_02949_));
 sg13g2_o21ai_1 _20101_ (.B1(_02954_),
    .Y(_00523_),
    .A1(_02949_),
    .A2(_02953_));
 sg13g2_nor2_1 _20102_ (.A(_12025_),
    .B(_02946_),
    .Y(_02955_));
 sg13g2_buf_2 _20103_ (.A(_02955_),
    .X(_02956_));
 sg13g2_buf_1 _20104_ (.A(_02956_),
    .X(_02957_));
 sg13g2_nor2_1 _20105_ (.A(net672),
    .B(_12033_),
    .Y(_02958_));
 sg13g2_buf_2 _20106_ (.A(_02958_),
    .X(_02959_));
 sg13g2_nor2b_1 _20107_ (.A(_02959_),
    .B_N(\cpu.dcache.r_data[7][10] ),
    .Y(_02960_));
 sg13g2_a21oi_1 _20108_ (.A1(net969),
    .A2(_02959_),
    .Y(_02961_),
    .B1(_02960_));
 sg13g2_nand2_1 _20109_ (.Y(_02962_),
    .A(_12042_),
    .B(_02957_));
 sg13g2_o21ai_1 _20110_ (.B1(_02962_),
    .Y(_00524_),
    .A1(net35),
    .A2(_02961_));
 sg13g2_buf_1 _20111_ (.A(_12046_),
    .X(_02963_));
 sg13g2_nor2b_1 _20112_ (.A(_02959_),
    .B_N(\cpu.dcache.r_data[7][11] ),
    .Y(_02964_));
 sg13g2_a21oi_1 _20113_ (.A1(net968),
    .A2(_02959_),
    .Y(_02965_),
    .B1(_02964_));
 sg13g2_nand2_1 _20114_ (.Y(_02966_),
    .A(_12051_),
    .B(net35));
 sg13g2_o21ai_1 _20115_ (.B1(_02966_),
    .Y(_00525_),
    .A1(_02957_),
    .A2(_02965_));
 sg13g2_nor2_1 _20116_ (.A(_09876_),
    .B(_12055_),
    .Y(_02967_));
 sg13g2_buf_2 _20117_ (.A(_02967_),
    .X(_02968_));
 sg13g2_nor2b_1 _20118_ (.A(_02968_),
    .B_N(\cpu.dcache.r_data[7][12] ),
    .Y(_02969_));
 sg13g2_a21oi_1 _20119_ (.A1(_02862_),
    .A2(_02968_),
    .Y(_02970_),
    .B1(_02969_));
 sg13g2_nand2_1 _20120_ (.Y(_02971_),
    .A(_12063_),
    .B(_02956_));
 sg13g2_o21ai_1 _20121_ (.B1(_02971_),
    .Y(_00526_),
    .A1(net35),
    .A2(_02970_));
 sg13g2_nor2b_1 _20122_ (.A(_02968_),
    .B_N(\cpu.dcache.r_data[7][13] ),
    .Y(_02972_));
 sg13g2_a21oi_1 _20123_ (.A1(_02875_),
    .A2(_02968_),
    .Y(_02973_),
    .B1(_02972_));
 sg13g2_nand2_1 _20124_ (.Y(_02974_),
    .A(_12073_),
    .B(_02956_));
 sg13g2_o21ai_1 _20125_ (.B1(_02974_),
    .Y(_00527_),
    .A1(net35),
    .A2(_02973_));
 sg13g2_nor2b_1 _20126_ (.A(_02968_),
    .B_N(\cpu.dcache.r_data[7][14] ),
    .Y(_02975_));
 sg13g2_a21oi_1 _20127_ (.A1(net969),
    .A2(_02968_),
    .Y(_02976_),
    .B1(_02975_));
 sg13g2_nand2_1 _20128_ (.Y(_02977_),
    .A(_12080_),
    .B(_02956_));
 sg13g2_o21ai_1 _20129_ (.B1(_02977_),
    .Y(_00528_),
    .A1(net35),
    .A2(_02976_));
 sg13g2_nor2b_1 _20130_ (.A(_02968_),
    .B_N(\cpu.dcache.r_data[7][15] ),
    .Y(_02978_));
 sg13g2_a21oi_1 _20131_ (.A1(net968),
    .A2(_02968_),
    .Y(_02979_),
    .B1(_02978_));
 sg13g2_nand2_1 _20132_ (.Y(_02980_),
    .A(_12087_),
    .B(_02956_));
 sg13g2_o21ai_1 _20133_ (.B1(_02980_),
    .Y(_00529_),
    .A1(net35),
    .A2(_02979_));
 sg13g2_nor2_1 _20134_ (.A(_12090_),
    .B(_02946_),
    .Y(_02981_));
 sg13g2_buf_1 _20135_ (.A(_02981_),
    .X(_02982_));
 sg13g2_buf_1 _20136_ (.A(_02982_),
    .X(_02983_));
 sg13g2_nor2_1 _20137_ (.A(net672),
    .B(_12096_),
    .Y(_02984_));
 sg13g2_buf_2 _20138_ (.A(_02984_),
    .X(_02985_));
 sg13g2_nor2b_1 _20139_ (.A(_02985_),
    .B_N(\cpu.dcache.r_data[7][16] ),
    .Y(_02986_));
 sg13g2_a21oi_1 _20140_ (.A1(net1075),
    .A2(_02985_),
    .Y(_02987_),
    .B1(_02986_));
 sg13g2_nand2_1 _20141_ (.Y(_02988_),
    .A(net970),
    .B(net34));
 sg13g2_o21ai_1 _20142_ (.B1(_02988_),
    .Y(_00530_),
    .A1(_02983_),
    .A2(_02987_));
 sg13g2_nor2b_1 _20143_ (.A(_02985_),
    .B_N(\cpu.dcache.r_data[7][17] ),
    .Y(_02989_));
 sg13g2_a21oi_1 _20144_ (.A1(net1074),
    .A2(_02985_),
    .Y(_02990_),
    .B1(_02989_));
 sg13g2_nand2_1 _20145_ (.Y(_02991_),
    .A(net850),
    .B(net34));
 sg13g2_o21ai_1 _20146_ (.B1(_02991_),
    .Y(_00531_),
    .A1(net34),
    .A2(_02990_));
 sg13g2_mux2_1 _20147_ (.A0(\cpu.dcache.r_data[7][18] ),
    .A1(net1084),
    .S(_02985_),
    .X(_02992_));
 sg13g2_nor2_1 _20148_ (.A(_02982_),
    .B(_02992_),
    .Y(_02993_));
 sg13g2_a21oi_1 _20149_ (.A1(net753),
    .A2(_02983_),
    .Y(_00532_),
    .B1(_02993_));
 sg13g2_mux2_1 _20150_ (.A0(\cpu.dcache.r_data[7][19] ),
    .A1(net1083),
    .S(_02985_),
    .X(_02994_));
 sg13g2_nor2_1 _20151_ (.A(_02982_),
    .B(_02994_),
    .Y(_02995_));
 sg13g2_a21oi_1 _20152_ (.A1(net721),
    .A2(net34),
    .Y(_00533_),
    .B1(_02995_));
 sg13g2_nor2b_1 _20153_ (.A(_02951_),
    .B_N(\cpu.dcache.r_data[7][1] ),
    .Y(_02996_));
 sg13g2_a21oi_1 _20154_ (.A1(net1074),
    .A2(_02951_),
    .Y(_02997_),
    .B1(_02996_));
 sg13g2_nand2_1 _20155_ (.Y(_02998_),
    .A(net1018),
    .B(net36));
 sg13g2_o21ai_1 _20156_ (.B1(_02998_),
    .Y(_00534_),
    .A1(net36),
    .A2(_02997_));
 sg13g2_or2_1 _20157_ (.X(_02999_),
    .B(_12125_),
    .A(net672));
 sg13g2_buf_1 _20158_ (.A(_02999_),
    .X(_03000_));
 sg13g2_mux2_1 _20159_ (.A0(net1079),
    .A1(\cpu.dcache.r_data[7][20] ),
    .S(_03000_),
    .X(_03001_));
 sg13g2_nor2_1 _20160_ (.A(_02982_),
    .B(_03001_),
    .Y(_03002_));
 sg13g2_a21oi_1 _20161_ (.A1(_02755_),
    .A2(net34),
    .Y(_00535_),
    .B1(_03002_));
 sg13g2_mux2_1 _20162_ (.A0(net1082),
    .A1(\cpu.dcache.r_data[7][21] ),
    .S(_03000_),
    .X(_03003_));
 sg13g2_mux2_1 _20163_ (.A0(_03003_),
    .A1(_12132_),
    .S(net34),
    .X(_00536_));
 sg13g2_mux2_1 _20164_ (.A0(net1081),
    .A1(\cpu.dcache.r_data[7][22] ),
    .S(_03000_),
    .X(_03004_));
 sg13g2_mux2_1 _20165_ (.A0(_03004_),
    .A1(net974),
    .S(net34),
    .X(_00537_));
 sg13g2_mux2_1 _20166_ (.A0(net1080),
    .A1(\cpu.dcache.r_data[7][23] ),
    .S(_03000_),
    .X(_03005_));
 sg13g2_nor2_1 _20167_ (.A(_02982_),
    .B(_03005_),
    .Y(_03006_));
 sg13g2_a21oi_1 _20168_ (.A1(net719),
    .A2(net34),
    .Y(_00538_),
    .B1(_03006_));
 sg13g2_nor2_1 _20169_ (.A(_12153_),
    .B(_02946_),
    .Y(_03007_));
 sg13g2_buf_2 _20170_ (.A(_03007_),
    .X(_03008_));
 sg13g2_buf_1 _20171_ (.A(_03008_),
    .X(_03009_));
 sg13g2_nor2_1 _20172_ (.A(net672),
    .B(_11995_),
    .Y(_03010_));
 sg13g2_buf_1 _20173_ (.A(_03010_),
    .X(_03011_));
 sg13g2_nor2b_1 _20174_ (.A(net514),
    .B_N(\cpu.dcache.r_data[7][24] ),
    .Y(_03012_));
 sg13g2_a21oi_1 _20175_ (.A1(net1075),
    .A2(net514),
    .Y(_03013_),
    .B1(_03012_));
 sg13g2_nand2_1 _20176_ (.Y(_03014_),
    .A(_12148_),
    .B(net33));
 sg13g2_o21ai_1 _20177_ (.B1(_03014_),
    .Y(_00539_),
    .A1(net33),
    .A2(_03013_));
 sg13g2_nor2b_1 _20178_ (.A(net514),
    .B_N(\cpu.dcache.r_data[7][25] ),
    .Y(_03015_));
 sg13g2_a21oi_1 _20179_ (.A1(net1074),
    .A2(net514),
    .Y(_03016_),
    .B1(_03015_));
 sg13g2_nand2_1 _20180_ (.Y(_03017_),
    .A(_12160_),
    .B(net33));
 sg13g2_o21ai_1 _20181_ (.B1(_03017_),
    .Y(_00540_),
    .A1(_03009_),
    .A2(_03016_));
 sg13g2_nor2b_1 _20182_ (.A(net514),
    .B_N(\cpu.dcache.r_data[7][26] ),
    .Y(_03018_));
 sg13g2_a21oi_1 _20183_ (.A1(net969),
    .A2(net514),
    .Y(_03019_),
    .B1(_03018_));
 sg13g2_nand2_1 _20184_ (.Y(_03020_),
    .A(_12042_),
    .B(_03008_));
 sg13g2_o21ai_1 _20185_ (.B1(_03020_),
    .Y(_00541_),
    .A1(_03009_),
    .A2(_03019_));
 sg13g2_nor2b_1 _20186_ (.A(net514),
    .B_N(\cpu.dcache.r_data[7][27] ),
    .Y(_03021_));
 sg13g2_a21oi_1 _20187_ (.A1(net968),
    .A2(net514),
    .Y(_03022_),
    .B1(_03021_));
 sg13g2_nand2_1 _20188_ (.Y(_03023_),
    .A(_12051_),
    .B(_03008_));
 sg13g2_o21ai_1 _20189_ (.B1(_03023_),
    .Y(_00542_),
    .A1(net33),
    .A2(_03022_));
 sg13g2_nor2_1 _20190_ (.A(_09876_),
    .B(_12166_),
    .Y(_03024_));
 sg13g2_buf_2 _20191_ (.A(_03024_),
    .X(_03025_));
 sg13g2_nor2b_1 _20192_ (.A(_03025_),
    .B_N(\cpu.dcache.r_data[7][28] ),
    .Y(_03026_));
 sg13g2_a21oi_1 _20193_ (.A1(net1075),
    .A2(_03025_),
    .Y(_03027_),
    .B1(_03026_));
 sg13g2_nand2_1 _20194_ (.Y(_03028_),
    .A(_12063_),
    .B(_03008_));
 sg13g2_o21ai_1 _20195_ (.B1(_03028_),
    .Y(_00543_),
    .A1(net33),
    .A2(_03027_));
 sg13g2_buf_2 _20196_ (.A(_12065_),
    .X(_03029_));
 sg13g2_nor2b_1 _20197_ (.A(_03025_),
    .B_N(\cpu.dcache.r_data[7][29] ),
    .Y(_03030_));
 sg13g2_a21oi_1 _20198_ (.A1(_03029_),
    .A2(_03025_),
    .Y(_03031_),
    .B1(_03030_));
 sg13g2_nand2_1 _20199_ (.Y(_03032_),
    .A(_12073_),
    .B(_03008_));
 sg13g2_o21ai_1 _20200_ (.B1(_03032_),
    .Y(_00544_),
    .A1(net33),
    .A2(_03031_));
 sg13g2_mux2_1 _20201_ (.A0(\cpu.dcache.r_data[7][2] ),
    .A1(net1084),
    .S(_02951_),
    .X(_03033_));
 sg13g2_nor2_1 _20202_ (.A(_02948_),
    .B(_03033_),
    .Y(_03034_));
 sg13g2_a21oi_1 _20203_ (.A1(_09884_),
    .A2(net36),
    .Y(_00545_),
    .B1(_03034_));
 sg13g2_nor2b_1 _20204_ (.A(_03025_),
    .B_N(\cpu.dcache.r_data[7][30] ),
    .Y(_03035_));
 sg13g2_a21oi_1 _20205_ (.A1(net969),
    .A2(_03025_),
    .Y(_03036_),
    .B1(_03035_));
 sg13g2_nand2_1 _20206_ (.Y(_03037_),
    .A(_12080_),
    .B(_03008_));
 sg13g2_o21ai_1 _20207_ (.B1(_03037_),
    .Y(_00546_),
    .A1(net33),
    .A2(_03036_));
 sg13g2_nor2b_1 _20208_ (.A(_03025_),
    .B_N(\cpu.dcache.r_data[7][31] ),
    .Y(_03038_));
 sg13g2_a21oi_1 _20209_ (.A1(net968),
    .A2(_03025_),
    .Y(_03039_),
    .B1(_03038_));
 sg13g2_nand2_1 _20210_ (.Y(_03040_),
    .A(_12087_),
    .B(_03008_));
 sg13g2_o21ai_1 _20211_ (.B1(_03040_),
    .Y(_00547_),
    .A1(net33),
    .A2(_03039_));
 sg13g2_mux2_1 _20212_ (.A0(\cpu.dcache.r_data[7][3] ),
    .A1(_12046_),
    .S(_02951_),
    .X(_03041_));
 sg13g2_nor2_1 _20213_ (.A(_02948_),
    .B(_03041_),
    .Y(_03042_));
 sg13g2_a21oi_1 _20214_ (.A1(net721),
    .A2(net36),
    .Y(_00548_),
    .B1(_03042_));
 sg13g2_or2_1 _20215_ (.X(_03043_),
    .B(_12190_),
    .A(net672));
 sg13g2_buf_1 _20216_ (.A(_03043_),
    .X(_03044_));
 sg13g2_mux2_1 _20217_ (.A0(_12122_),
    .A1(\cpu.dcache.r_data[7][4] ),
    .S(_03044_),
    .X(_03045_));
 sg13g2_nor2_1 _20218_ (.A(_02948_),
    .B(_03045_),
    .Y(_03046_));
 sg13g2_a21oi_1 _20219_ (.A1(net720),
    .A2(net36),
    .Y(_00549_),
    .B1(_03046_));
 sg13g2_mux2_1 _20220_ (.A0(net1082),
    .A1(\cpu.dcache.r_data[7][5] ),
    .S(_03044_),
    .X(_03047_));
 sg13g2_mux2_1 _20221_ (.A0(_03047_),
    .A1(net986),
    .S(net36),
    .X(_00550_));
 sg13g2_mux2_1 _20222_ (.A0(net1081),
    .A1(\cpu.dcache.r_data[7][6] ),
    .S(_03044_),
    .X(_03048_));
 sg13g2_mux2_1 _20223_ (.A0(_03048_),
    .A1(net974),
    .S(net36),
    .X(_00551_));
 sg13g2_mux2_1 _20224_ (.A0(net1080),
    .A1(\cpu.dcache.r_data[7][7] ),
    .S(_03044_),
    .X(_03049_));
 sg13g2_nor2_1 _20225_ (.A(_02948_),
    .B(_03049_),
    .Y(_03050_));
 sg13g2_a21oi_1 _20226_ (.A1(_02766_),
    .A2(net36),
    .Y(_00552_),
    .B1(_03050_));
 sg13g2_nor2b_1 _20227_ (.A(_02959_),
    .B_N(\cpu.dcache.r_data[7][8] ),
    .Y(_03051_));
 sg13g2_a21oi_1 _20228_ (.A1(_02862_),
    .A2(_02959_),
    .Y(_03052_),
    .B1(_03051_));
 sg13g2_nand2_1 _20229_ (.Y(_03053_),
    .A(_12148_),
    .B(_02956_));
 sg13g2_o21ai_1 _20230_ (.B1(_03053_),
    .Y(_00553_),
    .A1(net35),
    .A2(_03052_));
 sg13g2_nor2b_1 _20231_ (.A(_02959_),
    .B_N(\cpu.dcache.r_data[7][9] ),
    .Y(_03054_));
 sg13g2_a21oi_1 _20232_ (.A1(_03029_),
    .A2(_02959_),
    .Y(_03055_),
    .B1(_03054_));
 sg13g2_nand2_1 _20233_ (.Y(_03056_),
    .A(_12160_),
    .B(_02956_));
 sg13g2_o21ai_1 _20234_ (.B1(_03056_),
    .Y(_00554_),
    .A1(net35),
    .A2(_03055_));
 sg13g2_buf_1 _20235_ (.A(_08181_),
    .X(_03057_));
 sg13g2_buf_1 _20236_ (.A(\cpu.d_rstrobe_d ),
    .X(_03058_));
 sg13g2_nor2_1 _20237_ (.A(_03057_),
    .B(_03058_),
    .Y(_03059_));
 sg13g2_nand3_1 _20238_ (.B(_11996_),
    .C(_03059_),
    .A(_12009_),
    .Y(_03060_));
 sg13g2_o21ai_1 _20239_ (.B1(_03060_),
    .Y(_03061_),
    .A1(_11524_),
    .A2(_11997_));
 sg13g2_buf_2 _20240_ (.A(_03061_),
    .X(_03062_));
 sg13g2_xor2_1 _20241_ (.B(_12009_),
    .A(_03058_),
    .X(_03063_));
 sg13g2_nand3_1 _20242_ (.B(_11993_),
    .C(_03063_),
    .A(net987),
    .Y(_03064_));
 sg13g2_o21ai_1 _20243_ (.B1(_03064_),
    .Y(_03065_),
    .A1(_11524_),
    .A2(_11997_));
 sg13g2_buf_2 _20244_ (.A(_03065_),
    .X(_03066_));
 sg13g2_nor2b_1 _20245_ (.A(net519),
    .B_N(_03066_),
    .Y(_03067_));
 sg13g2_mux2_1 _20246_ (.A0(\cpu.dcache.r_dirty[0] ),
    .A1(_03062_),
    .S(_03067_),
    .X(_00555_));
 sg13g2_buf_1 _20247_ (.A(net605),
    .X(_03068_));
 sg13g2_buf_1 _20248_ (.A(net513),
    .X(_03069_));
 sg13g2_buf_1 _20249_ (.A(net455),
    .X(_03070_));
 sg13g2_nand2_1 _20250_ (.Y(_03071_),
    .A(_03070_),
    .B(_03066_));
 sg13g2_mux2_1 _20251_ (.A0(_03062_),
    .A1(\cpu.dcache.r_dirty[1] ),
    .S(_03071_),
    .X(_00556_));
 sg13g2_buf_1 _20252_ (.A(net602),
    .X(_03072_));
 sg13g2_buf_1 _20253_ (.A(net512),
    .X(_03073_));
 sg13g2_nand2_1 _20254_ (.Y(_03074_),
    .A(_03073_),
    .B(_03066_));
 sg13g2_mux2_1 _20255_ (.A0(_03062_),
    .A1(\cpu.dcache.r_dirty[2] ),
    .S(_03074_),
    .X(_00557_));
 sg13g2_buf_1 _20256_ (.A(net681),
    .X(_03075_));
 sg13g2_buf_1 _20257_ (.A(net582),
    .X(_03076_));
 sg13g2_nand2_1 _20258_ (.Y(_03077_),
    .A(_03076_),
    .B(_03066_));
 sg13g2_mux2_1 _20259_ (.A0(_03062_),
    .A1(\cpu.dcache.r_dirty[3] ),
    .S(_03077_),
    .X(_00558_));
 sg13g2_nand2_1 _20260_ (.Y(_03078_),
    .A(net463),
    .B(_03066_));
 sg13g2_mux2_1 _20261_ (.A0(_03062_),
    .A1(\cpu.dcache.r_dirty[4] ),
    .S(_03078_),
    .X(_00559_));
 sg13g2_buf_1 _20262_ (.A(_09273_),
    .X(_03079_));
 sg13g2_buf_1 _20263_ (.A(net581),
    .X(_03080_));
 sg13g2_buf_1 _20264_ (.A(_03080_),
    .X(_03081_));
 sg13g2_nand2_1 _20265_ (.Y(_03082_),
    .A(_03081_),
    .B(_03066_));
 sg13g2_mux2_1 _20266_ (.A0(_03062_),
    .A1(\cpu.dcache.r_dirty[5] ),
    .S(_03082_),
    .X(_00560_));
 sg13g2_buf_1 _20267_ (.A(_09420_),
    .X(_03083_));
 sg13g2_buf_1 _20268_ (.A(net580),
    .X(_03084_));
 sg13g2_nand2_1 _20269_ (.Y(_03085_),
    .A(_03084_),
    .B(_03066_));
 sg13g2_mux2_1 _20270_ (.A0(_03062_),
    .A1(\cpu.dcache.r_dirty[6] ),
    .S(_03085_),
    .X(_00561_));
 sg13g2_nand2_1 _20271_ (.Y(_03086_),
    .A(net530),
    .B(_03066_));
 sg13g2_mux2_1 _20272_ (.A0(_03062_),
    .A1(\cpu.dcache.r_dirty[7] ),
    .S(_03086_),
    .X(_00562_));
 sg13g2_buf_1 _20273_ (.A(_10473_),
    .X(_03087_));
 sg13g2_buf_1 _20274_ (.A(net848),
    .X(_03088_));
 sg13g2_buf_1 _20275_ (.A(_03088_),
    .X(_03089_));
 sg13g2_buf_1 _20276_ (.A(_12145_),
    .X(_03090_));
 sg13g2_buf_1 _20277_ (.A(_12145_),
    .X(_03091_));
 sg13g2_nand2_1 _20278_ (.Y(_03092_),
    .A(\cpu.dcache.r_tag[0][5] ),
    .B(net364));
 sg13g2_o21ai_1 _20279_ (.B1(_03092_),
    .Y(_00566_),
    .A1(_03089_),
    .A2(net365));
 sg13g2_mux2_1 _20280_ (.A0(net427),
    .A1(\cpu.dcache.r_tag[0][15] ),
    .S(net365),
    .X(_00567_));
 sg13g2_mux2_1 _20281_ (.A0(net432),
    .A1(\cpu.dcache.r_tag[0][16] ),
    .S(net365),
    .X(_00568_));
 sg13g2_mux2_1 _20282_ (.A0(net428),
    .A1(\cpu.dcache.r_tag[0][17] ),
    .S(_03090_),
    .X(_00569_));
 sg13g2_mux2_1 _20283_ (.A0(net431),
    .A1(\cpu.dcache.r_tag[0][18] ),
    .S(net365),
    .X(_00570_));
 sg13g2_mux2_1 _20284_ (.A0(net424),
    .A1(\cpu.dcache.r_tag[0][19] ),
    .S(net365),
    .X(_00571_));
 sg13g2_mux2_1 _20285_ (.A0(net425),
    .A1(\cpu.dcache.r_tag[0][20] ),
    .S(_03090_),
    .X(_00572_));
 sg13g2_mux2_1 _20286_ (.A0(net426),
    .A1(\cpu.dcache.r_tag[0][21] ),
    .S(net365),
    .X(_00573_));
 sg13g2_mux2_1 _20287_ (.A0(net430),
    .A1(\cpu.dcache.r_tag[0][22] ),
    .S(net365),
    .X(_00574_));
 sg13g2_mux2_1 _20288_ (.A0(_09687_),
    .A1(\cpu.dcache.r_tag[0][23] ),
    .S(net365),
    .X(_00575_));
 sg13g2_buf_2 _20289_ (.A(_09023_),
    .X(_03093_));
 sg13g2_buf_1 _20290_ (.A(net966),
    .X(_03094_));
 sg13g2_buf_1 _20291_ (.A(net847),
    .X(_03095_));
 sg13g2_mux2_1 _20292_ (.A0(net717),
    .A1(\cpu.dcache.r_tag[0][6] ),
    .S(_03091_),
    .X(_00576_));
 sg13g2_buf_2 _20293_ (.A(_09026_),
    .X(_03096_));
 sg13g2_buf_1 _20294_ (.A(net965),
    .X(_03097_));
 sg13g2_buf_1 _20295_ (.A(net846),
    .X(_03098_));
 sg13g2_mux2_1 _20296_ (.A0(net716),
    .A1(\cpu.dcache.r_tag[0][7] ),
    .S(net364),
    .X(_00577_));
 sg13g2_buf_1 _20297_ (.A(net1037),
    .X(_03099_));
 sg13g2_buf_1 _20298_ (.A(net845),
    .X(_03100_));
 sg13g2_mux2_1 _20299_ (.A0(net715),
    .A1(\cpu.dcache.r_tag[0][8] ),
    .S(net364),
    .X(_00578_));
 sg13g2_buf_1 _20300_ (.A(_10831_),
    .X(_03101_));
 sg13g2_buf_1 _20301_ (.A(net964),
    .X(_03102_));
 sg13g2_mux2_1 _20302_ (.A0(net844),
    .A1(\cpu.dcache.r_tag[0][9] ),
    .S(_03091_),
    .X(_00579_));
 sg13g2_buf_1 _20303_ (.A(net1095),
    .X(_03103_));
 sg13g2_buf_1 _20304_ (.A(net963),
    .X(_03104_));
 sg13g2_mux2_1 _20305_ (.A0(net843),
    .A1(\cpu.dcache.r_tag[0][10] ),
    .S(net364),
    .X(_00580_));
 sg13g2_buf_1 _20306_ (.A(_10907_),
    .X(_03105_));
 sg13g2_buf_1 _20307_ (.A(net962),
    .X(_03106_));
 sg13g2_mux2_1 _20308_ (.A0(net842),
    .A1(\cpu.dcache.r_tag[0][11] ),
    .S(net364),
    .X(_00581_));
 sg13g2_mux2_1 _20309_ (.A0(net376),
    .A1(\cpu.dcache.r_tag[0][12] ),
    .S(net364),
    .X(_00582_));
 sg13g2_mux2_1 _20310_ (.A0(net377),
    .A1(\cpu.dcache.r_tag[0][13] ),
    .S(net364),
    .X(_00583_));
 sg13g2_mux2_1 _20311_ (.A0(net429),
    .A1(\cpu.dcache.r_tag[0][14] ),
    .S(net364),
    .X(_00584_));
 sg13g2_buf_2 _20312_ (.A(net727),
    .X(_03107_));
 sg13g2_buf_2 _20313_ (.A(net640),
    .X(_03108_));
 sg13g2_buf_1 _20314_ (.A(net579),
    .X(_03109_));
 sg13g2_buf_1 _20315_ (.A(_12286_),
    .X(_03110_));
 sg13g2_mux2_1 _20316_ (.A0(\cpu.dcache.r_tag[1][5] ),
    .A1(net508),
    .S(net295),
    .X(_00585_));
 sg13g2_mux2_1 _20317_ (.A0(\cpu.dcache.r_tag[1][15] ),
    .A1(net427),
    .S(net295),
    .X(_00586_));
 sg13g2_mux2_1 _20318_ (.A0(\cpu.dcache.r_tag[1][16] ),
    .A1(net432),
    .S(net295),
    .X(_00587_));
 sg13g2_mux2_1 _20319_ (.A0(\cpu.dcache.r_tag[1][17] ),
    .A1(net428),
    .S(_03110_),
    .X(_00588_));
 sg13g2_mux2_1 _20320_ (.A0(\cpu.dcache.r_tag[1][18] ),
    .A1(net431),
    .S(net295),
    .X(_00589_));
 sg13g2_mux2_1 _20321_ (.A0(\cpu.dcache.r_tag[1][19] ),
    .A1(net424),
    .S(net295),
    .X(_00590_));
 sg13g2_mux2_1 _20322_ (.A0(\cpu.dcache.r_tag[1][20] ),
    .A1(net425),
    .S(_03110_),
    .X(_00591_));
 sg13g2_mux2_1 _20323_ (.A0(\cpu.dcache.r_tag[1][21] ),
    .A1(net426),
    .S(net295),
    .X(_00592_));
 sg13g2_mux2_1 _20324_ (.A0(\cpu.dcache.r_tag[1][22] ),
    .A1(net430),
    .S(net295),
    .X(_00593_));
 sg13g2_mux2_1 _20325_ (.A0(\cpu.dcache.r_tag[1][23] ),
    .A1(net375),
    .S(net295),
    .X(_00594_));
 sg13g2_buf_1 _20326_ (.A(net847),
    .X(_03111_));
 sg13g2_buf_1 _20327_ (.A(_12286_),
    .X(_03112_));
 sg13g2_mux2_1 _20328_ (.A0(\cpu.dcache.r_tag[1][6] ),
    .A1(net714),
    .S(net294),
    .X(_00595_));
 sg13g2_buf_1 _20329_ (.A(net846),
    .X(_03113_));
 sg13g2_mux2_1 _20330_ (.A0(\cpu.dcache.r_tag[1][7] ),
    .A1(net713),
    .S(net294),
    .X(_00596_));
 sg13g2_buf_1 _20331_ (.A(net845),
    .X(_03114_));
 sg13g2_mux2_1 _20332_ (.A0(\cpu.dcache.r_tag[1][8] ),
    .A1(net712),
    .S(net294),
    .X(_00597_));
 sg13g2_buf_1 _20333_ (.A(net964),
    .X(_03115_));
 sg13g2_mux2_1 _20334_ (.A0(\cpu.dcache.r_tag[1][9] ),
    .A1(net841),
    .S(net294),
    .X(_00598_));
 sg13g2_buf_1 _20335_ (.A(net963),
    .X(_03116_));
 sg13g2_mux2_1 _20336_ (.A0(\cpu.dcache.r_tag[1][10] ),
    .A1(net840),
    .S(_03112_),
    .X(_00599_));
 sg13g2_buf_1 _20337_ (.A(net962),
    .X(_03117_));
 sg13g2_mux2_1 _20338_ (.A0(\cpu.dcache.r_tag[1][11] ),
    .A1(net839),
    .S(_03112_),
    .X(_00600_));
 sg13g2_mux2_1 _20339_ (.A0(\cpu.dcache.r_tag[1][12] ),
    .A1(_09502_),
    .S(net294),
    .X(_00601_));
 sg13g2_mux2_1 _20340_ (.A0(\cpu.dcache.r_tag[1][13] ),
    .A1(net377),
    .S(net294),
    .X(_00602_));
 sg13g2_mux2_1 _20341_ (.A0(\cpu.dcache.r_tag[1][14] ),
    .A1(_09329_),
    .S(net294),
    .X(_00603_));
 sg13g2_buf_1 _20342_ (.A(_12409_),
    .X(_03118_));
 sg13g2_mux2_1 _20343_ (.A0(\cpu.dcache.r_tag[2][5] ),
    .A1(net508),
    .S(net363),
    .X(_00604_));
 sg13g2_mux2_1 _20344_ (.A0(\cpu.dcache.r_tag[2][15] ),
    .A1(net427),
    .S(_03118_),
    .X(_00605_));
 sg13g2_mux2_1 _20345_ (.A0(\cpu.dcache.r_tag[2][16] ),
    .A1(net432),
    .S(net363),
    .X(_00606_));
 sg13g2_mux2_1 _20346_ (.A0(\cpu.dcache.r_tag[2][17] ),
    .A1(net428),
    .S(_03118_),
    .X(_00607_));
 sg13g2_mux2_1 _20347_ (.A0(\cpu.dcache.r_tag[2][18] ),
    .A1(net431),
    .S(net363),
    .X(_00608_));
 sg13g2_mux2_1 _20348_ (.A0(\cpu.dcache.r_tag[2][19] ),
    .A1(net424),
    .S(net363),
    .X(_00609_));
 sg13g2_mux2_1 _20349_ (.A0(\cpu.dcache.r_tag[2][20] ),
    .A1(net425),
    .S(net363),
    .X(_00610_));
 sg13g2_mux2_1 _20350_ (.A0(\cpu.dcache.r_tag[2][21] ),
    .A1(net426),
    .S(net363),
    .X(_00611_));
 sg13g2_mux2_1 _20351_ (.A0(\cpu.dcache.r_tag[2][22] ),
    .A1(net430),
    .S(net363),
    .X(_00612_));
 sg13g2_mux2_1 _20352_ (.A0(\cpu.dcache.r_tag[2][23] ),
    .A1(net375),
    .S(net363),
    .X(_00613_));
 sg13g2_buf_1 _20353_ (.A(_12409_),
    .X(_03119_));
 sg13g2_mux2_1 _20354_ (.A0(\cpu.dcache.r_tag[2][6] ),
    .A1(net714),
    .S(net362),
    .X(_00614_));
 sg13g2_mux2_1 _20355_ (.A0(\cpu.dcache.r_tag[2][7] ),
    .A1(net713),
    .S(net362),
    .X(_00615_));
 sg13g2_mux2_1 _20356_ (.A0(\cpu.dcache.r_tag[2][8] ),
    .A1(net712),
    .S(net362),
    .X(_00616_));
 sg13g2_mux2_1 _20357_ (.A0(\cpu.dcache.r_tag[2][9] ),
    .A1(net841),
    .S(net362),
    .X(_00617_));
 sg13g2_mux2_1 _20358_ (.A0(\cpu.dcache.r_tag[2][10] ),
    .A1(net840),
    .S(net362),
    .X(_00618_));
 sg13g2_mux2_1 _20359_ (.A0(\cpu.dcache.r_tag[2][11] ),
    .A1(net839),
    .S(_03119_),
    .X(_00619_));
 sg13g2_mux2_1 _20360_ (.A0(\cpu.dcache.r_tag[2][12] ),
    .A1(net376),
    .S(net362),
    .X(_00620_));
 sg13g2_mux2_1 _20361_ (.A0(\cpu.dcache.r_tag[2][13] ),
    .A1(net377),
    .S(net362),
    .X(_00621_));
 sg13g2_mux2_1 _20362_ (.A0(\cpu.dcache.r_tag[2][14] ),
    .A1(net429),
    .S(_03119_),
    .X(_00622_));
 sg13g2_buf_1 _20363_ (.A(_12530_),
    .X(_03120_));
 sg13g2_mux2_1 _20364_ (.A0(\cpu.dcache.r_tag[3][5] ),
    .A1(net508),
    .S(_03120_),
    .X(_00623_));
 sg13g2_mux2_1 _20365_ (.A0(\cpu.dcache.r_tag[3][15] ),
    .A1(net427),
    .S(net222),
    .X(_00624_));
 sg13g2_mux2_1 _20366_ (.A0(\cpu.dcache.r_tag[3][16] ),
    .A1(net432),
    .S(_03120_),
    .X(_00625_));
 sg13g2_mux2_1 _20367_ (.A0(\cpu.dcache.r_tag[3][17] ),
    .A1(net428),
    .S(net222),
    .X(_00626_));
 sg13g2_mux2_1 _20368_ (.A0(\cpu.dcache.r_tag[3][18] ),
    .A1(net431),
    .S(net222),
    .X(_00627_));
 sg13g2_mux2_1 _20369_ (.A0(\cpu.dcache.r_tag[3][19] ),
    .A1(net424),
    .S(net222),
    .X(_00628_));
 sg13g2_mux2_1 _20370_ (.A0(\cpu.dcache.r_tag[3][20] ),
    .A1(net425),
    .S(net222),
    .X(_00629_));
 sg13g2_mux2_1 _20371_ (.A0(\cpu.dcache.r_tag[3][21] ),
    .A1(net426),
    .S(net222),
    .X(_00630_));
 sg13g2_mux2_1 _20372_ (.A0(\cpu.dcache.r_tag[3][22] ),
    .A1(net430),
    .S(net222),
    .X(_00631_));
 sg13g2_mux2_1 _20373_ (.A0(\cpu.dcache.r_tag[3][23] ),
    .A1(net375),
    .S(net222),
    .X(_00632_));
 sg13g2_buf_1 _20374_ (.A(_12530_),
    .X(_03121_));
 sg13g2_mux2_1 _20375_ (.A0(\cpu.dcache.r_tag[3][6] ),
    .A1(net714),
    .S(net221),
    .X(_00633_));
 sg13g2_mux2_1 _20376_ (.A0(\cpu.dcache.r_tag[3][7] ),
    .A1(net713),
    .S(net221),
    .X(_00634_));
 sg13g2_mux2_1 _20377_ (.A0(\cpu.dcache.r_tag[3][8] ),
    .A1(_03114_),
    .S(_03121_),
    .X(_00635_));
 sg13g2_mux2_1 _20378_ (.A0(\cpu.dcache.r_tag[3][9] ),
    .A1(net841),
    .S(net221),
    .X(_00636_));
 sg13g2_mux2_1 _20379_ (.A0(\cpu.dcache.r_tag[3][10] ),
    .A1(net840),
    .S(_03121_),
    .X(_00637_));
 sg13g2_mux2_1 _20380_ (.A0(\cpu.dcache.r_tag[3][11] ),
    .A1(net839),
    .S(net221),
    .X(_00638_));
 sg13g2_mux2_1 _20381_ (.A0(\cpu.dcache.r_tag[3][12] ),
    .A1(net376),
    .S(net221),
    .X(_00639_));
 sg13g2_mux2_1 _20382_ (.A0(\cpu.dcache.r_tag[3][13] ),
    .A1(net377),
    .S(net221),
    .X(_00640_));
 sg13g2_mux2_1 _20383_ (.A0(\cpu.dcache.r_tag[3][14] ),
    .A1(net429),
    .S(net221),
    .X(_00641_));
 sg13g2_buf_1 _20384_ (.A(_12646_),
    .X(_03122_));
 sg13g2_nand2_1 _20385_ (.Y(_03123_),
    .A(\cpu.dcache.r_tag[4][5] ),
    .B(_12646_));
 sg13g2_o21ai_1 _20386_ (.B1(_03123_),
    .Y(_00642_),
    .A1(_03089_),
    .A2(net412));
 sg13g2_mux2_1 _20387_ (.A0(_09399_),
    .A1(\cpu.dcache.r_tag[4][15] ),
    .S(net412),
    .X(_00643_));
 sg13g2_mux2_1 _20388_ (.A0(net432),
    .A1(\cpu.dcache.r_tag[4][16] ),
    .S(_03122_),
    .X(_00644_));
 sg13g2_mux2_1 _20389_ (.A0(_09362_),
    .A1(\cpu.dcache.r_tag[4][17] ),
    .S(_03122_),
    .X(_00645_));
 sg13g2_mux2_1 _20390_ (.A0(_09252_),
    .A1(\cpu.dcache.r_tag[4][18] ),
    .S(net412),
    .X(_00646_));
 sg13g2_mux2_1 _20391_ (.A0(net424),
    .A1(\cpu.dcache.r_tag[4][19] ),
    .S(net412),
    .X(_00647_));
 sg13g2_mux2_1 _20392_ (.A0(net425),
    .A1(\cpu.dcache.r_tag[4][20] ),
    .S(net412),
    .X(_00648_));
 sg13g2_mux2_1 _20393_ (.A0(net426),
    .A1(\cpu.dcache.r_tag[4][21] ),
    .S(net412),
    .X(_00649_));
 sg13g2_mux2_1 _20394_ (.A0(net430),
    .A1(\cpu.dcache.r_tag[4][22] ),
    .S(net412),
    .X(_00650_));
 sg13g2_buf_1 _20395_ (.A(_12646_),
    .X(_03124_));
 sg13g2_mux2_1 _20396_ (.A0(net375),
    .A1(\cpu.dcache.r_tag[4][23] ),
    .S(net411),
    .X(_00651_));
 sg13g2_mux2_1 _20397_ (.A0(net717),
    .A1(\cpu.dcache.r_tag[4][6] ),
    .S(net411),
    .X(_00652_));
 sg13g2_mux2_1 _20398_ (.A0(net716),
    .A1(\cpu.dcache.r_tag[4][7] ),
    .S(net411),
    .X(_00653_));
 sg13g2_mux2_1 _20399_ (.A0(net715),
    .A1(\cpu.dcache.r_tag[4][8] ),
    .S(net411),
    .X(_00654_));
 sg13g2_mux2_1 _20400_ (.A0(_03102_),
    .A1(\cpu.dcache.r_tag[4][9] ),
    .S(net411),
    .X(_00655_));
 sg13g2_mux2_1 _20401_ (.A0(net843),
    .A1(\cpu.dcache.r_tag[4][10] ),
    .S(net411),
    .X(_00656_));
 sg13g2_mux2_1 _20402_ (.A0(net842),
    .A1(\cpu.dcache.r_tag[4][11] ),
    .S(net411),
    .X(_00657_));
 sg13g2_mux2_1 _20403_ (.A0(net376),
    .A1(\cpu.dcache.r_tag[4][12] ),
    .S(_03124_),
    .X(_00658_));
 sg13g2_mux2_1 _20404_ (.A0(net377),
    .A1(\cpu.dcache.r_tag[4][13] ),
    .S(net411),
    .X(_00659_));
 sg13g2_mux2_1 _20405_ (.A0(_09329_),
    .A1(\cpu.dcache.r_tag[4][14] ),
    .S(_03124_),
    .X(_00660_));
 sg13g2_buf_1 _20406_ (.A(_02773_),
    .X(_03125_));
 sg13g2_mux2_1 _20407_ (.A0(\cpu.dcache.r_tag[5][5] ),
    .A1(net508),
    .S(net361),
    .X(_00661_));
 sg13g2_mux2_1 _20408_ (.A0(\cpu.dcache.r_tag[5][15] ),
    .A1(net427),
    .S(net361),
    .X(_00662_));
 sg13g2_mux2_1 _20409_ (.A0(\cpu.dcache.r_tag[5][16] ),
    .A1(net432),
    .S(_03125_),
    .X(_00663_));
 sg13g2_mux2_1 _20410_ (.A0(\cpu.dcache.r_tag[5][17] ),
    .A1(_09362_),
    .S(_03125_),
    .X(_00664_));
 sg13g2_mux2_1 _20411_ (.A0(\cpu.dcache.r_tag[5][18] ),
    .A1(net431),
    .S(net361),
    .X(_00665_));
 sg13g2_mux2_1 _20412_ (.A0(\cpu.dcache.r_tag[5][19] ),
    .A1(net424),
    .S(net361),
    .X(_00666_));
 sg13g2_mux2_1 _20413_ (.A0(\cpu.dcache.r_tag[5][20] ),
    .A1(net425),
    .S(net361),
    .X(_00667_));
 sg13g2_mux2_1 _20414_ (.A0(\cpu.dcache.r_tag[5][21] ),
    .A1(_09446_),
    .S(net361),
    .X(_00668_));
 sg13g2_mux2_1 _20415_ (.A0(\cpu.dcache.r_tag[5][22] ),
    .A1(net430),
    .S(net361),
    .X(_00669_));
 sg13g2_mux2_1 _20416_ (.A0(\cpu.dcache.r_tag[5][23] ),
    .A1(net375),
    .S(net361),
    .X(_00670_));
 sg13g2_buf_1 _20417_ (.A(_02773_),
    .X(_03126_));
 sg13g2_mux2_1 _20418_ (.A0(\cpu.dcache.r_tag[5][6] ),
    .A1(_03111_),
    .S(net360),
    .X(_00671_));
 sg13g2_mux2_1 _20419_ (.A0(\cpu.dcache.r_tag[5][7] ),
    .A1(_03113_),
    .S(_03126_),
    .X(_00672_));
 sg13g2_mux2_1 _20420_ (.A0(\cpu.dcache.r_tag[5][8] ),
    .A1(_03114_),
    .S(net360),
    .X(_00673_));
 sg13g2_mux2_1 _20421_ (.A0(\cpu.dcache.r_tag[5][9] ),
    .A1(_03115_),
    .S(_03126_),
    .X(_00674_));
 sg13g2_mux2_1 _20422_ (.A0(\cpu.dcache.r_tag[5][10] ),
    .A1(_03116_),
    .S(net360),
    .X(_00675_));
 sg13g2_mux2_1 _20423_ (.A0(\cpu.dcache.r_tag[5][11] ),
    .A1(net839),
    .S(net360),
    .X(_00676_));
 sg13g2_mux2_1 _20424_ (.A0(\cpu.dcache.r_tag[5][12] ),
    .A1(net376),
    .S(net360),
    .X(_00677_));
 sg13g2_mux2_1 _20425_ (.A0(\cpu.dcache.r_tag[5][13] ),
    .A1(net377),
    .S(net360),
    .X(_00678_));
 sg13g2_mux2_1 _20426_ (.A0(\cpu.dcache.r_tag[5][14] ),
    .A1(net429),
    .S(net360),
    .X(_00679_));
 sg13g2_buf_1 _20427_ (.A(_02895_),
    .X(_03127_));
 sg13g2_mux2_1 _20428_ (.A0(\cpu.dcache.r_tag[6][5] ),
    .A1(net508),
    .S(_03127_),
    .X(_00680_));
 sg13g2_mux2_1 _20429_ (.A0(\cpu.dcache.r_tag[6][15] ),
    .A1(_09399_),
    .S(net452),
    .X(_00681_));
 sg13g2_mux2_1 _20430_ (.A0(\cpu.dcache.r_tag[6][16] ),
    .A1(_09208_),
    .S(_03127_),
    .X(_00682_));
 sg13g2_mux2_1 _20431_ (.A0(\cpu.dcache.r_tag[6][17] ),
    .A1(net428),
    .S(net452),
    .X(_00683_));
 sg13g2_mux2_1 _20432_ (.A0(\cpu.dcache.r_tag[6][18] ),
    .A1(net431),
    .S(net452),
    .X(_00684_));
 sg13g2_mux2_1 _20433_ (.A0(\cpu.dcache.r_tag[6][19] ),
    .A1(net424),
    .S(net452),
    .X(_00685_));
 sg13g2_mux2_1 _20434_ (.A0(\cpu.dcache.r_tag[6][20] ),
    .A1(_09607_),
    .S(net452),
    .X(_00686_));
 sg13g2_mux2_1 _20435_ (.A0(\cpu.dcache.r_tag[6][21] ),
    .A1(net426),
    .S(net452),
    .X(_00687_));
 sg13g2_mux2_1 _20436_ (.A0(\cpu.dcache.r_tag[6][22] ),
    .A1(net430),
    .S(net452),
    .X(_00688_));
 sg13g2_buf_1 _20437_ (.A(_02894_),
    .X(_03128_));
 sg13g2_mux2_1 _20438_ (.A0(\cpu.dcache.r_tag[6][23] ),
    .A1(net375),
    .S(net507),
    .X(_00689_));
 sg13g2_mux2_1 _20439_ (.A0(\cpu.dcache.r_tag[6][6] ),
    .A1(_03111_),
    .S(net507),
    .X(_00690_));
 sg13g2_mux2_1 _20440_ (.A0(\cpu.dcache.r_tag[6][7] ),
    .A1(_03113_),
    .S(_03128_),
    .X(_00691_));
 sg13g2_mux2_1 _20441_ (.A0(\cpu.dcache.r_tag[6][8] ),
    .A1(net712),
    .S(net507),
    .X(_00692_));
 sg13g2_mux2_1 _20442_ (.A0(\cpu.dcache.r_tag[6][9] ),
    .A1(_03115_),
    .S(_03128_),
    .X(_00693_));
 sg13g2_mux2_1 _20443_ (.A0(\cpu.dcache.r_tag[6][10] ),
    .A1(_03116_),
    .S(net507),
    .X(_00694_));
 sg13g2_mux2_1 _20444_ (.A0(\cpu.dcache.r_tag[6][11] ),
    .A1(net839),
    .S(net507),
    .X(_00695_));
 sg13g2_mux2_1 _20445_ (.A0(\cpu.dcache.r_tag[6][12] ),
    .A1(net376),
    .S(net507),
    .X(_00696_));
 sg13g2_mux2_1 _20446_ (.A0(\cpu.dcache.r_tag[6][13] ),
    .A1(net377),
    .S(net507),
    .X(_00697_));
 sg13g2_nand2_1 _20447_ (.Y(_03129_),
    .A(net429),
    .B(net507));
 sg13g2_o21ai_1 _20448_ (.B1(_03129_),
    .Y(_00698_),
    .A1(_09338_),
    .A2(net452));
 sg13g2_buf_1 _20449_ (.A(_03011_),
    .X(_03130_));
 sg13g2_mux2_1 _20450_ (.A0(\cpu.dcache.r_tag[7][5] ),
    .A1(net508),
    .S(_03130_),
    .X(_00699_));
 sg13g2_mux2_1 _20451_ (.A0(\cpu.dcache.r_tag[7][15] ),
    .A1(net427),
    .S(net451),
    .X(_00700_));
 sg13g2_mux2_1 _20452_ (.A0(\cpu.dcache.r_tag[7][16] ),
    .A1(_09208_),
    .S(_03130_),
    .X(_00701_));
 sg13g2_mux2_1 _20453_ (.A0(\cpu.dcache.r_tag[7][17] ),
    .A1(net428),
    .S(net451),
    .X(_00702_));
 sg13g2_mux2_1 _20454_ (.A0(\cpu.dcache.r_tag[7][18] ),
    .A1(_09252_),
    .S(net451),
    .X(_00703_));
 sg13g2_mux2_1 _20455_ (.A0(\cpu.dcache.r_tag[7][19] ),
    .A1(net424),
    .S(net451),
    .X(_00704_));
 sg13g2_buf_1 _20456_ (.A(_03010_),
    .X(_03131_));
 sg13g2_nand2_1 _20457_ (.Y(_03132_),
    .A(net425),
    .B(net506));
 sg13g2_o21ai_1 _20458_ (.B1(_03132_),
    .Y(_00705_),
    .A1(_09614_),
    .A2(net451));
 sg13g2_mux2_1 _20459_ (.A0(\cpu.dcache.r_tag[7][21] ),
    .A1(net426),
    .S(net451),
    .X(_00706_));
 sg13g2_mux2_1 _20460_ (.A0(\cpu.dcache.r_tag[7][22] ),
    .A1(_09294_),
    .S(net451),
    .X(_00707_));
 sg13g2_mux2_1 _20461_ (.A0(\cpu.dcache.r_tag[7][23] ),
    .A1(_09687_),
    .S(net451),
    .X(_00708_));
 sg13g2_buf_2 _20462_ (.A(net847),
    .X(_03133_));
 sg13g2_mux2_1 _20463_ (.A0(\cpu.dcache.r_tag[7][6] ),
    .A1(net711),
    .S(net506),
    .X(_00709_));
 sg13g2_buf_1 _20464_ (.A(net846),
    .X(_03134_));
 sg13g2_mux2_1 _20465_ (.A0(\cpu.dcache.r_tag[7][7] ),
    .A1(_03134_),
    .S(net506),
    .X(_00710_));
 sg13g2_buf_1 _20466_ (.A(net845),
    .X(_03135_));
 sg13g2_mux2_1 _20467_ (.A0(\cpu.dcache.r_tag[7][8] ),
    .A1(_03135_),
    .S(net506),
    .X(_00711_));
 sg13g2_buf_1 _20468_ (.A(net964),
    .X(_03136_));
 sg13g2_mux2_1 _20469_ (.A0(\cpu.dcache.r_tag[7][9] ),
    .A1(_03136_),
    .S(net506),
    .X(_00712_));
 sg13g2_buf_1 _20470_ (.A(net963),
    .X(_03137_));
 sg13g2_mux2_1 _20471_ (.A0(\cpu.dcache.r_tag[7][10] ),
    .A1(_03137_),
    .S(_03131_),
    .X(_00713_));
 sg13g2_buf_1 _20472_ (.A(net962),
    .X(_03138_));
 sg13g2_mux2_1 _20473_ (.A0(\cpu.dcache.r_tag[7][11] ),
    .A1(_03138_),
    .S(_03131_),
    .X(_00714_));
 sg13g2_mux2_1 _20474_ (.A0(\cpu.dcache.r_tag[7][12] ),
    .A1(net376),
    .S(net506),
    .X(_00715_));
 sg13g2_mux2_1 _20475_ (.A0(\cpu.dcache.r_tag[7][13] ),
    .A1(net377),
    .S(net506),
    .X(_00716_));
 sg13g2_mux2_1 _20476_ (.A0(\cpu.dcache.r_tag[7][14] ),
    .A1(net429),
    .S(net506),
    .X(_00717_));
 sg13g2_buf_1 _20477_ (.A(net152),
    .X(_03139_));
 sg13g2_nor2_1 _20478_ (.A(_08945_),
    .B(net150),
    .Y(_03140_));
 sg13g2_buf_1 _20479_ (.A(_03140_),
    .X(_03141_));
 sg13g2_nor2_1 _20480_ (.A(net305),
    .B(net253),
    .Y(_03142_));
 sg13g2_buf_1 _20481_ (.A(_03142_),
    .X(_03143_));
 sg13g2_buf_1 _20482_ (.A(_08761_),
    .X(_03144_));
 sg13g2_nor2_1 _20483_ (.A(_08721_),
    .B(net220),
    .Y(_03145_));
 sg13g2_buf_1 _20484_ (.A(_03145_),
    .X(_03146_));
 sg13g2_a21oi_1 _20485_ (.A1(net186),
    .A2(_03143_),
    .Y(_03147_),
    .B1(_03146_));
 sg13g2_nor2_2 _20486_ (.A(net212),
    .B(_03147_),
    .Y(_03148_));
 sg13g2_a21oi_1 _20487_ (.A1(net151),
    .A2(_03141_),
    .Y(_03149_),
    .B1(_03148_));
 sg13g2_buf_1 _20488_ (.A(net187),
    .X(_03150_));
 sg13g2_nand2_1 _20489_ (.Y(_03151_),
    .A(_10120_),
    .B(net141));
 sg13g2_o21ai_1 _20490_ (.B1(_03151_),
    .Y(_00726_),
    .A1(net117),
    .A2(_03149_));
 sg13g2_nand2_1 _20491_ (.Y(_03152_),
    .A(net305),
    .B(_08802_));
 sg13g2_buf_1 _20492_ (.A(net186),
    .X(_03153_));
 sg13g2_buf_1 _20493_ (.A(net212),
    .X(_03154_));
 sg13g2_o21ai_1 _20494_ (.B1(net176),
    .Y(_03155_),
    .A1(net140),
    .A2(net211));
 sg13g2_buf_1 _20495_ (.A(net253),
    .X(_03156_));
 sg13g2_a21oi_1 _20496_ (.A1(_03152_),
    .A2(_03155_),
    .Y(_03157_),
    .B1(net219));
 sg13g2_buf_1 _20497_ (.A(_08935_),
    .X(_03158_));
 sg13g2_buf_1 _20498_ (.A(net218),
    .X(_03159_));
 sg13g2_buf_1 _20499_ (.A(net197),
    .X(_03160_));
 sg13g2_nor2_1 _20500_ (.A(net197),
    .B(net212),
    .Y(_03161_));
 sg13g2_nor2_1 _20501_ (.A(_08737_),
    .B(_08761_),
    .Y(_03162_));
 sg13g2_buf_1 _20502_ (.A(_03162_),
    .X(_03163_));
 sg13g2_nand2b_1 _20503_ (.Y(_03164_),
    .B(net196),
    .A_N(_03161_));
 sg13g2_o21ai_1 _20504_ (.B1(_03164_),
    .Y(_03165_),
    .A1(net175),
    .A2(_08947_));
 sg13g2_o21ai_1 _20505_ (.B1(net104),
    .Y(_03166_),
    .A1(_03157_),
    .A2(_03165_));
 sg13g2_o21ai_1 _20506_ (.B1(_03166_),
    .Y(_00727_),
    .A1(_11505_),
    .A2(_08926_));
 sg13g2_buf_1 _20507_ (.A(_08906_),
    .X(_03167_));
 sg13g2_nand3_1 _20508_ (.B(net116),
    .C(net177),
    .A(net121),
    .Y(_03168_));
 sg13g2_o21ai_1 _20509_ (.B1(_03168_),
    .Y(_00728_),
    .A1(_11888_),
    .A2(net105));
 sg13g2_buf_1 _20510_ (.A(net220),
    .X(_03169_));
 sg13g2_o21ai_1 _20511_ (.B1(net140),
    .Y(_03170_),
    .A1(net195),
    .A2(_03161_));
 sg13g2_nand2_1 _20512_ (.Y(_03171_),
    .A(\cpu.cond[2] ),
    .B(net141));
 sg13g2_o21ai_1 _20513_ (.B1(_03171_),
    .Y(_00729_),
    .A1(net117),
    .A2(_03170_));
 sg13g2_nand4_1 _20514_ (.B(net151),
    .C(net116),
    .A(_08925_),
    .Y(_03172_),
    .D(_08952_));
 sg13g2_o21ai_1 _20515_ (.B1(_03172_),
    .Y(_00730_),
    .A1(_09142_),
    .A2(net105));
 sg13g2_nor2_1 _20516_ (.A(_03158_),
    .B(_08762_),
    .Y(_03173_));
 sg13g2_buf_1 _20517_ (.A(_03173_),
    .X(_03174_));
 sg13g2_inv_1 _20518_ (.Y(_03175_),
    .A(_09714_));
 sg13g2_nor2_1 _20519_ (.A(_00153_),
    .B(net434),
    .Y(_03176_));
 sg13g2_mux2_1 _20520_ (.A0(\cpu.icache.r_data[5][24] ),
    .A1(\cpu.icache.r_data[7][24] ),
    .S(_08693_),
    .X(_03177_));
 sg13g2_a22oi_1 _20521_ (.Y(_03178_),
    .B1(_03177_),
    .B2(net793),
    .A2(_08582_),
    .A1(\cpu.icache.r_data[6][24] ));
 sg13g2_nor2_1 _20522_ (.A(net689),
    .B(_03178_),
    .Y(_03179_));
 sg13g2_a22oi_1 _20523_ (.Y(_03180_),
    .B1(net690),
    .B2(\cpu.icache.r_data[4][24] ),
    .A2(net468),
    .A1(\cpu.icache.r_data[2][24] ));
 sg13g2_a22oi_1 _20524_ (.Y(_03181_),
    .B1(net467),
    .B2(\cpu.icache.r_data[3][24] ),
    .A2(net535),
    .A1(\cpu.icache.r_data[1][24] ));
 sg13g2_nand2_1 _20525_ (.Y(_03182_),
    .A(_03180_),
    .B(_03181_));
 sg13g2_nor3_1 _20526_ (.A(_03176_),
    .B(_03179_),
    .C(_03182_),
    .Y(_03183_));
 sg13g2_nand2_1 _20527_ (.Y(_03184_),
    .A(_00152_),
    .B(net612));
 sg13g2_a22oi_1 _20528_ (.Y(_03185_),
    .B1(net611),
    .B2(\cpu.icache.r_data[5][8] ),
    .A2(net535),
    .A1(\cpu.icache.r_data[1][8] ));
 sg13g2_a22oi_1 _20529_ (.Y(_03186_),
    .B1(_08716_),
    .B2(\cpu.icache.r_data[3][8] ),
    .A2(_08700_),
    .A1(\cpu.icache.r_data[2][8] ));
 sg13g2_mux2_1 _20530_ (.A0(\cpu.icache.r_data[4][8] ),
    .A1(\cpu.icache.r_data[6][8] ),
    .S(net794),
    .X(_03187_));
 sg13g2_a22oi_1 _20531_ (.Y(_03188_),
    .B1(_03187_),
    .B2(net915),
    .A2(_08424_),
    .A1(\cpu.icache.r_data[7][8] ));
 sg13g2_or2_1 _20532_ (.X(_03189_),
    .B(_03188_),
    .A(net689));
 sg13g2_nand4_1 _20533_ (.B(_03185_),
    .C(_03186_),
    .A(_08689_),
    .Y(_03190_),
    .D(_03189_));
 sg13g2_a21oi_1 _20534_ (.A1(_03184_),
    .A2(_03190_),
    .Y(_03191_),
    .B1(_08707_));
 sg13g2_a21o_1 _20535_ (.A2(_03183_),
    .A1(net784),
    .B1(_03191_),
    .X(_03192_));
 sg13g2_buf_2 _20536_ (.A(_03192_),
    .X(_03193_));
 sg13g2_nor2_1 _20537_ (.A(_00155_),
    .B(net470),
    .Y(_03194_));
 sg13g2_mux2_1 _20538_ (.A0(\cpu.icache.r_data[5][25] ),
    .A1(\cpu.icache.r_data[7][25] ),
    .S(net794),
    .X(_03195_));
 sg13g2_a22oi_1 _20539_ (.Y(_03196_),
    .B1(_03195_),
    .B2(net793),
    .A2(_08742_),
    .A1(\cpu.icache.r_data[4][25] ));
 sg13g2_nor2_1 _20540_ (.A(net689),
    .B(_03196_),
    .Y(_03197_));
 sg13g2_a22oi_1 _20541_ (.Y(_03198_),
    .B1(net467),
    .B2(\cpu.icache.r_data[3][25] ),
    .A2(net534),
    .A1(\cpu.icache.r_data[6][25] ));
 sg13g2_a22oi_1 _20542_ (.Y(_03199_),
    .B1(_08785_),
    .B2(\cpu.icache.r_data[1][25] ),
    .A2(net465),
    .A1(\cpu.icache.r_data[2][25] ));
 sg13g2_nand2_1 _20543_ (.Y(_03200_),
    .A(_03198_),
    .B(_03199_));
 sg13g2_nor4_1 _20544_ (.A(net1044),
    .B(_03194_),
    .C(_03197_),
    .D(_03200_),
    .Y(_03201_));
 sg13g2_nand2_1 _20545_ (.Y(_03202_),
    .A(_00154_),
    .B(_08710_));
 sg13g2_nor2b_1 _20546_ (.A(net903),
    .B_N(\cpu.icache.r_data[4][9] ),
    .Y(_03203_));
 sg13g2_a21oi_1 _20547_ (.A1(_08325_),
    .A2(\cpu.icache.r_data[6][9] ),
    .Y(_03204_),
    .B1(_03203_));
 sg13g2_a22oi_1 _20548_ (.Y(_03205_),
    .B1(_08364_),
    .B2(\cpu.icache.r_data[7][9] ),
    .A2(_08752_),
    .A1(\cpu.icache.r_data[5][9] ));
 sg13g2_o21ai_1 _20549_ (.B1(_03205_),
    .Y(_03206_),
    .A1(net793),
    .A2(_03204_));
 sg13g2_nand2_1 _20550_ (.Y(_03207_),
    .A(net1050),
    .B(_03206_));
 sg13g2_nand2_1 _20551_ (.Y(_03208_),
    .A(\cpu.icache.r_data[1][9] ),
    .B(_08785_));
 sg13g2_a22oi_1 _20552_ (.Y(_03209_),
    .B1(net536),
    .B2(\cpu.icache.r_data[3][9] ),
    .A2(net465),
    .A1(\cpu.icache.r_data[2][9] ));
 sg13g2_nand4_1 _20553_ (.B(_03207_),
    .C(_03208_),
    .A(net470),
    .Y(_03210_),
    .D(_03209_));
 sg13g2_a21oi_1 _20554_ (.A1(_03202_),
    .A2(_03210_),
    .Y(_03211_),
    .B1(net902));
 sg13g2_or2_1 _20555_ (.X(_03212_),
    .B(_03211_),
    .A(_03201_));
 sg13g2_buf_1 _20556_ (.A(_03212_),
    .X(_03213_));
 sg13g2_a22oi_1 _20557_ (.Y(_03214_),
    .B1(net534),
    .B2(\cpu.icache.r_data[6][7] ),
    .A2(net533),
    .A1(\cpu.icache.r_data[1][7] ));
 sg13g2_a22oi_1 _20558_ (.Y(_03215_),
    .B1(net536),
    .B2(\cpu.icache.r_data[3][7] ),
    .A2(net465),
    .A1(\cpu.icache.r_data[2][7] ));
 sg13g2_mux2_1 _20559_ (.A0(\cpu.icache.r_data[5][7] ),
    .A1(\cpu.icache.r_data[7][7] ),
    .S(net903),
    .X(_03216_));
 sg13g2_a22oi_1 _20560_ (.Y(_03217_),
    .B1(_03216_),
    .B2(net912),
    .A2(_08742_),
    .A1(\cpu.icache.r_data[4][7] ));
 sg13g2_or2_1 _20561_ (.X(_03218_),
    .B(_03217_),
    .A(net785));
 sg13g2_and4_1 _20562_ (.A(net470),
    .B(_03214_),
    .C(_03215_),
    .D(_03218_),
    .X(_03219_));
 sg13g2_a21oi_1 _20563_ (.A1(_00150_),
    .A2(net612),
    .Y(_03220_),
    .B1(_03219_));
 sg13g2_nor2_1 _20564_ (.A(_00151_),
    .B(_08357_),
    .Y(_03221_));
 sg13g2_mux2_1 _20565_ (.A0(\cpu.icache.r_data[7][23] ),
    .A1(\cpu.icache.r_data[3][23] ),
    .S(net785),
    .X(_03222_));
 sg13g2_a22oi_1 _20566_ (.Y(_03223_),
    .B1(_03222_),
    .B2(_08693_),
    .A2(_08328_),
    .A1(\cpu.icache.r_data[5][23] ));
 sg13g2_nor2_1 _20567_ (.A(net915),
    .B(_03223_),
    .Y(_03224_));
 sg13g2_a22oi_1 _20568_ (.Y(_03225_),
    .B1(net534),
    .B2(\cpu.icache.r_data[6][23] ),
    .A2(net465),
    .A1(\cpu.icache.r_data[2][23] ));
 sg13g2_a22oi_1 _20569_ (.Y(_03226_),
    .B1(net533),
    .B2(\cpu.icache.r_data[1][23] ),
    .A2(net690),
    .A1(\cpu.icache.r_data[4][23] ));
 sg13g2_nand2_1 _20570_ (.Y(_03227_),
    .A(_03225_),
    .B(_03226_));
 sg13g2_or4_1 _20571_ (.A(net1044),
    .B(_03221_),
    .C(_03224_),
    .D(_03227_),
    .X(_03228_));
 sg13g2_o21ai_1 _20572_ (.B1(_03228_),
    .Y(_03229_),
    .A1(net902),
    .A2(_03220_));
 sg13g2_buf_1 _20573_ (.A(_03229_),
    .X(_03230_));
 sg13g2_and2_1 _20574_ (.A(net217),
    .B(_03230_),
    .X(_03231_));
 sg13g2_nand2_1 _20575_ (.Y(_03232_),
    .A(_03193_),
    .B(_03231_));
 sg13g2_nor3_1 _20576_ (.A(net211),
    .B(_03175_),
    .C(_03232_),
    .Y(_03233_));
 sg13g2_nand3_1 _20577_ (.B(_03174_),
    .C(_03233_),
    .A(net116),
    .Y(_03234_));
 sg13g2_inv_1 _20578_ (.Y(_03235_),
    .A(_00161_));
 sg13g2_nand2_1 _20579_ (.Y(_03236_),
    .A(\cpu.icache.r_data[2][20] ),
    .B(_08306_));
 sg13g2_a22oi_1 _20580_ (.Y(_03237_),
    .B1(net618),
    .B2(\cpu.icache.r_data[1][20] ),
    .A2(net699),
    .A1(\cpu.icache.r_data[4][20] ));
 sg13g2_a22oi_1 _20581_ (.Y(_03238_),
    .B1(net536),
    .B2(\cpu.icache.r_data[3][20] ),
    .A2(_08367_),
    .A1(\cpu.icache.r_data[7][20] ));
 sg13g2_a22oi_1 _20582_ (.Y(_03239_),
    .B1(net696),
    .B2(\cpu.icache.r_data[5][20] ),
    .A2(net538),
    .A1(\cpu.icache.r_data[6][20] ));
 sg13g2_nand4_1 _20583_ (.B(_03237_),
    .C(_03238_),
    .A(_03236_),
    .Y(_03240_),
    .D(_03239_));
 sg13g2_a21oi_1 _20584_ (.A1(_03235_),
    .A2(net612),
    .Y(_03241_),
    .B1(_03240_));
 sg13g2_nand2_1 _20585_ (.Y(_03242_),
    .A(_00160_),
    .B(net612));
 sg13g2_a22oi_1 _20586_ (.Y(_03243_),
    .B1(net538),
    .B2(\cpu.icache.r_data[6][4] ),
    .A2(net618),
    .A1(\cpu.icache.r_data[1][4] ));
 sg13g2_a22oi_1 _20587_ (.Y(_03244_),
    .B1(net536),
    .B2(\cpu.icache.r_data[3][4] ),
    .A2(_08306_),
    .A1(\cpu.icache.r_data[2][4] ));
 sg13g2_mux2_1 _20588_ (.A0(\cpu.icache.r_data[5][4] ),
    .A1(\cpu.icache.r_data[7][4] ),
    .S(net914),
    .X(_03245_));
 sg13g2_a22oi_1 _20589_ (.Y(_03246_),
    .B1(_03245_),
    .B2(_08331_),
    .A2(_08742_),
    .A1(\cpu.icache.r_data[4][4] ));
 sg13g2_or2_1 _20590_ (.X(_03247_),
    .B(_03246_),
    .A(net785));
 sg13g2_nand4_1 _20591_ (.B(_03243_),
    .C(_03244_),
    .A(_08300_),
    .Y(_03248_),
    .D(_03247_));
 sg13g2_nand3_1 _20592_ (.B(_03242_),
    .C(_03248_),
    .A(net1044),
    .Y(_03249_));
 sg13g2_o21ai_1 _20593_ (.B1(_03249_),
    .Y(_03250_),
    .A1(_08709_),
    .A2(_03241_));
 sg13g2_buf_2 _20594_ (.A(_03250_),
    .X(_03251_));
 sg13g2_buf_1 _20595_ (.A(_03251_),
    .X(_03252_));
 sg13g2_nor4_1 _20596_ (.A(net187),
    .B(_08951_),
    .C(_03234_),
    .D(net216),
    .Y(_03253_));
 sg13g2_a21o_1 _20597_ (.A2(net122),
    .A1(\cpu.dec.do_flush_all ),
    .B1(_03253_),
    .X(_00731_));
 sg13g2_nand2_1 _20598_ (.Y(_03254_),
    .A(net150),
    .B(_03143_));
 sg13g2_nor3_1 _20599_ (.A(net209),
    .B(net212),
    .C(_03254_),
    .Y(_03255_));
 sg13g2_mux2_1 _20600_ (.A0(_03255_),
    .A1(\cpu.dec.do_flush_write ),
    .S(net149),
    .X(_00732_));
 sg13g2_nor3_1 _20601_ (.A(net232),
    .B(_08947_),
    .C(net177),
    .Y(_03256_));
 sg13g2_buf_1 _20602_ (.A(_08945_),
    .X(_03257_));
 sg13g2_a22oi_1 _20603_ (.Y(_03258_),
    .B1(net196),
    .B2(_03252_),
    .A2(net254),
    .A1(net220));
 sg13g2_inv_1 _20604_ (.Y(_03259_),
    .A(_00156_));
 sg13g2_a22oi_1 _20605_ (.Y(_03260_),
    .B1(_08712_),
    .B2(\cpu.icache.r_data[5][2] ),
    .A2(_08315_),
    .A1(\cpu.icache.r_data[1][2] ));
 sg13g2_a22oi_1 _20606_ (.Y(_03261_),
    .B1(_08374_),
    .B2(\cpu.icache.r_data[3][2] ),
    .A2(net539),
    .A1(\cpu.icache.r_data[2][2] ));
 sg13g2_mux2_1 _20607_ (.A0(\cpu.icache.r_data[4][2] ),
    .A1(\cpu.icache.r_data[6][2] ),
    .S(_08605_),
    .X(_03262_));
 sg13g2_a22oi_1 _20608_ (.Y(_03263_),
    .B1(_03262_),
    .B2(_08302_),
    .A2(_08364_),
    .A1(\cpu.icache.r_data[7][2] ));
 sg13g2_or2_1 _20609_ (.X(_03264_),
    .B(_03263_),
    .A(_08691_));
 sg13g2_nand4_1 _20610_ (.B(_03260_),
    .C(_03261_),
    .A(_08357_),
    .Y(_03265_),
    .D(_03264_));
 sg13g2_o21ai_1 _20611_ (.B1(_03265_),
    .Y(_03266_),
    .A1(_03259_),
    .A2(_08298_));
 sg13g2_nand2_1 _20612_ (.Y(_03267_),
    .A(\cpu.icache.r_data[2][18] ),
    .B(_08784_));
 sg13g2_a22oi_1 _20613_ (.Y(_03268_),
    .B1(net533),
    .B2(\cpu.icache.r_data[1][18] ),
    .A2(_08310_),
    .A1(\cpu.icache.r_data[4][18] ));
 sg13g2_a22oi_1 _20614_ (.Y(_03269_),
    .B1(_08374_),
    .B2(\cpu.icache.r_data[3][18] ),
    .A2(_08367_),
    .A1(\cpu.icache.r_data[7][18] ));
 sg13g2_a22oi_1 _20615_ (.Y(_03270_),
    .B1(net611),
    .B2(\cpu.icache.r_data[5][18] ),
    .A2(_08321_),
    .A1(\cpu.icache.r_data[6][18] ));
 sg13g2_nand4_1 _20616_ (.B(_03268_),
    .C(_03269_),
    .A(_03267_),
    .Y(_03271_),
    .D(_03270_));
 sg13g2_nor2_1 _20617_ (.A(_00157_),
    .B(_08298_),
    .Y(_03272_));
 sg13g2_o21ai_1 _20618_ (.B1(net902),
    .Y(_03273_),
    .A1(_03271_),
    .A2(_03272_));
 sg13g2_o21ai_1 _20619_ (.B1(_03273_),
    .Y(_03274_),
    .A1(_08706_),
    .A2(_03266_));
 sg13g2_buf_1 _20620_ (.A(_03274_),
    .X(_03275_));
 sg13g2_buf_1 _20621_ (.A(_03275_),
    .X(_03276_));
 sg13g2_nand2_1 _20622_ (.Y(_03277_),
    .A(_09726_),
    .B(net194));
 sg13g2_o21ai_1 _20623_ (.B1(_03277_),
    .Y(_03278_),
    .A1(_09726_),
    .A2(net231));
 sg13g2_nand3_1 _20624_ (.B(_08906_),
    .C(_03278_),
    .A(net185),
    .Y(_03279_));
 sg13g2_o21ai_1 _20625_ (.B1(_03279_),
    .Y(_03280_),
    .A1(net174),
    .A2(_03258_));
 sg13g2_a21oi_1 _20626_ (.A1(net254),
    .A2(_03256_),
    .Y(_03281_),
    .B1(_03280_));
 sg13g2_nand3_1 _20627_ (.B(_03141_),
    .C(net196),
    .A(net254),
    .Y(_03282_));
 sg13g2_o21ai_1 _20628_ (.B1(_03282_),
    .Y(_03283_),
    .A1(_03141_),
    .A2(_03281_));
 sg13g2_mux2_1 _20629_ (.A0(_03283_),
    .A1(_10205_),
    .S(net149),
    .X(_00733_));
 sg13g2_inv_1 _20630_ (.Y(_03284_),
    .A(_03251_));
 sg13g2_nor2_1 _20631_ (.A(net218),
    .B(_08937_),
    .Y(_03285_));
 sg13g2_a21oi_1 _20632_ (.A1(_03284_),
    .A2(_03285_),
    .Y(_03286_),
    .B1(_08947_));
 sg13g2_buf_1 _20633_ (.A(_03286_),
    .X(_03287_));
 sg13g2_nand2_1 _20634_ (.Y(_03288_),
    .A(net232),
    .B(net220));
 sg13g2_buf_2 _20635_ (.A(_03288_),
    .X(_03289_));
 sg13g2_buf_1 _20636_ (.A(net305),
    .X(_03290_));
 sg13g2_nand2_1 _20637_ (.Y(_03291_),
    .A(net209),
    .B(_03290_));
 sg13g2_nand2_1 _20638_ (.Y(_03292_),
    .A(net211),
    .B(_03145_));
 sg13g2_buf_2 _20639_ (.A(_03292_),
    .X(_03293_));
 sg13g2_nand2_1 _20640_ (.Y(_03294_),
    .A(_03291_),
    .B(_03293_));
 sg13g2_inv_1 _20641_ (.Y(_03295_),
    .A(_03294_));
 sg13g2_o21ai_1 _20642_ (.B1(_03295_),
    .Y(_03296_),
    .A1(_03289_),
    .A2(_03193_));
 sg13g2_nand2_1 _20643_ (.Y(_03297_),
    .A(net116),
    .B(_09727_));
 sg13g2_nand2_1 _20644_ (.Y(_03298_),
    .A(_08947_),
    .B(_03297_));
 sg13g2_nor3_2 _20645_ (.A(_03158_),
    .B(net305),
    .C(net220),
    .Y(_03299_));
 sg13g2_nand2_1 _20646_ (.Y(_03300_),
    .A(net216),
    .B(_03299_));
 sg13g2_o21ai_1 _20647_ (.B1(_03300_),
    .Y(_03301_),
    .A1(_03293_),
    .A2(_03297_));
 sg13g2_inv_1 _20648_ (.Y(_03302_),
    .A(_03152_));
 sg13g2_nor3_1 _20649_ (.A(net218),
    .B(net305),
    .C(net186),
    .Y(_03303_));
 sg13g2_a21oi_1 _20650_ (.A1(net218),
    .A2(_03302_),
    .Y(_03304_),
    .B1(_03303_));
 sg13g2_nand2_1 _20651_ (.Y(_03305_),
    .A(_03144_),
    .B(_03251_));
 sg13g2_nor3_1 _20652_ (.A(net174),
    .B(_03304_),
    .C(_03305_),
    .Y(_03306_));
 sg13g2_buf_1 _20653_ (.A(_03306_),
    .X(_03307_));
 sg13g2_a221oi_1 _20654_ (.B2(_03301_),
    .C1(_03307_),
    .B1(_03298_),
    .A1(_03287_),
    .Y(_03308_),
    .A2(_03296_));
 sg13g2_nand2_1 _20655_ (.Y(_03309_),
    .A(\cpu.dec.imm[10] ),
    .B(net141));
 sg13g2_o21ai_1 _20656_ (.B1(_03309_),
    .Y(_00734_),
    .A1(net117),
    .A2(_03308_));
 sg13g2_nand2_1 _20657_ (.Y(_03310_),
    .A(_08945_),
    .B(_08804_));
 sg13g2_nor2_1 _20658_ (.A(_03310_),
    .B(_03174_),
    .Y(_03311_));
 sg13g2_buf_2 _20659_ (.A(_03311_),
    .X(_03312_));
 sg13g2_nand2_1 _20660_ (.Y(_03313_),
    .A(_08721_),
    .B(net196));
 sg13g2_buf_2 _20661_ (.A(_03313_),
    .X(_03314_));
 sg13g2_o21ai_1 _20662_ (.B1(_03293_),
    .Y(_03315_),
    .A1(net231),
    .A2(_03314_));
 sg13g2_a21oi_1 _20663_ (.A1(net784),
    .A2(_03183_),
    .Y(_03316_),
    .B1(_03191_));
 sg13g2_buf_1 _20664_ (.A(_03316_),
    .X(_03317_));
 sg13g2_nand3_1 _20665_ (.B(_03317_),
    .C(_03231_),
    .A(_08913_),
    .Y(_03318_));
 sg13g2_buf_1 _20666_ (.A(_03318_),
    .X(_03319_));
 sg13g2_o21ai_1 _20667_ (.B1(_03299_),
    .Y(_03320_),
    .A1(_03251_),
    .A2(net139));
 sg13g2_buf_1 _20668_ (.A(_03320_),
    .X(_03321_));
 sg13g2_and2_1 _20669_ (.A(net231),
    .B(net139),
    .X(_03322_));
 sg13g2_nor2_2 _20670_ (.A(net218),
    .B(net220),
    .Y(_03323_));
 sg13g2_o21ai_1 _20671_ (.B1(net232),
    .Y(_03324_),
    .A1(_08949_),
    .A2(_03323_));
 sg13g2_o21ai_1 _20672_ (.B1(_03159_),
    .Y(_03325_),
    .A1(net185),
    .A2(_08949_));
 sg13g2_nand2_1 _20673_ (.Y(_03326_),
    .A(_03324_),
    .B(_03325_));
 sg13g2_o21ai_1 _20674_ (.B1(_03326_),
    .Y(_03327_),
    .A1(_03321_),
    .A2(_03322_));
 sg13g2_a221oi_1 _20675_ (.B2(_03287_),
    .C1(_03307_),
    .B1(_03327_),
    .A1(_03312_),
    .Y(_03328_),
    .A2(_03315_));
 sg13g2_nand2_1 _20676_ (.Y(_03329_),
    .A(\cpu.dec.imm[11] ),
    .B(net141));
 sg13g2_o21ai_1 _20677_ (.B1(_03329_),
    .Y(_00735_),
    .A1(net117),
    .A2(_03328_));
 sg13g2_o21ai_1 _20678_ (.B1(_03293_),
    .Y(_03330_),
    .A1(_08929_),
    .A2(_03314_));
 sg13g2_and2_1 _20679_ (.A(_08929_),
    .B(net139),
    .X(_03331_));
 sg13g2_o21ai_1 _20680_ (.B1(_03326_),
    .Y(_03332_),
    .A1(_03321_),
    .A2(_03331_));
 sg13g2_a221oi_1 _20681_ (.B2(_03287_),
    .C1(_03307_),
    .B1(_03332_),
    .A1(_03312_),
    .Y(_03333_),
    .A2(_03330_));
 sg13g2_nand2_1 _20682_ (.Y(_03334_),
    .A(\cpu.dec.imm[12] ),
    .B(_03150_));
 sg13g2_o21ai_1 _20683_ (.B1(_03334_),
    .Y(_00736_),
    .A1(net117),
    .A2(_03333_));
 sg13g2_nand2_1 _20684_ (.Y(_03335_),
    .A(net218),
    .B(net253));
 sg13g2_buf_2 _20685_ (.A(_03335_),
    .X(_03336_));
 sg13g2_a21oi_1 _20686_ (.A1(_03336_),
    .A2(_03314_),
    .Y(_03337_),
    .B1(_08949_));
 sg13g2_and2_1 _20687_ (.A(_08949_),
    .B(net139),
    .X(_03338_));
 sg13g2_o21ai_1 _20688_ (.B1(_03326_),
    .Y(_03339_),
    .A1(_03321_),
    .A2(_03338_));
 sg13g2_a221oi_1 _20689_ (.B2(_03287_),
    .C1(_03307_),
    .B1(_03339_),
    .A1(_03312_),
    .Y(_03340_),
    .A2(_03337_));
 sg13g2_nand2_1 _20690_ (.Y(_03341_),
    .A(\cpu.dec.imm[13] ),
    .B(net141));
 sg13g2_o21ai_1 _20691_ (.B1(_03341_),
    .Y(_00737_),
    .A1(net117),
    .A2(_03340_));
 sg13g2_a22oi_1 _20692_ (.Y(_03342_),
    .B1(_03299_),
    .B2(net210),
    .A2(net177),
    .A1(net211));
 sg13g2_nor2b_1 _20693_ (.A(net210),
    .B_N(net139),
    .Y(_03343_));
 sg13g2_o21ai_1 _20694_ (.B1(_03326_),
    .Y(_03344_),
    .A1(_03321_),
    .A2(_03343_));
 sg13g2_a21oi_1 _20695_ (.A1(_03287_),
    .A2(_03344_),
    .Y(_03345_),
    .B1(_03307_));
 sg13g2_o21ai_1 _20696_ (.B1(_03345_),
    .Y(_03346_),
    .A1(_03297_),
    .A2(_03342_));
 sg13g2_mux2_1 _20697_ (.A0(_03346_),
    .A1(\cpu.dec.imm[14] ),
    .S(net149),
    .X(_00738_));
 sg13g2_o21ai_1 _20698_ (.B1(_03293_),
    .Y(_03347_),
    .A1(net210),
    .A2(_03314_));
 sg13g2_nand2_1 _20699_ (.Y(_03348_),
    .A(_03312_),
    .B(_03347_));
 sg13g2_a21oi_1 _20700_ (.A1(_03345_),
    .A2(_03348_),
    .Y(_03349_),
    .B1(net152));
 sg13g2_a21o_1 _20701_ (.A2(net122),
    .A1(\cpu.dec.imm[15] ),
    .B1(_03349_),
    .X(_00739_));
 sg13g2_buf_1 _20702_ (.A(net239),
    .X(_03350_));
 sg13g2_nor2_1 _20703_ (.A(net150),
    .B(_03319_),
    .Y(_03351_));
 sg13g2_o21ai_1 _20704_ (.B1(net219),
    .Y(_03352_),
    .A1(net215),
    .A2(_03351_));
 sg13g2_nand3_1 _20705_ (.B(_03254_),
    .C(_03352_),
    .A(_03152_),
    .Y(_03353_));
 sg13g2_nand2_1 _20706_ (.Y(_03354_),
    .A(net120),
    .B(net174));
 sg13g2_a21oi_1 _20707_ (.A1(net209),
    .A2(_03353_),
    .Y(_03355_),
    .B1(_03354_));
 sg13g2_nand2_1 _20708_ (.Y(_03356_),
    .A(_08783_),
    .B(net186));
 sg13g2_buf_1 _20709_ (.A(_03356_),
    .X(_03357_));
 sg13g2_nand2_1 _20710_ (.Y(_03358_),
    .A(net116),
    .B(_03174_));
 sg13g2_nand2b_1 _20711_ (.Y(_03359_),
    .B(_03358_),
    .A_N(_03148_));
 sg13g2_nor2_1 _20712_ (.A(_00159_),
    .B(_08297_),
    .Y(_03360_));
 sg13g2_mux2_1 _20713_ (.A0(\cpu.icache.r_data[5][19] ),
    .A1(\cpu.icache.r_data[7][19] ),
    .S(net794),
    .X(_03361_));
 sg13g2_a22oi_1 _20714_ (.Y(_03362_),
    .B1(_03361_),
    .B2(_08332_),
    .A2(_08582_),
    .A1(\cpu.icache.r_data[6][19] ));
 sg13g2_nor2_1 _20715_ (.A(_08739_),
    .B(_03362_),
    .Y(_03363_));
 sg13g2_a22oi_1 _20716_ (.Y(_03364_),
    .B1(_08310_),
    .B2(\cpu.icache.r_data[4][19] ),
    .A2(net539),
    .A1(\cpu.icache.r_data[2][19] ));
 sg13g2_a22oi_1 _20717_ (.Y(_03365_),
    .B1(net536),
    .B2(\cpu.icache.r_data[3][19] ),
    .A2(net613),
    .A1(\cpu.icache.r_data[1][19] ));
 sg13g2_nand2_1 _20718_ (.Y(_03366_),
    .A(_03364_),
    .B(_03365_));
 sg13g2_nor3_1 _20719_ (.A(_03360_),
    .B(_03363_),
    .C(_03366_),
    .Y(_03367_));
 sg13g2_nand2_1 _20720_ (.Y(_03368_),
    .A(_00158_),
    .B(_08658_));
 sg13g2_a22oi_1 _20721_ (.Y(_03369_),
    .B1(_08315_),
    .B2(\cpu.icache.r_data[1][3] ),
    .A2(net795),
    .A1(\cpu.icache.r_data[4][3] ));
 sg13g2_a22oi_1 _20722_ (.Y(_03370_),
    .B1(net536),
    .B2(\cpu.icache.r_data[3][3] ),
    .A2(_08358_),
    .A1(\cpu.icache.r_data[2][3] ));
 sg13g2_mux2_1 _20723_ (.A0(\cpu.icache.r_data[5][3] ),
    .A1(\cpu.icache.r_data[7][3] ),
    .S(net914),
    .X(_03371_));
 sg13g2_a22oi_1 _20724_ (.Y(_03372_),
    .B1(_03371_),
    .B2(_08331_),
    .A2(_08582_),
    .A1(\cpu.icache.r_data[6][3] ));
 sg13g2_or2_1 _20725_ (.X(_03373_),
    .B(_03372_),
    .A(net785));
 sg13g2_nand4_1 _20726_ (.B(_03369_),
    .C(_03370_),
    .A(_08300_),
    .Y(_03374_),
    .D(_03373_));
 sg13g2_a21oi_1 _20727_ (.A1(_03368_),
    .A2(_03374_),
    .Y(_03375_),
    .B1(_08705_));
 sg13g2_a21oi_1 _20728_ (.A1(net902),
    .A2(_03367_),
    .Y(_03376_),
    .B1(_03375_));
 sg13g2_buf_1 _20729_ (.A(_03376_),
    .X(_03377_));
 sg13g2_nand3_1 _20730_ (.B(_03359_),
    .C(net238),
    .A(net115),
    .Y(_03378_));
 sg13g2_o21ai_1 _20731_ (.B1(_03378_),
    .Y(_03379_),
    .A1(net233),
    .A2(_03355_));
 sg13g2_mux2_1 _20732_ (.A0(_03379_),
    .A1(_10327_),
    .S(net149),
    .X(_00740_));
 sg13g2_inv_1 _20733_ (.Y(_03380_),
    .A(_10458_));
 sg13g2_nor3_1 _20734_ (.A(net197),
    .B(net185),
    .C(net196),
    .Y(_03381_));
 sg13g2_a21o_1 _20735_ (.A2(_03367_),
    .A1(net688),
    .B1(_03375_),
    .X(_03382_));
 sg13g2_buf_1 _20736_ (.A(_03382_),
    .X(_03383_));
 sg13g2_nor2_1 _20737_ (.A(net120),
    .B(_03383_),
    .Y(_03384_));
 sg13g2_a221oi_1 _20738_ (.B2(net234),
    .C1(_03384_),
    .B1(_03381_),
    .A1(_03174_),
    .Y(_03385_),
    .A2(net216));
 sg13g2_nor2_1 _20739_ (.A(_03310_),
    .B(_03385_),
    .Y(_03386_));
 sg13g2_a21oi_1 _20740_ (.A1(_03148_),
    .A2(net216),
    .Y(_03387_),
    .B1(_03386_));
 sg13g2_nor2_1 _20741_ (.A(net218),
    .B(net305),
    .Y(_03388_));
 sg13g2_inv_1 _20742_ (.Y(_03389_),
    .A(_03388_));
 sg13g2_nor2_1 _20743_ (.A(net234),
    .B(_03389_),
    .Y(_03390_));
 sg13g2_nor3_1 _20744_ (.A(net186),
    .B(net238),
    .C(_03388_),
    .Y(_03391_));
 sg13g2_o21ai_1 _20745_ (.B1(_03169_),
    .Y(_03392_),
    .A1(_03390_),
    .A2(_03391_));
 sg13g2_nor3_1 _20746_ (.A(_03144_),
    .B(_08905_),
    .C(_08841_),
    .Y(_03393_));
 sg13g2_nor2_1 _20747_ (.A(net174),
    .B(_03393_),
    .Y(_03394_));
 sg13g2_a22oi_1 _20748_ (.Y(_03395_),
    .B1(_03392_),
    .B2(_03394_),
    .A2(_03285_),
    .A1(_03153_));
 sg13g2_a21oi_1 _20749_ (.A1(net140),
    .A2(_08913_),
    .Y(_03396_),
    .B1(_03395_));
 sg13g2_nand2_1 _20750_ (.Y(_03397_),
    .A(_08806_),
    .B(_03291_));
 sg13g2_nor2_2 _20751_ (.A(_03314_),
    .B(net139),
    .Y(_03398_));
 sg13g2_a21oi_1 _20752_ (.A1(net254),
    .A2(_03398_),
    .Y(_03399_),
    .B1(_03384_));
 sg13g2_nor2_1 _20753_ (.A(_03397_),
    .B(_03399_),
    .Y(_03400_));
 sg13g2_nor3_1 _20754_ (.A(net152),
    .B(_03396_),
    .C(_03400_),
    .Y(_03401_));
 sg13g2_a22oi_1 _20755_ (.Y(_00741_),
    .B1(_03387_),
    .B2(_03401_),
    .A2(_03139_),
    .A1(_03380_));
 sg13g2_nand2_1 _20756_ (.Y(_03402_),
    .A(_08764_),
    .B(_03251_));
 sg13g2_o21ai_1 _20757_ (.B1(_03402_),
    .Y(_03403_),
    .A1(_08913_),
    .A2(_03336_));
 sg13g2_a221oi_1 _20758_ (.B2(_08912_),
    .C1(_03403_),
    .B1(_03398_),
    .A1(_08928_),
    .Y(_03404_),
    .A2(_03143_));
 sg13g2_nor2_1 _20759_ (.A(net253),
    .B(net186),
    .Y(_03405_));
 sg13g2_o21ai_1 _20760_ (.B1(_03290_),
    .Y(_03406_),
    .A1(_08939_),
    .A2(net186));
 sg13g2_a21o_1 _20761_ (.A2(_03406_),
    .A1(_03254_),
    .B1(_03159_),
    .X(_03407_));
 sg13g2_o21ai_1 _20762_ (.B1(_03407_),
    .Y(_03408_),
    .A1(_03257_),
    .A2(_03405_));
 sg13g2_a21o_1 _20763_ (.A2(_03174_),
    .A1(_08928_),
    .B1(_03403_),
    .X(_03409_));
 sg13g2_nor3_1 _20764_ (.A(_09729_),
    .B(_03305_),
    .C(_03388_),
    .Y(_03410_));
 sg13g2_a221oi_1 _20765_ (.B2(_03167_),
    .C1(_03410_),
    .B1(_03409_),
    .A1(_08912_),
    .Y(_03411_),
    .A2(_03408_));
 sg13g2_o21ai_1 _20766_ (.B1(_03411_),
    .Y(_03412_),
    .A1(_03397_),
    .A2(_03404_));
 sg13g2_mux2_1 _20767_ (.A0(_03412_),
    .A1(_10427_),
    .S(_08960_),
    .X(_00742_));
 sg13g2_nand2b_1 _20768_ (.Y(_03413_),
    .B(_03398_),
    .A_N(_03397_));
 sg13g2_nor2_1 _20769_ (.A(net176),
    .B(_03256_),
    .Y(_03414_));
 sg13g2_nand3_1 _20770_ (.B(_03413_),
    .C(_03414_),
    .A(_08908_),
    .Y(_03415_));
 sg13g2_and2_1 _20771_ (.A(net210),
    .B(net115),
    .X(_03416_));
 sg13g2_a22oi_1 _20772_ (.Y(_03417_),
    .B1(_03416_),
    .B2(_03148_),
    .A2(_03415_),
    .A1(net211));
 sg13g2_nand2_1 _20773_ (.Y(_03418_),
    .A(\cpu.dec.imm[4] ),
    .B(net141));
 sg13g2_o21ai_1 _20774_ (.B1(_03418_),
    .Y(_00743_),
    .A1(net117),
    .A2(_03417_));
 sg13g2_nor3_1 _20775_ (.A(net151),
    .B(net231),
    .C(net196),
    .Y(_03419_));
 sg13g2_a21oi_1 _20776_ (.A1(net151),
    .A2(net194),
    .Y(_03420_),
    .B1(_03419_));
 sg13g2_and2_1 _20777_ (.A(_03299_),
    .B(_03319_),
    .X(_03421_));
 sg13g2_o21ai_1 _20778_ (.B1(net140),
    .Y(_03422_),
    .A1(net176),
    .A2(_03421_));
 sg13g2_nand3_1 _20779_ (.B(net116),
    .C(_03336_),
    .A(net120),
    .Y(_03423_));
 sg13g2_nand3_1 _20780_ (.B(_03422_),
    .C(_03423_),
    .A(_03276_),
    .Y(_03424_));
 sg13g2_o21ai_1 _20781_ (.B1(_03424_),
    .Y(_03425_),
    .A1(net115),
    .A2(_03420_));
 sg13g2_mux2_1 _20782_ (.A0(_03425_),
    .A1(\cpu.dec.imm[5] ),
    .S(net149),
    .X(_00744_));
 sg13g2_nor2_1 _20783_ (.A(_08945_),
    .B(_08905_),
    .Y(_03426_));
 sg13g2_buf_1 _20784_ (.A(_03426_),
    .X(_03427_));
 sg13g2_buf_1 _20785_ (.A(_03427_),
    .X(_03428_));
 sg13g2_o21ai_1 _20786_ (.B1(_03377_),
    .Y(_03429_),
    .A1(_03156_),
    .A2(_03388_));
 sg13g2_nand2_1 _20787_ (.Y(_03430_),
    .A(_03428_),
    .B(_03429_));
 sg13g2_o21ai_1 _20788_ (.B1(_03257_),
    .Y(_03431_),
    .A1(_09710_),
    .A2(_03336_));
 sg13g2_buf_1 _20789_ (.A(_03230_),
    .X(_03432_));
 sg13g2_nor3_1 _20790_ (.A(net212),
    .B(_03289_),
    .C(net193),
    .Y(_03433_));
 sg13g2_o21ai_1 _20791_ (.B1(net238),
    .Y(_03434_),
    .A1(_03285_),
    .A2(_03398_));
 sg13g2_nand2b_1 _20792_ (.Y(_03435_),
    .B(_03434_),
    .A_N(_03433_));
 sg13g2_a22oi_1 _20793_ (.Y(_03436_),
    .B1(_03435_),
    .B2(_03153_),
    .A2(_03431_),
    .A1(_03430_));
 sg13g2_nor3_1 _20794_ (.A(net219),
    .B(_08765_),
    .C(net193),
    .Y(_03437_));
 sg13g2_nor3_1 _20795_ (.A(net115),
    .B(_03384_),
    .C(_03437_),
    .Y(_03438_));
 sg13g2_nor3_1 _20796_ (.A(net152),
    .B(_03436_),
    .C(_03438_),
    .Y(_03439_));
 sg13g2_a21o_1 _20797_ (.A2(net122),
    .A1(\cpu.dec.imm[6] ),
    .B1(_03439_),
    .X(_00745_));
 sg13g2_inv_1 _20798_ (.Y(_03440_),
    .A(net233));
 sg13g2_a22oi_1 _20799_ (.Y(_03441_),
    .B1(_03161_),
    .B2(_03351_),
    .A2(_03427_),
    .A1(net215));
 sg13g2_a22oi_1 _20800_ (.Y(_03442_),
    .B1(_03427_),
    .B2(_03143_),
    .A2(_08806_),
    .A1(net239));
 sg13g2_or2_1 _20801_ (.X(_03443_),
    .B(_03442_),
    .A(_03160_));
 sg13g2_o21ai_1 _20802_ (.B1(_03443_),
    .Y(_03444_),
    .A1(net195),
    .A2(_03441_));
 sg13g2_nor2_1 _20803_ (.A(net253),
    .B(_08764_),
    .Y(_03445_));
 sg13g2_nand2_1 _20804_ (.Y(_03446_),
    .A(_03317_),
    .B(_03445_));
 sg13g2_a21oi_1 _20805_ (.A1(_03402_),
    .A2(_03446_),
    .Y(_03447_),
    .B1(net115));
 sg13g2_a221oi_1 _20806_ (.B2(_03444_),
    .C1(_03447_),
    .B1(net216),
    .A1(_03440_),
    .Y(_03448_),
    .A2(_03148_));
 sg13g2_buf_1 _20807_ (.A(net187),
    .X(_03449_));
 sg13g2_nand2_1 _20808_ (.Y(_03450_),
    .A(\cpu.dec.imm[7] ),
    .B(_03449_));
 sg13g2_o21ai_1 _20809_ (.B1(_03450_),
    .Y(_00746_),
    .A1(_03139_),
    .A2(_03448_));
 sg13g2_nor2_1 _20810_ (.A(net115),
    .B(net217),
    .Y(_03451_));
 sg13g2_inv_1 _20811_ (.Y(_03452_),
    .A(net194));
 sg13g2_o21ai_1 _20812_ (.B1(_03293_),
    .Y(_03453_),
    .A1(_03452_),
    .A2(_03314_));
 sg13g2_a221oi_1 _20813_ (.B2(_03312_),
    .C1(_03307_),
    .B1(_03453_),
    .A1(_03445_),
    .Y(_03454_),
    .A2(_03451_));
 sg13g2_a21oi_1 _20814_ (.A1(_03452_),
    .A2(net139),
    .Y(_03455_),
    .B1(_03321_));
 sg13g2_o21ai_1 _20815_ (.B1(_03295_),
    .Y(_03456_),
    .A1(_03289_),
    .A2(net217));
 sg13g2_o21ai_1 _20816_ (.B1(_03287_),
    .Y(_03457_),
    .A1(_03455_),
    .A2(_03456_));
 sg13g2_a21oi_1 _20817_ (.A1(_03454_),
    .A2(_03457_),
    .Y(_03458_),
    .B1(_08687_));
 sg13g2_a21o_1 _20818_ (.A2(net122),
    .A1(\cpu.dec.imm[8] ),
    .B1(_03458_),
    .X(_00747_));
 sg13g2_o21ai_1 _20819_ (.B1(_03293_),
    .Y(_03459_),
    .A1(_03314_),
    .A2(_03383_));
 sg13g2_a21oi_1 _20820_ (.A1(net139),
    .A2(_03383_),
    .Y(_03460_),
    .B1(_03321_));
 sg13g2_a21oi_1 _20821_ (.A1(net234),
    .A2(_03143_),
    .Y(_03461_),
    .B1(_03294_));
 sg13g2_nand2b_1 _20822_ (.Y(_03462_),
    .B(_03461_),
    .A_N(_03460_));
 sg13g2_a221oi_1 _20823_ (.B2(_03287_),
    .C1(_03307_),
    .B1(_03462_),
    .A1(_03312_),
    .Y(_03463_),
    .A2(_03459_));
 sg13g2_nand2_1 _20824_ (.Y(_03464_),
    .A(\cpu.dec.imm[9] ),
    .B(net138));
 sg13g2_o21ai_1 _20825_ (.B1(_03464_),
    .Y(_00748_),
    .A1(net117),
    .A2(_03463_));
 sg13g2_buf_1 _20826_ (.A(\cpu.dec.do_inv_mmu ),
    .X(_03465_));
 sg13g2_nor4_1 _20827_ (.A(net789),
    .B(net152),
    .C(net233),
    .D(_03234_),
    .Y(_03466_));
 sg13g2_a21o_1 _20828_ (.A2(net122),
    .A1(_03465_),
    .B1(_03466_),
    .X(_00749_));
 sg13g2_inv_1 _20829_ (.Y(_03467_),
    .A(\cpu.dec.io ));
 sg13g2_nand3_1 _20830_ (.B(net116),
    .C(_03381_),
    .A(net121),
    .Y(_03468_));
 sg13g2_o21ai_1 _20831_ (.B1(_03468_),
    .Y(_00750_),
    .A1(_03467_),
    .A2(net105));
 sg13g2_nor4_1 _20832_ (.A(_08843_),
    .B(_03251_),
    .C(_03275_),
    .D(net238),
    .Y(_03469_));
 sg13g2_buf_2 _20833_ (.A(_03469_),
    .X(_03470_));
 sg13g2_nand3_1 _20834_ (.B(net97),
    .C(_03470_),
    .A(net151),
    .Y(_03471_));
 sg13g2_nand2_1 _20835_ (.Y(_03472_),
    .A(_11508_),
    .B(net138));
 sg13g2_o21ai_1 _20836_ (.B1(_03472_),
    .Y(_00751_),
    .A1(_08688_),
    .A2(_03471_));
 sg13g2_inv_1 _20837_ (.Y(_03473_),
    .A(_11495_));
 sg13g2_nand2_1 _20838_ (.Y(_03474_),
    .A(net215),
    .B(net150));
 sg13g2_nand2_1 _20839_ (.Y(_03475_),
    .A(net174),
    .B(_03474_));
 sg13g2_nand3_1 _20840_ (.B(_03323_),
    .C(_03475_),
    .A(net121),
    .Y(_03476_));
 sg13g2_o21ai_1 _20841_ (.B1(_03476_),
    .Y(_00752_),
    .A1(_03473_),
    .A2(net105));
 sg13g2_nor4_1 _20842_ (.A(net187),
    .B(_08843_),
    .C(_08908_),
    .D(_08950_),
    .Y(_03477_));
 sg13g2_a21o_1 _20843_ (.A2(net122),
    .A1(\cpu.dec.mult ),
    .B1(_03477_),
    .X(_00753_));
 sg13g2_o21ai_1 _20844_ (.B1(_08954_),
    .Y(_03478_),
    .A1(net210),
    .A2(net211));
 sg13g2_nand3_1 _20845_ (.B(_03154_),
    .C(_08949_),
    .A(net209),
    .Y(_03479_));
 sg13g2_nand3_1 _20846_ (.B(net174),
    .C(_08879_),
    .A(_03160_),
    .Y(_03480_));
 sg13g2_nand4_1 _20847_ (.B(_03405_),
    .C(_03479_),
    .A(_03350_),
    .Y(_03481_),
    .D(_03480_));
 sg13g2_o21ai_1 _20848_ (.B1(_03481_),
    .Y(_03482_),
    .A1(_08807_),
    .A2(_03478_));
 sg13g2_nand2_1 _20849_ (.Y(_03483_),
    .A(net104),
    .B(_03482_));
 sg13g2_o21ai_1 _20850_ (.B1(_03483_),
    .Y(_00754_),
    .A1(_10131_),
    .A2(net105));
 sg13g2_nand2_1 _20851_ (.Y(_03484_),
    .A(net239),
    .B(net194));
 sg13g2_o21ai_1 _20852_ (.B1(_03484_),
    .Y(_03485_),
    .A1(net215),
    .A2(net193));
 sg13g2_nand2_1 _20853_ (.Y(_03486_),
    .A(_03323_),
    .B(_03485_));
 sg13g2_o21ai_1 _20854_ (.B1(_03486_),
    .Y(_03487_),
    .A1(net120),
    .A2(net193));
 sg13g2_nand2_1 _20855_ (.Y(_03488_),
    .A(net175),
    .B(_08762_));
 sg13g2_a21oi_1 _20856_ (.A1(_03289_),
    .A2(net194),
    .Y(_03489_),
    .B1(net175));
 sg13g2_a21o_1 _20857_ (.A2(net193),
    .A1(_03289_),
    .B1(_08947_),
    .X(_03490_));
 sg13g2_o21ai_1 _20858_ (.B1(_03490_),
    .Y(_03491_),
    .A1(_03357_),
    .A2(_03489_));
 sg13g2_nand3_1 _20859_ (.B(net211),
    .C(_03470_),
    .A(net197),
    .Y(_03492_));
 sg13g2_o21ai_1 _20860_ (.B1(_03492_),
    .Y(_03493_),
    .A1(_03432_),
    .A2(_03470_));
 sg13g2_nor2_1 _20861_ (.A(net197),
    .B(_03432_),
    .Y(_03494_));
 sg13g2_a21oi_1 _20862_ (.A1(_03289_),
    .A2(_03493_),
    .Y(_03495_),
    .B1(_03494_));
 sg13g2_nor3_1 _20863_ (.A(_09729_),
    .B(_03146_),
    .C(_03495_),
    .Y(_03496_));
 sg13g2_a221oi_1 _20864_ (.B2(_03491_),
    .C1(_03496_),
    .B1(_03488_),
    .A1(_03167_),
    .Y(_03497_),
    .A2(_03487_));
 sg13g2_nand2_1 _20865_ (.Y(_03498_),
    .A(\cpu.dec.r_rd[0] ),
    .B(net138));
 sg13g2_o21ai_1 _20866_ (.B1(_03498_),
    .Y(_00755_),
    .A1(net123),
    .A2(_03497_));
 sg13g2_o21ai_1 _20867_ (.B1(_08947_),
    .Y(_03499_),
    .A1(_09729_),
    .A2(_03470_));
 sg13g2_o21ai_1 _20868_ (.B1(_09729_),
    .Y(_03500_),
    .A1(net220),
    .A2(_08947_));
 sg13g2_a22oi_1 _20869_ (.Y(_03501_),
    .B1(_03500_),
    .B2(net209),
    .A2(_03499_),
    .A1(_08941_));
 sg13g2_inv_1 _20870_ (.Y(_03502_),
    .A(_03501_));
 sg13g2_nor3_1 _20871_ (.A(net197),
    .B(_03143_),
    .C(_03357_),
    .Y(_03503_));
 sg13g2_o21ai_1 _20872_ (.B1(net209),
    .Y(_03504_),
    .A1(net220),
    .A2(net238));
 sg13g2_o21ai_1 _20873_ (.B1(_03504_),
    .Y(_03505_),
    .A1(net219),
    .A2(_03193_));
 sg13g2_nor2_1 _20874_ (.A(net215),
    .B(_03193_),
    .Y(_03506_));
 sg13g2_a22oi_1 _20875_ (.Y(_03507_),
    .B1(_03506_),
    .B2(_03323_),
    .A2(_03505_),
    .A1(net215));
 sg13g2_nand4_1 _20876_ (.B(_08842_),
    .C(_03233_),
    .A(_08824_),
    .Y(_03508_),
    .D(_03251_));
 sg13g2_nor3_1 _20877_ (.A(net194),
    .B(_03383_),
    .C(_03508_),
    .Y(_03509_));
 sg13g2_nor2_1 _20878_ (.A(_09727_),
    .B(_03509_),
    .Y(_03510_));
 sg13g2_nor3_1 _20879_ (.A(_03310_),
    .B(_03507_),
    .C(_03510_),
    .Y(_03511_));
 sg13g2_a221oi_1 _20880_ (.B2(net238),
    .C1(_03511_),
    .B1(_03503_),
    .A1(_03317_),
    .Y(_03512_),
    .A2(_03502_));
 sg13g2_nand2_1 _20881_ (.Y(_03513_),
    .A(\cpu.dec.r_rd[1] ),
    .B(_03449_));
 sg13g2_o21ai_1 _20882_ (.B1(_03513_),
    .Y(_00756_),
    .A1(net123),
    .A2(_03512_));
 sg13g2_nand2_1 _20883_ (.Y(_03514_),
    .A(net239),
    .B(_03252_));
 sg13g2_o21ai_1 _20884_ (.B1(_03514_),
    .Y(_03515_),
    .A1(net239),
    .A2(net217));
 sg13g2_nand2_1 _20885_ (.Y(_03516_),
    .A(_03323_),
    .B(_03515_));
 sg13g2_o21ai_1 _20886_ (.B1(_03516_),
    .Y(_03517_),
    .A1(net120),
    .A2(_03213_));
 sg13g2_a22oi_1 _20887_ (.Y(_03518_),
    .B1(_03517_),
    .B2(_03312_),
    .A2(_03503_),
    .A1(net216));
 sg13g2_o21ai_1 _20888_ (.B1(_03518_),
    .Y(_03519_),
    .A1(_03213_),
    .A2(_03501_));
 sg13g2_mux2_1 _20889_ (.A0(_03519_),
    .A1(\cpu.dec.r_rd[2] ),
    .S(_08960_),
    .X(_00757_));
 sg13g2_a21oi_1 _20890_ (.A1(net219),
    .A2(net234),
    .Y(_03520_),
    .B1(net185));
 sg13g2_nand3b_1 _20891_ (.B(net234),
    .C(net185),
    .Y(_03521_),
    .A_N(_03470_));
 sg13g2_o21ai_1 _20892_ (.B1(_03521_),
    .Y(_03522_),
    .A1(net175),
    .A2(_03520_));
 sg13g2_o21ai_1 _20893_ (.B1(net115),
    .Y(_03523_),
    .A1(net212),
    .A2(_08913_));
 sg13g2_o21ai_1 _20894_ (.B1(net150),
    .Y(_03524_),
    .A1(net195),
    .A2(net176));
 sg13g2_a22oi_1 _20895_ (.Y(_03525_),
    .B1(_03524_),
    .B2(net215),
    .A2(_03523_),
    .A1(net219));
 sg13g2_nor2_1 _20896_ (.A(net175),
    .B(_03525_),
    .Y(_03526_));
 sg13g2_a221oi_1 _20897_ (.B2(_03522_),
    .C1(_03526_),
    .B1(net97),
    .A1(net151),
    .Y(_03527_),
    .A2(net174));
 sg13g2_nand2_1 _20898_ (.Y(_03528_),
    .A(\cpu.dec.r_rd[3] ),
    .B(net138));
 sg13g2_o21ai_1 _20899_ (.B1(_03528_),
    .Y(_00758_),
    .A1(net123),
    .A2(_03527_));
 sg13g2_or2_1 _20900_ (.X(_03529_),
    .B(net193),
    .A(net195));
 sg13g2_a21oi_1 _20901_ (.A1(net120),
    .A2(_03529_),
    .Y(_03530_),
    .B1(net115));
 sg13g2_nand2_1 _20902_ (.Y(_03531_),
    .A(_08762_),
    .B(_03336_));
 sg13g2_nor2_1 _20903_ (.A(_08902_),
    .B(_03470_),
    .Y(_03532_));
 sg13g2_nor2_1 _20904_ (.A(net120),
    .B(_03532_),
    .Y(_03533_));
 sg13g2_or2_1 _20905_ (.X(_03534_),
    .B(_03533_),
    .A(_03445_));
 sg13g2_a22oi_1 _20906_ (.Y(_03535_),
    .B1(_03534_),
    .B2(_03427_),
    .A2(_03531_),
    .A1(_08806_));
 sg13g2_nand2_1 _20907_ (.Y(_03536_),
    .A(_03312_),
    .B(_03314_));
 sg13g2_a21oi_1 _20908_ (.A1(_03535_),
    .A2(_03536_),
    .Y(_03537_),
    .B1(net193));
 sg13g2_o21ai_1 _20909_ (.B1(net104),
    .Y(_03538_),
    .A1(_03530_),
    .A2(_03537_));
 sg13g2_o21ai_1 _20910_ (.B1(_03538_),
    .Y(_00759_),
    .A1(_10101_),
    .A2(net104));
 sg13g2_o21ai_1 _20911_ (.B1(net195),
    .Y(_03539_),
    .A1(net239),
    .A2(net150));
 sg13g2_nand3_1 _20912_ (.B(_03474_),
    .C(_03539_),
    .A(_03336_),
    .Y(_03540_));
 sg13g2_a22oi_1 _20913_ (.Y(_03541_),
    .B1(_03351_),
    .B2(_03163_),
    .A2(_03405_),
    .A1(net215));
 sg13g2_nor2_1 _20914_ (.A(net175),
    .B(_03541_),
    .Y(_03542_));
 sg13g2_a21oi_1 _20915_ (.A1(_03317_),
    .A2(_03540_),
    .Y(_03543_),
    .B1(_03542_));
 sg13g2_o21ai_1 _20916_ (.B1(_08943_),
    .Y(_03544_),
    .A1(net195),
    .A2(_03317_));
 sg13g2_a221oi_1 _20917_ (.B2(net151),
    .C1(net174),
    .B1(_03532_),
    .A1(_03193_),
    .Y(_03545_),
    .A2(_03405_));
 sg13g2_a21oi_1 _20918_ (.A1(net140),
    .A2(_03398_),
    .Y(_03546_),
    .B1(_03545_));
 sg13g2_a21o_1 _20919_ (.A2(_03544_),
    .A1(net140),
    .B1(_03546_),
    .X(_03547_));
 sg13g2_o21ai_1 _20920_ (.B1(_03547_),
    .Y(_03548_),
    .A1(net176),
    .A2(_03543_));
 sg13g2_mux2_1 _20921_ (.A0(_03548_),
    .A1(_10052_),
    .S(_03150_),
    .X(_00760_));
 sg13g2_nand2_1 _20922_ (.Y(_03549_),
    .A(net219),
    .B(_03141_));
 sg13g2_a21oi_1 _20923_ (.A1(_03535_),
    .A2(_03549_),
    .Y(_03550_),
    .B1(net217));
 sg13g2_a221oi_1 _20924_ (.B2(_09727_),
    .C1(_03310_),
    .B1(net217),
    .A1(net209),
    .Y(_03551_),
    .A2(net196));
 sg13g2_o21ai_1 _20925_ (.B1(net104),
    .Y(_03552_),
    .A1(_03550_),
    .A2(_03551_));
 sg13g2_o21ai_1 _20926_ (.B1(_03552_),
    .Y(_00761_),
    .A1(_10099_),
    .A2(net104));
 sg13g2_nand2_1 _20927_ (.Y(_03553_),
    .A(net218),
    .B(net239));
 sg13g2_nand2_1 _20928_ (.Y(_03554_),
    .A(net234),
    .B(_03533_));
 sg13g2_nand2b_1 _20929_ (.Y(_03555_),
    .B(_03554_),
    .A_N(_03553_));
 sg13g2_nand2_1 _20930_ (.Y(_03556_),
    .A(net150),
    .B(_03555_));
 sg13g2_nand2_1 _20931_ (.Y(_03557_),
    .A(_03350_),
    .B(_08906_));
 sg13g2_nand2_1 _20932_ (.Y(_03558_),
    .A(net232),
    .B(_03154_));
 sg13g2_a21oi_1 _20933_ (.A1(_03557_),
    .A2(_03558_),
    .Y(_03559_),
    .B1(net175));
 sg13g2_a221oi_1 _20934_ (.B2(net176),
    .C1(_03559_),
    .B1(_03556_),
    .A1(_08937_),
    .Y(_03560_),
    .A2(net140));
 sg13g2_a221oi_1 _20935_ (.B2(net97),
    .C1(net195),
    .B1(_03554_),
    .A1(_03161_),
    .Y(_03561_),
    .A2(_03474_));
 sg13g2_a21oi_1 _20936_ (.A1(net195),
    .A2(_03560_),
    .Y(_03562_),
    .B1(_03561_));
 sg13g2_nand2_1 _20937_ (.Y(_03563_),
    .A(_10248_),
    .B(net138));
 sg13g2_o21ai_1 _20938_ (.B1(_03563_),
    .Y(_00762_),
    .A1(net123),
    .A2(_03562_));
 sg13g2_nor2_1 _20939_ (.A(net177),
    .B(net194),
    .Y(_03564_));
 sg13g2_a21oi_1 _20940_ (.A1(net177),
    .A2(net193),
    .Y(_03565_),
    .B1(_03564_));
 sg13g2_nor2_1 _20941_ (.A(net233),
    .B(_08904_),
    .Y(_03566_));
 sg13g2_o21ai_1 _20942_ (.B1(_03389_),
    .Y(_03567_),
    .A1(_03553_),
    .A2(_03566_));
 sg13g2_a21oi_2 _20943_ (.B1(net140),
    .Y(_03568_),
    .A2(_03567_),
    .A1(_03169_));
 sg13g2_nor3_1 _20944_ (.A(net97),
    .B(_03452_),
    .C(_03568_),
    .Y(_03569_));
 sg13g2_a21oi_1 _20945_ (.A1(net97),
    .A2(_03565_),
    .Y(_03570_),
    .B1(_03569_));
 sg13g2_nand2_1 _20946_ (.Y(_03571_),
    .A(_11049_),
    .B(net138));
 sg13g2_o21ai_1 _20947_ (.B1(_03571_),
    .Y(_00763_),
    .A1(net123),
    .A2(_03570_));
 sg13g2_nor2_1 _20948_ (.A(_03336_),
    .B(_03317_),
    .Y(_03572_));
 sg13g2_a21oi_1 _20949_ (.A1(_03336_),
    .A2(_03383_),
    .Y(_03573_),
    .B1(_03572_));
 sg13g2_nor3_1 _20950_ (.A(net97),
    .B(_03383_),
    .C(_03568_),
    .Y(_03574_));
 sg13g2_a21oi_1 _20951_ (.A1(net97),
    .A2(_03573_),
    .Y(_03575_),
    .B1(_03574_));
 sg13g2_nand2_1 _20952_ (.Y(_03576_),
    .A(net592),
    .B(net138));
 sg13g2_o21ai_1 _20953_ (.B1(_03576_),
    .Y(_00764_),
    .A1(net123),
    .A2(_03575_));
 sg13g2_nor2_1 _20954_ (.A(net177),
    .B(net216),
    .Y(_03577_));
 sg13g2_a21oi_1 _20955_ (.A1(net177),
    .A2(net217),
    .Y(_03578_),
    .B1(_03577_));
 sg13g2_o21ai_1 _20956_ (.B1(_09729_),
    .Y(_03579_),
    .A1(_03284_),
    .A2(_03568_));
 sg13g2_o21ai_1 _20957_ (.B1(_03579_),
    .Y(_03580_),
    .A1(_09729_),
    .A2(_03578_));
 sg13g2_nand2_1 _20958_ (.Y(_03581_),
    .A(_10897_),
    .B(net138));
 sg13g2_o21ai_1 _20959_ (.B1(_03581_),
    .Y(_00765_),
    .A1(net123),
    .A2(_03580_));
 sg13g2_nand2_1 _20960_ (.Y(_03582_),
    .A(_09729_),
    .B(_03568_));
 sg13g2_a22oi_1 _20961_ (.Y(_03583_),
    .B1(_08913_),
    .B2(net219),
    .A2(_09710_),
    .A1(net185));
 sg13g2_nand3b_1 _20962_ (.B(net97),
    .C(net175),
    .Y(_03584_),
    .A_N(_03583_));
 sg13g2_nand3_1 _20963_ (.B(_03582_),
    .C(_03584_),
    .A(net121),
    .Y(_03585_));
 sg13g2_o21ai_1 _20964_ (.B1(_03585_),
    .Y(_00766_),
    .A1(net737),
    .A2(net104));
 sg13g2_nor4_1 _20965_ (.A(net187),
    .B(_08904_),
    .C(_08908_),
    .D(_08951_),
    .Y(_03586_));
 sg13g2_a21o_1 _20966_ (.A2(net122),
    .A1(_10642_),
    .B1(_03586_),
    .X(_00767_));
 sg13g2_nor4_1 _20967_ (.A(_08686_),
    .B(_08807_),
    .C(_03440_),
    .D(_08904_),
    .Y(_03587_));
 sg13g2_a21o_1 _20968_ (.A2(_08883_),
    .A1(\cpu.dec.r_set_cc ),
    .B1(_03587_),
    .X(_00768_));
 sg13g2_nand2_1 _20969_ (.Y(_03588_),
    .A(net176),
    .B(net177));
 sg13g2_o21ai_1 _20970_ (.B1(_03588_),
    .Y(_03589_),
    .A1(net176),
    .A2(_03254_));
 sg13g2_buf_1 _20971_ (.A(\cpu.dec.r_store ),
    .X(_03590_));
 sg13g2_mux2_1 _20972_ (.A0(_03589_),
    .A1(_03590_),
    .S(net141),
    .X(_00769_));
 sg13g2_nand2b_1 _20973_ (.Y(_03591_),
    .B(_03509_),
    .A_N(_03358_));
 sg13g2_nand2_1 _20974_ (.Y(_03592_),
    .A(\cpu.dec.r_swapsp ),
    .B(net152));
 sg13g2_o21ai_1 _20975_ (.B1(_03592_),
    .Y(_00770_),
    .A1(net123),
    .A2(_03591_));
 sg13g2_nor4_1 _20976_ (.A(_03358_),
    .B(_03452_),
    .C(net238),
    .D(_03508_),
    .Y(_03593_));
 sg13g2_mux2_1 _20977_ (.A0(_03593_),
    .A1(\cpu.dec.r_sys_call ),
    .S(net141),
    .X(_00771_));
 sg13g2_o21ai_1 _20978_ (.B1(_08765_),
    .Y(_03594_),
    .A1(net254),
    .A2(_03232_));
 sg13g2_nor2_1 _20979_ (.A(_03175_),
    .B(_03232_),
    .Y(_03595_));
 sg13g2_nand3_1 _20980_ (.B(_03470_),
    .C(_03595_),
    .A(_03174_),
    .Y(_03596_));
 sg13g2_nand4_1 _20981_ (.B(_03141_),
    .C(_03594_),
    .A(_03289_),
    .Y(_03597_),
    .D(_03596_));
 sg13g2_buf_1 _20982_ (.A(_08222_),
    .X(_03598_));
 sg13g2_or2_1 _20983_ (.X(_03599_),
    .B(_10753_),
    .A(_03598_));
 sg13g2_nand2_1 _20984_ (.Y(_03600_),
    .A(net232),
    .B(_03599_));
 sg13g2_o21ai_1 _20985_ (.B1(net253),
    .Y(_03601_),
    .A1(net232),
    .A2(_03599_));
 sg13g2_nor2_1 _20986_ (.A(_03193_),
    .B(_03230_),
    .Y(_03602_));
 sg13g2_xor2_1 _20987_ (.B(_03602_),
    .A(net217),
    .X(_03603_));
 sg13g2_nor3_2 _20988_ (.A(net961),
    .B(net234),
    .C(_03603_),
    .Y(_03604_));
 sg13g2_a22oi_1 _20989_ (.Y(_03605_),
    .B1(_03604_),
    .B2(net196),
    .A2(_03601_),
    .A1(_03600_));
 sg13g2_or2_1 _20990_ (.X(_03606_),
    .B(net210),
    .A(_08762_));
 sg13g2_o21ai_1 _20991_ (.B1(_03606_),
    .Y(_03607_),
    .A1(net197),
    .A2(_03605_));
 sg13g2_nand4_1 _20992_ (.B(_08949_),
    .C(_09714_),
    .A(net961),
    .Y(_03608_),
    .D(_03470_));
 sg13g2_a22oi_1 _20993_ (.Y(_03609_),
    .B1(_03608_),
    .B2(_03255_),
    .A2(_03607_),
    .A1(net116));
 sg13g2_o21ai_1 _20994_ (.B1(net233),
    .Y(_03610_),
    .A1(net231),
    .A2(net216));
 sg13g2_a21oi_1 _20995_ (.A1(_03233_),
    .A2(_03610_),
    .Y(_03611_),
    .B1(_03509_));
 sg13g2_nor3_1 _20996_ (.A(net789),
    .B(_09727_),
    .C(_03611_),
    .Y(_03612_));
 sg13g2_nor2_1 _20997_ (.A(net961),
    .B(_03603_),
    .Y(_03613_));
 sg13g2_nor2_1 _20998_ (.A(_08132_),
    .B(_08901_),
    .Y(_03614_));
 sg13g2_a21oi_1 _20999_ (.A1(net961),
    .A2(_08902_),
    .Y(_03615_),
    .B1(_03614_));
 sg13g2_nand2_1 _21000_ (.Y(_03616_),
    .A(net231),
    .B(_03615_));
 sg13g2_nand2_1 _21001_ (.Y(_03617_),
    .A(_03276_),
    .B(net238));
 sg13g2_xnor2_1 _21002_ (.Y(_03618_),
    .A(_03284_),
    .B(_03617_));
 sg13g2_o21ai_1 _21003_ (.B1(net239),
    .Y(_03619_),
    .A1(_03616_),
    .A2(_03618_));
 sg13g2_a22oi_1 _21004_ (.Y(_03620_),
    .B1(_03619_),
    .B2(net197),
    .A2(_03613_),
    .A1(net232));
 sg13g2_o21ai_1 _21005_ (.B1(_03604_),
    .Y(_03621_),
    .A1(net253),
    .A2(_03533_));
 sg13g2_o21ai_1 _21006_ (.B1(_03621_),
    .Y(_03622_),
    .A1(_03156_),
    .A2(_03620_));
 sg13g2_mux2_1 _21007_ (.A0(_08843_),
    .A1(net194),
    .S(_08949_),
    .X(_03623_));
 sg13g2_nor2b_1 _21008_ (.A(_08860_),
    .B_N(_03623_),
    .Y(_03624_));
 sg13g2_o21ai_1 _21009_ (.B1(_08948_),
    .Y(_03625_),
    .A1(_03566_),
    .A2(_03624_));
 sg13g2_a21oi_1 _21010_ (.A1(_09730_),
    .A2(_03623_),
    .Y(_03626_),
    .B1(_03141_));
 sg13g2_nand3_1 _21011_ (.B(_03421_),
    .C(_03604_),
    .A(_08806_),
    .Y(_03627_));
 sg13g2_nand3_1 _21012_ (.B(_03626_),
    .C(_03627_),
    .A(_03625_),
    .Y(_03628_));
 sg13g2_a21oi_1 _21013_ (.A1(_03428_),
    .A2(_03622_),
    .Y(_03629_),
    .B1(_03628_));
 sg13g2_o21ai_1 _21014_ (.B1(_03629_),
    .Y(_03630_),
    .A1(_03609_),
    .A2(_03612_));
 sg13g2_nand3_1 _21015_ (.B(_03597_),
    .C(_03630_),
    .A(_08925_),
    .Y(_03631_));
 sg13g2_o21ai_1 _21016_ (.B1(_03631_),
    .Y(_00772_),
    .A1(_10260_),
    .A2(net104));
 sg13g2_buf_1 _21017_ (.A(net1118),
    .X(_03632_));
 sg13g2_buf_1 _21018_ (.A(net960),
    .X(_03633_));
 sg13g2_nand2b_1 _21019_ (.Y(_03634_),
    .B(net1102),
    .A_N(net1015));
 sg13g2_buf_1 _21020_ (.A(_03634_),
    .X(_03635_));
 sg13g2_inv_1 _21021_ (.Y(_03636_),
    .A(_10021_));
 sg13g2_nand3_1 _21022_ (.B(_03636_),
    .C(_10017_),
    .A(net1103),
    .Y(_03637_));
 sg13g2_buf_1 _21023_ (.A(_03637_),
    .X(_03638_));
 sg13g2_nor2_1 _21024_ (.A(_03635_),
    .B(_03638_),
    .Y(_03639_));
 sg13g2_buf_1 _21025_ (.A(_03639_),
    .X(_03640_));
 sg13g2_buf_1 _21026_ (.A(net578),
    .X(_03641_));
 sg13g2_mux2_1 _21027_ (.A0(\cpu.ex.r_10[0] ),
    .A1(net835),
    .S(net505),
    .X(_00777_));
 sg13g2_mux2_1 _21028_ (.A0(\cpu.ex.r_10[10] ),
    .A1(net837),
    .S(net505),
    .X(_00778_));
 sg13g2_mux2_1 _21029_ (.A0(\cpu.ex.r_10[11] ),
    .A1(net836),
    .S(net505),
    .X(_00779_));
 sg13g2_buf_1 _21030_ (.A(net589),
    .X(_03642_));
 sg13g2_buf_1 _21031_ (.A(_03642_),
    .X(_03643_));
 sg13g2_mux2_1 _21032_ (.A0(\cpu.ex.r_10[12] ),
    .A1(net450),
    .S(net505),
    .X(_00780_));
 sg13g2_buf_1 _21033_ (.A(net601),
    .X(_03644_));
 sg13g2_buf_1 _21034_ (.A(net503),
    .X(_03645_));
 sg13g2_mux2_1 _21035_ (.A0(\cpu.ex.r_10[13] ),
    .A1(net449),
    .S(net505),
    .X(_00781_));
 sg13g2_buf_1 _21036_ (.A(net732),
    .X(_03646_));
 sg13g2_buf_1 _21037_ (.A(net639),
    .X(_03647_));
 sg13g2_mux2_1 _21038_ (.A0(\cpu.ex.r_10[14] ),
    .A1(net577),
    .S(net505),
    .X(_00782_));
 sg13g2_buf_1 _21039_ (.A(net731),
    .X(_03648_));
 sg13g2_buf_1 _21040_ (.A(net638),
    .X(_03649_));
 sg13g2_mux2_1 _21041_ (.A0(\cpu.ex.r_10[15] ),
    .A1(net576),
    .S(net505),
    .X(_00783_));
 sg13g2_buf_1 _21042_ (.A(net755),
    .X(_03650_));
 sg13g2_buf_2 _21043_ (.A(net637),
    .X(_03651_));
 sg13g2_buf_1 _21044_ (.A(net575),
    .X(_03652_));
 sg13g2_mux2_1 _21045_ (.A0(\cpu.ex.r_10[1] ),
    .A1(net502),
    .S(_03641_),
    .X(_00784_));
 sg13g2_buf_2 _21046_ (.A(net456),
    .X(_03653_));
 sg13g2_nand2_1 _21047_ (.Y(_03654_),
    .A(net410),
    .B(net578));
 sg13g2_o21ai_1 _21048_ (.B1(_03654_),
    .Y(_00785_),
    .A1(_10442_),
    .A2(net505));
 sg13g2_buf_1 _21049_ (.A(net464),
    .X(_03655_));
 sg13g2_mux2_1 _21050_ (.A0(\cpu.ex.r_10[3] ),
    .A1(net409),
    .S(net578),
    .X(_00786_));
 sg13g2_buf_1 _21051_ (.A(net585),
    .X(_03656_));
 sg13g2_buf_2 _21052_ (.A(_03656_),
    .X(_03657_));
 sg13g2_buf_1 _21053_ (.A(_03657_),
    .X(_03658_));
 sg13g2_mux2_1 _21054_ (.A0(\cpu.ex.r_10[4] ),
    .A1(net408),
    .S(net578),
    .X(_00787_));
 sg13g2_nand2_1 _21055_ (.Y(_03659_),
    .A(net579),
    .B(_03640_));
 sg13g2_o21ai_1 _21056_ (.B1(_03659_),
    .Y(_00788_),
    .A1(_10515_),
    .A2(_03641_));
 sg13g2_mux2_1 _21057_ (.A0(\cpu.ex.r_10[6] ),
    .A1(net711),
    .S(net578),
    .X(_00789_));
 sg13g2_mux2_1 _21058_ (.A0(\cpu.ex.r_10[7] ),
    .A1(net710),
    .S(net578),
    .X(_00790_));
 sg13g2_mux2_1 _21059_ (.A0(\cpu.ex.r_10[8] ),
    .A1(net709),
    .S(net578),
    .X(_00791_));
 sg13g2_mux2_1 _21060_ (.A0(\cpu.ex.r_10[9] ),
    .A1(net838),
    .S(net578),
    .X(_00792_));
 sg13g2_nor2_1 _21061_ (.A(_10026_),
    .B(_03638_),
    .Y(_03660_));
 sg13g2_buf_2 _21062_ (.A(_03660_),
    .X(_03661_));
 sg13g2_buf_1 _21063_ (.A(_03661_),
    .X(_03662_));
 sg13g2_mux2_1 _21064_ (.A0(\cpu.ex.r_11[0] ),
    .A1(net835),
    .S(_03662_),
    .X(_00793_));
 sg13g2_mux2_1 _21065_ (.A0(\cpu.ex.r_11[10] ),
    .A1(net837),
    .S(net500),
    .X(_00794_));
 sg13g2_mux2_1 _21066_ (.A0(\cpu.ex.r_11[11] ),
    .A1(net836),
    .S(net500),
    .X(_00795_));
 sg13g2_mux2_1 _21067_ (.A0(\cpu.ex.r_11[12] ),
    .A1(net450),
    .S(net500),
    .X(_00796_));
 sg13g2_mux2_1 _21068_ (.A0(\cpu.ex.r_11[13] ),
    .A1(net449),
    .S(net500),
    .X(_00797_));
 sg13g2_mux2_1 _21069_ (.A0(\cpu.ex.r_11[14] ),
    .A1(net577),
    .S(net500),
    .X(_00798_));
 sg13g2_mux2_1 _21070_ (.A0(\cpu.ex.r_11[15] ),
    .A1(net576),
    .S(net500),
    .X(_00799_));
 sg13g2_mux2_1 _21071_ (.A0(\cpu.ex.r_11[1] ),
    .A1(net502),
    .S(_03662_),
    .X(_00800_));
 sg13g2_buf_1 _21072_ (.A(net410),
    .X(_03663_));
 sg13g2_mux2_1 _21073_ (.A0(\cpu.ex.r_11[2] ),
    .A1(_03663_),
    .S(net500),
    .X(_00801_));
 sg13g2_mux2_1 _21074_ (.A0(\cpu.ex.r_11[3] ),
    .A1(net409),
    .S(net500),
    .X(_00802_));
 sg13g2_mux2_1 _21075_ (.A0(\cpu.ex.r_11[4] ),
    .A1(net408),
    .S(_03661_),
    .X(_00803_));
 sg13g2_mux2_1 _21076_ (.A0(\cpu.ex.r_11[5] ),
    .A1(net508),
    .S(_03661_),
    .X(_00804_));
 sg13g2_mux2_1 _21077_ (.A0(\cpu.ex.r_11[6] ),
    .A1(net711),
    .S(_03661_),
    .X(_00805_));
 sg13g2_mux2_1 _21078_ (.A0(\cpu.ex.r_11[7] ),
    .A1(net710),
    .S(_03661_),
    .X(_00806_));
 sg13g2_mux2_1 _21079_ (.A0(\cpu.ex.r_11[8] ),
    .A1(net709),
    .S(_03661_),
    .X(_00807_));
 sg13g2_mux2_1 _21080_ (.A0(\cpu.ex.r_11[9] ),
    .A1(net838),
    .S(_03661_),
    .X(_00808_));
 sg13g2_nand3_1 _21081_ (.B(_10021_),
    .C(_10017_),
    .A(net1103),
    .Y(_03664_));
 sg13g2_buf_1 _21082_ (.A(_03664_),
    .X(_03665_));
 sg13g2_nor3_1 _21083_ (.A(net1102),
    .B(net1015),
    .C(_03665_),
    .Y(_03666_));
 sg13g2_buf_4 _21084_ (.X(_03667_),
    .A(_03666_));
 sg13g2_buf_1 _21085_ (.A(_03667_),
    .X(_03668_));
 sg13g2_mux2_1 _21086_ (.A0(\cpu.ex.r_12[0] ),
    .A1(net835),
    .S(net574),
    .X(_00809_));
 sg13g2_mux2_1 _21087_ (.A0(\cpu.ex.r_12[10] ),
    .A1(net837),
    .S(net574),
    .X(_00810_));
 sg13g2_mux2_1 _21088_ (.A0(\cpu.ex.r_12[11] ),
    .A1(net836),
    .S(net574),
    .X(_00811_));
 sg13g2_mux2_1 _21089_ (.A0(\cpu.ex.r_12[12] ),
    .A1(net450),
    .S(net574),
    .X(_00812_));
 sg13g2_mux2_1 _21090_ (.A0(\cpu.ex.r_12[13] ),
    .A1(net449),
    .S(net574),
    .X(_00813_));
 sg13g2_mux2_1 _21091_ (.A0(\cpu.ex.r_12[14] ),
    .A1(net577),
    .S(net574),
    .X(_00814_));
 sg13g2_mux2_1 _21092_ (.A0(\cpu.ex.r_12[15] ),
    .A1(net576),
    .S(net574),
    .X(_00815_));
 sg13g2_mux2_1 _21093_ (.A0(\cpu.ex.r_12[1] ),
    .A1(net502),
    .S(_03668_),
    .X(_00816_));
 sg13g2_mux2_1 _21094_ (.A0(\cpu.ex.r_12[2] ),
    .A1(net359),
    .S(_03668_),
    .X(_00817_));
 sg13g2_mux2_1 _21095_ (.A0(\cpu.ex.r_12[3] ),
    .A1(net409),
    .S(_03667_),
    .X(_00818_));
 sg13g2_mux2_1 _21096_ (.A0(\cpu.ex.r_12[4] ),
    .A1(_03658_),
    .S(_03667_),
    .X(_00819_));
 sg13g2_mux2_1 _21097_ (.A0(\cpu.ex.r_12[5] ),
    .A1(net508),
    .S(_03667_),
    .X(_00820_));
 sg13g2_nand2_1 _21098_ (.Y(_03669_),
    .A(net847),
    .B(_03667_));
 sg13g2_o21ai_1 _21099_ (.B1(_03669_),
    .Y(_00821_),
    .A1(_10691_),
    .A2(net574));
 sg13g2_mux2_1 _21100_ (.A0(\cpu.ex.r_12[7] ),
    .A1(net710),
    .S(_03667_),
    .X(_00822_));
 sg13g2_mux2_1 _21101_ (.A0(\cpu.ex.r_12[8] ),
    .A1(net709),
    .S(_03667_),
    .X(_00823_));
 sg13g2_mux2_1 _21102_ (.A0(\cpu.ex.r_12[9] ),
    .A1(net838),
    .S(_03667_),
    .X(_00824_));
 sg13g2_inv_1 _21103_ (.Y(_03670_),
    .A(net1102));
 sg13g2_nand2_1 _21104_ (.Y(_03671_),
    .A(_03670_),
    .B(net1015));
 sg13g2_nor2_1 _21105_ (.A(_03665_),
    .B(_03671_),
    .Y(_03672_));
 sg13g2_buf_1 _21106_ (.A(_03672_),
    .X(_03673_));
 sg13g2_buf_1 _21107_ (.A(net636),
    .X(_03674_));
 sg13g2_mux2_1 _21108_ (.A0(\cpu.ex.r_13[0] ),
    .A1(net835),
    .S(net573),
    .X(_00825_));
 sg13g2_nand2_1 _21109_ (.Y(_03675_),
    .A(net963),
    .B(net636));
 sg13g2_o21ai_1 _21110_ (.B1(_03675_),
    .Y(_00826_),
    .A1(_10949_),
    .A2(net573));
 sg13g2_nand2_1 _21111_ (.Y(_03676_),
    .A(net962),
    .B(net636));
 sg13g2_o21ai_1 _21112_ (.B1(_03676_),
    .Y(_00827_),
    .A1(_10922_),
    .A2(net573));
 sg13g2_mux2_1 _21113_ (.A0(\cpu.ex.r_13[12] ),
    .A1(net450),
    .S(_03674_),
    .X(_00828_));
 sg13g2_mux2_1 _21114_ (.A0(\cpu.ex.r_13[13] ),
    .A1(net449),
    .S(_03674_),
    .X(_00829_));
 sg13g2_mux2_1 _21115_ (.A0(\cpu.ex.r_13[14] ),
    .A1(net577),
    .S(net573),
    .X(_00830_));
 sg13g2_mux2_1 _21116_ (.A0(\cpu.ex.r_13[15] ),
    .A1(net576),
    .S(net573),
    .X(_00831_));
 sg13g2_mux2_1 _21117_ (.A0(\cpu.ex.r_13[1] ),
    .A1(net502),
    .S(net573),
    .X(_00832_));
 sg13g2_mux2_1 _21118_ (.A0(\cpu.ex.r_13[2] ),
    .A1(net359),
    .S(net573),
    .X(_00833_));
 sg13g2_mux2_1 _21119_ (.A0(\cpu.ex.r_13[3] ),
    .A1(net409),
    .S(net636),
    .X(_00834_));
 sg13g2_mux2_1 _21120_ (.A0(\cpu.ex.r_13[4] ),
    .A1(net408),
    .S(_03673_),
    .X(_00835_));
 sg13g2_mux2_1 _21121_ (.A0(\cpu.ex.r_13[5] ),
    .A1(_03109_),
    .S(_03673_),
    .X(_00836_));
 sg13g2_inv_1 _21122_ (.Y(_03677_),
    .A(\cpu.ex.r_13[6] ));
 sg13g2_nand2_1 _21123_ (.Y(_03678_),
    .A(net847),
    .B(net636));
 sg13g2_o21ai_1 _21124_ (.B1(_03678_),
    .Y(_00837_),
    .A1(_03677_),
    .A2(net573));
 sg13g2_mux2_1 _21125_ (.A0(\cpu.ex.r_13[7] ),
    .A1(net710),
    .S(net636),
    .X(_00838_));
 sg13g2_mux2_1 _21126_ (.A0(\cpu.ex.r_13[8] ),
    .A1(net709),
    .S(net636),
    .X(_00839_));
 sg13g2_mux2_1 _21127_ (.A0(\cpu.ex.r_13[9] ),
    .A1(net838),
    .S(net636),
    .X(_00840_));
 sg13g2_nor2_1 _21128_ (.A(_03635_),
    .B(_03665_),
    .Y(_03679_));
 sg13g2_buf_1 _21129_ (.A(_03679_),
    .X(_03680_));
 sg13g2_buf_1 _21130_ (.A(net572),
    .X(_03681_));
 sg13g2_mux2_1 _21131_ (.A0(\cpu.ex.r_14[0] ),
    .A1(net835),
    .S(net499),
    .X(_00841_));
 sg13g2_mux2_1 _21132_ (.A0(\cpu.ex.r_14[10] ),
    .A1(net837),
    .S(net499),
    .X(_00842_));
 sg13g2_mux2_1 _21133_ (.A0(\cpu.ex.r_14[11] ),
    .A1(_03138_),
    .S(net499),
    .X(_00843_));
 sg13g2_mux2_1 _21134_ (.A0(\cpu.ex.r_14[12] ),
    .A1(net450),
    .S(_03681_),
    .X(_00844_));
 sg13g2_mux2_1 _21135_ (.A0(\cpu.ex.r_14[13] ),
    .A1(net449),
    .S(net499),
    .X(_00845_));
 sg13g2_nand2_1 _21136_ (.Y(_03682_),
    .A(net639),
    .B(net572));
 sg13g2_o21ai_1 _21137_ (.B1(_03682_),
    .Y(_00846_),
    .A1(_11061_),
    .A2(_03681_));
 sg13g2_nand2_1 _21138_ (.Y(_03683_),
    .A(net638),
    .B(_03680_));
 sg13g2_o21ai_1 _21139_ (.B1(_03683_),
    .Y(_00847_),
    .A1(_11187_),
    .A2(net499));
 sg13g2_mux2_1 _21140_ (.A0(\cpu.ex.r_14[1] ),
    .A1(net502),
    .S(net499),
    .X(_00848_));
 sg13g2_mux2_1 _21141_ (.A0(\cpu.ex.r_14[2] ),
    .A1(net359),
    .S(net499),
    .X(_00849_));
 sg13g2_mux2_1 _21142_ (.A0(\cpu.ex.r_14[3] ),
    .A1(_03655_),
    .S(net572),
    .X(_00850_));
 sg13g2_mux2_1 _21143_ (.A0(\cpu.ex.r_14[4] ),
    .A1(net408),
    .S(net572),
    .X(_00851_));
 sg13g2_mux2_1 _21144_ (.A0(\cpu.ex.r_14[5] ),
    .A1(_03109_),
    .S(net572),
    .X(_00852_));
 sg13g2_mux2_1 _21145_ (.A0(\cpu.ex.r_14[6] ),
    .A1(net711),
    .S(net572),
    .X(_00853_));
 sg13g2_nand2_1 _21146_ (.Y(_03684_),
    .A(net846),
    .B(net572));
 sg13g2_o21ai_1 _21147_ (.B1(_03684_),
    .Y(_00854_),
    .A1(_10784_),
    .A2(net499));
 sg13g2_mux2_1 _21148_ (.A0(\cpu.ex.r_14[8] ),
    .A1(net709),
    .S(net572),
    .X(_00855_));
 sg13g2_mux2_1 _21149_ (.A0(\cpu.ex.r_14[9] ),
    .A1(net838),
    .S(_03680_),
    .X(_00856_));
 sg13g2_nor2_1 _21150_ (.A(_10026_),
    .B(_03665_),
    .Y(_03685_));
 sg13g2_buf_2 _21151_ (.A(_03685_),
    .X(_03686_));
 sg13g2_buf_1 _21152_ (.A(_03686_),
    .X(_03687_));
 sg13g2_mux2_1 _21153_ (.A0(\cpu.ex.r_15[0] ),
    .A1(net835),
    .S(net571),
    .X(_00857_));
 sg13g2_mux2_1 _21154_ (.A0(\cpu.ex.r_15[10] ),
    .A1(net837),
    .S(net571),
    .X(_00858_));
 sg13g2_mux2_1 _21155_ (.A0(\cpu.ex.r_15[11] ),
    .A1(net836),
    .S(net571),
    .X(_00859_));
 sg13g2_mux2_1 _21156_ (.A0(\cpu.ex.r_15[12] ),
    .A1(net450),
    .S(net571),
    .X(_00860_));
 sg13g2_mux2_1 _21157_ (.A0(\cpu.ex.r_15[13] ),
    .A1(net449),
    .S(net571),
    .X(_00861_));
 sg13g2_mux2_1 _21158_ (.A0(\cpu.ex.r_15[14] ),
    .A1(net577),
    .S(net571),
    .X(_00862_));
 sg13g2_mux2_1 _21159_ (.A0(\cpu.ex.r_15[15] ),
    .A1(net576),
    .S(net571),
    .X(_00863_));
 sg13g2_mux2_1 _21160_ (.A0(\cpu.ex.r_15[1] ),
    .A1(net502),
    .S(_03687_),
    .X(_00864_));
 sg13g2_mux2_1 _21161_ (.A0(\cpu.ex.r_15[2] ),
    .A1(net359),
    .S(_03687_),
    .X(_00865_));
 sg13g2_mux2_1 _21162_ (.A0(\cpu.ex.r_15[3] ),
    .A1(net409),
    .S(net571),
    .X(_00866_));
 sg13g2_mux2_1 _21163_ (.A0(\cpu.ex.r_15[4] ),
    .A1(net408),
    .S(_03686_),
    .X(_00867_));
 sg13g2_buf_1 _21164_ (.A(_03107_),
    .X(_03688_));
 sg13g2_mux2_1 _21165_ (.A0(\cpu.ex.r_15[5] ),
    .A1(net570),
    .S(_03686_),
    .X(_00868_));
 sg13g2_mux2_1 _21166_ (.A0(\cpu.ex.r_15[6] ),
    .A1(net711),
    .S(_03686_),
    .X(_00869_));
 sg13g2_mux2_1 _21167_ (.A0(\cpu.ex.r_15[7] ),
    .A1(net710),
    .S(_03686_),
    .X(_00870_));
 sg13g2_mux2_1 _21168_ (.A0(\cpu.ex.r_15[8] ),
    .A1(net709),
    .S(_03686_),
    .X(_00871_));
 sg13g2_mux2_1 _21169_ (.A0(\cpu.ex.r_15[9] ),
    .A1(net838),
    .S(_03686_),
    .X(_00872_));
 sg13g2_nor3_1 _21170_ (.A(net1102),
    .B(net1015),
    .C(_03638_),
    .Y(_03689_));
 sg13g2_buf_4 _21171_ (.X(_03690_),
    .A(_03689_));
 sg13g2_buf_1 _21172_ (.A(_03690_),
    .X(_03691_));
 sg13g2_nand2_1 _21173_ (.Y(_03692_),
    .A(_03633_),
    .B(_03690_));
 sg13g2_o21ai_1 _21174_ (.B1(_03692_),
    .Y(_00873_),
    .A1(_10164_),
    .A2(_03691_));
 sg13g2_mux2_1 _21175_ (.A0(\cpu.ex.r_8[10] ),
    .A1(net837),
    .S(net498),
    .X(_00874_));
 sg13g2_mux2_1 _21176_ (.A0(\cpu.ex.r_8[11] ),
    .A1(net836),
    .S(net498),
    .X(_00875_));
 sg13g2_mux2_1 _21177_ (.A0(\cpu.ex.r_8[12] ),
    .A1(net450),
    .S(net498),
    .X(_00876_));
 sg13g2_mux2_1 _21178_ (.A0(\cpu.ex.r_8[13] ),
    .A1(net449),
    .S(_03691_),
    .X(_00877_));
 sg13g2_mux2_1 _21179_ (.A0(\cpu.ex.r_8[14] ),
    .A1(_03647_),
    .S(net498),
    .X(_00878_));
 sg13g2_mux2_1 _21180_ (.A0(\cpu.ex.r_8[15] ),
    .A1(_03649_),
    .S(net498),
    .X(_00879_));
 sg13g2_mux2_1 _21181_ (.A0(\cpu.ex.r_8[1] ),
    .A1(_03652_),
    .S(net498),
    .X(_00880_));
 sg13g2_mux2_1 _21182_ (.A0(\cpu.ex.r_8[2] ),
    .A1(net359),
    .S(net498),
    .X(_00881_));
 sg13g2_mux2_1 _21183_ (.A0(\cpu.ex.r_8[3] ),
    .A1(net409),
    .S(net498),
    .X(_00882_));
 sg13g2_mux2_1 _21184_ (.A0(\cpu.ex.r_8[4] ),
    .A1(net408),
    .S(_03690_),
    .X(_00883_));
 sg13g2_mux2_1 _21185_ (.A0(\cpu.ex.r_8[5] ),
    .A1(net570),
    .S(_03690_),
    .X(_00884_));
 sg13g2_mux2_1 _21186_ (.A0(\cpu.ex.r_8[6] ),
    .A1(net711),
    .S(_03690_),
    .X(_00885_));
 sg13g2_mux2_1 _21187_ (.A0(\cpu.ex.r_8[7] ),
    .A1(net710),
    .S(_03690_),
    .X(_00886_));
 sg13g2_mux2_1 _21188_ (.A0(\cpu.ex.r_8[8] ),
    .A1(_03135_),
    .S(_03690_),
    .X(_00887_));
 sg13g2_mux2_1 _21189_ (.A0(\cpu.ex.r_8[9] ),
    .A1(_03136_),
    .S(_03690_),
    .X(_00888_));
 sg13g2_nor2_1 _21190_ (.A(_03638_),
    .B(_03671_),
    .Y(_03693_));
 sg13g2_buf_4 _21191_ (.X(_03694_),
    .A(_03693_));
 sg13g2_buf_1 _21192_ (.A(_03694_),
    .X(_03695_));
 sg13g2_mux2_1 _21193_ (.A0(\cpu.ex.r_9[0] ),
    .A1(net835),
    .S(net497),
    .X(_00889_));
 sg13g2_mux2_1 _21194_ (.A0(\cpu.ex.r_9[10] ),
    .A1(net837),
    .S(net497),
    .X(_00890_));
 sg13g2_mux2_1 _21195_ (.A0(\cpu.ex.r_9[11] ),
    .A1(net836),
    .S(net497),
    .X(_00891_));
 sg13g2_buf_1 _21196_ (.A(net589),
    .X(_03696_));
 sg13g2_mux2_1 _21197_ (.A0(\cpu.ex.r_9[12] ),
    .A1(net496),
    .S(net497),
    .X(_00892_));
 sg13g2_buf_1 _21198_ (.A(net503),
    .X(_03697_));
 sg13g2_mux2_1 _21199_ (.A0(\cpu.ex.r_9[13] ),
    .A1(net447),
    .S(net497),
    .X(_00893_));
 sg13g2_mux2_1 _21200_ (.A0(\cpu.ex.r_9[14] ),
    .A1(_03647_),
    .S(_03695_),
    .X(_00894_));
 sg13g2_mux2_1 _21201_ (.A0(\cpu.ex.r_9[15] ),
    .A1(_03649_),
    .S(net497),
    .X(_00895_));
 sg13g2_mux2_1 _21202_ (.A0(\cpu.ex.r_9[1] ),
    .A1(net502),
    .S(_03695_),
    .X(_00896_));
 sg13g2_mux2_1 _21203_ (.A0(\cpu.ex.r_9[2] ),
    .A1(net359),
    .S(net497),
    .X(_00897_));
 sg13g2_mux2_1 _21204_ (.A0(\cpu.ex.r_9[3] ),
    .A1(net409),
    .S(_03694_),
    .X(_00898_));
 sg13g2_mux2_1 _21205_ (.A0(\cpu.ex.r_9[4] ),
    .A1(net408),
    .S(_03694_),
    .X(_00899_));
 sg13g2_mux2_1 _21206_ (.A0(\cpu.ex.r_9[5] ),
    .A1(net570),
    .S(_03694_),
    .X(_00900_));
 sg13g2_nand2_1 _21207_ (.Y(_03698_),
    .A(net847),
    .B(_03694_));
 sg13g2_o21ai_1 _21208_ (.B1(_03698_),
    .Y(_00901_),
    .A1(_10683_),
    .A2(net497));
 sg13g2_mux2_1 _21209_ (.A0(\cpu.ex.r_9[7] ),
    .A1(net710),
    .S(_03694_),
    .X(_00902_));
 sg13g2_mux2_1 _21210_ (.A0(\cpu.ex.r_9[8] ),
    .A1(net709),
    .S(_03694_),
    .X(_00903_));
 sg13g2_mux2_1 _21211_ (.A0(\cpu.ex.r_9[9] ),
    .A1(net838),
    .S(_03694_),
    .X(_00904_));
 sg13g2_nor2_1 _21212_ (.A(net1103),
    .B(_10021_),
    .Y(_03699_));
 sg13g2_nand4_1 _21213_ (.B(net1015),
    .C(_10017_),
    .A(net1102),
    .Y(_03700_),
    .D(_03699_));
 sg13g2_nor2_1 _21214_ (.A(_08132_),
    .B(_03700_),
    .Y(_03701_));
 sg13g2_buf_2 _21215_ (.A(_03701_),
    .X(_03702_));
 sg13g2_buf_1 _21216_ (.A(_03702_),
    .X(_03703_));
 sg13g2_mux2_1 _21217_ (.A0(\cpu.ex.r_epc[1] ),
    .A1(_03652_),
    .S(_03703_),
    .X(_00906_));
 sg13g2_mux2_1 _21218_ (.A0(\cpu.ex.r_epc[11] ),
    .A1(net836),
    .S(net569),
    .X(_00907_));
 sg13g2_mux2_1 _21219_ (.A0(\cpu.ex.r_epc[12] ),
    .A1(net496),
    .S(net569),
    .X(_00908_));
 sg13g2_mux2_1 _21220_ (.A0(\cpu.ex.r_epc[13] ),
    .A1(net447),
    .S(net569),
    .X(_00909_));
 sg13g2_nand2_1 _21221_ (.Y(_03704_),
    .A(net639),
    .B(_03702_));
 sg13g2_o21ai_1 _21222_ (.B1(_03704_),
    .Y(_00910_),
    .A1(_11074_),
    .A2(net569));
 sg13g2_buf_1 _21223_ (.A(net731),
    .X(_03705_));
 sg13g2_mux2_1 _21224_ (.A0(\cpu.ex.r_epc[15] ),
    .A1(net635),
    .S(_03703_),
    .X(_00911_));
 sg13g2_mux2_1 _21225_ (.A0(\cpu.ex.r_epc[2] ),
    .A1(net359),
    .S(net569),
    .X(_00912_));
 sg13g2_mux2_1 _21226_ (.A0(\cpu.ex.r_epc[3] ),
    .A1(_03655_),
    .S(net569),
    .X(_00913_));
 sg13g2_mux2_1 _21227_ (.A0(\cpu.ex.r_epc[4] ),
    .A1(_03658_),
    .S(net569),
    .X(_00914_));
 sg13g2_mux2_1 _21228_ (.A0(\cpu.ex.r_epc[5] ),
    .A1(net570),
    .S(net569),
    .X(_00915_));
 sg13g2_mux2_1 _21229_ (.A0(\cpu.ex.r_epc[6] ),
    .A1(net711),
    .S(_03702_),
    .X(_00916_));
 sg13g2_mux2_1 _21230_ (.A0(\cpu.ex.r_epc[7] ),
    .A1(net710),
    .S(_03702_),
    .X(_00917_));
 sg13g2_mux2_1 _21231_ (.A0(\cpu.ex.r_epc[8] ),
    .A1(net709),
    .S(_03702_),
    .X(_00918_));
 sg13g2_mux2_1 _21232_ (.A0(\cpu.ex.r_epc[9] ),
    .A1(net838),
    .S(_03702_),
    .X(_00919_));
 sg13g2_mux2_1 _21233_ (.A0(\cpu.ex.r_epc[10] ),
    .A1(net837),
    .S(_03702_),
    .X(_00920_));
 sg13g2_nand4_1 _21234_ (.B(net1015),
    .C(_10017_),
    .A(_03670_),
    .Y(_03706_),
    .D(_03699_));
 sg13g2_buf_1 _21235_ (.A(_03706_),
    .X(_03707_));
 sg13g2_buf_1 _21236_ (.A(_03707_),
    .X(_03708_));
 sg13g2_buf_1 _21237_ (.A(_03707_),
    .X(_03709_));
 sg13g2_nand2_1 _21238_ (.Y(_03710_),
    .A(\cpu.ex.r_lr[1] ),
    .B(net633));
 sg13g2_o21ai_1 _21239_ (.B1(_03710_),
    .Y(_00926_),
    .A1(net673),
    .A2(net634));
 sg13g2_mux2_1 _21240_ (.A0(net842),
    .A1(\cpu.ex.r_lr[11] ),
    .S(net634),
    .X(_00927_));
 sg13g2_buf_1 _21241_ (.A(net504),
    .X(_03711_));
 sg13g2_mux2_1 _21242_ (.A0(net446),
    .A1(\cpu.ex.r_lr[12] ),
    .S(net634),
    .X(_00928_));
 sg13g2_buf_1 _21243_ (.A(net503),
    .X(_03712_));
 sg13g2_mux2_1 _21244_ (.A0(_03712_),
    .A1(\cpu.ex.r_lr[13] ),
    .S(net634),
    .X(_00929_));
 sg13g2_buf_1 _21245_ (.A(net639),
    .X(_03713_));
 sg13g2_mux2_1 _21246_ (.A0(_03713_),
    .A1(\cpu.ex.r_lr[14] ),
    .S(net634),
    .X(_00930_));
 sg13g2_buf_1 _21247_ (.A(net638),
    .X(_03714_));
 sg13g2_mux2_1 _21248_ (.A0(net567),
    .A1(\cpu.ex.r_lr[15] ),
    .S(net634),
    .X(_00931_));
 sg13g2_nand2_1 _21249_ (.Y(_03715_),
    .A(\cpu.ex.r_lr[2] ),
    .B(_03709_));
 sg13g2_o21ai_1 _21250_ (.B1(_03715_),
    .Y(_00932_),
    .A1(net644),
    .A2(_03708_));
 sg13g2_nand2_1 _21251_ (.Y(_03716_),
    .A(\cpu.ex.r_lr[3] ),
    .B(_03709_));
 sg13g2_o21ai_1 _21252_ (.B1(_03716_),
    .Y(_00933_),
    .A1(net781),
    .A2(_03708_));
 sg13g2_buf_1 _21253_ (.A(net645),
    .X(_03717_));
 sg13g2_buf_1 _21254_ (.A(net566),
    .X(_03718_));
 sg13g2_nand2_1 _21255_ (.Y(_03719_),
    .A(\cpu.ex.r_lr[4] ),
    .B(net633));
 sg13g2_o21ai_1 _21256_ (.B1(_03719_),
    .Y(_00934_),
    .A1(_03718_),
    .A2(net634));
 sg13g2_nand2_1 _21257_ (.Y(_03720_),
    .A(\cpu.ex.r_lr[5] ),
    .B(net633));
 sg13g2_o21ai_1 _21258_ (.B1(_03720_),
    .Y(_00935_),
    .A1(net641),
    .A2(net634));
 sg13g2_mux2_1 _21259_ (.A0(_03095_),
    .A1(\cpu.ex.r_lr[6] ),
    .S(net633),
    .X(_00936_));
 sg13g2_mux2_1 _21260_ (.A0(net716),
    .A1(\cpu.ex.r_lr[7] ),
    .S(net633),
    .X(_00937_));
 sg13g2_mux2_1 _21261_ (.A0(net715),
    .A1(\cpu.ex.r_lr[8] ),
    .S(net633),
    .X(_00938_));
 sg13g2_mux2_1 _21262_ (.A0(_03102_),
    .A1(\cpu.ex.r_lr[9] ),
    .S(net633),
    .X(_00939_));
 sg13g2_mux2_1 _21263_ (.A0(net843),
    .A1(\cpu.ex.r_lr[10] ),
    .S(net633),
    .X(_00940_));
 sg13g2_buf_1 _21264_ (.A(_10348_),
    .X(_03721_));
 sg13g2_buf_8 _21265_ (.A(_11462_),
    .X(_03722_));
 sg13g2_nor2_1 _21266_ (.A(net293),
    .B(_03722_),
    .Y(_03723_));
 sg13g2_xnor2_1 _21267_ (.Y(_03724_),
    .A(net72),
    .B(_03723_));
 sg13g2_nor2_1 _21268_ (.A(net202),
    .B(_11071_),
    .Y(_03725_));
 sg13g2_nor2_1 _21269_ (.A(_11860_),
    .B(_11840_),
    .Y(_03726_));
 sg13g2_o21ai_1 _21270_ (.B1(_03726_),
    .Y(_03727_),
    .A1(net78),
    .A2(_03725_));
 sg13g2_mux2_1 _21271_ (.A0(_11860_),
    .A1(_11862_),
    .S(net199),
    .X(_03728_));
 sg13g2_a221oi_1 _21272_ (.B2(_11847_),
    .C1(_11072_),
    .B1(_03728_),
    .A1(_11323_),
    .Y(_03729_),
    .A2(_11213_));
 sg13g2_nand3_1 _21273_ (.B(_11213_),
    .C(_11855_),
    .A(_11860_),
    .Y(_03730_));
 sg13g2_nand2_1 _21274_ (.Y(_03731_),
    .A(_11072_),
    .B(_03730_));
 sg13g2_nand3b_1 _21275_ (.B(_03731_),
    .C(_11470_),
    .Y(_03732_),
    .A_N(_03729_));
 sg13g2_nand2_1 _21276_ (.Y(_03733_),
    .A(_03727_),
    .B(_03732_));
 sg13g2_nand2_1 _21277_ (.Y(_03734_),
    .A(\cpu.ex.r_mult[15] ),
    .B(net683));
 sg13g2_or2_1 _21278_ (.X(_03735_),
    .B(_03734_),
    .A(net78));
 sg13g2_nor3_1 _21279_ (.A(_11836_),
    .B(_11837_),
    .C(_03735_),
    .Y(_03736_));
 sg13g2_a21oi_1 _21280_ (.A1(_03727_),
    .A2(_03732_),
    .Y(_03737_),
    .B1(_03734_));
 sg13g2_nand2_1 _21281_ (.Y(_03738_),
    .A(_11794_),
    .B(_11071_));
 sg13g2_a21oi_1 _21282_ (.A1(_11860_),
    .A2(net199),
    .Y(_03739_),
    .B1(_03738_));
 sg13g2_nor2_1 _21283_ (.A(_11860_),
    .B(net199),
    .Y(_03740_));
 sg13g2_o21ai_1 _21284_ (.B1(net587),
    .Y(_03741_),
    .A1(_03739_),
    .A2(_03740_));
 sg13g2_nor2_1 _21285_ (.A(_03741_),
    .B(_03735_),
    .Y(_03742_));
 sg13g2_a221oi_1 _21286_ (.B2(_11834_),
    .C1(_03742_),
    .B1(_03737_),
    .A1(_03733_),
    .Y(_03743_),
    .A2(_03736_));
 sg13g2_buf_8 _21287_ (.A(_03743_),
    .X(_03744_));
 sg13g2_o21ai_1 _21288_ (.B1(_03733_),
    .Y(_03745_),
    .A1(_11834_),
    .A2(_11838_));
 sg13g2_inv_1 _21289_ (.Y(_03746_),
    .A(_03741_));
 sg13g2_a22oi_1 _21290_ (.Y(_03747_),
    .B1(net73),
    .B2(_03746_),
    .A2(_11546_),
    .A1(\cpu.ex.r_mult[15] ));
 sg13g2_a21oi_1 _21291_ (.A1(_03745_),
    .A2(_03747_),
    .Y(_03748_),
    .B1(_11475_));
 sg13g2_a22oi_1 _21292_ (.Y(_03749_),
    .B1(_03744_),
    .B2(_03748_),
    .A2(_11621_),
    .A1(_10153_));
 sg13g2_nand2_1 _21293_ (.Y(_03750_),
    .A(net835),
    .B(net597));
 sg13g2_o21ai_1 _21294_ (.B1(_03750_),
    .Y(_03751_),
    .A1(_11465_),
    .A2(_03749_));
 sg13g2_a21o_1 _21295_ (.A2(_03724_),
    .A1(_11661_),
    .B1(_03751_),
    .X(_00941_));
 sg13g2_buf_1 _21296_ (.A(_10349_),
    .X(_03752_));
 sg13g2_buf_1 _21297_ (.A(net292),
    .X(_03753_));
 sg13g2_nor3_1 _21298_ (.A(net293),
    .B(net73),
    .C(_03753_),
    .Y(_03754_));
 sg13g2_a21oi_1 _21299_ (.A1(net245),
    .A2(net72),
    .Y(_03755_),
    .B1(net244));
 sg13g2_nor3_1 _21300_ (.A(_11462_),
    .B(_03754_),
    .C(_03755_),
    .Y(_03756_));
 sg13g2_xnor2_1 _21301_ (.Y(_03757_),
    .A(_11370_),
    .B(_03756_));
 sg13g2_inv_1 _21302_ (.Y(_03758_),
    .A(_10153_));
 sg13g2_and2_1 _21303_ (.A(_03758_),
    .B(_03744_),
    .X(_03759_));
 sg13g2_nor2_1 _21304_ (.A(_03758_),
    .B(_03744_),
    .Y(_03760_));
 sg13g2_nor3_1 _21305_ (.A(_11633_),
    .B(_03759_),
    .C(_03760_),
    .Y(_03761_));
 sg13g2_a221oi_1 _21306_ (.B2(net79),
    .C1(_03761_),
    .B1(_03757_),
    .A1(net1000),
    .Y(_03762_),
    .A2(_11621_));
 sg13g2_buf_1 _21307_ (.A(net597),
    .X(_03763_));
 sg13g2_nand2_1 _21308_ (.Y(_03764_),
    .A(net575),
    .B(net494));
 sg13g2_o21ai_1 _21309_ (.B1(_03764_),
    .Y(_00942_),
    .A1(net458),
    .A2(_03762_));
 sg13g2_and2_1 _21310_ (.A(_11394_),
    .B(net241),
    .X(_03765_));
 sg13g2_nor2_1 _21311_ (.A(_11394_),
    .B(net241),
    .Y(_03766_));
 sg13g2_nor3_1 _21312_ (.A(net29),
    .B(_03765_),
    .C(_03766_),
    .Y(_03767_));
 sg13g2_xor2_1 _21313_ (.B(_03767_),
    .A(_11396_),
    .X(_03768_));
 sg13g2_buf_1 _21314_ (.A(_11557_),
    .X(_03769_));
 sg13g2_xnor2_1 _21315_ (.Y(_03770_),
    .A(net1000),
    .B(_03760_));
 sg13g2_nor2_1 _21316_ (.A(_11817_),
    .B(_03770_),
    .Y(_03771_));
 sg13g2_a221oi_1 _21317_ (.B2(net999),
    .C1(_03771_),
    .B1(_03769_),
    .A1(net410),
    .Y(_03772_),
    .A2(_03763_));
 sg13g2_o21ai_1 _21318_ (.B1(_03772_),
    .Y(_00943_),
    .A1(_11818_),
    .A2(_03768_));
 sg13g2_nand2_1 _21319_ (.Y(_03773_),
    .A(net464),
    .B(net597));
 sg13g2_nand2_1 _21320_ (.Y(_03774_),
    .A(net999),
    .B(_11418_));
 sg13g2_o21ai_1 _21321_ (.B1(net1000),
    .Y(_03775_),
    .A1(_11394_),
    .A2(net241));
 sg13g2_a21oi_1 _21322_ (.A1(_11394_),
    .A2(net241),
    .Y(_03776_),
    .B1(net1000));
 sg13g2_o21ai_1 _21323_ (.B1(net999),
    .Y(_03777_),
    .A1(_03766_),
    .A2(_03776_));
 sg13g2_o21ai_1 _21324_ (.B1(_03777_),
    .Y(_03778_),
    .A1(net999),
    .A2(_03775_));
 sg13g2_a22oi_1 _21325_ (.Y(_03779_),
    .B1(_03778_),
    .B2(net523),
    .A2(_03765_),
    .A1(_03774_));
 sg13g2_xnor2_1 _21326_ (.Y(_03780_),
    .A(_11584_),
    .B(_03779_));
 sg13g2_nand2_1 _21327_ (.Y(_03781_),
    .A(_11402_),
    .B(net29));
 sg13g2_o21ai_1 _21328_ (.B1(_03781_),
    .Y(_03782_),
    .A1(net29),
    .A2(_03780_));
 sg13g2_inv_1 _21329_ (.Y(_03783_),
    .A(net1000));
 sg13g2_nor3_1 _21330_ (.A(_03758_),
    .B(_03783_),
    .C(_03744_),
    .Y(_03784_));
 sg13g2_xnor2_1 _21331_ (.Y(_03785_),
    .A(net999),
    .B(_03784_));
 sg13g2_o21ai_1 _21332_ (.B1(_11556_),
    .Y(_03786_),
    .A1(_11633_),
    .A2(_03785_));
 sg13g2_a21oi_1 _21333_ (.A1(net79),
    .A2(_03782_),
    .Y(_03787_),
    .B1(_03786_));
 sg13g2_and2_1 _21334_ (.A(net458),
    .B(_03773_),
    .X(_03788_));
 sg13g2_a221oi_1 _21335_ (.B2(_03787_),
    .C1(_03788_),
    .B1(_03773_),
    .A1(_11297_),
    .Y(_00944_),
    .A2(net358));
 sg13g2_inv_1 _21336_ (.Y(_03789_),
    .A(net1002));
 sg13g2_o21ai_1 _21337_ (.B1(_11394_),
    .Y(_03790_),
    .A1(_11411_),
    .A2(_11407_));
 sg13g2_buf_1 _21338_ (.A(_03790_),
    .X(_03791_));
 sg13g2_nand2_1 _21339_ (.Y(_03792_),
    .A(_03791_),
    .B(_11414_));
 sg13g2_nor2_1 _21340_ (.A(net302),
    .B(_03792_),
    .Y(_03793_));
 sg13g2_a21oi_1 _21341_ (.A1(_03791_),
    .A2(_11414_),
    .Y(_03794_),
    .B1(net247));
 sg13g2_nor3_1 _21342_ (.A(net29),
    .B(_03793_),
    .C(_03794_),
    .Y(_03795_));
 sg13g2_nand2_1 _21343_ (.Y(_03796_),
    .A(net1001),
    .B(_11418_));
 sg13g2_xnor2_1 _21344_ (.Y(_03797_),
    .A(_03795_),
    .B(_03796_));
 sg13g2_nand2_1 _21345_ (.Y(_03798_),
    .A(net71),
    .B(_03797_));
 sg13g2_nor2_1 _21346_ (.A(net458),
    .B(_11633_),
    .Y(_03799_));
 sg13g2_nand3_1 _21347_ (.B(net1000),
    .C(net999),
    .A(_10153_),
    .Y(_03800_));
 sg13g2_buf_1 _21348_ (.A(_03800_),
    .X(_03801_));
 sg13g2_nor2_1 _21349_ (.A(_03744_),
    .B(_03801_),
    .Y(_03802_));
 sg13g2_xnor2_1 _21350_ (.Y(_03803_),
    .A(_11297_),
    .B(_03802_));
 sg13g2_a221oi_1 _21351_ (.B2(_03803_),
    .C1(net358),
    .B1(_03799_),
    .A1(net448),
    .Y(_03804_),
    .A2(net597));
 sg13g2_a22oi_1 _21352_ (.Y(_00945_),
    .B1(_03798_),
    .B2(_03804_),
    .A2(net358),
    .A1(_03789_));
 sg13g2_nand2_1 _21353_ (.Y(_03805_),
    .A(net1001),
    .B(_03802_));
 sg13g2_xnor2_1 _21354_ (.Y(_03806_),
    .A(net1002),
    .B(_03805_));
 sg13g2_a22oi_1 _21355_ (.Y(_03807_),
    .B1(_11815_),
    .B2(_03806_),
    .A2(_11621_),
    .A1(net1003));
 sg13g2_nor2_1 _21356_ (.A(_11297_),
    .B(_10576_),
    .Y(_03808_));
 sg13g2_nand2_1 _21357_ (.Y(_03809_),
    .A(_10240_),
    .B(_11404_));
 sg13g2_nor2_1 _21358_ (.A(_03758_),
    .B(net370),
    .Y(_03810_));
 sg13g2_o21ai_1 _21359_ (.B1(_03810_),
    .Y(_03811_),
    .A1(_10240_),
    .A2(_11404_));
 sg13g2_a21oi_1 _21360_ (.A1(_03809_),
    .A2(_03811_),
    .Y(_03812_),
    .B1(net301));
 sg13g2_nor2_1 _21361_ (.A(net1001),
    .B(net302),
    .Y(_03813_));
 sg13g2_nor2_1 _21362_ (.A(_09153_),
    .B(_03813_),
    .Y(_03814_));
 sg13g2_a21oi_1 _21363_ (.A1(_10240_),
    .A2(net299),
    .Y(_03815_),
    .B1(net372));
 sg13g2_o21ai_1 _21364_ (.B1(_11402_),
    .Y(_03816_),
    .A1(_11275_),
    .A2(net302));
 sg13g2_a21oi_1 _21365_ (.A1(_03811_),
    .A2(_03815_),
    .Y(_03817_),
    .B1(_03816_));
 sg13g2_a221oi_1 _21366_ (.B2(_03814_),
    .C1(_03817_),
    .B1(_03812_),
    .A1(net652),
    .Y(_03818_),
    .A2(_03808_));
 sg13g2_and4_1 _21367_ (.A(net374),
    .B(_11468_),
    .C(_11391_),
    .D(_03818_),
    .X(_03819_));
 sg13g2_buf_1 _21368_ (.A(_03819_),
    .X(_03820_));
 sg13g2_o21ai_1 _21369_ (.B1(_09146_),
    .Y(_03821_),
    .A1(_11395_),
    .A2(net1001));
 sg13g2_and3_1 _21370_ (.X(_03822_),
    .A(net302),
    .B(net299),
    .C(_03821_));
 sg13g2_xnor2_1 _21371_ (.Y(_03823_),
    .A(_11395_),
    .B(net299));
 sg13g2_nor4_1 _21372_ (.A(_03808_),
    .B(_03813_),
    .C(_03821_),
    .D(_03823_),
    .Y(_03824_));
 sg13g2_or2_1 _21373_ (.X(_03825_),
    .B(_03824_),
    .A(_03822_));
 sg13g2_xnor2_1 _21374_ (.Y(_03826_),
    .A(net999),
    .B(net301));
 sg13g2_nor2_1 _21375_ (.A(_03758_),
    .B(net292),
    .Y(_03827_));
 sg13g2_and4_1 _21376_ (.A(_03758_),
    .B(_11409_),
    .C(_10349_),
    .D(net301),
    .X(_03828_));
 sg13g2_a21oi_1 _21377_ (.A1(_03826_),
    .A2(_03827_),
    .Y(_03829_),
    .B1(_03828_));
 sg13g2_o21ai_1 _21378_ (.B1(_11248_),
    .Y(_03830_),
    .A1(_10153_),
    .A2(_11409_));
 sg13g2_nand3_1 _21379_ (.B(net372),
    .C(_03830_),
    .A(net292),
    .Y(_03831_));
 sg13g2_o21ai_1 _21380_ (.B1(_03831_),
    .Y(_03832_),
    .A1(_09153_),
    .A2(_03829_));
 sg13g2_a21o_1 _21381_ (.A2(_03808_),
    .A1(net652),
    .B1(_03817_),
    .X(_03833_));
 sg13g2_a221oi_1 _21382_ (.B2(_03832_),
    .C1(_03833_),
    .B1(_03825_),
    .A1(_03812_),
    .Y(_03834_),
    .A2(_03814_));
 sg13g2_and3_1 _21383_ (.X(_03835_),
    .A(_11466_),
    .B(_11368_),
    .C(_03818_));
 sg13g2_buf_1 _21384_ (.A(_03835_),
    .X(_03836_));
 sg13g2_nor3_2 _21385_ (.A(_03820_),
    .B(_03834_),
    .C(_03836_),
    .Y(_03837_));
 sg13g2_nor2_1 _21386_ (.A(net246),
    .B(_03837_),
    .Y(_03838_));
 sg13g2_nor4_2 _21387_ (.A(net230),
    .B(_03820_),
    .C(_03834_),
    .Y(_03839_),
    .D(_03836_));
 sg13g2_nor3_1 _21388_ (.A(_11462_),
    .B(_03838_),
    .C(_03839_),
    .Y(_03840_));
 sg13g2_nand2_1 _21389_ (.Y(_03841_),
    .A(net1002),
    .B(net588));
 sg13g2_xnor2_1 _21390_ (.Y(_03842_),
    .A(_03840_),
    .B(_03841_));
 sg13g2_a21oi_1 _21391_ (.A1(net79),
    .A2(_03842_),
    .Y(_03843_),
    .B1(net494));
 sg13g2_a221oi_1 _21392_ (.B2(_03843_),
    .C1(_10031_),
    .B1(_03807_),
    .A1(net718),
    .Y(_00946_),
    .A2(net494));
 sg13g2_o21ai_1 _21393_ (.B1(_11270_),
    .Y(_03844_),
    .A1(net246),
    .A2(_03794_));
 sg13g2_nand3_1 _21394_ (.B(_03791_),
    .C(_11414_),
    .A(net247),
    .Y(_03845_));
 sg13g2_nor2_1 _21395_ (.A(_11272_),
    .B(_03796_),
    .Y(_03846_));
 sg13g2_a22oi_1 _21396_ (.Y(_03847_),
    .B1(_03845_),
    .B2(_03846_),
    .A2(_03792_),
    .A1(_11300_));
 sg13g2_o21ai_1 _21397_ (.B1(_03847_),
    .Y(_03848_),
    .A1(net651),
    .A2(_03844_));
 sg13g2_xnor2_1 _21398_ (.Y(_03849_),
    .A(net198),
    .B(_03848_));
 sg13g2_nor2_1 _21399_ (.A(net29),
    .B(_03849_),
    .Y(_03850_));
 sg13g2_nor2_1 _21400_ (.A(_11286_),
    .B(net651),
    .Y(_03851_));
 sg13g2_xnor2_1 _21401_ (.Y(_03852_),
    .A(_03850_),
    .B(_03851_));
 sg13g2_nor4_1 _21402_ (.A(_11297_),
    .B(_03789_),
    .C(_03744_),
    .D(_03801_),
    .Y(_03853_));
 sg13g2_buf_2 _21403_ (.A(_03853_),
    .X(_03854_));
 sg13g2_xnor2_1 _21404_ (.Y(_03855_),
    .A(net1003),
    .B(_03854_));
 sg13g2_nor2_1 _21405_ (.A(_11817_),
    .B(_03855_),
    .Y(_03856_));
 sg13g2_a221oi_1 _21406_ (.B2(net1096),
    .C1(_03856_),
    .B1(net358),
    .A1(_03094_),
    .Y(_03857_),
    .A2(net494));
 sg13g2_o21ai_1 _21407_ (.B1(_03857_),
    .Y(_00947_),
    .A1(_11818_),
    .A2(_03852_));
 sg13g2_a22oi_1 _21408_ (.Y(_03858_),
    .B1(net358),
    .B2(net1004),
    .A2(net494),
    .A1(net846));
 sg13g2_nand2_1 _21409_ (.Y(_03859_),
    .A(net1003),
    .B(_03854_));
 sg13g2_xnor2_1 _21410_ (.Y(_03860_),
    .A(net1096),
    .B(_03859_));
 sg13g2_nand2_1 _21411_ (.Y(_03861_),
    .A(net1096),
    .B(net523));
 sg13g2_nand2_1 _21412_ (.Y(_03862_),
    .A(net198),
    .B(_03839_));
 sg13g2_nor2_1 _21413_ (.A(net201),
    .B(_03841_),
    .Y(_03863_));
 sg13g2_a22oi_1 _21414_ (.Y(_03864_),
    .B1(_03863_),
    .B2(_03837_),
    .A2(_03851_),
    .A1(_03839_));
 sg13g2_nor3_1 _21415_ (.A(_03789_),
    .B(_11286_),
    .C(net651),
    .Y(_03865_));
 sg13g2_nand2_1 _21416_ (.Y(_03866_),
    .A(net224),
    .B(net246));
 sg13g2_a22oi_1 _21417_ (.Y(_03867_),
    .B1(_03865_),
    .B2(net246),
    .A2(_03851_),
    .A1(net224));
 sg13g2_o21ai_1 _21418_ (.B1(_03867_),
    .Y(_03868_),
    .A1(_03841_),
    .A2(_03866_));
 sg13g2_a21oi_1 _21419_ (.A1(_03837_),
    .A2(_03865_),
    .Y(_03869_),
    .B1(_03868_));
 sg13g2_nand3_1 _21420_ (.B(_03864_),
    .C(_03869_),
    .A(_03862_),
    .Y(_03870_));
 sg13g2_xnor2_1 _21421_ (.Y(_03871_),
    .A(net228),
    .B(_03870_));
 sg13g2_nor2_1 _21422_ (.A(net29),
    .B(_03871_),
    .Y(_03872_));
 sg13g2_xnor2_1 _21423_ (.Y(_03873_),
    .A(_03861_),
    .B(_03872_));
 sg13g2_a22oi_1 _21424_ (.Y(_03874_),
    .B1(_03873_),
    .B2(net71),
    .A2(_03860_),
    .A1(_03799_));
 sg13g2_nand2_1 _21425_ (.Y(_00948_),
    .A(_03858_),
    .B(_03874_));
 sg13g2_nand2_1 _21426_ (.Y(_03875_),
    .A(net1004),
    .B(net521));
 sg13g2_nand2_1 _21427_ (.Y(_03876_),
    .A(_10725_),
    .B(net587));
 sg13g2_nand3_1 _21428_ (.B(net1002),
    .C(net1003),
    .A(net1001),
    .Y(_03877_));
 sg13g2_nor4_2 _21429_ (.A(_03744_),
    .B(_03801_),
    .C(_03876_),
    .Y(_03878_),
    .D(_03877_));
 sg13g2_nand2_1 _21430_ (.Y(_03879_),
    .A(_11308_),
    .B(_03878_));
 sg13g2_o21ai_1 _21431_ (.B1(_03879_),
    .Y(_03880_),
    .A1(_03875_),
    .A2(_03878_));
 sg13g2_a21oi_1 _21432_ (.A1(_03791_),
    .A2(_11414_),
    .Y(_03881_),
    .B1(_11303_));
 sg13g2_nor2_1 _21433_ (.A(_11320_),
    .B(_03881_),
    .Y(_03882_));
 sg13g2_xnor2_1 _21434_ (.Y(_03883_),
    .A(net226),
    .B(_03882_));
 sg13g2_nor2_1 _21435_ (.A(_11462_),
    .B(_03883_),
    .Y(_03884_));
 sg13g2_nand2_1 _21436_ (.Y(_03885_),
    .A(net1004),
    .B(net588));
 sg13g2_xnor2_1 _21437_ (.Y(_03886_),
    .A(_03884_),
    .B(_03885_));
 sg13g2_nor2_1 _21438_ (.A(_11306_),
    .B(_11556_),
    .Y(_03887_));
 sg13g2_a221oi_1 _21439_ (.B2(net79),
    .C1(_03887_),
    .B1(_03886_),
    .A1(net997),
    .Y(_03888_),
    .A2(_03880_));
 sg13g2_nand2_1 _21440_ (.Y(_03889_),
    .A(net845),
    .B(net494));
 sg13g2_o21ai_1 _21441_ (.B1(_03889_),
    .Y(_00949_),
    .A1(net458),
    .A2(_03888_));
 sg13g2_nand2b_1 _21442_ (.Y(_03890_),
    .B(net228),
    .A_N(_03861_));
 sg13g2_nand4_1 _21443_ (.B(_03864_),
    .C(_03869_),
    .A(_03862_),
    .Y(_03891_),
    .D(_03890_));
 sg13g2_buf_2 _21444_ (.A(_03891_),
    .X(_03892_));
 sg13g2_nor2_1 _21445_ (.A(_11243_),
    .B(net205),
    .Y(_03893_));
 sg13g2_nor2_1 _21446_ (.A(_03861_),
    .B(_03893_),
    .Y(_03894_));
 sg13g2_o21ai_1 _21447_ (.B1(_11270_),
    .Y(_03895_),
    .A1(net1003),
    .A2(net198));
 sg13g2_inv_1 _21448_ (.Y(_03896_),
    .A(_03895_));
 sg13g2_o21ai_1 _21449_ (.B1(_03896_),
    .Y(_03897_),
    .A1(net246),
    .A2(_03837_));
 sg13g2_nand2_1 _21450_ (.Y(_03898_),
    .A(net1003),
    .B(net198));
 sg13g2_o21ai_1 _21451_ (.B1(_03839_),
    .Y(_03899_),
    .A1(net1003),
    .A2(net198));
 sg13g2_nand3_1 _21452_ (.B(_03898_),
    .C(_03899_),
    .A(_03897_),
    .Y(_03900_));
 sg13g2_nor2_1 _21453_ (.A(net223),
    .B(_03885_),
    .Y(_03901_));
 sg13g2_a22oi_1 _21454_ (.Y(_03902_),
    .B1(_03900_),
    .B2(_03901_),
    .A2(_03894_),
    .A1(_03892_));
 sg13g2_inv_1 _21455_ (.Y(_03903_),
    .A(_03885_));
 sg13g2_nor2_1 _21456_ (.A(net226),
    .B(net223),
    .Y(_03904_));
 sg13g2_a22oi_1 _21457_ (.Y(_03905_),
    .B1(_03892_),
    .B2(_03904_),
    .A2(_03903_),
    .A1(net205));
 sg13g2_a21o_1 _21458_ (.A2(_03905_),
    .A1(_03902_),
    .B1(net225),
    .X(_03906_));
 sg13g2_nand3_1 _21459_ (.B(_03902_),
    .C(_03905_),
    .A(net225),
    .Y(_03907_));
 sg13g2_and2_1 _21460_ (.A(_03906_),
    .B(_03907_),
    .X(_03908_));
 sg13g2_inv_1 _21461_ (.Y(_03909_),
    .A(_11462_));
 sg13g2_nand2_1 _21462_ (.Y(_03910_),
    .A(net1097),
    .B(net588));
 sg13g2_and3_1 _21463_ (.X(_03911_),
    .A(_03909_),
    .B(net79),
    .C(_03910_));
 sg13g2_nor2_1 _21464_ (.A(_11634_),
    .B(_03910_),
    .Y(_03912_));
 sg13g2_nand3_1 _21465_ (.B(_03906_),
    .C(_03907_),
    .A(_03909_),
    .Y(_03913_));
 sg13g2_nand2_1 _21466_ (.Y(_03914_),
    .A(_10835_),
    .B(_11621_));
 sg13g2_nand2_1 _21467_ (.Y(_03915_),
    .A(net1097),
    .B(net521));
 sg13g2_nand4_1 _21468_ (.B(_09158_),
    .C(_03878_),
    .A(net1004),
    .Y(_03916_),
    .D(_03915_));
 sg13g2_or3_1 _21469_ (.A(_11475_),
    .B(_03878_),
    .C(_03915_),
    .X(_03917_));
 sg13g2_nand4_1 _21470_ (.B(_11308_),
    .C(net1097),
    .A(net997),
    .Y(_03918_),
    .D(net521));
 sg13g2_nand4_1 _21471_ (.B(_03916_),
    .C(_03917_),
    .A(_03914_),
    .Y(_03919_),
    .D(_03918_));
 sg13g2_a221oi_1 _21472_ (.B2(_03913_),
    .C1(_03919_),
    .B1(_03912_),
    .A1(_03908_),
    .Y(_03920_),
    .A2(_03911_));
 sg13g2_nand2_1 _21473_ (.Y(_03921_),
    .A(net964),
    .B(net494));
 sg13g2_o21ai_1 _21474_ (.B1(_03921_),
    .Y(_00950_),
    .A1(net458),
    .A2(_03920_));
 sg13g2_nor2_1 _21475_ (.A(_11253_),
    .B(net651),
    .Y(_03922_));
 sg13g2_nor2_1 _21476_ (.A(net523),
    .B(_03904_),
    .Y(_03923_));
 sg13g2_xnor2_1 _21477_ (.Y(_03924_),
    .A(net225),
    .B(_03910_));
 sg13g2_o21ai_1 _21478_ (.B1(_11268_),
    .Y(_03925_),
    .A1(net226),
    .A2(_03885_));
 sg13g2_or3_1 _21479_ (.A(_03923_),
    .B(_03924_),
    .C(_03925_),
    .X(_03926_));
 sg13g2_buf_1 _21480_ (.A(_03926_),
    .X(_03927_));
 sg13g2_nor2_1 _21481_ (.A(_03893_),
    .B(_03927_),
    .Y(_03928_));
 sg13g2_a21oi_1 _21482_ (.A1(_03892_),
    .A2(_03928_),
    .Y(_03929_),
    .B1(_11315_));
 sg13g2_xnor2_1 _21483_ (.Y(_03930_),
    .A(net145),
    .B(_03929_));
 sg13g2_nand2_1 _21484_ (.Y(_03931_),
    .A(_03909_),
    .B(_03930_));
 sg13g2_xnor2_1 _21485_ (.Y(_03932_),
    .A(_03922_),
    .B(_03931_));
 sg13g2_nand3_1 _21486_ (.B(net1097),
    .C(_03878_),
    .A(net1004),
    .Y(_03933_));
 sg13g2_xnor2_1 _21487_ (.Y(_03934_),
    .A(_11253_),
    .B(_03933_));
 sg13g2_a22oi_1 _21488_ (.Y(_03935_),
    .B1(net358),
    .B2(_10947_),
    .A2(net597),
    .A1(net1095));
 sg13g2_o21ai_1 _21489_ (.B1(_03935_),
    .Y(_03936_),
    .A1(_11817_),
    .A2(_03934_));
 sg13g2_a21o_1 _21490_ (.A2(_03932_),
    .A1(net71),
    .B1(_03936_),
    .X(_00951_));
 sg13g2_nor4_1 _21491_ (.A(_11253_),
    .B(net651),
    .C(_03893_),
    .D(_03927_),
    .Y(_03937_));
 sg13g2_nor3_1 _21492_ (.A(net182),
    .B(_03893_),
    .C(_03927_),
    .Y(_03938_));
 sg13g2_o21ai_1 _21493_ (.B1(_03892_),
    .Y(_03939_),
    .A1(_03937_),
    .A2(_03938_));
 sg13g2_o21ai_1 _21494_ (.B1(_11315_),
    .Y(_03940_),
    .A1(net145),
    .A2(_03922_));
 sg13g2_inv_1 _21495_ (.Y(_03941_),
    .A(_03940_));
 sg13g2_a21oi_1 _21496_ (.A1(net145),
    .A2(_03922_),
    .Y(_03942_),
    .B1(_03941_));
 sg13g2_and3_1 _21497_ (.X(_03943_),
    .A(net181),
    .B(_03939_),
    .C(_03942_));
 sg13g2_a21oi_1 _21498_ (.A1(_03939_),
    .A2(_03942_),
    .Y(_03944_),
    .B1(net181));
 sg13g2_o21ai_1 _21499_ (.B1(_03909_),
    .Y(_03945_),
    .A1(_03943_),
    .A2(_03944_));
 sg13g2_nor2_1 _21500_ (.A(_11241_),
    .B(net651),
    .Y(_03946_));
 sg13g2_xnor2_1 _21501_ (.Y(_03947_),
    .A(_03945_),
    .B(_03946_));
 sg13g2_nand3_1 _21502_ (.B(net1097),
    .C(_10835_),
    .A(net1004),
    .Y(_03948_));
 sg13g2_nor2_1 _21503_ (.A(_03876_),
    .B(_03948_),
    .Y(_03949_));
 sg13g2_nand3_1 _21504_ (.B(_03854_),
    .C(_03949_),
    .A(net1003),
    .Y(_03950_));
 sg13g2_xnor2_1 _21505_ (.Y(_03951_),
    .A(_11241_),
    .B(_03950_));
 sg13g2_a22oi_1 _21506_ (.Y(_03952_),
    .B1(net358),
    .B2(net998),
    .A2(net597),
    .A1(_10907_));
 sg13g2_o21ai_1 _21507_ (.B1(_03952_),
    .Y(_03953_),
    .A1(_11817_),
    .A2(_03951_));
 sg13g2_a21o_1 _21508_ (.A2(_03947_),
    .A1(net71),
    .B1(_03953_),
    .X(_00952_));
 sg13g2_a22oi_1 _21509_ (.Y(_03954_),
    .B1(_03769_),
    .B2(_11014_),
    .A2(_03763_),
    .A1(net504));
 sg13g2_nor4_2 _21510_ (.A(_11286_),
    .B(_11241_),
    .C(_03876_),
    .Y(_03955_),
    .D(_03948_));
 sg13g2_and2_1 _21511_ (.A(_03854_),
    .B(_03955_),
    .X(_03956_));
 sg13g2_xor2_1 _21512_ (.B(_03956_),
    .A(net998),
    .X(_03957_));
 sg13g2_nand2_1 _21513_ (.Y(_03958_),
    .A(_11431_),
    .B(net523));
 sg13g2_nor2_1 _21514_ (.A(_11319_),
    .B(_11417_),
    .Y(_03959_));
 sg13g2_xnor2_1 _21515_ (.Y(_03960_),
    .A(net203),
    .B(_03959_));
 sg13g2_nor2_1 _21516_ (.A(net29),
    .B(_03960_),
    .Y(_03961_));
 sg13g2_xnor2_1 _21517_ (.Y(_03962_),
    .A(_03958_),
    .B(_03961_));
 sg13g2_a22oi_1 _21518_ (.Y(_03963_),
    .B1(_03962_),
    .B2(net71),
    .A2(_03957_),
    .A1(_03799_));
 sg13g2_nand2_1 _21519_ (.Y(_00953_),
    .A(_03954_),
    .B(_03963_));
 sg13g2_nand2_1 _21520_ (.Y(_03964_),
    .A(_11014_),
    .B(net523));
 sg13g2_nand2_1 _21521_ (.Y(_03965_),
    .A(net203),
    .B(_03959_));
 sg13g2_o21ai_1 _21522_ (.B1(net178),
    .Y(_03966_),
    .A1(_11319_),
    .A2(_11417_));
 sg13g2_nand2b_1 _21523_ (.Y(_03967_),
    .B(_03966_),
    .A_N(_03958_));
 sg13g2_a21o_1 _21524_ (.A2(_03967_),
    .A1(_03965_),
    .B1(net143),
    .X(_03968_));
 sg13g2_nand3_1 _21525_ (.B(_03965_),
    .C(_03967_),
    .A(net143),
    .Y(_03969_));
 sg13g2_a21oi_1 _21526_ (.A1(_03968_),
    .A2(_03969_),
    .Y(_03970_),
    .B1(net29));
 sg13g2_xnor2_1 _21527_ (.Y(_03971_),
    .A(_03964_),
    .B(_03970_));
 sg13g2_nand3_1 _21528_ (.B(_03854_),
    .C(_03955_),
    .A(net998),
    .Y(_03972_));
 sg13g2_xnor2_1 _21529_ (.Y(_03973_),
    .A(_11420_),
    .B(_03972_));
 sg13g2_a22oi_1 _21530_ (.Y(_03974_),
    .B1(net358),
    .B2(_11112_),
    .A2(net597),
    .A1(net601));
 sg13g2_o21ai_1 _21531_ (.B1(_03974_),
    .Y(_03975_),
    .A1(_11817_),
    .A2(_03973_));
 sg13g2_a21o_1 _21532_ (.A2(_03971_),
    .A1(net71),
    .B1(_03975_),
    .X(_00954_));
 sg13g2_nand2_1 _21533_ (.Y(_03976_),
    .A(net732),
    .B(net597));
 sg13g2_o21ai_1 _21534_ (.B1(net522),
    .Y(_03977_),
    .A1(_11047_),
    .A2(_11556_));
 sg13g2_and2_1 _21535_ (.A(_11556_),
    .B(_03976_),
    .X(_03978_));
 sg13g2_and2_1 _21536_ (.A(net998),
    .B(_11014_),
    .X(_03979_));
 sg13g2_nand3_1 _21537_ (.B(_03955_),
    .C(_03979_),
    .A(_03854_),
    .Y(_03980_));
 sg13g2_xnor2_1 _21538_ (.Y(_03981_),
    .A(_11112_),
    .B(_03980_));
 sg13g2_o21ai_1 _21539_ (.B1(net178),
    .Y(_03982_),
    .A1(_11420_),
    .A2(_11846_));
 sg13g2_or2_1 _21540_ (.X(_03983_),
    .B(_11454_),
    .A(net998));
 sg13g2_a22oi_1 _21541_ (.Y(_03984_),
    .B1(_03982_),
    .B2(_03983_),
    .A2(_11447_),
    .A1(_11446_));
 sg13g2_or2_1 _21542_ (.X(_03985_),
    .B(net203),
    .A(net998));
 sg13g2_o21ai_1 _21543_ (.B1(_11452_),
    .Y(_03986_),
    .A1(_11454_),
    .A2(_03985_));
 sg13g2_o21ai_1 _21544_ (.B1(net147),
    .Y(_03987_),
    .A1(_03984_),
    .A2(_03986_));
 sg13g2_or3_1 _21545_ (.A(net147),
    .B(_03984_),
    .C(_03986_),
    .X(_03988_));
 sg13g2_a21oi_1 _21546_ (.A1(_03987_),
    .A2(_03988_),
    .Y(_03989_),
    .B1(_03722_));
 sg13g2_xnor2_1 _21547_ (.Y(_03990_),
    .A(_11439_),
    .B(_03989_));
 sg13g2_a22oi_1 _21548_ (.Y(_03991_),
    .B1(_03990_),
    .B2(net79),
    .A2(_03981_),
    .A1(_11815_));
 sg13g2_a22oi_1 _21549_ (.Y(_00955_),
    .B1(_03978_),
    .B2(_03991_),
    .A2(_03977_),
    .A1(_03976_));
 sg13g2_nand4_1 _21550_ (.B(_03854_),
    .C(_03955_),
    .A(_11112_),
    .Y(_03992_),
    .D(_03979_));
 sg13g2_xnor2_1 _21551_ (.Y(_03993_),
    .A(_11047_),
    .B(_03992_));
 sg13g2_nand2_1 _21552_ (.Y(_03994_),
    .A(_03959_),
    .B(_11441_));
 sg13g2_nand2_1 _21553_ (.Y(_03995_),
    .A(_11459_),
    .B(_03994_));
 sg13g2_xnor2_1 _21554_ (.Y(_03996_),
    .A(net199),
    .B(_03995_));
 sg13g2_nor2_1 _21555_ (.A(_11449_),
    .B(_11634_),
    .Y(_03997_));
 sg13g2_a221oi_1 _21556_ (.B2(_03997_),
    .C1(_11621_),
    .B1(_03996_),
    .A1(_11815_),
    .Y(_03998_),
    .A2(_03993_));
 sg13g2_o21ai_1 _21557_ (.B1(net522),
    .Y(_03999_),
    .A1(\cpu.ex.r_mult[31] ),
    .A2(_11556_));
 sg13g2_nand2_1 _21558_ (.Y(_04000_),
    .A(net638),
    .B(net494));
 sg13g2_o21ai_1 _21559_ (.B1(_04000_),
    .Y(_00956_),
    .A1(_03998_),
    .A2(_03999_));
 sg13g2_a221oi_1 _21560_ (.B2(_11536_),
    .C1(_11500_),
    .B1(_11535_),
    .A1(_11532_),
    .Y(_04001_),
    .A2(_11534_));
 sg13g2_buf_2 _21561_ (.A(_04001_),
    .X(_04002_));
 sg13g2_nand2_1 _21562_ (.Y(_04003_),
    .A(_10260_),
    .B(_10261_));
 sg13g2_nor2_1 _21563_ (.A(_11496_),
    .B(_04003_),
    .Y(_04004_));
 sg13g2_buf_1 _21564_ (.A(_04004_),
    .X(_04005_));
 sg13g2_nor2b_1 _21565_ (.A(_11503_),
    .B_N(net1119),
    .Y(_04006_));
 sg13g2_mux2_1 _21566_ (.A0(_04006_),
    .A1(_09018_),
    .S(_11898_),
    .X(_04007_));
 sg13g2_nand3_1 _21567_ (.B(net214),
    .C(_04007_),
    .A(net729),
    .Y(_04008_));
 sg13g2_buf_2 _21568_ (.A(_04008_),
    .X(_04009_));
 sg13g2_and2_1 _21569_ (.A(net1042),
    .B(_11234_),
    .X(_04010_));
 sg13g2_buf_1 _21570_ (.A(_04010_),
    .X(_04011_));
 sg13g2_nand2_2 _21571_ (.Y(_04012_),
    .A(net374),
    .B(net370));
 sg13g2_nand2_1 _21572_ (.Y(_04013_),
    .A(net301),
    .B(net296));
 sg13g2_buf_2 _21573_ (.A(_04013_),
    .X(_04014_));
 sg13g2_o21ai_1 _21574_ (.B1(_11482_),
    .Y(_04015_),
    .A1(_04012_),
    .A2(_04014_));
 sg13g2_buf_1 _21575_ (.A(_10939_),
    .X(_04016_));
 sg13g2_nor2_1 _21576_ (.A(net300),
    .B(net296),
    .Y(_04017_));
 sg13g2_nor2_1 _21577_ (.A(net300),
    .B(net299),
    .Y(_04018_));
 sg13g2_buf_2 _21578_ (.A(_04018_),
    .X(_04019_));
 sg13g2_a22oi_1 _21579_ (.Y(_04020_),
    .B1(_04019_),
    .B2(net146),
    .A2(_04017_),
    .A1(_04016_));
 sg13g2_a21o_1 _21580_ (.A2(_11124_),
    .A1(net227),
    .B1(_11126_),
    .X(_04021_));
 sg13g2_buf_1 _21581_ (.A(_04021_),
    .X(_04022_));
 sg13g2_buf_1 _21582_ (.A(_04022_),
    .X(_04023_));
 sg13g2_nand3_1 _21583_ (.B(net114),
    .C(_04019_),
    .A(net237),
    .Y(_04024_));
 sg13g2_o21ai_1 _21584_ (.B1(_04024_),
    .Y(_04025_),
    .A1(net237),
    .A2(_04020_));
 sg13g2_nand2_1 _21585_ (.Y(_04026_),
    .A(net293),
    .B(_04025_));
 sg13g2_nand2_1 _21586_ (.Y(_04027_),
    .A(_10431_),
    .B(net371));
 sg13g2_buf_2 _21587_ (.A(_04027_),
    .X(_04028_));
 sg13g2_nor2_1 _21588_ (.A(_04012_),
    .B(_04028_),
    .Y(_04029_));
 sg13g2_buf_1 _21589_ (.A(_04029_),
    .X(_04030_));
 sg13g2_buf_1 _21590_ (.A(_04030_),
    .X(_04031_));
 sg13g2_nand2_1 _21591_ (.Y(_04032_),
    .A(net374),
    .B(net292));
 sg13g2_buf_2 _21592_ (.A(_04032_),
    .X(_04033_));
 sg13g2_nand2_1 _21593_ (.Y(_04034_),
    .A(_11399_),
    .B(net299));
 sg13g2_buf_1 _21594_ (.A(_04034_),
    .X(_04035_));
 sg13g2_nor2_1 _21595_ (.A(_04033_),
    .B(_04035_),
    .Y(_04036_));
 sg13g2_buf_1 _21596_ (.A(_04036_),
    .X(_04037_));
 sg13g2_nand2_2 _21597_ (.Y(_04038_),
    .A(_10348_),
    .B(net292));
 sg13g2_nor2_1 _21598_ (.A(_04038_),
    .B(_04035_),
    .Y(_04039_));
 sg13g2_buf_1 _21599_ (.A(_04039_),
    .X(_04040_));
 sg13g2_and2_1 _21600_ (.A(_11351_),
    .B(net171),
    .X(_04041_));
 sg13g2_a221oi_1 _21601_ (.B2(net204),
    .C1(_04041_),
    .B1(net172),
    .A1(_10678_),
    .Y(_04042_),
    .A2(net173));
 sg13g2_inv_1 _21602_ (.Y(_04043_),
    .A(_00175_));
 sg13g2_mux2_1 _21603_ (.A0(_04043_),
    .A1(_11893_),
    .S(net250),
    .X(_04044_));
 sg13g2_buf_1 _21604_ (.A(_04044_),
    .X(_04045_));
 sg13g2_buf_1 _21605_ (.A(_04045_),
    .X(_04046_));
 sg13g2_nand2_1 _21606_ (.Y(_04047_),
    .A(_10348_),
    .B(net370));
 sg13g2_buf_2 _21607_ (.A(_04047_),
    .X(_04048_));
 sg13g2_nor3_1 _21608_ (.A(_11399_),
    .B(net371),
    .C(_04048_),
    .Y(_04049_));
 sg13g2_buf_1 _21609_ (.A(_04049_),
    .X(_04050_));
 sg13g2_buf_1 _21610_ (.A(net192),
    .X(_04051_));
 sg13g2_nor2_1 _21611_ (.A(_04033_),
    .B(_04028_),
    .Y(_04052_));
 sg13g2_buf_2 _21612_ (.A(_04052_),
    .X(_04053_));
 sg13g2_buf_1 _21613_ (.A(_04053_),
    .X(_04054_));
 sg13g2_buf_1 _21614_ (.A(net206),
    .X(_04055_));
 sg13g2_a22oi_1 _21615_ (.Y(_04056_),
    .B1(net136),
    .B2(net168),
    .A2(net169),
    .A1(net170));
 sg13g2_buf_1 _21616_ (.A(net207),
    .X(_04057_));
 sg13g2_nor2_1 _21617_ (.A(_04028_),
    .B(_04048_),
    .Y(_04058_));
 sg13g2_buf_1 _21618_ (.A(_04058_),
    .X(_04059_));
 sg13g2_buf_1 _21619_ (.A(_04059_),
    .X(_04060_));
 sg13g2_nand2_1 _21620_ (.Y(_04061_),
    .A(net167),
    .B(net166));
 sg13g2_buf_1 _21621_ (.A(_10505_),
    .X(_04062_));
 sg13g2_nor2_1 _21622_ (.A(_04038_),
    .B(_04028_),
    .Y(_04063_));
 sg13g2_buf_1 _21623_ (.A(_04063_),
    .X(_04064_));
 sg13g2_buf_1 _21624_ (.A(_04064_),
    .X(_04065_));
 sg13g2_nand2_1 _21625_ (.Y(_04066_),
    .A(net191),
    .B(net165));
 sg13g2_and2_1 _21626_ (.A(_04061_),
    .B(_04066_),
    .X(_04067_));
 sg13g2_buf_1 _21627_ (.A(_11157_),
    .X(_04068_));
 sg13g2_nor2_1 _21628_ (.A(_04012_),
    .B(_04035_),
    .Y(_04069_));
 sg13g2_buf_1 _21629_ (.A(_04069_),
    .X(_04070_));
 sg13g2_nor2_1 _21630_ (.A(_04033_),
    .B(_04014_),
    .Y(_04071_));
 sg13g2_buf_1 _21631_ (.A(_11098_),
    .X(_04072_));
 sg13g2_and2_1 _21632_ (.A(_10579_),
    .B(_10609_),
    .X(_04073_));
 sg13g2_buf_1 _21633_ (.A(_04073_),
    .X(_04074_));
 sg13g2_nand2_1 _21634_ (.Y(_04075_),
    .A(_11480_),
    .B(_10350_));
 sg13g2_nor2_1 _21635_ (.A(_10348_),
    .B(net370),
    .Y(_04076_));
 sg13g2_nand2_1 _21636_ (.Y(_04077_),
    .A(_11480_),
    .B(_04076_));
 sg13g2_buf_1 _21637_ (.A(_04077_),
    .X(_04078_));
 sg13g2_o21ai_1 _21638_ (.B1(net164),
    .Y(_04079_),
    .A1(net213),
    .A2(_04075_));
 sg13g2_a221oi_1 _21639_ (.B2(net135),
    .C1(_04079_),
    .B1(_04071_),
    .A1(net113),
    .Y(_04080_),
    .A2(_04070_));
 sg13g2_and4_1 _21640_ (.A(_04042_),
    .B(_04056_),
    .C(_04067_),
    .D(_04080_),
    .X(_04081_));
 sg13g2_nor2_1 _21641_ (.A(_08910_),
    .B(_09712_),
    .Y(_04082_));
 sg13g2_buf_1 _21642_ (.A(_04082_),
    .X(_04083_));
 sg13g2_a21oi_1 _21643_ (.A1(_04026_),
    .A2(_04081_),
    .Y(_04084_),
    .B1(net834));
 sg13g2_a21o_1 _21644_ (.A2(_04015_),
    .A1(_04011_),
    .B1(_04084_),
    .X(_04085_));
 sg13g2_and2_1 _21645_ (.A(_11480_),
    .B(_04076_),
    .X(_04086_));
 sg13g2_buf_1 _21646_ (.A(_04086_),
    .X(_04087_));
 sg13g2_buf_1 _21647_ (.A(_04087_),
    .X(_04088_));
 sg13g2_buf_1 _21648_ (.A(net134),
    .X(_04089_));
 sg13g2_buf_1 _21649_ (.A(net112),
    .X(_04090_));
 sg13g2_nand2_1 _21650_ (.Y(_04091_),
    .A(_11389_),
    .B(_04090_));
 sg13g2_inv_1 _21651_ (.Y(_04092_),
    .A(net200));
 sg13g2_buf_1 _21652_ (.A(_04092_),
    .X(_04093_));
 sg13g2_nand3_1 _21653_ (.B(net133),
    .C(_04090_),
    .A(_09732_),
    .Y(_04094_));
 sg13g2_nor2_1 _21654_ (.A(net897),
    .B(_09151_),
    .Y(_04095_));
 sg13g2_nor2_1 _21655_ (.A(_11554_),
    .B(_04095_),
    .Y(_04096_));
 sg13g2_buf_1 _21656_ (.A(_04096_),
    .X(_04097_));
 sg13g2_buf_1 _21657_ (.A(_04097_),
    .X(_04098_));
 sg13g2_a21oi_1 _21658_ (.A1(_08882_),
    .A2(_11256_),
    .Y(_04099_),
    .B1(net291));
 sg13g2_a21o_1 _21659_ (.A2(_10258_),
    .A1(_10826_),
    .B1(_10352_),
    .X(_04100_));
 sg13g2_buf_1 _21660_ (.A(_04100_),
    .X(_04101_));
 sg13g2_buf_1 _21661_ (.A(_04101_),
    .X(_04102_));
 sg13g2_nand2_1 _21662_ (.Y(_04103_),
    .A(net132),
    .B(_11369_));
 sg13g2_nand2_1 _21663_ (.Y(_04104_),
    .A(_11383_),
    .B(net292));
 sg13g2_nand2_1 _21664_ (.Y(_04105_),
    .A(_04103_),
    .B(_04104_));
 sg13g2_nor2_1 _21665_ (.A(\cpu.dec.r_op[7] ),
    .B(_09708_),
    .Y(_04106_));
 sg13g2_nor2_1 _21666_ (.A(net1123),
    .B(_08932_),
    .Y(_04107_));
 sg13g2_nor4_1 _21667_ (.A(_08881_),
    .B(net1113),
    .C(_09718_),
    .D(_09731_),
    .Y(_04108_));
 sg13g2_nand4_1 _21668_ (.B(_04082_),
    .C(_04107_),
    .A(_04106_),
    .Y(_04109_),
    .D(_04108_));
 sg13g2_buf_2 _21669_ (.A(_04109_),
    .X(_04110_));
 sg13g2_and2_1 _21670_ (.A(_04106_),
    .B(_04110_),
    .X(_04111_));
 sg13g2_buf_1 _21671_ (.A(_04111_),
    .X(_04112_));
 sg13g2_a21oi_1 _21672_ (.A1(net200),
    .A2(_04105_),
    .Y(_04113_),
    .B1(_04112_));
 sg13g2_nand2_1 _21673_ (.Y(_04114_),
    .A(_04106_),
    .B(_04110_));
 sg13g2_buf_1 _21674_ (.A(_04114_),
    .X(_04115_));
 sg13g2_o21ai_1 _21675_ (.B1(net245),
    .Y(_04116_),
    .A1(net200),
    .A2(_04115_));
 sg13g2_nand2_1 _21676_ (.Y(_04117_),
    .A(net200),
    .B(_04115_));
 sg13g2_o21ai_1 _21677_ (.B1(_04117_),
    .Y(_04118_),
    .A1(_11533_),
    .A2(_11385_));
 sg13g2_nor3_1 _21678_ (.A(_03721_),
    .B(_04105_),
    .C(_04118_),
    .Y(_04119_));
 sg13g2_a21oi_1 _21679_ (.A1(_04105_),
    .A2(_04116_),
    .Y(_04120_),
    .B1(_04119_));
 sg13g2_o21ai_1 _21680_ (.B1(_04120_),
    .Y(_04121_),
    .A1(net1123),
    .A2(_04113_));
 sg13g2_mux2_1 _21681_ (.A0(_08959_),
    .A1(_08933_),
    .S(_04103_),
    .X(_04122_));
 sg13g2_o21ai_1 _21682_ (.B1(_04104_),
    .Y(_04123_),
    .A1(_09719_),
    .A2(_04122_));
 sg13g2_nand4_1 _21683_ (.B(_04099_),
    .C(_04121_),
    .A(_04094_),
    .Y(_04124_),
    .D(_04123_));
 sg13g2_a21oi_1 _21684_ (.A1(_04085_),
    .A2(_04091_),
    .Y(_04125_),
    .B1(_04124_));
 sg13g2_or2_1 _21685_ (.X(_04126_),
    .B(_04125_),
    .A(_04009_));
 sg13g2_a21oi_1 _21686_ (.A1(_11562_),
    .A2(_04002_),
    .Y(_04127_),
    .B1(_04126_));
 sg13g2_nand2_1 _21687_ (.Y(_04128_),
    .A(_08186_),
    .B(net729));
 sg13g2_nor4_1 _21688_ (.A(_11508_),
    .B(net373),
    .C(_04128_),
    .D(_11898_),
    .Y(_04129_));
 sg13g2_buf_1 _21689_ (.A(_04129_),
    .X(_04130_));
 sg13g2_nand2_1 _21690_ (.Y(_04131_),
    .A(\cpu.dec.iready ),
    .B(_00183_));
 sg13g2_nor2_2 _21691_ (.A(\cpu.ex.r_branch_stall ),
    .B(_04131_),
    .Y(_04132_));
 sg13g2_nor2_1 _21692_ (.A(net387),
    .B(_04132_),
    .Y(_04133_));
 sg13g2_nor3_1 _21693_ (.A(_10260_),
    .B(_11496_),
    .C(net1031),
    .Y(_04134_));
 sg13g2_o21ai_1 _21694_ (.B1(_09018_),
    .Y(_04135_),
    .A1(_04133_),
    .A2(_04134_));
 sg13g2_nor3_1 _21695_ (.A(_09013_),
    .B(_10261_),
    .C(_04128_),
    .Y(_04136_));
 sg13g2_a21oi_1 _21696_ (.A1(net387),
    .A2(_04136_),
    .Y(_04137_),
    .B1(net897));
 sg13g2_nand3b_1 _21697_ (.B(_04135_),
    .C(_04137_),
    .Y(_04138_),
    .A_N(net95));
 sg13g2_nor2b_1 _21698_ (.A(_04138_),
    .B_N(_04009_),
    .Y(_04139_));
 sg13g2_buf_1 _21699_ (.A(_04139_),
    .X(_04140_));
 sg13g2_buf_1 _21700_ (.A(_04140_),
    .X(_04141_));
 sg13g2_a22oi_1 _21701_ (.Y(_04142_),
    .B1(_04141_),
    .B2(net688),
    .A2(net95),
    .A1(_10326_));
 sg13g2_nand2b_1 _21702_ (.Y(_00957_),
    .B(_04142_),
    .A_N(_04127_));
 sg13g2_buf_1 _21703_ (.A(_04009_),
    .X(_04143_));
 sg13g2_nand2_1 _21704_ (.Y(_04144_),
    .A(net183),
    .B(_11034_));
 sg13g2_nand2_1 _21705_ (.Y(_04145_),
    .A(net181),
    .B(_10939_));
 sg13g2_nand2_1 _21706_ (.Y(_04146_),
    .A(_04144_),
    .B(_04145_));
 sg13g2_o21ai_1 _21707_ (.B1(_11036_),
    .Y(_04147_),
    .A1(_10807_),
    .A2(_10881_));
 sg13g2_buf_1 _21708_ (.A(_04147_),
    .X(_04148_));
 sg13g2_nor2_1 _21709_ (.A(_10339_),
    .B(_11889_),
    .Y(_04149_));
 sg13g2_a21oi_1 _21710_ (.A1(_10941_),
    .A2(_10339_),
    .Y(_04150_),
    .B1(_04149_));
 sg13g2_buf_2 _21711_ (.A(_04150_),
    .X(_04151_));
 sg13g2_o21ai_1 _21712_ (.B1(_04151_),
    .Y(_04152_),
    .A1(net145),
    .A2(_04148_));
 sg13g2_nand2_1 _21713_ (.Y(_04153_),
    .A(net145),
    .B(_04148_));
 sg13g2_nand2_1 _21714_ (.Y(_04154_),
    .A(_04152_),
    .B(_04153_));
 sg13g2_xor2_1 _21715_ (.B(_04154_),
    .A(_04146_),
    .X(_04155_));
 sg13g2_nand2_1 _21716_ (.Y(_04156_),
    .A(_11277_),
    .B(_10738_));
 sg13g2_xnor2_1 _21717_ (.Y(_04157_),
    .A(net207),
    .B(net249));
 sg13g2_buf_2 _21718_ (.A(_04157_),
    .X(_04158_));
 sg13g2_nand3_1 _21719_ (.B(_04156_),
    .C(_04158_),
    .A(_10671_),
    .Y(_04159_));
 sg13g2_nor2_1 _21720_ (.A(_11389_),
    .B(net371),
    .Y(_04160_));
 sg13g2_nand2b_1 _21721_ (.Y(_04161_),
    .B(_10258_),
    .A_N(_10334_));
 sg13g2_or2_1 _21722_ (.X(_04162_),
    .B(_10334_),
    .A(_10326_));
 sg13g2_mux2_1 _21723_ (.A0(_04161_),
    .A1(_04162_),
    .S(_10338_),
    .X(_04163_));
 sg13g2_a221oi_1 _21724_ (.B2(net250),
    .C1(_10348_),
    .B1(_10291_),
    .A1(_10259_),
    .Y(_04164_),
    .A2(_10264_));
 sg13g2_a221oi_1 _21725_ (.B2(net250),
    .C1(_10349_),
    .B1(_10258_),
    .A1(_11380_),
    .Y(_04165_),
    .A2(_11381_));
 sg13g2_a221oi_1 _21726_ (.B2(_04164_),
    .C1(_04165_),
    .B1(_04163_),
    .A1(_11389_),
    .Y(_04166_),
    .A2(_10463_));
 sg13g2_a21oi_1 _21727_ (.A1(_10472_),
    .A2(_10503_),
    .Y(_04167_),
    .B1(net230));
 sg13g2_a21oi_2 _21728_ (.B1(_10576_),
    .Y(_04168_),
    .A2(_10609_),
    .A1(_10579_));
 sg13g2_a21o_1 _21729_ (.A2(_10431_),
    .A1(_04045_),
    .B1(_04168_),
    .X(_04169_));
 sg13g2_nor4_2 _21730_ (.A(_04160_),
    .B(_04166_),
    .C(_04167_),
    .Y(_04170_),
    .D(_04169_));
 sg13g2_and3_1 _21731_ (.X(_04171_),
    .A(_10472_),
    .B(_10503_),
    .C(net230));
 sg13g2_a221oi_1 _21732_ (.B2(_10576_),
    .C1(_04171_),
    .B1(net213),
    .A1(_10390_),
    .Y(_04172_),
    .A2(_11398_));
 sg13g2_nand3_1 _21733_ (.B(_10503_),
    .C(_10540_),
    .A(_10472_),
    .Y(_04173_));
 sg13g2_a21oi_1 _21734_ (.A1(_04168_),
    .A2(_04173_),
    .Y(_04174_),
    .B1(_04167_));
 sg13g2_nor2b_1 _21735_ (.A(_04172_),
    .B_N(_04174_),
    .Y(_04175_));
 sg13g2_buf_1 _21736_ (.A(_04175_),
    .X(_04176_));
 sg13g2_or3_1 _21737_ (.A(_04159_),
    .B(_04170_),
    .C(_04176_),
    .X(_04177_));
 sg13g2_buf_1 _21738_ (.A(_04177_),
    .X(_04178_));
 sg13g2_a21oi_1 _21739_ (.A1(net224),
    .A2(net206),
    .Y(_04179_),
    .B1(net228));
 sg13g2_a21oi_1 _21740_ (.A1(_11290_),
    .A2(net206),
    .Y(_04180_),
    .B1(net207));
 sg13g2_o21ai_1 _21741_ (.B1(_10679_),
    .Y(_04181_),
    .A1(_04179_),
    .A2(_04180_));
 sg13g2_nand2_1 _21742_ (.Y(_04182_),
    .A(_10671_),
    .B(_04181_));
 sg13g2_a21oi_1 _21743_ (.A1(_04178_),
    .A2(_04182_),
    .Y(_04183_),
    .B1(_11256_));
 sg13g2_a21oi_1 _21744_ (.A1(_10671_),
    .A2(_04181_),
    .Y(_04184_),
    .B1(_10878_));
 sg13g2_a21oi_1 _21745_ (.A1(_04178_),
    .A2(_04184_),
    .Y(_04185_),
    .B1(_10856_));
 sg13g2_nand2_1 _21746_ (.Y(_04186_),
    .A(_04151_),
    .B(_10996_));
 sg13g2_o21ai_1 _21747_ (.B1(_04186_),
    .Y(_04187_),
    .A1(_04183_),
    .A2(_04185_));
 sg13g2_nand2_1 _21748_ (.Y(_04188_),
    .A(net204),
    .B(_11255_));
 sg13g2_nand2_1 _21749_ (.Y(_04189_),
    .A(_04187_),
    .B(_04188_));
 sg13g2_xnor2_1 _21750_ (.Y(_04190_),
    .A(_04146_),
    .B(_04189_));
 sg13g2_buf_1 _21751_ (.A(_10738_),
    .X(_04191_));
 sg13g2_nand3_1 _21752_ (.B(_11284_),
    .C(net163),
    .A(_09708_),
    .Y(_04192_));
 sg13g2_nand4_1 _21753_ (.B(net201),
    .C(net206),
    .A(_09708_),
    .Y(_04193_),
    .D(_04158_));
 sg13g2_o21ai_1 _21754_ (.B1(_04193_),
    .Y(_04194_),
    .A1(_04158_),
    .A2(_04192_));
 sg13g2_buf_1 _21755_ (.A(_04194_),
    .X(_04195_));
 sg13g2_nand2_1 _21756_ (.Y(_04196_),
    .A(net207),
    .B(net223));
 sg13g2_and2_1 _21757_ (.A(_10801_),
    .B(_04196_),
    .X(_04197_));
 sg13g2_nand3_1 _21758_ (.B(net163),
    .C(_04197_),
    .A(_09708_),
    .Y(_04198_));
 sg13g2_nand3_1 _21759_ (.B(net198),
    .C(_04197_),
    .A(_09708_),
    .Y(_04199_));
 sg13g2_inv_1 _21760_ (.Y(_04200_),
    .A(_10805_));
 sg13g2_a21oi_2 _21761_ (.B1(_04200_),
    .Y(_04201_),
    .A2(_10613_),
    .A1(_10468_));
 sg13g2_a21oi_1 _21762_ (.A1(_04198_),
    .A2(_04199_),
    .Y(_04202_),
    .B1(_04201_));
 sg13g2_nand3_1 _21763_ (.B(net206),
    .C(_04158_),
    .A(_09708_),
    .Y(_04203_));
 sg13g2_nand3_1 _21764_ (.B(net201),
    .C(_04158_),
    .A(_09708_),
    .Y(_04204_));
 sg13g2_a21o_1 _21765_ (.A2(_10613_),
    .A1(_10468_),
    .B1(_04200_),
    .X(_04205_));
 sg13g2_a21oi_1 _21766_ (.A1(_04203_),
    .A2(_04204_),
    .Y(_04206_),
    .B1(_04205_));
 sg13g2_nor4_1 _21767_ (.A(_04097_),
    .B(_04195_),
    .C(_04202_),
    .D(_04206_),
    .Y(_04207_));
 sg13g2_buf_1 _21768_ (.A(_04207_),
    .X(_04208_));
 sg13g2_mux2_1 _21769_ (.A0(net1041),
    .A1(net1040),
    .S(_11035_),
    .X(_04209_));
 sg13g2_nand2_1 _21770_ (.Y(_04210_),
    .A(_11033_),
    .B(_11034_));
 sg13g2_o21ai_1 _21771_ (.B1(_04210_),
    .Y(_04211_),
    .A1(net1027),
    .A2(_04209_));
 sg13g2_nand2_1 _21772_ (.Y(_04212_),
    .A(net297),
    .B(_11480_));
 sg13g2_and2_1 _21773_ (.A(_09712_),
    .B(net146),
    .X(_04213_));
 sg13g2_nor2_1 _21774_ (.A(net119),
    .B(_04075_),
    .Y(_04214_));
 sg13g2_a221oi_1 _21775_ (.B2(net165),
    .C1(_04214_),
    .B1(_04213_),
    .A1(_04011_),
    .Y(_04215_),
    .A2(_04212_));
 sg13g2_buf_1 _21776_ (.A(_11480_),
    .X(_04216_));
 sg13g2_buf_1 _21777_ (.A(_11127_),
    .X(_04217_));
 sg13g2_o21ai_1 _21778_ (.B1(_04033_),
    .Y(_04218_),
    .A1(_04217_),
    .A2(_04048_));
 sg13g2_nand2_1 _21779_ (.Y(_04219_),
    .A(net190),
    .B(_04218_));
 sg13g2_a221oi_1 _21780_ (.B2(_04219_),
    .C1(net834),
    .B1(_04215_),
    .A1(_11028_),
    .Y(_04220_),
    .A2(net112));
 sg13g2_a21oi_1 _21781_ (.A1(net1043),
    .A2(net242),
    .Y(_04221_),
    .B1(_04220_));
 sg13g2_nor2_1 _21782_ (.A(net242),
    .B(_11405_),
    .Y(_04222_));
 sg13g2_nand2_1 _21783_ (.Y(_04223_),
    .A(_11481_),
    .B(_04222_));
 sg13g2_nor2_1 _21784_ (.A(_10770_),
    .B(_04223_),
    .Y(_04224_));
 sg13g2_and2_1 _21785_ (.A(_11351_),
    .B(_04050_),
    .X(_04225_));
 sg13g2_nor2_1 _21786_ (.A(_04224_),
    .B(_04225_),
    .Y(_04226_));
 sg13g2_a22oi_1 _21787_ (.Y(_04227_),
    .B1(_04054_),
    .B2(net168),
    .A2(net173),
    .A1(net229));
 sg13g2_a221oi_1 _21788_ (.B2(net133),
    .C1(net112),
    .B1(_04070_),
    .A1(_04062_),
    .Y(_04228_),
    .A2(net166));
 sg13g2_buf_1 _21789_ (.A(_10128_),
    .X(_04229_));
 sg13g2_a22oi_1 _21790_ (.Y(_04230_),
    .B1(_04037_),
    .B2(net162),
    .A2(net171),
    .A1(net170));
 sg13g2_nor3_2 _21791_ (.A(net242),
    .B(net296),
    .C(_04012_),
    .Y(_04231_));
 sg13g2_buf_1 _21792_ (.A(_04231_),
    .X(_04232_));
 sg13g2_nor2_1 _21793_ (.A(_04035_),
    .B(_04048_),
    .Y(_04233_));
 sg13g2_buf_1 _21794_ (.A(_04233_),
    .X(_04234_));
 sg13g2_a22oi_1 _21795_ (.Y(_04235_),
    .B1(net161),
    .B2(_04102_),
    .A2(net189),
    .A1(_10678_));
 sg13g2_and2_1 _21796_ (.A(_04230_),
    .B(_04235_),
    .X(_04236_));
 sg13g2_nand4_1 _21797_ (.B(_04227_),
    .C(_04228_),
    .A(_04226_),
    .Y(_04237_),
    .D(_04236_));
 sg13g2_nand2_1 _21798_ (.Y(_04238_),
    .A(_04151_),
    .B(net96));
 sg13g2_nand3_1 _21799_ (.B(_04237_),
    .C(_04238_),
    .A(net1026),
    .Y(_04239_));
 sg13g2_nand4_1 _21800_ (.B(_04211_),
    .C(_04221_),
    .A(_04208_),
    .Y(_04240_),
    .D(_04239_));
 sg13g2_a21oi_1 _21801_ (.A1(net1063),
    .A2(_04190_),
    .Y(_04241_),
    .B1(_04240_));
 sg13g2_o21ai_1 _21802_ (.B1(_04241_),
    .Y(_04242_),
    .A1(_04110_),
    .A2(_04155_));
 sg13g2_o21ai_1 _21803_ (.B1(_04242_),
    .Y(_04243_),
    .A1(_11500_),
    .A2(\cpu.ex.c_mult[11] ));
 sg13g2_buf_1 _21804_ (.A(_08629_),
    .X(_04244_));
 sg13g2_inv_1 _21805_ (.Y(_04245_),
    .A(_08656_));
 sg13g2_and2_1 _21806_ (.A(_08705_),
    .B(net788),
    .X(_04246_));
 sg13g2_buf_1 _21807_ (.A(_04246_),
    .X(_04247_));
 sg13g2_nand3_1 _21808_ (.B(_08673_),
    .C(_04247_),
    .A(net1046),
    .Y(_04248_));
 sg13g2_nor2_1 _21809_ (.A(_08648_),
    .B(_04248_),
    .Y(_04249_));
 sg13g2_nand3_1 _21810_ (.B(_08620_),
    .C(_04249_),
    .A(_08611_),
    .Y(_04250_));
 sg13g2_nor2_1 _21811_ (.A(net958),
    .B(_04250_),
    .Y(_04251_));
 sg13g2_nand2_1 _21812_ (.Y(_04252_),
    .A(_08639_),
    .B(_04251_));
 sg13g2_xnor2_1 _21813_ (.Y(_04253_),
    .A(_10882_),
    .B(_04252_));
 sg13g2_buf_1 _21814_ (.A(net95),
    .X(_04254_));
 sg13g2_a22oi_1 _21815_ (.Y(_04255_),
    .B1(_04253_),
    .B2(net83),
    .A2(net32),
    .A1(net959));
 sg13g2_o21ai_1 _21816_ (.B1(_04255_),
    .Y(_00958_),
    .A1(_04143_),
    .A2(_04243_));
 sg13g2_xnor2_1 _21817_ (.Y(_04256_),
    .A(net178),
    .B(net113));
 sg13g2_and3_1 _21818_ (.X(_04257_),
    .A(_10878_),
    .B(_10671_),
    .C(_04181_));
 sg13g2_nand4_1 _21819_ (.B(_10671_),
    .C(_04156_),
    .A(_10878_),
    .Y(_04258_),
    .D(_04158_));
 sg13g2_nor3_1 _21820_ (.A(_04170_),
    .B(_04176_),
    .C(_04258_),
    .Y(_04259_));
 sg13g2_nand2_1 _21821_ (.Y(_04260_),
    .A(_04145_),
    .B(_04188_));
 sg13g2_or3_1 _21822_ (.A(_04257_),
    .B(_04259_),
    .C(_04260_),
    .X(_04261_));
 sg13g2_nor2_1 _21823_ (.A(net204),
    .B(_11263_),
    .Y(_04262_));
 sg13g2_inv_1 _21824_ (.Y(_04263_),
    .A(_04144_));
 sg13g2_a21oi_1 _21825_ (.A1(_04145_),
    .A2(_04262_),
    .Y(_04264_),
    .B1(_04263_));
 sg13g2_o21ai_1 _21826_ (.B1(_04264_),
    .Y(_04265_),
    .A1(_04185_),
    .A2(_04261_));
 sg13g2_xnor2_1 _21827_ (.Y(_04266_),
    .A(_04256_),
    .B(_04265_));
 sg13g2_nand2b_1 _21828_ (.Y(_04267_),
    .B(_11001_),
    .A_N(_11040_));
 sg13g2_xor2_1 _21829_ (.B(_04256_),
    .A(_04267_),
    .X(_04268_));
 sg13g2_and4_1 _21830_ (.A(_04106_),
    .B(_04083_),
    .C(_04107_),
    .D(_04108_),
    .X(_04269_));
 sg13g2_buf_1 _21831_ (.A(_04269_),
    .X(_04270_));
 sg13g2_nand2_1 _21832_ (.Y(_04271_),
    .A(_11485_),
    .B(net113));
 sg13g2_mux2_1 _21833_ (.A0(net1040),
    .A1(net1041),
    .S(_04271_),
    .X(_04272_));
 sg13g2_nand2_1 _21834_ (.Y(_04273_),
    .A(net203),
    .B(_11028_));
 sg13g2_o21ai_1 _21835_ (.B1(_04273_),
    .Y(_04274_),
    .A1(net1027),
    .A2(_04272_));
 sg13g2_o21ai_1 _21836_ (.B1(_04033_),
    .Y(_04275_),
    .A1(net119),
    .A2(_04048_));
 sg13g2_a22oi_1 _21837_ (.Y(_04276_),
    .B1(_04212_),
    .B2(net1042),
    .A2(net190),
    .A1(net298));
 sg13g2_inv_1 _21838_ (.Y(_04277_),
    .A(_04276_));
 sg13g2_a22oi_1 _21839_ (.Y(_04278_),
    .B1(_04277_),
    .B2(net118),
    .A2(_04275_),
    .A1(net190));
 sg13g2_nand2_1 _21840_ (.Y(_04279_),
    .A(_04217_),
    .B(net134));
 sg13g2_inv_1 _21841_ (.Y(_04280_),
    .A(_04279_));
 sg13g2_nor3_1 _21842_ (.A(net834),
    .B(_04278_),
    .C(_04280_),
    .Y(_04281_));
 sg13g2_a21oi_1 _21843_ (.A1(net1043),
    .A2(net247),
    .Y(_04282_),
    .B1(_04281_));
 sg13g2_nand2_1 _21844_ (.Y(_04283_),
    .A(net204),
    .B(net192));
 sg13g2_and2_1 _21845_ (.A(net164),
    .B(_04283_),
    .X(_04284_));
 sg13g2_nor2_2 _21846_ (.A(_04038_),
    .B(_04014_),
    .Y(_04285_));
 sg13g2_a22oi_1 _21847_ (.Y(_04286_),
    .B1(_04285_),
    .B2(net133),
    .A2(net161),
    .A1(net162));
 sg13g2_a22oi_1 _21848_ (.Y(_04287_),
    .B1(_04232_),
    .B2(_11351_),
    .A2(_04060_),
    .A1(net168));
 sg13g2_a22oi_1 _21849_ (.Y(_04288_),
    .B1(net173),
    .B2(_04062_),
    .A2(_04040_),
    .A1(net229));
 sg13g2_and4_1 _21850_ (.A(_04284_),
    .B(_04286_),
    .C(_04287_),
    .D(_04288_),
    .X(_04289_));
 sg13g2_buf_1 _21851_ (.A(_10669_),
    .X(_04290_));
 sg13g2_nand2_1 _21852_ (.Y(_04291_),
    .A(net170),
    .B(net172));
 sg13g2_o21ai_1 _21853_ (.B1(_04291_),
    .Y(_04292_),
    .A1(net160),
    .A2(_04223_));
 sg13g2_a221oi_1 _21854_ (.B2(net132),
    .C1(_04292_),
    .B1(_04070_),
    .A1(net167),
    .Y(_04293_),
    .A2(net136));
 sg13g2_o21ai_1 _21855_ (.B1(_09731_),
    .Y(_04294_),
    .A1(net137),
    .A2(net164));
 sg13g2_a21o_1 _21856_ (.A2(_04293_),
    .A1(_04289_),
    .B1(_04294_),
    .X(_04295_));
 sg13g2_nand4_1 _21857_ (.B(_04274_),
    .C(_04282_),
    .A(_04208_),
    .Y(_04296_),
    .D(_04295_));
 sg13g2_a221oi_1 _21858_ (.B2(net632),
    .C1(_04296_),
    .B1(_04268_),
    .A1(net1063),
    .Y(_04297_),
    .A2(_04266_));
 sg13g2_a21o_1 _21859_ (.A2(_04002_),
    .A1(_11793_),
    .B1(_04297_),
    .X(_04298_));
 sg13g2_nand3_1 _21860_ (.B(_08629_),
    .C(_04251_),
    .A(_08639_),
    .Y(_04299_));
 sg13g2_xnor2_1 _21861_ (.Y(_04300_),
    .A(_11002_),
    .B(_04299_));
 sg13g2_a22oi_1 _21862_ (.Y(_04301_),
    .B1(_04300_),
    .B2(net83),
    .A2(net32),
    .A1(_08464_));
 sg13g2_o21ai_1 _21863_ (.B1(_04301_),
    .Y(_00959_),
    .A1(net77),
    .A2(_04298_));
 sg13g2_a21o_1 _21864_ (.A2(_11041_),
    .A1(_11001_),
    .B1(_11178_),
    .X(_04302_));
 sg13g2_buf_1 _21865_ (.A(_04302_),
    .X(_04303_));
 sg13g2_xnor2_1 _21866_ (.Y(_04304_),
    .A(net142),
    .B(net131));
 sg13g2_xor2_1 _21867_ (.B(_04304_),
    .A(_04303_),
    .X(_04305_));
 sg13g2_nor2_1 _21868_ (.A(net203),
    .B(_04260_),
    .Y(_04306_));
 sg13g2_a21oi_1 _21869_ (.A1(_11157_),
    .A2(_04144_),
    .Y(_04307_),
    .B1(_11177_));
 sg13g2_a221oi_1 _21870_ (.B2(_04187_),
    .C1(_04307_),
    .B1(_04306_),
    .A1(_11028_),
    .Y(_04308_),
    .A2(_04265_));
 sg13g2_buf_1 _21871_ (.A(_04308_),
    .X(_04309_));
 sg13g2_xnor2_1 _21872_ (.Y(_04310_),
    .A(_04304_),
    .B(net30));
 sg13g2_a22oi_1 _21873_ (.Y(_04311_),
    .B1(_04051_),
    .B2(net118),
    .A2(net134),
    .A1(net135));
 sg13g2_o21ai_1 _21874_ (.B1(net1042),
    .Y(_04312_),
    .A1(net146),
    .A2(net134));
 sg13g2_nand2_1 _21875_ (.Y(_04313_),
    .A(_11100_),
    .B(net134));
 sg13g2_nand2b_1 _21876_ (.Y(_04314_),
    .B(_04313_),
    .A_N(_04312_));
 sg13g2_o21ai_1 _21877_ (.B1(_04314_),
    .Y(_04315_),
    .A1(_09713_),
    .A2(_04311_));
 sg13g2_a21oi_1 _21878_ (.A1(net1043),
    .A2(_10541_),
    .Y(_04316_),
    .B1(_04315_));
 sg13g2_nor2_1 _21879_ (.A(net143),
    .B(net131),
    .Y(_04317_));
 sg13g2_mux2_1 _21880_ (.A0(net1041),
    .A1(net1040),
    .S(_04317_),
    .X(_04318_));
 sg13g2_o21ai_1 _21881_ (.B1(_11182_),
    .Y(_04319_),
    .A1(net1027),
    .A2(_04318_));
 sg13g2_nand2_1 _21882_ (.Y(_04320_),
    .A(_11028_),
    .B(net96));
 sg13g2_nor2_1 _21883_ (.A(_10128_),
    .B(_03752_),
    .Y(_04321_));
 sg13g2_a21oi_1 _21884_ (.A1(_03753_),
    .A2(net213),
    .Y(_04322_),
    .B1(_04321_));
 sg13g2_a22oi_1 _21885_ (.Y(_04323_),
    .B1(_04322_),
    .B2(net245),
    .A2(_11481_),
    .A1(net191));
 sg13g2_a21oi_1 _21886_ (.A1(net137),
    .A2(net192),
    .Y(_04324_),
    .B1(net134));
 sg13g2_nand2_1 _21887_ (.Y(_04325_),
    .A(_11351_),
    .B(_04064_));
 sg13g2_nand3_1 _21888_ (.B(_04324_),
    .C(_04325_),
    .A(_04061_),
    .Y(_04326_));
 sg13g2_nor2_1 _21889_ (.A(net242),
    .B(net160),
    .Y(_04327_));
 sg13g2_a21oi_1 _21890_ (.A1(net133),
    .A2(net242),
    .Y(_04328_),
    .B1(_04327_));
 sg13g2_nor3_1 _21891_ (.A(net241),
    .B(_04033_),
    .C(_04328_),
    .Y(_04329_));
 sg13g2_a22oi_1 _21892_ (.Y(_04330_),
    .B1(_04285_),
    .B2(net132),
    .A2(_04233_),
    .A1(_04045_));
 sg13g2_nand2_1 _21893_ (.Y(_04331_),
    .A(_10817_),
    .B(net173));
 sg13g2_nand2_1 _21894_ (.Y(_04332_),
    .A(net204),
    .B(_04231_));
 sg13g2_nand3_1 _21895_ (.B(_04331_),
    .C(_04332_),
    .A(_04330_),
    .Y(_04333_));
 sg13g2_nor3_1 _21896_ (.A(_04326_),
    .B(_04329_),
    .C(_04333_),
    .Y(_04334_));
 sg13g2_o21ai_1 _21897_ (.B1(_04334_),
    .Y(_04335_),
    .A1(_04035_),
    .A2(_04323_));
 sg13g2_nand3_1 _21898_ (.B(_04320_),
    .C(_04335_),
    .A(net1026),
    .Y(_04336_));
 sg13g2_nand4_1 _21899_ (.B(_04316_),
    .C(_04319_),
    .A(_04208_),
    .Y(_04337_),
    .D(_04336_));
 sg13g2_a221oi_1 _21900_ (.B2(net1063),
    .C1(_04337_),
    .B1(_04310_),
    .A1(net632),
    .Y(_04338_),
    .A2(_04305_));
 sg13g2_a21o_1 _21901_ (.A2(_04002_),
    .A1(_11823_),
    .B1(_04338_),
    .X(_04339_));
 sg13g2_nor2_1 _21902_ (.A(_08229_),
    .B(_04299_),
    .Y(_04340_));
 sg13g2_xnor2_1 _21903_ (.Y(_04341_),
    .A(_11125_),
    .B(_04340_));
 sg13g2_a22oi_1 _21904_ (.Y(_04342_),
    .B1(_04341_),
    .B2(net83),
    .A2(net32),
    .A1(net616));
 sg13g2_o21ai_1 _21905_ (.B1(_04342_),
    .Y(_00960_),
    .A1(net77),
    .A2(_04339_));
 sg13g2_nand2_1 _21906_ (.Y(_04343_),
    .A(_11845_),
    .B(_04002_));
 sg13g2_nand2_1 _21907_ (.Y(_04344_),
    .A(net179),
    .B(net119));
 sg13g2_nand2_2 _21908_ (.Y(_04345_),
    .A(_11073_),
    .B(_11098_));
 sg13g2_and2_1 _21909_ (.A(_04344_),
    .B(_04345_),
    .X(_04346_));
 sg13g2_buf_1 _21910_ (.A(_04346_),
    .X(_04347_));
 sg13g2_nor2_1 _21911_ (.A(net142),
    .B(net131),
    .Y(_04348_));
 sg13g2_or2_1 _21912_ (.X(_04349_),
    .B(net30),
    .A(_04348_));
 sg13g2_nand2_1 _21913_ (.Y(_04350_),
    .A(_04344_),
    .B(_04345_));
 sg13g2_mux2_1 _21914_ (.A0(_04350_),
    .A1(net131),
    .S(net30),
    .X(_04351_));
 sg13g2_nand2_1 _21915_ (.Y(_04352_),
    .A(net131),
    .B(_04350_));
 sg13g2_o21ai_1 _21916_ (.B1(net1063),
    .Y(_04353_),
    .A1(net30),
    .A2(_04352_));
 sg13g2_a221oi_1 _21917_ (.B2(net142),
    .C1(_04353_),
    .B1(_04351_),
    .A1(_04347_),
    .Y(_04354_),
    .A2(_04349_));
 sg13g2_a22oi_1 _21918_ (.Y(_04355_),
    .B1(_04019_),
    .B2(net133),
    .A2(net113),
    .A1(net190));
 sg13g2_nor2_1 _21919_ (.A(_04048_),
    .B(_04355_),
    .Y(_04356_));
 sg13g2_a22oi_1 _21920_ (.Y(_04357_),
    .B1(_04019_),
    .B2(net132),
    .A2(_04017_),
    .A1(net191));
 sg13g2_nor2_1 _21921_ (.A(_04033_),
    .B(_04357_),
    .Y(_04358_));
 sg13g2_a22oi_1 _21922_ (.Y(_04359_),
    .B1(_04285_),
    .B2(net162),
    .A2(net166),
    .A1(_10678_));
 sg13g2_nand2_1 _21923_ (.Y(_04360_),
    .A(_04046_),
    .B(_04070_));
 sg13g2_nand2_1 _21924_ (.Y(_04361_),
    .A(net137),
    .B(_04231_));
 sg13g2_nand3_1 _21925_ (.B(_04360_),
    .C(_04361_),
    .A(_04359_),
    .Y(_04362_));
 sg13g2_nor3_1 _21926_ (.A(_04356_),
    .B(_04358_),
    .C(_04362_),
    .Y(_04363_));
 sg13g2_nor2_1 _21927_ (.A(_04151_),
    .B(_04223_),
    .Y(_04364_));
 sg13g2_a21oi_1 _21928_ (.A1(net229),
    .A2(net161),
    .Y(_04365_),
    .B1(_04364_));
 sg13g2_a21oi_1 _21929_ (.A1(net167),
    .A2(net173),
    .Y(_04366_),
    .B1(net112));
 sg13g2_a22oi_1 _21930_ (.Y(_04367_),
    .B1(_04054_),
    .B2(_11351_),
    .A2(net171),
    .A1(net168));
 sg13g2_nand4_1 _21931_ (.B(_04365_),
    .C(_04366_),
    .A(_04363_),
    .Y(_04368_),
    .D(_04367_));
 sg13g2_nand3_1 _21932_ (.B(_04279_),
    .C(_04368_),
    .A(net1026),
    .Y(_04369_));
 sg13g2_nand2_1 _21933_ (.Y(_04370_),
    .A(_04317_),
    .B(_04347_));
 sg13g2_o21ai_1 _21934_ (.B1(_04370_),
    .Y(_04371_),
    .A1(_11182_),
    .A2(_04347_));
 sg13g2_nand2_1 _21935_ (.Y(_04372_),
    .A(net1041),
    .B(_04350_));
 sg13g2_nand4_1 _21936_ (.B(net142),
    .C(net131),
    .A(net1123),
    .Y(_04373_),
    .D(_04347_));
 sg13g2_a22oi_1 _21937_ (.Y(_04374_),
    .B1(_11181_),
    .B2(net1040),
    .A2(net201),
    .A1(net1114));
 sg13g2_nand2_1 _21938_ (.Y(_04375_),
    .A(net147),
    .B(net119));
 sg13g2_a22oi_1 _21939_ (.Y(_04376_),
    .B1(net96),
    .B2(_04213_),
    .A2(_04375_),
    .A1(_09718_));
 sg13g2_nand4_1 _21940_ (.B(_04373_),
    .C(_04374_),
    .A(_04372_),
    .Y(_04377_),
    .D(_04376_));
 sg13g2_a21oi_1 _21941_ (.A1(net632),
    .A2(_04371_),
    .Y(_04378_),
    .B1(_04377_));
 sg13g2_nand2_1 _21942_ (.Y(_04379_),
    .A(_04369_),
    .B(_04378_));
 sg13g2_nand2_1 _21943_ (.Y(_04380_),
    .A(net1042),
    .B(_11234_));
 sg13g2_buf_2 _21944_ (.A(_04380_),
    .X(_04381_));
 sg13g2_nand2_1 _21945_ (.Y(_04382_),
    .A(_04381_),
    .B(_04208_));
 sg13g2_nand3_1 _21946_ (.B(net632),
    .C(_04347_),
    .A(_11182_),
    .Y(_04383_));
 sg13g2_nor3_1 _21947_ (.A(_04110_),
    .B(_04317_),
    .C(_04347_),
    .Y(_04384_));
 sg13g2_nor2_1 _21948_ (.A(_04303_),
    .B(_04384_),
    .Y(_04385_));
 sg13g2_a21oi_1 _21949_ (.A1(_04303_),
    .A2(_04383_),
    .Y(_04386_),
    .B1(_04385_));
 sg13g2_or4_1 _21950_ (.A(_04354_),
    .B(_04379_),
    .C(_04382_),
    .D(_04386_),
    .X(_04387_));
 sg13g2_nand2_1 _21951_ (.Y(_04388_),
    .A(_04343_),
    .B(_04387_));
 sg13g2_nand2_1 _21952_ (.Y(_04389_),
    .A(net616),
    .B(_04340_));
 sg13g2_xnor2_1 _21953_ (.Y(_04390_),
    .A(_11068_),
    .B(_04389_));
 sg13g2_a22oi_1 _21954_ (.Y(_04391_),
    .B1(_04390_),
    .B2(net83),
    .A2(net32),
    .A1(_08438_));
 sg13g2_o21ai_1 _21955_ (.B1(_04391_),
    .Y(_00961_),
    .A1(net77),
    .A2(_04388_));
 sg13g2_nor3_1 _21956_ (.A(net143),
    .B(net30),
    .C(_04345_),
    .Y(_04392_));
 sg13g2_xnor2_1 _21957_ (.Y(_04393_),
    .A(_11445_),
    .B(net146));
 sg13g2_buf_2 _21958_ (.A(_04393_),
    .X(_04394_));
 sg13g2_nor3_1 _21959_ (.A(net179),
    .B(net131),
    .C(_04394_),
    .Y(_04395_));
 sg13g2_o21ai_1 _21960_ (.B1(_04395_),
    .Y(_04396_),
    .A1(net143),
    .A2(net30));
 sg13g2_nor2b_1 _21961_ (.A(_04392_),
    .B_N(_04396_),
    .Y(_04397_));
 sg13g2_o21ai_1 _21962_ (.B1(_04344_),
    .Y(_04398_),
    .A1(net143),
    .A2(net30));
 sg13g2_nand2_1 _21963_ (.Y(_04399_),
    .A(net143),
    .B(net30));
 sg13g2_nor2b_1 _21964_ (.A(_04394_),
    .B_N(_04345_),
    .Y(_04400_));
 sg13g2_nor2_1 _21965_ (.A(net114),
    .B(_04400_),
    .Y(_04401_));
 sg13g2_a22oi_1 _21966_ (.Y(_04402_),
    .B1(_04344_),
    .B2(net143),
    .A2(net114),
    .A1(net135));
 sg13g2_nor2_1 _21967_ (.A(_04394_),
    .B(_04402_),
    .Y(_04403_));
 sg13g2_nand2_1 _21968_ (.Y(_04404_),
    .A(net135),
    .B(_04348_));
 sg13g2_o21ai_1 _21969_ (.B1(net1123),
    .Y(_04405_),
    .A1(_04394_),
    .A2(_04404_));
 sg13g2_a21o_1 _21970_ (.A2(_04403_),
    .A1(_04309_),
    .B1(_04405_),
    .X(_04406_));
 sg13g2_a221oi_1 _21971_ (.B2(_04401_),
    .C1(_04406_),
    .B1(_04399_),
    .A1(_04394_),
    .Y(_04407_),
    .A2(_04398_));
 sg13g2_xnor2_1 _21972_ (.Y(_04408_),
    .A(_11185_),
    .B(_04394_));
 sg13g2_nor2_1 _21973_ (.A(net298),
    .B(net292),
    .Y(_04409_));
 sg13g2_nand2_1 _21974_ (.Y(_04410_),
    .A(_11351_),
    .B(_04409_));
 sg13g2_nor2_1 _21975_ (.A(_04151_),
    .B(net297),
    .Y(_04411_));
 sg13g2_nor2_1 _21976_ (.A(net237),
    .B(net160),
    .Y(_04412_));
 sg13g2_o21ai_1 _21977_ (.B1(net245),
    .Y(_04413_),
    .A1(_04411_),
    .A2(_04412_));
 sg13g2_a21oi_1 _21978_ (.A1(_04410_),
    .A2(_04413_),
    .Y(_04414_),
    .B1(_04028_));
 sg13g2_nor2_1 _21979_ (.A(_10128_),
    .B(_11369_),
    .Y(_04415_));
 sg13g2_a21oi_1 _21980_ (.A1(net200),
    .A2(_11542_),
    .Y(_04416_),
    .B1(_04415_));
 sg13g2_nand2_1 _21981_ (.Y(_04417_),
    .A(_10348_),
    .B(_04103_));
 sg13g2_o21ai_1 _21982_ (.B1(_04417_),
    .Y(_04418_),
    .A1(net293),
    .A2(_04416_));
 sg13g2_a21oi_1 _21983_ (.A1(_10939_),
    .A2(_04064_),
    .Y(_04419_),
    .B1(_04087_));
 sg13g2_a22oi_1 _21984_ (.Y(_04420_),
    .B1(net192),
    .B2(net114),
    .A2(net171),
    .A1(net167));
 sg13g2_nand2_1 _21985_ (.Y(_04421_),
    .A(net168),
    .B(net172));
 sg13g2_a22oi_1 _21986_ (.Y(_04422_),
    .B1(_04285_),
    .B2(_04045_),
    .A2(_04070_),
    .A1(net229));
 sg13g2_nand4_1 _21987_ (.B(_04420_),
    .C(_04421_),
    .A(_04419_),
    .Y(_04423_),
    .D(_04422_));
 sg13g2_a221oi_1 _21988_ (.B2(net191),
    .C1(_04423_),
    .B1(net161),
    .A1(net113),
    .Y(_04424_),
    .A2(net189));
 sg13g2_o21ai_1 _21989_ (.B1(_04424_),
    .Y(_04425_),
    .A1(_04014_),
    .A2(_04418_));
 sg13g2_and2_1 _21990_ (.A(net1026),
    .B(_04313_),
    .X(_04426_));
 sg13g2_o21ai_1 _21991_ (.B1(_04426_),
    .Y(_04427_),
    .A1(_04414_),
    .A2(_04425_));
 sg13g2_nor2_1 _21992_ (.A(_11533_),
    .B(_04345_),
    .Y(_04428_));
 sg13g2_mux2_1 _21993_ (.A0(net1113),
    .A1(_08932_),
    .S(_11238_),
    .X(_04429_));
 sg13g2_nor2_1 _21994_ (.A(_09718_),
    .B(_04429_),
    .Y(_04430_));
 sg13g2_nor2_1 _21995_ (.A(_11237_),
    .B(_04430_),
    .Y(_04431_));
 sg13g2_a221oi_1 _21996_ (.B2(_04428_),
    .C1(_04431_),
    .B1(_04394_),
    .A1(net1043),
    .Y(_04432_),
    .A2(net223));
 sg13g2_nand4_1 _21997_ (.B(_04208_),
    .C(_04427_),
    .A(_04381_),
    .Y(_04433_),
    .D(_04432_));
 sg13g2_a221oi_1 _21998_ (.B2(net632),
    .C1(_04433_),
    .B1(_04408_),
    .A1(_04397_),
    .Y(_04434_),
    .A2(_04407_));
 sg13g2_a21o_1 _21999_ (.A2(_04002_),
    .A1(_11881_),
    .B1(_04434_),
    .X(_04435_));
 sg13g2_nand3_1 _22000_ (.B(net906),
    .C(_04340_),
    .A(_08339_),
    .Y(_04436_));
 sg13g2_xnor2_1 _22001_ (.Y(_04437_),
    .A(_11214_),
    .B(_04436_));
 sg13g2_a22oi_1 _22002_ (.Y(_04438_),
    .B1(_04437_),
    .B2(net83),
    .A2(net32),
    .A1(_08231_));
 sg13g2_o21ai_1 _22003_ (.B1(_04438_),
    .Y(_00962_),
    .A1(net77),
    .A2(_04435_));
 sg13g2_buf_1 _22004_ (.A(net387),
    .X(_04439_));
 sg13g2_nor4_1 _22005_ (.A(net1122),
    .B(_10260_),
    .C(net897),
    .D(net1031),
    .Y(_04440_));
 sg13g2_nand2_1 _22006_ (.Y(_04441_),
    .A(net290),
    .B(_04440_));
 sg13g2_a21oi_1 _22007_ (.A1(net1044),
    .A2(net95),
    .Y(_04442_),
    .B1(_04140_));
 sg13g2_a21oi_1 _22008_ (.A1(net688),
    .A2(net95),
    .Y(_04443_),
    .B1(net691));
 sg13g2_a21o_1 _22009_ (.A2(_04442_),
    .A1(net691),
    .B1(_04443_),
    .X(_04444_));
 sg13g2_nand2_2 _22010_ (.Y(_04445_),
    .A(net291),
    .B(_11538_));
 sg13g2_nand2_1 _22011_ (.Y(_04446_),
    .A(_10505_),
    .B(_04231_));
 sg13g2_a22oi_1 _22012_ (.Y(_04447_),
    .B1(net161),
    .B2(net113),
    .A2(net165),
    .A1(net168));
 sg13g2_nor2_1 _22013_ (.A(net213),
    .B(_04048_),
    .Y(_04448_));
 sg13g2_a21oi_1 _22014_ (.A1(net293),
    .A2(_04381_),
    .Y(_04449_),
    .B1(net244));
 sg13g2_o21ai_1 _22015_ (.B1(_04216_),
    .Y(_04450_),
    .A1(_04448_),
    .A2(_04449_));
 sg13g2_nand2_1 _22016_ (.Y(_04451_),
    .A(_04057_),
    .B(net292));
 sg13g2_o21ai_1 _22017_ (.B1(_04451_),
    .Y(_04452_),
    .A1(_10856_),
    .A2(net237));
 sg13g2_nor2_1 _22018_ (.A(net160),
    .B(_04048_),
    .Y(_04453_));
 sg13g2_a21o_1 _22019_ (.A2(_04452_),
    .A1(net245),
    .B1(_04453_),
    .X(_04454_));
 sg13g2_nand2_1 _22020_ (.Y(_04455_),
    .A(net237),
    .B(net137));
 sg13g2_o21ai_1 _22021_ (.B1(_04455_),
    .Y(_04456_),
    .A1(net237),
    .A2(net131));
 sg13g2_mux2_1 _22022_ (.A0(_04411_),
    .A1(_04456_),
    .S(net298),
    .X(_04457_));
 sg13g2_nand3_1 _22023_ (.B(net244),
    .C(net118),
    .A(_08911_),
    .Y(_04458_));
 sg13g2_nand2_1 _22024_ (.Y(_04459_),
    .A(net298),
    .B(_11234_));
 sg13g2_o21ai_1 _22025_ (.B1(_04459_),
    .Y(_04460_),
    .A1(net298),
    .A2(_11100_));
 sg13g2_nand2_1 _22026_ (.Y(_04461_),
    .A(net237),
    .B(_04460_));
 sg13g2_a21oi_1 _22027_ (.A1(_04458_),
    .A2(_04461_),
    .Y(_04462_),
    .B1(_04014_));
 sg13g2_a221oi_1 _22028_ (.B2(_04017_),
    .C1(_04462_),
    .B1(_04457_),
    .A1(_04222_),
    .Y(_04463_),
    .A2(_04454_));
 sg13g2_nand4_1 _22029_ (.B(_04447_),
    .C(_04450_),
    .A(_04446_),
    .Y(_04464_),
    .D(_04463_));
 sg13g2_nor2_1 _22030_ (.A(net170),
    .B(net164),
    .Y(_04465_));
 sg13g2_nor2_1 _22031_ (.A(net834),
    .B(_04465_),
    .Y(_04466_));
 sg13g2_o21ai_1 _22032_ (.B1(_04163_),
    .Y(_04467_),
    .A1(_04165_),
    .A2(_04164_));
 sg13g2_xnor2_1 _22033_ (.Y(_04468_),
    .A(net162),
    .B(net241));
 sg13g2_xnor2_1 _22034_ (.Y(_04469_),
    .A(_04467_),
    .B(_04468_));
 sg13g2_a22oi_1 _22035_ (.Y(_04470_),
    .B1(_04051_),
    .B2(_04093_),
    .A2(net112),
    .A1(net132));
 sg13g2_inv_1 _22036_ (.Y(_04471_),
    .A(_04470_));
 sg13g2_a221oi_1 _22037_ (.B2(_09732_),
    .C1(net291),
    .B1(_04471_),
    .A1(net1043),
    .Y(_04472_),
    .A2(_10996_));
 sg13g2_inv_1 _22038_ (.Y(_04473_),
    .A(_09718_));
 sg13g2_o21ai_1 _22039_ (.B1(net1041),
    .Y(_04474_),
    .A1(_11389_),
    .A2(net241));
 sg13g2_nand3_1 _22040_ (.B(net162),
    .C(_11565_),
    .A(_08959_),
    .Y(_04475_));
 sg13g2_nand3_1 _22041_ (.B(_04474_),
    .C(_04475_),
    .A(_04473_),
    .Y(_04476_));
 sg13g2_nand2b_1 _22042_ (.Y(_04477_),
    .B(_04476_),
    .A_N(_10465_));
 sg13g2_nor3_1 _22043_ (.A(_10340_),
    .B(_10351_),
    .C(_10355_),
    .Y(_04478_));
 sg13g2_xnor2_1 _22044_ (.Y(_04479_),
    .A(_04478_),
    .B(_04468_));
 sg13g2_nand2_1 _22045_ (.Y(_04480_),
    .A(_04115_),
    .B(_04479_));
 sg13g2_nand3_1 _22046_ (.B(_04477_),
    .C(_04480_),
    .A(_04472_),
    .Y(_04481_));
 sg13g2_a221oi_1 _22047_ (.B2(_08122_),
    .C1(_04481_),
    .B1(_04469_),
    .A1(_04464_),
    .Y(_04482_),
    .A2(_04466_));
 sg13g2_nor2_1 _22048_ (.A(_04009_),
    .B(_04482_),
    .Y(_04483_));
 sg13g2_o21ai_1 _22049_ (.B1(_04483_),
    .Y(_04484_),
    .A1(_11579_),
    .A2(_04445_));
 sg13g2_nand3_1 _22050_ (.B(_04444_),
    .C(_04484_),
    .A(_04441_),
    .Y(_00963_));
 sg13g2_nor2b_1 _22051_ (.A(_00253_),
    .B_N(_04440_),
    .Y(_04485_));
 sg13g2_o21ai_1 _22052_ (.B1(net290),
    .Y(_04486_),
    .A1(_04136_),
    .A2(_04485_));
 sg13g2_nand3_1 _22053_ (.B(net688),
    .C(_04130_),
    .A(net691),
    .Y(_04487_));
 sg13g2_nand2_1 _22054_ (.Y(_04488_),
    .A(net691),
    .B(net688));
 sg13g2_a21oi_1 _22055_ (.A1(net95),
    .A2(_04488_),
    .Y(_04489_),
    .B1(_04140_));
 sg13g2_mux2_1 _22056_ (.A0(_04487_),
    .A1(_04489_),
    .S(net692),
    .X(_04490_));
 sg13g2_nor2_1 _22057_ (.A(_11586_),
    .B(_04478_),
    .Y(_04491_));
 sg13g2_a21oi_1 _22058_ (.A1(_10432_),
    .A2(_10464_),
    .Y(_04492_),
    .B1(_11389_));
 sg13g2_nor2_1 _22059_ (.A(_04491_),
    .B(_04492_),
    .Y(_04493_));
 sg13g2_xnor2_1 _22060_ (.Y(_04494_),
    .A(_10390_),
    .B(net300));
 sg13g2_xnor2_1 _22061_ (.Y(_04495_),
    .A(_04493_),
    .B(_04494_));
 sg13g2_a21oi_1 _22062_ (.A1(net244),
    .A2(net163),
    .Y(_04496_),
    .B1(net293));
 sg13g2_nor2_1 _22063_ (.A(net244),
    .B(_04381_),
    .Y(_04497_));
 sg13g2_o21ai_1 _22064_ (.B1(net190),
    .Y(_04498_),
    .A1(_04496_),
    .A2(_04497_));
 sg13g2_nor2_1 _22065_ (.A(net297),
    .B(_04290_),
    .Y(_04499_));
 sg13g2_nor2_1 _22066_ (.A(_04151_),
    .B(_03752_),
    .Y(_04500_));
 sg13g2_o21ai_1 _22067_ (.B1(net298),
    .Y(_04501_),
    .A1(_04499_),
    .A2(_04500_));
 sg13g2_a21oi_1 _22068_ (.A1(_04410_),
    .A2(_04501_),
    .Y(_04502_),
    .B1(_04028_));
 sg13g2_nand3_1 _22069_ (.B(_04019_),
    .C(_04011_),
    .A(_04038_),
    .Y(_04503_));
 sg13g2_a221oi_1 _22070_ (.B2(net146),
    .C1(_04224_),
    .B1(_04285_),
    .A1(net135),
    .Y(_04504_),
    .A2(_04070_));
 sg13g2_a22oi_1 _22071_ (.Y(_04505_),
    .B1(net161),
    .B2(net114),
    .A2(net171),
    .A1(net137));
 sg13g2_a22oi_1 _22072_ (.Y(_04506_),
    .B1(net192),
    .B2(net191),
    .A2(net172),
    .A1(net113));
 sg13g2_nand4_1 _22073_ (.B(_04504_),
    .C(_04505_),
    .A(_04503_),
    .Y(_04507_),
    .D(_04506_));
 sg13g2_nor2_1 _22074_ (.A(_04502_),
    .B(_04507_),
    .Y(_04508_));
 sg13g2_a221oi_1 _22075_ (.B2(_04508_),
    .C1(net834),
    .B1(_04498_),
    .A1(net213),
    .Y(_04509_),
    .A2(net96));
 sg13g2_or2_1 _22076_ (.X(_04510_),
    .B(_04166_),
    .A(_04160_));
 sg13g2_buf_1 _22077_ (.A(_04510_),
    .X(_04511_));
 sg13g2_xor2_1 _22078_ (.B(_04494_),
    .A(_04511_),
    .X(_04512_));
 sg13g2_mux2_1 _22079_ (.A0(_08932_),
    .A1(_08958_),
    .S(_10467_),
    .X(_04513_));
 sg13g2_or2_1 _22080_ (.X(_04514_),
    .B(_04513_),
    .A(_09718_));
 sg13g2_nand2_1 _22081_ (.Y(_04515_),
    .A(_10390_),
    .B(net300));
 sg13g2_nand2_1 _22082_ (.Y(_04516_),
    .A(_09731_),
    .B(net190));
 sg13g2_a21oi_1 _22083_ (.A1(net1114),
    .A2(net183),
    .Y(_04517_),
    .B1(_04097_));
 sg13g2_o21ai_1 _22084_ (.B1(_04517_),
    .Y(_04518_),
    .A1(_04418_),
    .A2(_04516_));
 sg13g2_a221oi_1 _22085_ (.B2(_04515_),
    .C1(_04518_),
    .B1(_04514_),
    .A1(_08121_),
    .Y(_04519_),
    .A2(_04512_));
 sg13g2_nor2b_1 _22086_ (.A(_04509_),
    .B_N(_04519_),
    .Y(_04520_));
 sg13g2_o21ai_1 _22087_ (.B1(_04520_),
    .Y(_04521_),
    .A1(_04112_),
    .A2(_04495_));
 sg13g2_nor2b_1 _22088_ (.A(_04009_),
    .B_N(_04521_),
    .Y(_04522_));
 sg13g2_o21ai_1 _22089_ (.B1(_04522_),
    .Y(_04523_),
    .A1(_11606_),
    .A2(_04445_));
 sg13g2_nand3_1 _22090_ (.B(_04490_),
    .C(_04523_),
    .A(_04486_),
    .Y(_00964_));
 sg13g2_a21o_1 _22091_ (.A2(_10466_),
    .A1(_10356_),
    .B1(_10467_),
    .X(_04524_));
 sg13g2_nand2_1 _22092_ (.Y(_04525_),
    .A(net247),
    .B(net213));
 sg13g2_nor2b_1 _22093_ (.A(_04168_),
    .B_N(_04525_),
    .Y(_04526_));
 sg13g2_xnor2_1 _22094_ (.Y(_04527_),
    .A(_04524_),
    .B(_04526_));
 sg13g2_nor2_1 _22095_ (.A(_11400_),
    .B(_04511_),
    .Y(_04528_));
 sg13g2_nand2_1 _22096_ (.Y(_04529_),
    .A(_11400_),
    .B(_04511_));
 sg13g2_o21ai_1 _22097_ (.B1(_04529_),
    .Y(_04530_),
    .A1(_10390_),
    .A2(_04528_));
 sg13g2_xor2_1 _22098_ (.B(_04530_),
    .A(_04526_),
    .X(_04531_));
 sg13g2_nor2_1 _22099_ (.A(net302),
    .B(net213),
    .Y(_04532_));
 sg13g2_mux2_1 _22100_ (.A0(_08933_),
    .A1(net1040),
    .S(_04532_),
    .X(_04533_));
 sg13g2_nand2_1 _22101_ (.Y(_04534_),
    .A(_11274_),
    .B(net213));
 sg13g2_o21ai_1 _22102_ (.B1(_04534_),
    .Y(_04535_),
    .A1(net1027),
    .A2(_04533_));
 sg13g2_a221oi_1 _22103_ (.B2(_04093_),
    .C1(_04089_),
    .B1(net165),
    .A1(net162),
    .Y(_04536_),
    .A2(net169));
 sg13g2_o21ai_1 _22104_ (.B1(_04536_),
    .Y(_04537_),
    .A1(_11383_),
    .A2(_04075_));
 sg13g2_nand3b_1 _22105_ (.B(_04537_),
    .C(net1026),
    .Y(_04538_),
    .A_N(_04465_));
 sg13g2_a21oi_1 _22106_ (.A1(net1043),
    .A2(_11485_),
    .Y(_04539_),
    .B1(net291));
 sg13g2_a22oi_1 _22107_ (.Y(_04540_),
    .B1(net169),
    .B2(net168),
    .A2(_04040_),
    .A1(_04068_));
 sg13g2_a21oi_1 _22108_ (.A1(_11482_),
    .A2(_04014_),
    .Y(_04541_),
    .B1(_04381_));
 sg13g2_a221oi_1 _22109_ (.B2(net118),
    .C1(_04541_),
    .B1(_04070_),
    .A1(_04016_),
    .Y(_04542_),
    .A2(_04031_));
 sg13g2_a21oi_1 _22110_ (.A1(_04057_),
    .A2(net189),
    .Y(_04543_),
    .B1(_04088_));
 sg13g2_a22oi_1 _22111_ (.Y(_04544_),
    .B1(net161),
    .B2(net135),
    .A2(net172),
    .A1(net114));
 sg13g2_nand4_1 _22112_ (.B(_04542_),
    .C(_04543_),
    .A(_04540_),
    .Y(_04545_),
    .D(_04544_));
 sg13g2_nor2_1 _22113_ (.A(_10856_),
    .B(net297),
    .Y(_04546_));
 sg13g2_nor2_1 _22114_ (.A(net293),
    .B(_04546_),
    .Y(_04547_));
 sg13g2_nor3_1 _22115_ (.A(net245),
    .B(_04499_),
    .C(_04500_),
    .Y(_04548_));
 sg13g2_nor3_1 _22116_ (.A(_04028_),
    .B(_04547_),
    .C(_04548_),
    .Y(_04549_));
 sg13g2_a21oi_1 _22117_ (.A1(_11377_),
    .A2(net96),
    .Y(_04550_),
    .B1(net834));
 sg13g2_o21ai_1 _22118_ (.B1(_04550_),
    .Y(_04551_),
    .A1(_04545_),
    .A2(_04549_));
 sg13g2_nand4_1 _22119_ (.B(_04538_),
    .C(_04539_),
    .A(_04535_),
    .Y(_04552_),
    .D(_04551_));
 sg13g2_a221oi_1 _22120_ (.B2(net1063),
    .C1(_04552_),
    .B1(_04531_),
    .A1(_04115_),
    .Y(_04553_),
    .A2(_04527_));
 sg13g2_inv_1 _22121_ (.Y(_04554_),
    .A(_04553_));
 sg13g2_o21ai_1 _22122_ (.B1(_04554_),
    .Y(_04555_),
    .A1(_11500_),
    .A2(\cpu.ex.c_mult[4] ));
 sg13g2_nand2_1 _22123_ (.Y(_04556_),
    .A(net688),
    .B(net788));
 sg13g2_a21o_1 _22124_ (.A2(_04556_),
    .A1(_04130_),
    .B1(_04140_),
    .X(_04557_));
 sg13g2_nor2_1 _22125_ (.A(net1046),
    .B(_04556_),
    .Y(_04558_));
 sg13g2_nor4_1 _22126_ (.A(net1122),
    .B(net387),
    .C(_09123_),
    .D(_04132_),
    .Y(_04559_));
 sg13g2_a221oi_1 _22127_ (.B2(net95),
    .C1(_04559_),
    .B1(_04558_),
    .A1(net1046),
    .Y(_04560_),
    .A2(_04557_));
 sg13g2_o21ai_1 _22128_ (.B1(_04560_),
    .Y(_00965_),
    .A1(net77),
    .A2(_04555_));
 sg13g2_buf_1 _22129_ (.A(_08673_),
    .X(_04561_));
 sg13g2_nand2_1 _22130_ (.Y(_04562_),
    .A(net1046),
    .B(_04247_));
 sg13g2_xor2_1 _22131_ (.B(_04562_),
    .A(_10469_),
    .X(_04563_));
 sg13g2_a22oi_1 _22132_ (.Y(_04564_),
    .B1(_04563_),
    .B2(net83),
    .A2(net32),
    .A1(net957));
 sg13g2_nand2b_1 _22133_ (.Y(_04565_),
    .B(_04173_),
    .A_N(_04167_));
 sg13g2_o21ai_1 _22134_ (.B1(_04525_),
    .Y(_04566_),
    .A1(_04168_),
    .A2(_04530_));
 sg13g2_xor2_1 _22135_ (.B(_04566_),
    .A(_04565_),
    .X(_04567_));
 sg13g2_a21oi_1 _22136_ (.A1(_04524_),
    .A2(_04534_),
    .Y(_04568_),
    .B1(_04532_));
 sg13g2_xnor2_1 _22137_ (.Y(_04569_),
    .A(_04565_),
    .B(_04568_));
 sg13g2_nand2b_1 _22138_ (.Y(_04570_),
    .B(_10802_),
    .A_N(_08932_));
 sg13g2_o21ai_1 _22139_ (.B1(_04570_),
    .Y(_04571_),
    .A1(net1113),
    .A2(_10802_));
 sg13g2_a21o_1 _22140_ (.A2(_04571_),
    .A1(_04473_),
    .B1(_10804_),
    .X(_04572_));
 sg13g2_a22oi_1 _22141_ (.Y(_04573_),
    .B1(net189),
    .B2(net162),
    .A2(net169),
    .A1(net170));
 sg13g2_a221oi_1 _22142_ (.B2(net132),
    .C1(_04089_),
    .B1(net165),
    .A1(net133),
    .Y(_04574_),
    .A2(net136));
 sg13g2_o21ai_1 _22143_ (.B1(_09731_),
    .Y(_04575_),
    .A1(net229),
    .A2(net164));
 sg13g2_a21o_1 _22144_ (.A2(_04574_),
    .A1(_04573_),
    .B1(_04575_),
    .X(_04576_));
 sg13g2_a21oi_1 _22145_ (.A1(net1114),
    .A2(_11846_),
    .Y(_04577_),
    .B1(_04097_));
 sg13g2_nand2_1 _22146_ (.Y(_04578_),
    .A(_11586_),
    .B(_04012_));
 sg13g2_a22oi_1 _22147_ (.Y(_04579_),
    .B1(_04578_),
    .B2(net242),
    .A2(net190),
    .A1(net237));
 sg13g2_nand2_1 _22148_ (.Y(_04580_),
    .A(net297),
    .B(_04290_));
 sg13g2_nand3_1 _22149_ (.B(net190),
    .C(_04580_),
    .A(net298),
    .Y(_04581_));
 sg13g2_o21ai_1 _22150_ (.B1(_04581_),
    .Y(_04582_),
    .A1(_04381_),
    .A2(_04579_));
 sg13g2_nand2_1 _22151_ (.Y(_04583_),
    .A(net167),
    .B(net192));
 sg13g2_a22oi_1 _22152_ (.Y(_04584_),
    .B1(net166),
    .B2(net137),
    .A2(net172),
    .A1(net135));
 sg13g2_and2_1 _22153_ (.A(_10967_),
    .B(_04053_),
    .X(_04585_));
 sg13g2_a21o_1 _22154_ (.A2(_04039_),
    .A1(net114),
    .B1(_04585_),
    .X(_04586_));
 sg13g2_a221oi_1 _22155_ (.B2(net146),
    .C1(_04586_),
    .B1(net161),
    .A1(net113),
    .Y(_04587_),
    .A2(net173));
 sg13g2_nand4_1 _22156_ (.B(_04583_),
    .C(_04584_),
    .A(_04325_),
    .Y(_04588_),
    .D(_04587_));
 sg13g2_a21oi_1 _22157_ (.A1(_04191_),
    .A2(net112),
    .Y(_04589_),
    .B1(net834));
 sg13g2_o21ai_1 _22158_ (.B1(_04589_),
    .Y(_04590_),
    .A1(_04582_),
    .A2(_04588_));
 sg13g2_nand4_1 _22159_ (.B(_04576_),
    .C(_04577_),
    .A(_04572_),
    .Y(_04591_),
    .D(_04590_));
 sg13g2_a221oi_1 _22160_ (.B2(_04115_),
    .C1(_04591_),
    .B1(_04569_),
    .A1(net1063),
    .Y(_04592_),
    .A2(_04567_));
 sg13g2_nor2_1 _22161_ (.A(_04009_),
    .B(_04592_),
    .Y(_04593_));
 sg13g2_o21ai_1 _22162_ (.B1(_04593_),
    .Y(_04594_),
    .A1(_11639_),
    .A2(_04445_));
 sg13g2_nand2_1 _22163_ (.Y(_00966_),
    .A(_04564_),
    .B(_04594_));
 sg13g2_xnor2_1 _22164_ (.Y(_04595_),
    .A(_10814_),
    .B(_04248_));
 sg13g2_a22oi_1 _22165_ (.Y(_04596_),
    .B1(_04595_),
    .B2(net83),
    .A2(net32),
    .A1(\cpu.ex.pc[6] ));
 sg13g2_xnor2_1 _22166_ (.Y(_04597_),
    .A(_10739_),
    .B(_04201_));
 sg13g2_a22oi_1 _22167_ (.Y(_04598_),
    .B1(net172),
    .B2(_11235_),
    .A2(net171),
    .A1(net135));
 sg13g2_a21oi_1 _22168_ (.A1(_04023_),
    .A2(net173),
    .Y(_04599_),
    .B1(_04364_));
 sg13g2_a22oi_1 _22169_ (.Y(_04600_),
    .B1(net166),
    .B2(_11157_),
    .A2(net136),
    .A1(net137));
 sg13g2_a21oi_1 _22170_ (.A1(_10856_),
    .A2(_11542_),
    .Y(_04601_),
    .B1(_10348_));
 sg13g2_o21ai_1 _22171_ (.B1(_04216_),
    .Y(_04602_),
    .A1(_04453_),
    .A2(_04601_));
 sg13g2_nand4_1 _22172_ (.B(_04599_),
    .C(_04600_),
    .A(_04598_),
    .Y(_04603_),
    .D(_04602_));
 sg13g2_a21o_1 _22173_ (.A2(_04603_),
    .A1(_09712_),
    .B1(net1042),
    .X(_04604_));
 sg13g2_o21ai_1 _22174_ (.B1(_11584_),
    .Y(_04605_),
    .A1(net297),
    .A2(_11565_));
 sg13g2_nand2_1 _22175_ (.Y(_04606_),
    .A(_11482_),
    .B(_04605_));
 sg13g2_a21oi_1 _22176_ (.A1(net118),
    .A2(_04606_),
    .Y(_04607_),
    .B1(_04603_));
 sg13g2_a21oi_1 _22177_ (.A1(_10770_),
    .A2(net96),
    .Y(_04608_),
    .B1(_04607_));
 sg13g2_or2_1 _22178_ (.X(_04609_),
    .B(_04176_),
    .A(_04170_));
 sg13g2_xor2_1 _22179_ (.B(_04609_),
    .A(_10739_),
    .X(_04610_));
 sg13g2_nand2_1 _22180_ (.Y(_04611_),
    .A(_11377_),
    .B(net112));
 sg13g2_a21oi_1 _22181_ (.A1(net162),
    .A2(net165),
    .Y(_04612_),
    .B1(_04088_));
 sg13g2_a22oi_1 _22182_ (.Y(_04613_),
    .B1(_04232_),
    .B2(net170),
    .A2(net166),
    .A1(net133));
 sg13g2_a22oi_1 _22183_ (.Y(_04614_),
    .B1(net136),
    .B2(net132),
    .A2(net169),
    .A1(_10611_));
 sg13g2_nand3_1 _22184_ (.B(_04613_),
    .C(_04614_),
    .A(_04612_),
    .Y(_04615_));
 sg13g2_nand3_1 _22185_ (.B(_04611_),
    .C(_04615_),
    .A(_09731_),
    .Y(_04616_));
 sg13g2_nor2_1 _22186_ (.A(net198),
    .B(net163),
    .Y(_04617_));
 sg13g2_mux2_1 _22187_ (.A0(_08932_),
    .A1(net1113),
    .S(_04617_),
    .X(_04618_));
 sg13g2_nand2_1 _22188_ (.Y(_04619_),
    .A(net224),
    .B(net163));
 sg13g2_o21ai_1 _22189_ (.B1(_04619_),
    .Y(_04620_),
    .A1(_09718_),
    .A2(_04618_));
 sg13g2_a21oi_1 _22190_ (.A1(net1114),
    .A2(net179),
    .Y(_04621_),
    .B1(_04097_));
 sg13g2_nand3_1 _22191_ (.B(_04620_),
    .C(_04621_),
    .A(_04616_),
    .Y(_04622_));
 sg13g2_a221oi_1 _22192_ (.B2(net1123),
    .C1(_04622_),
    .B1(_04610_),
    .A1(_04604_),
    .Y(_04623_),
    .A2(_04608_));
 sg13g2_o21ai_1 _22193_ (.B1(_04623_),
    .Y(_04624_),
    .A1(_04112_),
    .A2(_04597_));
 sg13g2_nor2b_1 _22194_ (.A(_04009_),
    .B_N(_04624_),
    .Y(_04625_));
 sg13g2_o21ai_1 _22195_ (.B1(_04625_),
    .Y(_04626_),
    .A1(_11663_),
    .A2(_04445_));
 sg13g2_nand2_1 _22196_ (.Y(_00967_),
    .A(_04596_),
    .B(_04626_));
 sg13g2_inv_1 _22197_ (.Y(_04627_),
    .A(_11682_));
 sg13g2_nor2_1 _22198_ (.A(_04627_),
    .B(_04445_),
    .Y(_04628_));
 sg13g2_o21ai_1 _22199_ (.B1(_04055_),
    .Y(_04629_),
    .A1(_11277_),
    .A2(_04201_));
 sg13g2_o21ai_1 _22200_ (.B1(_04629_),
    .Y(_04630_),
    .A1(_11652_),
    .A2(_04205_));
 sg13g2_xnor2_1 _22201_ (.Y(_04631_),
    .A(_04158_),
    .B(_04630_));
 sg13g2_o21ai_1 _22202_ (.B1(net163),
    .Y(_04632_),
    .A1(_04170_),
    .A2(_04176_));
 sg13g2_nor3_1 _22203_ (.A(net163),
    .B(_04170_),
    .C(_04176_),
    .Y(_04633_));
 sg13g2_a21oi_1 _22204_ (.A1(_11652_),
    .A2(_04632_),
    .Y(_04634_),
    .B1(_04633_));
 sg13g2_xnor2_1 _22205_ (.Y(_04635_),
    .A(_04158_),
    .B(_04634_));
 sg13g2_mux2_1 _22206_ (.A0(net1040),
    .A1(net1041),
    .S(_04196_),
    .X(_04636_));
 sg13g2_o21ai_1 _22207_ (.B1(_10801_),
    .Y(_04637_),
    .A1(net1027),
    .A2(_04636_));
 sg13g2_a21oi_1 _22208_ (.A1(net1114),
    .A2(net202),
    .Y(_04638_),
    .B1(net291));
 sg13g2_nand2_1 _22209_ (.Y(_04639_),
    .A(_04191_),
    .B(net112));
 sg13g2_a221oi_1 _22210_ (.B2(net170),
    .C1(_04079_),
    .B1(_04065_),
    .A1(net191),
    .Y(_04640_),
    .A2(net169));
 sg13g2_o21ai_1 _22211_ (.B1(_04640_),
    .Y(_04641_),
    .A1(_04028_),
    .A2(_04418_));
 sg13g2_nand3_1 _22212_ (.B(_04639_),
    .C(_04641_),
    .A(net1026),
    .Y(_04642_));
 sg13g2_nand2_1 _22213_ (.Y(_04643_),
    .A(net160),
    .B(net134));
 sg13g2_a22oi_1 _22214_ (.Y(_04644_),
    .B1(_04059_),
    .B2(_04022_),
    .A2(_04053_),
    .A1(_11157_));
 sg13g2_a21oi_1 _22215_ (.A1(_11098_),
    .A2(_04030_),
    .Y(_04645_),
    .B1(_04225_));
 sg13g2_nand4_1 _22216_ (.B(_04419_),
    .C(_04644_),
    .A(_04332_),
    .Y(_04646_),
    .D(_04645_));
 sg13g2_a21oi_1 _22217_ (.A1(net118),
    .A2(net171),
    .Y(_04647_),
    .B1(_04646_));
 sg13g2_a21oi_1 _22218_ (.A1(net1042),
    .A2(_04646_),
    .Y(_04648_),
    .B1(_09712_));
 sg13g2_a21oi_1 _22219_ (.A1(_11405_),
    .A2(_11481_),
    .Y(_04649_),
    .B1(net242));
 sg13g2_nand2b_1 _22220_ (.Y(_04650_),
    .B(_04011_),
    .A_N(_04649_));
 sg13g2_o21ai_1 _22221_ (.B1(_04650_),
    .Y(_04651_),
    .A1(_04647_),
    .A2(_04648_));
 sg13g2_nand2_1 _22222_ (.Y(_04652_),
    .A(_04643_),
    .B(_04651_));
 sg13g2_nand4_1 _22223_ (.B(_04638_),
    .C(_04642_),
    .A(_04637_),
    .Y(_04653_),
    .D(_04652_));
 sg13g2_a221oi_1 _22224_ (.B2(net1063),
    .C1(_04653_),
    .B1(_04635_),
    .A1(_04115_),
    .Y(_04654_),
    .A2(_04631_));
 sg13g2_or2_1 _22225_ (.X(_04655_),
    .B(_04654_),
    .A(net77));
 sg13g2_buf_1 _22226_ (.A(_08611_),
    .X(_04656_));
 sg13g2_xnor2_1 _22227_ (.Y(_04657_),
    .A(_10740_),
    .B(_04249_));
 sg13g2_a22oi_1 _22228_ (.Y(_04658_),
    .B1(_04657_),
    .B2(_04254_),
    .A2(_04141_),
    .A1(net956));
 sg13g2_o21ai_1 _22229_ (.B1(_04658_),
    .Y(_00968_),
    .A1(_04628_),
    .A2(_04655_));
 sg13g2_a221oi_1 _22230_ (.B2(net201),
    .C1(_04201_),
    .B1(net206),
    .A1(net167),
    .Y(_04659_),
    .A2(net223));
 sg13g2_buf_1 _22231_ (.A(_04659_),
    .X(_04660_));
 sg13g2_a21oi_1 _22232_ (.A1(_11665_),
    .A2(_04619_),
    .Y(_04661_),
    .B1(net167));
 sg13g2_a21o_1 _22233_ (.A2(net163),
    .A1(_11290_),
    .B1(_04661_),
    .X(_04662_));
 sg13g2_buf_1 _22234_ (.A(_04662_),
    .X(_04663_));
 sg13g2_o21ai_1 _22235_ (.B1(net632),
    .Y(_04664_),
    .A1(_04660_),
    .A2(_04663_));
 sg13g2_a21oi_1 _22236_ (.A1(_10770_),
    .A2(_11665_),
    .Y(_04665_),
    .B1(_04634_));
 sg13g2_a21oi_1 _22237_ (.A1(net167),
    .A2(net228),
    .Y(_04666_),
    .B1(_04665_));
 sg13g2_a221oi_1 _22238_ (.B2(_04045_),
    .C1(_04087_),
    .B1(_04053_),
    .A1(_04092_),
    .Y(_04667_),
    .A2(_04039_));
 sg13g2_a22oi_1 _22239_ (.Y(_04668_),
    .B1(_04059_),
    .B2(_10128_),
    .A2(_04030_),
    .A1(_04101_));
 sg13g2_a22oi_1 _22240_ (.Y(_04669_),
    .B1(_04064_),
    .B2(net229),
    .A2(net192),
    .A1(_10817_));
 sg13g2_nand4_1 _22241_ (.B(_04667_),
    .C(_04668_),
    .A(_04446_),
    .Y(_04670_),
    .D(_04669_));
 sg13g2_o21ai_1 _22242_ (.B1(_09731_),
    .Y(_04671_),
    .A1(_10769_),
    .A2(net164));
 sg13g2_inv_1 _22243_ (.Y(_04672_),
    .A(_04671_));
 sg13g2_o21ai_1 _22244_ (.B1(_08932_),
    .Y(_04673_),
    .A1(net205),
    .A2(_10669_));
 sg13g2_nand3_1 _22245_ (.B(_11244_),
    .C(_10678_),
    .A(net1113),
    .Y(_04674_));
 sg13g2_and2_1 _22246_ (.A(_04673_),
    .B(_04674_),
    .X(_04675_));
 sg13g2_a22oi_1 _22247_ (.Y(_04676_),
    .B1(_04675_),
    .B2(_04473_),
    .A2(net160),
    .A1(net205));
 sg13g2_a221oi_1 _22248_ (.B2(_04672_),
    .C1(_04676_),
    .B1(_04670_),
    .A1(net1114),
    .Y(_04677_),
    .A2(_11466_));
 sg13g2_a22oi_1 _22249_ (.Y(_04678_),
    .B1(_04059_),
    .B2(_11098_),
    .A2(_04030_),
    .A1(_11234_));
 sg13g2_nand4_1 _22250_ (.B(_04283_),
    .C(_04650_),
    .A(net164),
    .Y(_04679_),
    .D(_04678_));
 sg13g2_a22oi_1 _22251_ (.Y(_04680_),
    .B1(_04064_),
    .B2(_11157_),
    .A2(_04053_),
    .A1(_04022_));
 sg13g2_nand2_1 _22252_ (.Y(_04681_),
    .A(_04361_),
    .B(_04680_));
 sg13g2_a21oi_1 _22253_ (.A1(_10856_),
    .A2(net134),
    .Y(_04682_),
    .B1(net834));
 sg13g2_o21ai_1 _22254_ (.B1(_04682_),
    .Y(_04683_),
    .A1(_04679_),
    .A2(_04681_));
 sg13g2_nand3_1 _22255_ (.B(_04677_),
    .C(_04683_),
    .A(_04110_),
    .Y(_04684_));
 sg13g2_nor4_2 _22256_ (.A(_04195_),
    .B(_04202_),
    .C(_04206_),
    .Y(_04685_),
    .D(_04684_));
 sg13g2_nand2b_1 _22257_ (.Y(_04686_),
    .B(_04685_),
    .A_N(_04666_));
 sg13g2_a21oi_1 _22258_ (.A1(_04664_),
    .A2(_04686_),
    .Y(_04687_),
    .B1(_10680_));
 sg13g2_nor3_1 _22259_ (.A(_04110_),
    .B(_04660_),
    .C(_04663_),
    .Y(_04688_));
 sg13g2_a21o_1 _22260_ (.A2(_04666_),
    .A1(_04685_),
    .B1(_04688_),
    .X(_04689_));
 sg13g2_a22oi_1 _22261_ (.Y(_04690_),
    .B1(_04689_),
    .B2(_10680_),
    .A2(_04685_),
    .A1(_11533_));
 sg13g2_nand2b_1 _22262_ (.Y(_04691_),
    .B(_04690_),
    .A_N(_04687_));
 sg13g2_mux2_1 _22263_ (.A0(_11703_),
    .A1(_04691_),
    .S(_11500_),
    .X(_04692_));
 sg13g2_buf_1 _22264_ (.A(_08620_),
    .X(_04693_));
 sg13g2_nand2_1 _22265_ (.Y(_04694_),
    .A(_08611_),
    .B(_04249_));
 sg13g2_xnor2_1 _22266_ (.Y(_04695_),
    .A(_10643_),
    .B(_04694_));
 sg13g2_a22oi_1 _22267_ (.Y(_04696_),
    .B1(_04695_),
    .B2(net83),
    .A2(_04140_),
    .A1(net955));
 sg13g2_o21ai_1 _22268_ (.B1(_04696_),
    .Y(_00969_),
    .A1(net77),
    .A2(_04692_));
 sg13g2_or3_1 _22269_ (.A(_10820_),
    .B(_04660_),
    .C(_04663_),
    .X(_04697_));
 sg13g2_nand2_1 _22270_ (.Y(_04698_),
    .A(net160),
    .B(_04697_));
 sg13g2_o21ai_1 _22271_ (.B1(_10820_),
    .Y(_04699_),
    .A1(_04660_),
    .A2(_04663_));
 sg13g2_xnor2_1 _22272_ (.Y(_04700_),
    .A(_10856_),
    .B(_10878_));
 sg13g2_nor2_1 _22273_ (.A(_04110_),
    .B(_04700_),
    .Y(_04701_));
 sg13g2_and2_1 _22274_ (.A(_04699_),
    .B(_04701_),
    .X(_04702_));
 sg13g2_and3_1 _22275_ (.X(_04703_),
    .A(net160),
    .B(net632),
    .C(_04700_));
 sg13g2_nand2_1 _22276_ (.Y(_04704_),
    .A(_04270_),
    .B(_04700_));
 sg13g2_nor2_1 _22277_ (.A(_04699_),
    .B(_04704_),
    .Y(_04705_));
 sg13g2_a221oi_1 _22278_ (.B2(_04697_),
    .C1(_04705_),
    .B1(_04703_),
    .A1(_04698_),
    .Y(_04706_),
    .A2(_04702_));
 sg13g2_nor4_1 _22279_ (.A(_04270_),
    .B(_04195_),
    .C(_04202_),
    .D(_04206_),
    .Y(_04707_));
 sg13g2_inv_1 _22280_ (.Y(_04708_),
    .A(net1042));
 sg13g2_nand2b_1 _22281_ (.Y(_04709_),
    .B(_04649_),
    .A_N(net173));
 sg13g2_a22oi_1 _22282_ (.Y(_04710_),
    .B1(net189),
    .B2(_11157_),
    .A2(net165),
    .A1(net114));
 sg13g2_a22oi_1 _22283_ (.Y(_04711_),
    .B1(net166),
    .B2(_11234_),
    .A2(_04053_),
    .A1(_04072_));
 sg13g2_nand3_1 _22284_ (.B(_04710_),
    .C(_04711_),
    .A(_04324_),
    .Y(_04712_));
 sg13g2_a21oi_1 _22285_ (.A1(_11236_),
    .A2(_04709_),
    .Y(_04713_),
    .B1(_04712_));
 sg13g2_nand2_1 _22286_ (.Y(_04714_),
    .A(_09712_),
    .B(_04712_));
 sg13g2_o21ai_1 _22287_ (.B1(_04714_),
    .Y(_04715_),
    .A1(_04708_),
    .A2(_04713_));
 sg13g2_nand2_1 _22288_ (.Y(_04716_),
    .A(_04178_),
    .B(_04182_));
 sg13g2_xor2_1 _22289_ (.B(_04700_),
    .A(_04716_),
    .X(_04717_));
 sg13g2_mux2_1 _22290_ (.A0(_08932_),
    .A1(net1113),
    .S(_10879_),
    .X(_04718_));
 sg13g2_o21ai_1 _22291_ (.B1(_11036_),
    .Y(_04719_),
    .A1(_09718_),
    .A2(_04718_));
 sg13g2_a22oi_1 _22292_ (.Y(_04720_),
    .B1(net189),
    .B2(net206),
    .A2(net136),
    .A1(net229));
 sg13g2_a221oi_1 _22293_ (.B2(_04045_),
    .C1(_04087_),
    .B1(_04059_),
    .A1(_04092_),
    .Y(_04721_),
    .A2(net172));
 sg13g2_a22oi_1 _22294_ (.Y(_04722_),
    .B1(_04030_),
    .B2(_10128_),
    .A2(_04039_),
    .A1(net132));
 sg13g2_and2_1 _22295_ (.A(_04721_),
    .B(_04722_),
    .X(_04723_));
 sg13g2_nand4_1 _22296_ (.B(_04583_),
    .C(_04720_),
    .A(_04066_),
    .Y(_04724_),
    .D(_04723_));
 sg13g2_nand3_1 _22297_ (.B(_04643_),
    .C(_04724_),
    .A(_09731_),
    .Y(_04725_));
 sg13g2_nand2_1 _22298_ (.Y(_04726_),
    .A(net1114),
    .B(net244));
 sg13g2_nand3_1 _22299_ (.B(_04725_),
    .C(_04726_),
    .A(_04719_),
    .Y(_04727_));
 sg13g2_a221oi_1 _22300_ (.B2(net1123),
    .C1(_04727_),
    .B1(_04717_),
    .A1(_04238_),
    .Y(_04728_),
    .A2(_04715_));
 sg13g2_a21oi_1 _22301_ (.A1(_04707_),
    .A2(_04728_),
    .Y(_04729_),
    .B1(_04098_));
 sg13g2_a21oi_1 _22302_ (.A1(_11538_),
    .A2(_11722_),
    .Y(_04730_),
    .B1(_11500_));
 sg13g2_a21oi_1 _22303_ (.A1(_04706_),
    .A2(_04729_),
    .Y(_04731_),
    .B1(_04730_));
 sg13g2_xnor2_1 _22304_ (.Y(_04732_),
    .A(_10874_),
    .B(_04250_));
 sg13g2_a22oi_1 _22305_ (.Y(_04733_),
    .B1(_04732_),
    .B2(net95),
    .A2(_04140_),
    .A1(_08656_));
 sg13g2_o21ai_1 _22306_ (.B1(_04733_),
    .Y(_00970_),
    .A1(net77),
    .A2(_04731_));
 sg13g2_and2_1 _22307_ (.A(_04186_),
    .B(_04188_),
    .X(_04734_));
 sg13g2_xor2_1 _22308_ (.B(_04734_),
    .A(_04148_),
    .X(_04735_));
 sg13g2_nor2_1 _22309_ (.A(_04183_),
    .B(_04185_),
    .Y(_04736_));
 sg13g2_xnor2_1 _22310_ (.Y(_04737_),
    .A(_04736_),
    .B(_04734_));
 sg13g2_a22oi_1 _22311_ (.Y(_04738_),
    .B1(net189),
    .B2(_04022_),
    .A2(_04053_),
    .A1(_11234_));
 sg13g2_a22oi_1 _22312_ (.Y(_04739_),
    .B1(net165),
    .B2(_11098_),
    .A2(net192),
    .A1(_11157_));
 sg13g2_nand3_1 _22313_ (.B(_04738_),
    .C(_04739_),
    .A(net164),
    .Y(_04740_));
 sg13g2_nand3_1 _22314_ (.B(_11235_),
    .C(_04222_),
    .A(net244),
    .Y(_04741_));
 sg13g2_nand2b_1 _22315_ (.Y(_04742_),
    .B(_04741_),
    .A_N(_04740_));
 sg13g2_nor2_1 _22316_ (.A(_04381_),
    .B(_04649_),
    .Y(_04743_));
 sg13g2_a221oi_1 _22317_ (.B2(net1042),
    .C1(_04743_),
    .B1(_04742_),
    .A1(_09712_),
    .Y(_04744_),
    .A2(_04740_));
 sg13g2_a21o_1 _22318_ (.A2(net96),
    .A1(_11034_),
    .B1(_04744_),
    .X(_04745_));
 sg13g2_nand2_1 _22319_ (.Y(_04746_),
    .A(net1043),
    .B(net296));
 sg13g2_mux2_1 _22320_ (.A0(net1040),
    .A1(net1041),
    .S(_10997_),
    .X(_04747_));
 sg13g2_nand2_1 _22321_ (.Y(_04748_),
    .A(_04151_),
    .B(_11263_));
 sg13g2_o21ai_1 _22322_ (.B1(_04748_),
    .Y(_04749_),
    .A1(net1027),
    .A2(_04747_));
 sg13g2_a22oi_1 _22323_ (.Y(_04750_),
    .B1(_04065_),
    .B2(_04055_),
    .A2(net171),
    .A1(_04229_));
 sg13g2_a22oi_1 _22324_ (.Y(_04751_),
    .B1(net136),
    .B2(net191),
    .A2(net169),
    .A1(_10678_));
 sg13g2_and2_1 _22325_ (.A(_04750_),
    .B(_04751_),
    .X(_04752_));
 sg13g2_a22oi_1 _22326_ (.Y(_04753_),
    .B1(_04037_),
    .B2(_04102_),
    .A2(_04031_),
    .A1(_04046_));
 sg13g2_nand2_1 _22327_ (.Y(_04754_),
    .A(_04543_),
    .B(_04753_));
 sg13g2_a221oi_1 _22328_ (.B2(net133),
    .C1(_04754_),
    .B1(_04234_),
    .A1(_10611_),
    .Y(_04755_),
    .A2(_04060_));
 sg13g2_o21ai_1 _22329_ (.B1(net1026),
    .Y(_04756_),
    .A1(_11351_),
    .A2(_04078_));
 sg13g2_a21o_1 _22330_ (.A2(_04755_),
    .A1(_04752_),
    .B1(_04756_),
    .X(_04757_));
 sg13g2_nand4_1 _22331_ (.B(_04746_),
    .C(_04749_),
    .A(_04745_),
    .Y(_04758_),
    .D(_04757_));
 sg13g2_a221oi_1 _22332_ (.B2(net1063),
    .C1(_04758_),
    .B1(_04737_),
    .A1(net632),
    .Y(_04759_),
    .A2(_04735_));
 sg13g2_a22oi_1 _22333_ (.Y(_04760_),
    .B1(_04208_),
    .B2(_04759_),
    .A2(_04002_),
    .A1(_11747_));
 sg13g2_nand2b_1 _22334_ (.Y(_04761_),
    .B(_04760_),
    .A_N(_04143_));
 sg13g2_buf_1 _22335_ (.A(_08639_),
    .X(_04762_));
 sg13g2_xnor2_1 _22336_ (.Y(_04763_),
    .A(_00272_),
    .B(_04251_));
 sg13g2_a22oi_1 _22337_ (.Y(_04764_),
    .B1(_04763_),
    .B2(_04254_),
    .A2(net32),
    .A1(net954));
 sg13g2_nand2_1 _22338_ (.Y(_00971_),
    .A(_04761_),
    .B(_04764_));
 sg13g2_buf_1 _22339_ (.A(_00234_),
    .X(_04765_));
 sg13g2_nor4_1 _22340_ (.A(net1103),
    .B(_10021_),
    .C(_04765_),
    .D(_03635_),
    .Y(_04766_));
 sg13g2_buf_2 _22341_ (.A(_04766_),
    .X(_04767_));
 sg13g2_buf_1 _22342_ (.A(_04767_),
    .X(_04768_));
 sg13g2_mux2_1 _22343_ (.A0(_10223_),
    .A1(net502),
    .S(net493),
    .X(_00974_));
 sg13g2_mux2_1 _22344_ (.A0(_10898_),
    .A1(net836),
    .S(net493),
    .X(_00975_));
 sg13g2_mux2_1 _22345_ (.A0(_11018_),
    .A1(net496),
    .S(net493),
    .X(_00976_));
 sg13g2_mux2_1 _22346_ (.A0(_11105_),
    .A1(net447),
    .S(_04768_),
    .X(_00977_));
 sg13g2_buf_1 _22347_ (.A(net639),
    .X(_04769_));
 sg13g2_mux2_1 _22348_ (.A0(_11052_),
    .A1(_04769_),
    .S(net493),
    .X(_00978_));
 sg13g2_mux2_1 _22349_ (.A0(_11191_),
    .A1(net635),
    .S(net493),
    .X(_00979_));
 sg13g2_mux2_1 _22350_ (.A0(_10093_),
    .A1(net359),
    .S(net493),
    .X(_00980_));
 sg13g2_mux2_1 _22351_ (.A0(_10359_),
    .A1(net409),
    .S(_04768_),
    .X(_00981_));
 sg13g2_mux2_1 _22352_ (.A0(_10558_),
    .A1(net408),
    .S(net493),
    .X(_00982_));
 sg13g2_mux2_1 _22353_ (.A0(_10485_),
    .A1(net570),
    .S(net493),
    .X(_00983_));
 sg13g2_mux2_1 _22354_ (.A0(_10695_),
    .A1(net711),
    .S(_04767_),
    .X(_00984_));
 sg13g2_mux2_1 _22355_ (.A0(_10755_),
    .A1(_03134_),
    .S(_04767_),
    .X(_00985_));
 sg13g2_buf_1 _22356_ (.A(net1037),
    .X(_04770_));
 sg13g2_mux2_1 _22357_ (.A0(_10631_),
    .A1(_04770_),
    .S(_04767_),
    .X(_00986_));
 sg13g2_buf_1 _22358_ (.A(_10831_),
    .X(_04771_));
 sg13g2_mux2_1 _22359_ (.A0(_10839_),
    .A1(_04771_),
    .S(_04767_),
    .X(_00987_));
 sg13g2_mux2_1 _22360_ (.A0(_10957_),
    .A1(_03137_),
    .S(_04767_),
    .X(_00988_));
 sg13g2_or2_1 _22361_ (.X(_04772_),
    .B(_03635_),
    .A(_10022_));
 sg13g2_buf_1 _22362_ (.A(_04772_),
    .X(_04773_));
 sg13g2_buf_1 _22363_ (.A(_04773_),
    .X(_04774_));
 sg13g2_nor2_1 _22364_ (.A(_08397_),
    .B(_04765_),
    .Y(_04775_));
 sg13g2_nand2_1 _22365_ (.Y(_04776_),
    .A(_03633_),
    .B(_04775_));
 sg13g2_nor2_1 _22366_ (.A(_08397_),
    .B(_03636_),
    .Y(_04777_));
 sg13g2_a21oi_1 _22367_ (.A1(_03636_),
    .A2(\cpu.ex.r_wb_swapsp ),
    .Y(_04778_),
    .B1(_04777_));
 sg13g2_or4_1 _22368_ (.A(net1103),
    .B(_04765_),
    .C(_03635_),
    .D(_04778_),
    .X(_04779_));
 sg13g2_buf_1 _22369_ (.A(_04779_),
    .X(_04780_));
 sg13g2_buf_1 _22370_ (.A(_04780_),
    .X(_04781_));
 sg13g2_nand2_1 _22371_ (.Y(_04782_),
    .A(\cpu.ex.r_stmp[0] ),
    .B(_04781_));
 sg13g2_o21ai_1 _22372_ (.B1(_04782_),
    .Y(_00989_),
    .A1(net492),
    .A2(_04776_));
 sg13g2_mux2_1 _22373_ (.A0(net1095),
    .A1(_10957_),
    .S(net492),
    .X(_04783_));
 sg13g2_buf_1 _22374_ (.A(_04780_),
    .X(_04784_));
 sg13g2_mux2_1 _22375_ (.A0(_04783_),
    .A1(\cpu.ex.r_stmp[10] ),
    .S(_04784_),
    .X(_00990_));
 sg13g2_mux2_1 _22376_ (.A0(_10907_),
    .A1(_10898_),
    .S(net492),
    .X(_04785_));
 sg13g2_mux2_1 _22377_ (.A0(_04785_),
    .A1(\cpu.ex.r_stmp[11] ),
    .S(net406),
    .X(_00991_));
 sg13g2_mux2_1 _22378_ (.A0(net589),
    .A1(_11018_),
    .S(_04774_),
    .X(_04786_));
 sg13g2_mux2_1 _22379_ (.A0(_04786_),
    .A1(\cpu.ex.r_stmp[12] ),
    .S(net406),
    .X(_00992_));
 sg13g2_mux2_1 _22380_ (.A0(_09483_),
    .A1(_11105_),
    .S(net492),
    .X(_04787_));
 sg13g2_mux2_1 _22381_ (.A0(_04787_),
    .A1(\cpu.ex.r_stmp[13] ),
    .S(net406),
    .X(_00993_));
 sg13g2_buf_1 _22382_ (.A(_04773_),
    .X(_04788_));
 sg13g2_mux2_1 _22383_ (.A0(_11042_),
    .A1(_11052_),
    .S(net491),
    .X(_04789_));
 sg13g2_mux2_1 _22384_ (.A0(_04789_),
    .A1(\cpu.ex.r_stmp[14] ),
    .S(net406),
    .X(_00994_));
 sg13g2_mux2_1 _22385_ (.A0(net731),
    .A1(_11191_),
    .S(_04788_),
    .X(_04790_));
 sg13g2_mux2_1 _22386_ (.A0(_04790_),
    .A1(\cpu.ex.r_stmp[15] ),
    .S(net407),
    .X(_00995_));
 sg13g2_nor2_1 _22387_ (.A(net673),
    .B(net491),
    .Y(_04791_));
 sg13g2_a21oi_1 _22388_ (.A1(_10223_),
    .A2(net492),
    .Y(_04792_),
    .B1(_04791_));
 sg13g2_nand2_1 _22389_ (.Y(_04793_),
    .A(\cpu.ex.r_stmp[1] ),
    .B(net407));
 sg13g2_o21ai_1 _22390_ (.B1(_04793_),
    .Y(_00996_),
    .A1(net406),
    .A2(_04792_));
 sg13g2_nor2_1 _22391_ (.A(_11988_),
    .B(_04788_),
    .Y(_04794_));
 sg13g2_a21oi_1 _22392_ (.A1(_10093_),
    .A2(net492),
    .Y(_04795_),
    .B1(_04794_));
 sg13g2_nand2_1 _22393_ (.Y(_04796_),
    .A(\cpu.ex.r_stmp[2] ),
    .B(net407));
 sg13g2_o21ai_1 _22394_ (.B1(_04796_),
    .Y(_00997_),
    .A1(net406),
    .A2(_04795_));
 sg13g2_nor2_1 _22395_ (.A(_09052_),
    .B(net491),
    .Y(_04797_));
 sg13g2_a21oi_1 _22396_ (.A1(_10359_),
    .A2(_04774_),
    .Y(_04798_),
    .B1(_04797_));
 sg13g2_nand2_1 _22397_ (.Y(_04799_),
    .A(\cpu.ex.r_stmp[3] ),
    .B(_04781_));
 sg13g2_o21ai_1 _22398_ (.B1(_04799_),
    .Y(_00998_),
    .A1(_04784_),
    .A2(_04798_));
 sg13g2_nor2_1 _22399_ (.A(net566),
    .B(net491),
    .Y(_04800_));
 sg13g2_a21oi_1 _22400_ (.A1(_10558_),
    .A2(net492),
    .Y(_04801_),
    .B1(_04800_));
 sg13g2_nand2_1 _22401_ (.Y(_04802_),
    .A(\cpu.ex.r_stmp[4] ),
    .B(net407));
 sg13g2_o21ai_1 _22402_ (.B1(_04802_),
    .Y(_00999_),
    .A1(net406),
    .A2(_04801_));
 sg13g2_nor2_1 _22403_ (.A(net718),
    .B(_04773_),
    .Y(_04803_));
 sg13g2_a21oi_1 _22404_ (.A1(_10485_),
    .A2(net492),
    .Y(_04804_),
    .B1(_04803_));
 sg13g2_nand2_1 _22405_ (.Y(_04805_),
    .A(\cpu.ex.r_stmp[5] ),
    .B(_04780_));
 sg13g2_o21ai_1 _22406_ (.B1(_04805_),
    .Y(_01000_),
    .A1(net406),
    .A2(_04804_));
 sg13g2_mux2_1 _22407_ (.A0(_03093_),
    .A1(_10695_),
    .S(net491),
    .X(_04806_));
 sg13g2_mux2_1 _22408_ (.A0(_04806_),
    .A1(\cpu.ex.r_stmp[6] ),
    .S(net407),
    .X(_01001_));
 sg13g2_mux2_1 _22409_ (.A0(net965),
    .A1(_10755_),
    .S(net491),
    .X(_04807_));
 sg13g2_mux2_1 _22410_ (.A0(_04807_),
    .A1(\cpu.ex.r_stmp[7] ),
    .S(net407),
    .X(_01002_));
 sg13g2_mux2_1 _22411_ (.A0(net1037),
    .A1(_10631_),
    .S(net491),
    .X(_04808_));
 sg13g2_mux2_1 _22412_ (.A0(_04808_),
    .A1(\cpu.ex.r_stmp[8] ),
    .S(net407),
    .X(_01003_));
 sg13g2_mux2_1 _22413_ (.A0(_10831_),
    .A1(_10839_),
    .S(net491),
    .X(_04809_));
 sg13g2_mux2_1 _22414_ (.A0(_04809_),
    .A1(\cpu.ex.r_stmp[9] ),
    .S(net407),
    .X(_01004_));
 sg13g2_buf_1 _22415_ (.A(_11515_),
    .X(_04810_));
 sg13g2_a21oi_1 _22416_ (.A1(_11503_),
    .A2(_11504_),
    .Y(_04811_),
    .B1(_11505_));
 sg13g2_nor2_1 _22417_ (.A(net373),
    .B(_04811_),
    .Y(_04812_));
 sg13g2_nand2_1 _22418_ (.Y(_04813_),
    .A(net191),
    .B(net136));
 sg13g2_o21ai_1 _22419_ (.B1(_04813_),
    .Y(_04814_),
    .A1(_04074_),
    .A2(_04223_));
 sg13g2_a221oi_1 _22420_ (.B2(_10967_),
    .C1(_04814_),
    .B1(_04234_),
    .A1(net168),
    .Y(_04815_),
    .A2(net166));
 sg13g2_a22oi_1 _22421_ (.Y(_04816_),
    .B1(net189),
    .B2(net170),
    .A2(net169),
    .A1(_04229_));
 sg13g2_nand2b_1 _22422_ (.Y(_04817_),
    .B(_04011_),
    .A_N(_11482_));
 sg13g2_and4_1 _22423_ (.A(_04366_),
    .B(_04815_),
    .C(_04816_),
    .D(_04817_),
    .X(_04818_));
 sg13g2_mux4_1 _22424_ (.S0(_11543_),
    .A0(_04068_),
    .A1(_04072_),
    .A2(_04023_),
    .A3(_11236_),
    .S1(net245),
    .X(_04819_));
 sg13g2_a21oi_1 _22425_ (.A1(_11543_),
    .A2(net137),
    .Y(_04820_),
    .B1(_04546_));
 sg13g2_o21ai_1 _22426_ (.B1(_04017_),
    .Y(_04821_),
    .A1(_11467_),
    .A2(_04499_));
 sg13g2_a21oi_1 _22427_ (.A1(_11467_),
    .A2(_04820_),
    .Y(_04822_),
    .B1(_04821_));
 sg13g2_a21oi_1 _22428_ (.A1(_04019_),
    .A2(_04819_),
    .Y(_04823_),
    .B1(_04822_));
 sg13g2_a221oi_1 _22429_ (.B2(_04823_),
    .C1(_04083_),
    .B1(_04818_),
    .A1(_11383_),
    .Y(_04824_),
    .A2(net96));
 sg13g2_and2_1 _22430_ (.A(_04107_),
    .B(_04112_),
    .X(_04825_));
 sg13g2_nor3_1 _22431_ (.A(net1113),
    .B(net293),
    .C(net200),
    .Y(_04826_));
 sg13g2_a21oi_1 _22432_ (.A1(net200),
    .A2(_04825_),
    .Y(_04827_),
    .B1(_04826_));
 sg13g2_or2_1 _22433_ (.X(_04828_),
    .B(_04827_),
    .A(net1027));
 sg13g2_nor2b_1 _22434_ (.A(_09719_),
    .B_N(_04825_),
    .Y(_04829_));
 sg13g2_o21ai_1 _22435_ (.B1(_03721_),
    .Y(_04830_),
    .A1(net200),
    .A2(_04829_));
 sg13g2_a221oi_1 _22436_ (.B2(_04830_),
    .C1(_04098_),
    .B1(_04828_),
    .A1(_08882_),
    .Y(_04831_),
    .A2(_11244_));
 sg13g2_nor2b_1 _22437_ (.A(_04824_),
    .B_N(_04831_),
    .Y(_04832_));
 sg13g2_nor2_1 _22438_ (.A(net961),
    .B(_04812_),
    .Y(_04833_));
 sg13g2_a21oi_1 _22439_ (.A1(_04812_),
    .A2(_04832_),
    .Y(_04834_),
    .B1(_04833_));
 sg13g2_nand2_1 _22440_ (.Y(_04835_),
    .A(net111),
    .B(_04834_));
 sg13g2_a22oi_1 _22441_ (.Y(_04836_),
    .B1(net681),
    .B2(\cpu.dcache.r_data[3][16] ),
    .A2(net675),
    .A1(\cpu.dcache.r_data[7][16] ));
 sg13g2_a22oi_1 _22442_ (.Y(_04837_),
    .B1(net580),
    .B2(\cpu.dcache.r_data[6][16] ),
    .A2(net581),
    .A1(\cpu.dcache.r_data[5][16] ));
 sg13g2_a22oi_1 _22443_ (.Y(_04838_),
    .B1(net604),
    .B2(\cpu.dcache.r_data[4][16] ),
    .A2(net602),
    .A1(\cpu.dcache.r_data[2][16] ));
 sg13g2_nand3_1 _22444_ (.B(_04837_),
    .C(_04838_),
    .A(_04836_),
    .Y(_04839_));
 sg13g2_nand2b_1 _22445_ (.Y(_04840_),
    .B(net758),
    .A_N(\cpu.dcache.r_data[0][16] ));
 sg13g2_o21ai_1 _22446_ (.B1(_04840_),
    .Y(_04841_),
    .A1(net758),
    .A2(_04839_));
 sg13g2_o21ai_1 _22447_ (.B1(net455),
    .Y(_04842_),
    .A1(\cpu.dcache.r_data[1][16] ),
    .A2(_04839_));
 sg13g2_o21ai_1 _22448_ (.B1(_04842_),
    .Y(_04843_),
    .A1(net413),
    .A2(_04841_));
 sg13g2_inv_2 _22449_ (.Y(_04844_),
    .A(_11984_));
 sg13g2_nand2_1 _22450_ (.Y(_04845_),
    .A(net1122),
    .B(net896));
 sg13g2_a21o_1 _22451_ (.A2(net1038),
    .A1(_08190_),
    .B1(_04845_),
    .X(_04846_));
 sg13g2_buf_2 _22452_ (.A(_04846_),
    .X(_04847_));
 sg13g2_nor3_1 _22453_ (.A(net1038),
    .B(net1119),
    .C(_04845_),
    .Y(_04848_));
 sg13g2_buf_1 _22454_ (.A(_04848_),
    .X(_04849_));
 sg13g2_a21oi_1 _22455_ (.A1(_04844_),
    .A2(_04847_),
    .Y(_04850_),
    .B1(net564));
 sg13g2_a21oi_1 _22456_ (.A1(net637),
    .A2(_04843_),
    .Y(_04851_),
    .B1(_04850_));
 sg13g2_buf_1 _22457_ (.A(net754),
    .X(_04852_));
 sg13g2_mux2_1 _22458_ (.A0(\cpu.dcache.r_data[5][8] ),
    .A1(\cpu.dcache.r_data[7][8] ),
    .S(net608),
    .X(_04853_));
 sg13g2_a22oi_1 _22459_ (.Y(_04854_),
    .B1(_04853_),
    .B2(_12460_),
    .A2(_09426_),
    .A1(\cpu.dcache.r_data[4][8] ));
 sg13g2_buf_1 _22460_ (.A(_09464_),
    .X(_04855_));
 sg13g2_a22oi_1 _22461_ (.Y(_04856_),
    .B1(net580),
    .B2(\cpu.dcache.r_data[6][8] ),
    .A2(net681),
    .A1(\cpu.dcache.r_data[3][8] ));
 sg13g2_o21ai_1 _22462_ (.B1(_04856_),
    .Y(_04857_),
    .A1(_00279_),
    .A2(net490));
 sg13g2_a221oi_1 _22463_ (.B2(\cpu.dcache.r_data[2][8] ),
    .C1(_04857_),
    .B1(net512),
    .A1(\cpu.dcache.r_data[1][8] ),
    .Y(_04858_),
    .A2(_03068_));
 sg13g2_o21ai_1 _22464_ (.B1(_04858_),
    .Y(_04859_),
    .A1(_09174_),
    .A2(_04854_));
 sg13g2_inv_1 _22465_ (.Y(_04860_),
    .A(_00278_));
 sg13g2_a22oi_1 _22466_ (.Y(_04861_),
    .B1(_09447_),
    .B2(_04860_),
    .A2(net510),
    .A1(\cpu.dcache.r_data[5][24] ));
 sg13g2_buf_1 _22467_ (.A(net580),
    .X(_04862_));
 sg13g2_a22oi_1 _22468_ (.Y(_04863_),
    .B1(net489),
    .B2(\cpu.dcache.r_data[6][24] ),
    .A2(net513),
    .A1(\cpu.dcache.r_data[1][24] ));
 sg13g2_a22oi_1 _22469_ (.Y(_04864_),
    .B1(net529),
    .B2(\cpu.dcache.r_data[4][24] ),
    .A2(net512),
    .A1(\cpu.dcache.r_data[2][24] ));
 sg13g2_a22oi_1 _22470_ (.Y(_04865_),
    .B1(net582),
    .B2(\cpu.dcache.r_data[3][24] ),
    .A2(net599),
    .A1(\cpu.dcache.r_data[7][24] ));
 sg13g2_nand4_1 _22471_ (.B(_04863_),
    .C(_04864_),
    .A(_04861_),
    .Y(_04866_),
    .D(_04865_));
 sg13g2_a221oi_1 _22472_ (.B2(_04844_),
    .C1(_04847_),
    .B1(_04866_),
    .A1(_04852_),
    .Y(_04867_),
    .A2(_04859_));
 sg13g2_mux2_1 _22473_ (.A0(\cpu.dcache.r_data[1][0] ),
    .A1(\cpu.dcache.r_data[3][0] ),
    .S(net608),
    .X(_04868_));
 sg13g2_a22oi_1 _22474_ (.Y(_04869_),
    .B1(_04868_),
    .B2(net517),
    .A2(net680),
    .A1(\cpu.dcache.r_data[2][0] ));
 sg13g2_inv_1 _22475_ (.Y(_04870_),
    .A(_04869_));
 sg13g2_mux4_1 _22476_ (.S0(net517),
    .A0(\cpu.dcache.r_data[4][0] ),
    .A1(\cpu.dcache.r_data[5][0] ),
    .A2(\cpu.dcache.r_data[6][0] ),
    .A3(\cpu.dcache.r_data[7][0] ),
    .S1(net532),
    .X(_04871_));
 sg13g2_a22oi_1 _22477_ (.Y(_04872_),
    .B1(_04871_),
    .B2(_11939_),
    .A2(_04870_),
    .A1(net1028));
 sg13g2_nor2_1 _22478_ (.A(\cpu.dcache.r_data[0][0] ),
    .B(net490),
    .Y(_04873_));
 sg13g2_a21oi_1 _22479_ (.A1(net490),
    .A2(_04872_),
    .Y(_04874_),
    .B1(_04873_));
 sg13g2_nand2_1 _22480_ (.Y(_04875_),
    .A(_11984_),
    .B(_04847_));
 sg13g2_nor2_1 _22481_ (.A(_04874_),
    .B(_04875_),
    .Y(_04876_));
 sg13g2_nor3_1 _22482_ (.A(_04851_),
    .B(_04867_),
    .C(_04876_),
    .Y(_04877_));
 sg13g2_nand2_1 _22483_ (.Y(_04878_),
    .A(net673),
    .B(_04874_));
 sg13g2_or3_1 _22484_ (.A(net1038),
    .B(net1119),
    .C(_04845_),
    .X(_04879_));
 sg13g2_buf_1 _22485_ (.A(_04879_),
    .X(_04880_));
 sg13g2_a21oi_1 _22486_ (.A1(_04851_),
    .A2(_04878_),
    .Y(_04881_),
    .B1(_04880_));
 sg13g2_nor3_1 _22487_ (.A(net967),
    .B(_04877_),
    .C(_04881_),
    .Y(_04882_));
 sg13g2_nand2b_1 _22488_ (.Y(_04883_),
    .B(net674),
    .A_N(_09028_));
 sg13g2_buf_2 _22489_ (.A(_04883_),
    .X(_04884_));
 sg13g2_o21ai_1 _22490_ (.B1(net777),
    .Y(_04885_),
    .A1(_09297_),
    .A2(_09367_));
 sg13g2_buf_2 _22491_ (.A(_04885_),
    .X(_04886_));
 sg13g2_nor2_1 _22492_ (.A(net763),
    .B(_09051_),
    .Y(_04887_));
 sg13g2_and2_1 _22493_ (.A(_09039_),
    .B(_04887_),
    .X(_04888_));
 sg13g2_buf_1 _22494_ (.A(_04888_),
    .X(_04889_));
 sg13g2_buf_1 _22495_ (.A(net405),
    .X(_04890_));
 sg13g2_nand2_2 _22496_ (.Y(_04891_),
    .A(net609),
    .B(net1111));
 sg13g2_nor2_1 _22497_ (.A(net676),
    .B(_04891_),
    .Y(_04892_));
 sg13g2_buf_1 _22498_ (.A(_04892_),
    .X(_04893_));
 sg13g2_a22oi_1 _22499_ (.Y(_04894_),
    .B1(net404),
    .B2(\cpu.uart.r_x_invert ),
    .A2(net357),
    .A1(\cpu.uart.r_div_value[0] ));
 sg13g2_nand2_1 _22500_ (.Y(_04895_),
    .A(net609),
    .B(_09872_));
 sg13g2_buf_2 _22501_ (.A(_04895_),
    .X(_04896_));
 sg13g2_nor2_1 _22502_ (.A(net676),
    .B(_04896_),
    .Y(_04897_));
 sg13g2_buf_1 _22503_ (.A(_04897_),
    .X(_04898_));
 sg13g2_nand2_1 _22504_ (.Y(_04899_),
    .A(net777),
    .B(net608));
 sg13g2_nor2_1 _22505_ (.A(net598),
    .B(_04899_),
    .Y(_04900_));
 sg13g2_buf_1 _22506_ (.A(_04900_),
    .X(_04901_));
 sg13g2_buf_1 _22507_ (.A(_04901_),
    .X(_04902_));
 sg13g2_a22oi_1 _22508_ (.Y(_04903_),
    .B1(net355),
    .B2(\cpu.uart.r_div_value[8] ),
    .A2(_04898_),
    .A1(_08972_));
 sg13g2_nand2_1 _22509_ (.Y(_04904_),
    .A(_04894_),
    .B(_04903_));
 sg13g2_a21oi_1 _22510_ (.A1(\cpu.uart.r_in[0] ),
    .A2(_04886_),
    .Y(_04905_),
    .B1(_04904_));
 sg13g2_o21ai_1 _22511_ (.B1(net967),
    .Y(_04906_),
    .A1(_04884_),
    .A2(_04905_));
 sg13g2_nand2_1 _22512_ (.Y(_04907_),
    .A(_09872_),
    .B(net677));
 sg13g2_buf_2 _22513_ (.A(_04907_),
    .X(_04908_));
 sg13g2_nor2_1 _22514_ (.A(net1025),
    .B(_09616_),
    .Y(_04909_));
 sg13g2_buf_1 _22515_ (.A(_04909_),
    .X(_04910_));
 sg13g2_a22oi_1 _22516_ (.Y(_04911_),
    .B1(_04910_),
    .B2(\cpu.intr.r_timer_reload[0] ),
    .A2(net528),
    .A1(_09930_));
 sg13g2_o21ai_1 _22517_ (.B1(_04911_),
    .Y(_04912_),
    .A1(_00264_),
    .A2(_04908_));
 sg13g2_nand2_1 _22518_ (.Y(_04913_),
    .A(net881),
    .B(net646));
 sg13g2_mux2_1 _22519_ (.A0(\cpu.intr.r_clock_cmp[16] ),
    .A1(\cpu.intr.r_timer_reload[16] ),
    .S(net464),
    .X(_04914_));
 sg13g2_a22oi_1 _22520_ (.Y(_04915_),
    .B1(_04914_),
    .B2(net456),
    .A2(net680),
    .A1(_09792_));
 sg13g2_buf_1 _22521_ (.A(\cpu.intr.r_clock_count[16] ),
    .X(_04916_));
 sg13g2_nor2_1 _22522_ (.A(net1025),
    .B(_02697_),
    .Y(_04917_));
 sg13g2_buf_2 _22523_ (.A(_04917_),
    .X(_04918_));
 sg13g2_nor2_1 _22524_ (.A(_08972_),
    .B(_08973_),
    .Y(_04919_));
 sg13g2_nor3_1 _22525_ (.A(_04919_),
    .B(net676),
    .C(net598),
    .Y(_04920_));
 sg13g2_a221oi_1 _22526_ (.B2(\cpu.intr.r_clock_cmp[0] ),
    .C1(_04920_),
    .B1(_04918_),
    .A1(_04916_),
    .Y(_04921_),
    .A2(net461));
 sg13g2_o21ai_1 _22527_ (.B1(_04921_),
    .Y(_04922_),
    .A1(_04913_),
    .A2(_04915_));
 sg13g2_nor2_1 _22528_ (.A(_04912_),
    .B(_04922_),
    .Y(_04923_));
 sg13g2_buf_1 _22529_ (.A(net356),
    .X(_04924_));
 sg13g2_and2_1 _22530_ (.A(net598),
    .B(_04896_),
    .X(_04925_));
 sg13g2_nor2_1 _22531_ (.A(net608),
    .B(_04925_),
    .Y(_04926_));
 sg13g2_nor3_1 _22532_ (.A(net646),
    .B(_04919_),
    .C(_04926_),
    .Y(_04927_));
 sg13g2_o21ai_1 _22533_ (.B1(\cpu.intr.r_enable[0] ),
    .Y(_04928_),
    .A1(net289),
    .A2(_04927_));
 sg13g2_a21oi_1 _22534_ (.A1(_04923_),
    .A2(_04928_),
    .Y(_04929_),
    .B1(net674));
 sg13g2_nand2_1 _22535_ (.Y(_04930_),
    .A(net763),
    .B(net883));
 sg13g2_a21oi_1 _22536_ (.A1(net685),
    .A2(_04930_),
    .Y(_04931_),
    .B1(net609));
 sg13g2_inv_1 _22537_ (.Y(_04932_),
    .A(_09031_));
 sg13g2_nand2_1 _22538_ (.Y(_04933_),
    .A(net777),
    .B(_09542_));
 sg13g2_nor2_1 _22539_ (.A(_09037_),
    .B(_04933_),
    .Y(_04934_));
 sg13g2_a21oi_1 _22540_ (.A1(_09051_),
    .A2(_04932_),
    .Y(_04935_),
    .B1(_04934_));
 sg13g2_nor3_1 _22541_ (.A(net1111),
    .B(_09261_),
    .C(_09379_),
    .Y(_04936_));
 sg13g2_a21oi_1 _22542_ (.A1(net1111),
    .A2(_04935_),
    .Y(_04937_),
    .B1(_04936_));
 sg13g2_nor2_1 _22543_ (.A(_04931_),
    .B(_04937_),
    .Y(_04938_));
 sg13g2_nand2b_1 _22544_ (.Y(_04939_),
    .B(_04887_),
    .A_N(net598));
 sg13g2_buf_1 _22545_ (.A(_04939_),
    .X(_04940_));
 sg13g2_a21oi_1 _22546_ (.A1(_04940_),
    .A2(_04908_),
    .Y(_04941_),
    .B1(_09781_));
 sg13g2_nor2_1 _22547_ (.A(_04938_),
    .B(_04941_),
    .Y(_04942_));
 sg13g2_buf_2 _22548_ (.A(_04942_),
    .X(_04943_));
 sg13g2_a22oi_1 _22549_ (.Y(_04944_),
    .B1(\cpu.spi.r_timeout[0] ),
    .B2(net464),
    .A2(_09031_),
    .A1(_08976_));
 sg13g2_nand3_1 _22550_ (.B(net781),
    .C(\cpu.spi.r_ready ),
    .A(net754),
    .Y(_04945_));
 sg13g2_o21ai_1 _22551_ (.B1(_04945_),
    .Y(_04946_),
    .A1(net754),
    .A2(_04944_));
 sg13g2_nor2_1 _22552_ (.A(net1111),
    .B(_09340_),
    .Y(_04947_));
 sg13g2_buf_2 _22553_ (.A(_04947_),
    .X(_04948_));
 sg13g2_nand2b_1 _22554_ (.Y(_04949_),
    .B(net405),
    .A_N(_00203_));
 sg13g2_o21ai_1 _22555_ (.B1(_04949_),
    .Y(_04950_),
    .A1(_00281_),
    .A2(_04940_));
 sg13g2_a21oi_1 _22556_ (.A1(\cpu.spi.r_mode[1][0] ),
    .A2(_04948_),
    .Y(_04951_),
    .B1(_04950_));
 sg13g2_and2_1 _22557_ (.A(net994),
    .B(net405),
    .X(_04952_));
 sg13g2_buf_1 _22558_ (.A(_04952_),
    .X(_04953_));
 sg13g2_buf_1 _22559_ (.A(_09542_),
    .X(_04954_));
 sg13g2_nor2_1 _22560_ (.A(_04954_),
    .B(_04940_),
    .Y(_04955_));
 sg13g2_buf_2 _22561_ (.A(_04955_),
    .X(_04956_));
 sg13g2_buf_1 _22562_ (.A(\cpu.spi.r_clk_count[2][0] ),
    .X(_04957_));
 sg13g2_nand3_1 _22563_ (.B(_09542_),
    .C(net677),
    .A(net1111),
    .Y(_04958_));
 sg13g2_buf_2 _22564_ (.A(_04958_),
    .X(_04959_));
 sg13g2_nor2_1 _22565_ (.A(_00280_),
    .B(_04959_),
    .Y(_04960_));
 sg13g2_a221oi_1 _22566_ (.B2(_04957_),
    .C1(_04960_),
    .B1(_04956_),
    .A1(\cpu.spi.r_mode[2][0] ),
    .Y(_04961_),
    .A2(_04953_));
 sg13g2_o21ai_1 _22567_ (.B1(_04961_),
    .Y(_04962_),
    .A1(net857),
    .A2(_04951_));
 sg13g2_a221oi_1 _22568_ (.B2(net456),
    .C1(_04962_),
    .B1(_04946_),
    .A1(_09073_),
    .Y(_04963_),
    .A2(_04943_));
 sg13g2_nor2_1 _22569_ (.A(_09030_),
    .B(_04963_),
    .Y(_04964_));
 sg13g2_buf_2 _22570_ (.A(\cpu.gpio.r_spi_miso_src[0][0] ),
    .X(_04965_));
 sg13g2_nor3_2 _22571_ (.A(net879),
    .B(net883),
    .C(_02697_),
    .Y(_04966_));
 sg13g2_buf_2 _22572_ (.A(\cpu.gpio.r_uart_rx_src[0] ),
    .X(_04967_));
 sg13g2_inv_1 _22573_ (.Y(_04968_),
    .A(_04967_));
 sg13g2_a22oi_1 _22574_ (.Y(_04969_),
    .B1(net356),
    .B2(_08991_),
    .A2(_04889_),
    .A1(_08990_));
 sg13g2_o21ai_1 _22575_ (.B1(_04969_),
    .Y(_04970_),
    .A1(_04968_),
    .A2(_04908_));
 sg13g2_buf_2 _22576_ (.A(\cpu.gpio.r_src_io[4][0] ),
    .X(_04971_));
 sg13g2_nor3_1 _22577_ (.A(_09542_),
    .B(_04899_),
    .C(_04896_),
    .Y(_04972_));
 sg13g2_buf_1 _22578_ (.A(_04972_),
    .X(_04973_));
 sg13g2_nor3_2 _22579_ (.A(net952),
    .B(_04899_),
    .C(_04891_),
    .Y(_04974_));
 sg13g2_buf_2 _22580_ (.A(\cpu.gpio.r_src_io[6][0] ),
    .X(_04975_));
 sg13g2_a22oi_1 _22581_ (.Y(_04976_),
    .B1(_04974_),
    .B2(_04975_),
    .A2(net354),
    .A1(_04971_));
 sg13g2_buf_2 _22582_ (.A(\cpu.gpio.r_src_o[6][0] ),
    .X(_04977_));
 sg13g2_nand2_1 _22583_ (.Y(_04978_),
    .A(net994),
    .B(_04892_));
 sg13g2_buf_1 _22584_ (.A(_04978_),
    .X(_04979_));
 sg13g2_inv_1 _22585_ (.Y(_04980_),
    .A(_04979_));
 sg13g2_nor3_2 _22586_ (.A(net952),
    .B(net676),
    .C(_04896_),
    .Y(_04981_));
 sg13g2_buf_2 _22587_ (.A(\cpu.gpio.r_src_o[4][0] ),
    .X(_04982_));
 sg13g2_a22oi_1 _22588_ (.Y(_04983_),
    .B1(_04981_),
    .B2(_04982_),
    .A2(_04980_),
    .A1(_04977_));
 sg13g2_nand2_1 _22589_ (.Y(_04984_),
    .A(_04976_),
    .B(_04983_));
 sg13g2_a221oi_1 _22590_ (.B2(net848),
    .C1(_04984_),
    .B1(_04970_),
    .A1(_04965_),
    .Y(_04985_),
    .A2(_04966_));
 sg13g2_o21ai_1 _22591_ (.B1(_09542_),
    .Y(_04986_),
    .A1(net1111),
    .A2(net763));
 sg13g2_nor2_1 _22592_ (.A(_09781_),
    .B(net685),
    .Y(_04987_));
 sg13g2_nor2_1 _22593_ (.A(_10473_),
    .B(net781),
    .Y(_04988_));
 sg13g2_a21oi_1 _22594_ (.A1(_04986_),
    .A2(_04987_),
    .Y(_04989_),
    .B1(_04988_));
 sg13g2_o21ai_1 _22595_ (.B1(_04930_),
    .Y(_04990_),
    .A1(net781),
    .A2(net883));
 sg13g2_o21ai_1 _22596_ (.B1(_04930_),
    .Y(_04991_),
    .A1(_04896_),
    .A2(_04933_));
 sg13g2_a22oi_1 _22597_ (.Y(_04992_),
    .B1(net883),
    .B2(_04987_),
    .A2(net685),
    .A1(net763));
 sg13g2_nor2_1 _22598_ (.A(net879),
    .B(_04992_),
    .Y(_04993_));
 sg13g2_a221oi_1 _22599_ (.B2(_09781_),
    .C1(_04993_),
    .B1(_04991_),
    .A1(_09037_),
    .Y(_04994_),
    .A2(_04990_));
 sg13g2_o21ai_1 _22600_ (.B1(_04994_),
    .Y(_04995_),
    .A1(net609),
    .A2(_04989_));
 sg13g2_buf_2 _22601_ (.A(_04995_),
    .X(_04996_));
 sg13g2_nand3_1 _22602_ (.B(_08991_),
    .C(_04996_),
    .A(_08990_),
    .Y(_04997_));
 sg13g2_nand2b_1 _22603_ (.Y(_04998_),
    .B(_09028_),
    .A_N(net966));
 sg13g2_buf_1 _22604_ (.A(_04998_),
    .X(_04999_));
 sg13g2_a21oi_1 _22605_ (.A1(_04985_),
    .A2(_04997_),
    .Y(_05000_),
    .B1(_04999_));
 sg13g2_nor4_1 _22606_ (.A(_04906_),
    .B(_04929_),
    .C(_04964_),
    .D(_05000_),
    .Y(_05001_));
 sg13g2_nand2_1 _22607_ (.Y(_05002_),
    .A(net1122),
    .B(_11528_));
 sg13g2_buf_2 _22608_ (.A(_05002_),
    .X(_05003_));
 sg13g2_buf_1 _22609_ (.A(_05003_),
    .X(_05004_));
 sg13g2_nor3_1 _22610_ (.A(_04882_),
    .B(_05001_),
    .C(net68),
    .Y(_05005_));
 sg13g2_a21oi_1 _22611_ (.A1(net1122),
    .A2(_11526_),
    .Y(_05006_),
    .B1(_08190_));
 sg13g2_o21ai_1 _22612_ (.B1(net144),
    .Y(_05007_),
    .A1(_05005_),
    .A2(_05006_));
 sg13g2_nand2_1 _22613_ (.Y(_05008_),
    .A(net291),
    .B(net649));
 sg13g2_nand2_1 _22614_ (.Y(_05009_),
    .A(net214),
    .B(_11515_));
 sg13g2_buf_2 _22615_ (.A(_05009_),
    .X(_05010_));
 sg13g2_nor2_1 _22616_ (.A(_05008_),
    .B(_05010_),
    .Y(_05011_));
 sg13g2_a22oi_1 _22617_ (.Y(_01005_),
    .B1(_05011_),
    .B2(_11494_),
    .A2(_05007_),
    .A1(_04835_));
 sg13g2_nand2_1 _22618_ (.Y(_05012_),
    .A(net649),
    .B(_04760_));
 sg13g2_buf_1 _22619_ (.A(_04811_),
    .X(_05013_));
 sg13g2_buf_1 _22620_ (.A(net630),
    .X(_05014_));
 sg13g2_a21oi_1 _22621_ (.A1(_05014_),
    .A2(_04763_),
    .Y(_05015_),
    .B1(_05010_));
 sg13g2_buf_1 _22622_ (.A(net373),
    .X(_05016_));
 sg13g2_nand2_2 _22623_ (.Y(_05017_),
    .A(net288),
    .B(_11515_));
 sg13g2_buf_1 _22624_ (.A(net1038),
    .X(_05018_));
 sg13g2_nor2_1 _22625_ (.A(net763),
    .B(_04926_),
    .Y(_05019_));
 sg13g2_buf_2 _22626_ (.A(_05019_),
    .X(_05020_));
 sg13g2_nor3_1 _22627_ (.A(net896),
    .B(net674),
    .C(_05020_),
    .Y(_05021_));
 sg13g2_buf_2 _22628_ (.A(_05021_),
    .X(_05022_));
 sg13g2_buf_1 _22629_ (.A(_04910_),
    .X(_05023_));
 sg13g2_buf_1 _22630_ (.A(_04918_),
    .X(_05024_));
 sg13g2_a22oi_1 _22631_ (.Y(_05025_),
    .B1(net403),
    .B2(\cpu.intr.r_clock_cmp[10] ),
    .A2(net488),
    .A1(\cpu.intr.r_timer_reload[10] ));
 sg13g2_nor2_1 _22632_ (.A(net879),
    .B(_02697_),
    .Y(_05026_));
 sg13g2_buf_1 _22633_ (.A(_05026_),
    .X(_05027_));
 sg13g2_a22oi_1 _22634_ (.Y(_05028_),
    .B1(net444),
    .B2(\cpu.intr.r_clock_cmp[26] ),
    .A2(net462),
    .A1(_09987_));
 sg13g2_buf_1 _22635_ (.A(\cpu.intr.r_clock_count[26] ),
    .X(_05029_));
 sg13g2_buf_1 _22636_ (.A(_04948_),
    .X(_05030_));
 sg13g2_a22oi_1 _22637_ (.Y(_05031_),
    .B1(net487),
    .B2(_09794_),
    .A2(net423),
    .A1(_05029_));
 sg13g2_nand3_1 _22638_ (.B(_05028_),
    .C(_05031_),
    .A(_05025_),
    .Y(_05032_));
 sg13g2_buf_1 _22639_ (.A(net603),
    .X(_05033_));
 sg13g2_inv_1 _22640_ (.Y(_05034_),
    .A(_00092_));
 sg13g2_a22oi_1 _22641_ (.Y(_05035_),
    .B1(net486),
    .B2(_05034_),
    .A2(net511),
    .A1(\cpu.dcache.r_data[3][26] ));
 sg13g2_a22oi_1 _22642_ (.Y(_05036_),
    .B1(net529),
    .B2(\cpu.dcache.r_data[4][26] ),
    .A2(_03069_),
    .A1(\cpu.dcache.r_data[1][26] ));
 sg13g2_a22oi_1 _22643_ (.Y(_05037_),
    .B1(net510),
    .B2(\cpu.dcache.r_data[5][26] ),
    .A2(net599),
    .A1(\cpu.dcache.r_data[7][26] ));
 sg13g2_a22oi_1 _22644_ (.Y(_05038_),
    .B1(net489),
    .B2(\cpu.dcache.r_data[6][26] ),
    .A2(net512),
    .A1(\cpu.dcache.r_data[2][26] ));
 sg13g2_nand4_1 _22645_ (.B(_05036_),
    .C(_05037_),
    .A(_05035_),
    .Y(_05039_),
    .D(_05038_));
 sg13g2_a22oi_1 _22646_ (.Y(_05040_),
    .B1(_03083_),
    .B2(\cpu.dcache.r_data[6][10] ),
    .A2(net581),
    .A1(\cpu.dcache.r_data[5][10] ));
 sg13g2_a22oi_1 _22647_ (.Y(_05041_),
    .B1(net604),
    .B2(\cpu.dcache.r_data[4][10] ),
    .A2(net681),
    .A1(\cpu.dcache.r_data[3][10] ));
 sg13g2_nand2_1 _22648_ (.Y(_05042_),
    .A(_05040_),
    .B(_05041_));
 sg13g2_a221oi_1 _22649_ (.B2(\cpu.dcache.r_data[2][10] ),
    .C1(_05042_),
    .B1(net512),
    .A1(\cpu.dcache.r_data[7][10] ),
    .Y(_05043_),
    .A2(net675));
 sg13g2_mux2_1 _22650_ (.A0(_00093_),
    .A1(_05043_),
    .S(net676),
    .X(_05044_));
 sg13g2_nor2_1 _22651_ (.A(\cpu.dcache.r_data[1][10] ),
    .B(net531),
    .Y(_05045_));
 sg13g2_a22oi_1 _22652_ (.Y(_05046_),
    .B1(_05045_),
    .B2(_05043_),
    .A2(_05044_),
    .A1(net531));
 sg13g2_mux2_1 _22653_ (.A0(_05039_),
    .A1(_05046_),
    .S(net631),
    .X(_05047_));
 sg13g2_buf_1 _22654_ (.A(_04849_),
    .X(_05048_));
 sg13g2_a22oi_1 _22655_ (.Y(_05049_),
    .B1(_05047_),
    .B2(net485),
    .A2(_05032_),
    .A1(_05022_));
 sg13g2_inv_2 _22656_ (.Y(_05050_),
    .A(_04847_));
 sg13g2_inv_1 _22657_ (.Y(_05051_),
    .A(_00140_));
 sg13g2_a22oi_1 _22658_ (.Y(_05052_),
    .B1(net603),
    .B2(_05051_),
    .A2(net681),
    .A1(\cpu.dcache.r_data[3][31] ));
 sg13g2_a22oi_1 _22659_ (.Y(_05053_),
    .B1(net604),
    .B2(\cpu.dcache.r_data[4][31] ),
    .A2(net513),
    .A1(\cpu.dcache.r_data[1][31] ));
 sg13g2_a22oi_1 _22660_ (.Y(_05054_),
    .B1(_09420_),
    .B2(\cpu.dcache.r_data[6][31] ),
    .A2(net769),
    .A1(\cpu.dcache.r_data[7][31] ));
 sg13g2_a22oi_1 _22661_ (.Y(_05055_),
    .B1(net581),
    .B2(\cpu.dcache.r_data[5][31] ),
    .A2(net602),
    .A1(\cpu.dcache.r_data[2][31] ));
 sg13g2_nand4_1 _22662_ (.B(_05053_),
    .C(_05054_),
    .A(_05052_),
    .Y(_05056_),
    .D(_05055_));
 sg13g2_inv_1 _22663_ (.Y(_05057_),
    .A(_00139_));
 sg13g2_a22oi_1 _22664_ (.Y(_05058_),
    .B1(net603),
    .B2(_05057_),
    .A2(net681),
    .A1(\cpu.dcache.r_data[3][23] ));
 sg13g2_a22oi_1 _22665_ (.Y(_05059_),
    .B1(net769),
    .B2(\cpu.dcache.r_data[7][23] ),
    .A2(net513),
    .A1(\cpu.dcache.r_data[1][23] ));
 sg13g2_a22oi_1 _22666_ (.Y(_05060_),
    .B1(_09273_),
    .B2(\cpu.dcache.r_data[5][23] ),
    .A2(net604),
    .A1(\cpu.dcache.r_data[4][23] ));
 sg13g2_a22oi_1 _22667_ (.Y(_05061_),
    .B1(net677),
    .B2(\cpu.dcache.r_data[6][23] ),
    .A2(net602),
    .A1(\cpu.dcache.r_data[2][23] ));
 sg13g2_nand4_1 _22668_ (.B(_05059_),
    .C(_05060_),
    .A(_05058_),
    .Y(_05062_),
    .D(_05061_));
 sg13g2_nor2_2 _22669_ (.A(_09873_),
    .B(_05050_),
    .Y(_05063_));
 sg13g2_a22oi_1 _22670_ (.Y(_05064_),
    .B1(_05062_),
    .B2(_05063_),
    .A2(_05056_),
    .A1(_05050_));
 sg13g2_inv_1 _22671_ (.Y(_05065_),
    .A(_00141_));
 sg13g2_a22oi_1 _22672_ (.Y(_05066_),
    .B1(net603),
    .B2(_05065_),
    .A2(net681),
    .A1(\cpu.dcache.r_data[3][15] ));
 sg13g2_a22oi_1 _22673_ (.Y(_05067_),
    .B1(net604),
    .B2(\cpu.dcache.r_data[4][15] ),
    .A2(_03068_),
    .A1(\cpu.dcache.r_data[1][15] ));
 sg13g2_a22oi_1 _22674_ (.Y(_05068_),
    .B1(net580),
    .B2(\cpu.dcache.r_data[6][15] ),
    .A2(net675),
    .A1(\cpu.dcache.r_data[7][15] ));
 sg13g2_a22oi_1 _22675_ (.Y(_05069_),
    .B1(net581),
    .B2(\cpu.dcache.r_data[5][15] ),
    .A2(net602),
    .A1(\cpu.dcache.r_data[2][15] ));
 sg13g2_nand4_1 _22676_ (.B(_05067_),
    .C(_05068_),
    .A(_05066_),
    .Y(_05070_),
    .D(_05069_));
 sg13g2_nor2_1 _22677_ (.A(_09775_),
    .B(_04847_),
    .Y(_05071_));
 sg13g2_mux2_1 _22678_ (.A0(\cpu.dcache.r_data[5][7] ),
    .A1(\cpu.dcache.r_data[7][7] ),
    .S(net685),
    .X(_05072_));
 sg13g2_a22oi_1 _22679_ (.Y(_05073_),
    .B1(_05072_),
    .B2(net609),
    .A2(net680),
    .A1(\cpu.dcache.r_data[6][7] ));
 sg13g2_nor2_1 _22680_ (.A(net777),
    .B(_05073_),
    .Y(_05074_));
 sg13g2_mux2_1 _22681_ (.A0(\cpu.dcache.r_data[1][7] ),
    .A1(\cpu.dcache.r_data[3][7] ),
    .S(net608),
    .X(_05075_));
 sg13g2_a22oi_1 _22682_ (.Y(_05076_),
    .B1(_05075_),
    .B2(net609),
    .A2(net680),
    .A1(\cpu.dcache.r_data[2][7] ));
 sg13g2_nor2_1 _22683_ (.A(_09305_),
    .B(_05076_),
    .Y(_05077_));
 sg13g2_nand2_1 _22684_ (.Y(_05078_),
    .A(\cpu.dcache.r_data[4][7] ),
    .B(net604));
 sg13g2_o21ai_1 _22685_ (.B1(_05078_),
    .Y(_05079_),
    .A1(_00138_),
    .A2(net490));
 sg13g2_nor3_2 _22686_ (.A(_05074_),
    .B(_05077_),
    .C(_05079_),
    .Y(_05080_));
 sg13g2_nor2_1 _22687_ (.A(_04875_),
    .B(_05080_),
    .Y(_05081_));
 sg13g2_a21oi_1 _22688_ (.A1(_05070_),
    .A2(_05071_),
    .Y(_05082_),
    .B1(_05081_));
 sg13g2_o21ai_1 _22689_ (.B1(_05082_),
    .Y(_05083_),
    .A1(_11984_),
    .A2(_05064_));
 sg13g2_inv_1 _22690_ (.Y(_05084_),
    .A(_05062_));
 sg13g2_mux2_1 _22691_ (.A0(_05084_),
    .A1(_05080_),
    .S(net879),
    .X(_05085_));
 sg13g2_nand2_1 _22692_ (.Y(_05086_),
    .A(net564),
    .B(_05085_));
 sg13g2_o21ai_1 _22693_ (.B1(_05086_),
    .Y(_05087_),
    .A1(net564),
    .A2(_05083_));
 sg13g2_and2_1 _22694_ (.A(_10473_),
    .B(_04889_),
    .X(_05088_));
 sg13g2_buf_2 _22695_ (.A(_05088_),
    .X(_05089_));
 sg13g2_a21o_1 _22696_ (.A2(_04996_),
    .A1(_08987_),
    .B1(_05089_),
    .X(_05090_));
 sg13g2_nor3_1 _22697_ (.A(net879),
    .B(_00148_),
    .C(_02697_),
    .Y(_05091_));
 sg13g2_a22oi_1 _22698_ (.Y(_05092_),
    .B1(_09273_),
    .B2(net10),
    .A2(_09300_),
    .A1(\cpu.gpio.genblk1[7].srcs_o[0] ));
 sg13g2_nor2_1 _22699_ (.A(net676),
    .B(net598),
    .Y(_05093_));
 sg13g2_buf_1 _22700_ (.A(_05093_),
    .X(_05094_));
 sg13g2_a21oi_1 _22701_ (.A1(_08992_),
    .A2(_05094_),
    .Y(_05095_),
    .B1(net404));
 sg13g2_nand2b_1 _22702_ (.Y(_05096_),
    .B(_08993_),
    .A_N(_05095_));
 sg13g2_o21ai_1 _22703_ (.B1(_05096_),
    .Y(_05097_),
    .A1(net1025),
    .A2(_05092_));
 sg13g2_or2_1 _22704_ (.X(_05098_),
    .B(_05097_),
    .A(_05091_));
 sg13g2_and2_1 _22705_ (.A(net952),
    .B(\cpu.gpio.genblk2[7].srcs_io[0] ),
    .X(_05099_));
 sg13g2_nor2_1 _22706_ (.A(net952),
    .B(_00146_),
    .Y(_05100_));
 sg13g2_a22oi_1 _22707_ (.Y(_05101_),
    .B1(_05100_),
    .B2(_04897_),
    .A2(_05099_),
    .A1(_09964_));
 sg13g2_nor2_1 _22708_ (.A(_10473_),
    .B(_00147_),
    .Y(_05102_));
 sg13g2_nor2b_1 _22709_ (.A(net994),
    .B_N(_08987_),
    .Y(_05103_));
 sg13g2_a22oi_1 _22710_ (.Y(_05104_),
    .B1(_05103_),
    .B2(_04897_),
    .A2(_05102_),
    .A1(_05094_));
 sg13g2_buf_1 _22711_ (.A(\cpu.gpio.r_src_io[5][3] ),
    .X(_05105_));
 sg13g2_inv_1 _22712_ (.Y(_05106_),
    .A(_00144_));
 sg13g2_a22oi_1 _22713_ (.Y(_05107_),
    .B1(_04974_),
    .B2(_05106_),
    .A2(net354),
    .A1(_05105_));
 sg13g2_inv_1 _22714_ (.Y(_05108_),
    .A(_00145_));
 sg13g2_nor2_1 _22715_ (.A(net994),
    .B(_04940_),
    .Y(_05109_));
 sg13g2_buf_1 _22716_ (.A(_05109_),
    .X(_05110_));
 sg13g2_a22oi_1 _22717_ (.Y(_05111_),
    .B1(_05110_),
    .B2(_08992_),
    .A2(_04980_),
    .A1(_05108_));
 sg13g2_nand4_1 _22718_ (.B(_05104_),
    .C(_05107_),
    .A(_05101_),
    .Y(_05112_),
    .D(_05111_));
 sg13g2_a221oi_1 _22719_ (.B2(_04954_),
    .C1(_05112_),
    .B1(_05098_),
    .A1(\cpu.gpio.r_enable_in[7] ),
    .Y(_05113_),
    .A2(_05090_));
 sg13g2_nor2_1 _22720_ (.A(net674),
    .B(_05020_),
    .Y(_05114_));
 sg13g2_buf_2 _22721_ (.A(\cpu.intr.r_clock_count[23] ),
    .X(_05115_));
 sg13g2_mux2_1 _22722_ (.A0(\cpu.intr.r_clock_cmp[7] ),
    .A1(\cpu.intr.r_clock_cmp[23] ),
    .S(net1025),
    .X(_05116_));
 sg13g2_a22oi_1 _22723_ (.Y(_05117_),
    .B1(_05116_),
    .B2(net581),
    .A2(_09964_),
    .A1(_05115_));
 sg13g2_nand2_1 _22724_ (.Y(_05118_),
    .A(\cpu.intr.r_timer_reload[7] ),
    .B(_04910_));
 sg13g2_a22oi_1 _22725_ (.Y(_05119_),
    .B1(net677),
    .B2(_09815_),
    .A2(net769),
    .A1(\cpu.intr.r_timer_reload[23] ));
 sg13g2_nand2b_1 _22726_ (.Y(_05120_),
    .B(net1025),
    .A_N(_05119_));
 sg13g2_a22oi_1 _22727_ (.Y(_05121_),
    .B1(_04948_),
    .B2(_09795_),
    .A2(_09921_),
    .A1(_09970_));
 sg13g2_nand4_1 _22728_ (.B(_05118_),
    .C(_05120_),
    .A(_05117_),
    .Y(_05122_),
    .D(_05121_));
 sg13g2_buf_1 _22729_ (.A(\cpu.spi.r_clk_count[2][7] ),
    .X(_05123_));
 sg13g2_inv_1 _22730_ (.Y(_05124_),
    .A(_00143_));
 sg13g2_a22oi_1 _22731_ (.Y(_05125_),
    .B1(_05110_),
    .B2(_05124_),
    .A2(_04956_),
    .A1(_05123_));
 sg13g2_nor2_1 _22732_ (.A(net781),
    .B(_04891_),
    .Y(_05126_));
 sg13g2_buf_2 _22733_ (.A(_05126_),
    .X(_05127_));
 sg13g2_nor2_1 _22734_ (.A(_00142_),
    .B(_04959_),
    .Y(_05128_));
 sg13g2_a21oi_1 _22735_ (.A1(\cpu.spi.r_timeout[7] ),
    .A2(_05127_),
    .Y(_05129_),
    .B1(_05128_));
 sg13g2_nand2b_1 _22736_ (.Y(_05130_),
    .B(_04943_),
    .A_N(_00200_));
 sg13g2_nand3_1 _22737_ (.B(_05129_),
    .C(_05130_),
    .A(_05125_),
    .Y(_05131_));
 sg13g2_and2_1 _22738_ (.A(_09023_),
    .B(_09028_),
    .X(_05132_));
 sg13g2_buf_1 _22739_ (.A(_05132_),
    .X(_05133_));
 sg13g2_a22oi_1 _22740_ (.Y(_05134_),
    .B1(_04886_),
    .B2(\cpu.uart.r_in[7] ),
    .A2(net405),
    .A1(\cpu.uart.r_div_value[7] ));
 sg13g2_nor2_1 _22741_ (.A(_04884_),
    .B(_05134_),
    .Y(_05135_));
 sg13g2_a221oi_1 _22742_ (.B2(_05133_),
    .C1(_05135_),
    .B1(_05131_),
    .A1(_05114_),
    .Y(_05136_),
    .A2(_05122_));
 sg13g2_o21ai_1 _22743_ (.B1(_05136_),
    .Y(_05137_),
    .A1(_04999_),
    .A2(_05113_));
 sg13g2_nor2_1 _22744_ (.A(net896),
    .B(_05137_),
    .Y(_05138_));
 sg13g2_a21oi_1 _22745_ (.A1(net896),
    .A2(_05087_),
    .Y(_05139_),
    .B1(_05138_));
 sg13g2_a21oi_1 _22746_ (.A1(net1038),
    .A2(_05139_),
    .Y(_05140_),
    .B1(_11515_));
 sg13g2_buf_2 _22747_ (.A(_05140_),
    .X(_05141_));
 sg13g2_o21ai_1 _22748_ (.B1(_05141_),
    .Y(_05142_),
    .A1(net832),
    .A2(_05049_));
 sg13g2_a21oi_1 _22749_ (.A1(net1122),
    .A2(_11528_),
    .Y(_05143_),
    .B1(_11515_));
 sg13g2_buf_2 _22750_ (.A(_05143_),
    .X(_05144_));
 sg13g2_mux2_1 _22751_ (.A0(_05142_),
    .A1(net1095),
    .S(_05144_),
    .X(_05145_));
 sg13g2_o21ai_1 _22752_ (.B1(_05145_),
    .Y(_05146_),
    .A1(net954),
    .A2(_05017_));
 sg13g2_a21oi_1 _22753_ (.A1(_05012_),
    .A2(_05015_),
    .Y(_01006_),
    .B1(_05146_));
 sg13g2_buf_1 _22754_ (.A(net111),
    .X(_05147_));
 sg13g2_or3_1 _22755_ (.A(net373),
    .B(net649),
    .C(_04253_),
    .X(_05148_));
 sg13g2_o21ai_1 _22756_ (.B1(_05148_),
    .Y(_05149_),
    .A1(net959),
    .A2(net214));
 sg13g2_nor2_1 _22757_ (.A(net563),
    .B(_05010_),
    .Y(_05150_));
 sg13g2_buf_1 _22758_ (.A(net1038),
    .X(_05151_));
 sg13g2_a22oi_1 _22759_ (.Y(_05152_),
    .B1(net444),
    .B2(\cpu.intr.r_clock_cmp[27] ),
    .A2(net488),
    .A1(\cpu.intr.r_timer_reload[11] ));
 sg13g2_a22oi_1 _22760_ (.Y(_05153_),
    .B1(net487),
    .B2(_09793_),
    .A2(net462),
    .A1(_09992_));
 sg13g2_buf_2 _22761_ (.A(\cpu.intr.r_clock_count[27] ),
    .X(_05154_));
 sg13g2_a22oi_1 _22762_ (.Y(_05155_),
    .B1(net403),
    .B2(\cpu.intr.r_clock_cmp[11] ),
    .A2(net423),
    .A1(_05154_));
 sg13g2_nand3_1 _22763_ (.B(_05153_),
    .C(_05155_),
    .A(_05152_),
    .Y(_05156_));
 sg13g2_mux2_1 _22764_ (.A0(\cpu.dcache.r_data[1][27] ),
    .A1(\cpu.dcache.r_data[3][27] ),
    .S(net532),
    .X(_05157_));
 sg13g2_a22oi_1 _22765_ (.Y(_05158_),
    .B1(_05157_),
    .B2(net456),
    .A2(net680),
    .A1(\cpu.dcache.r_data[2][27] ));
 sg13g2_inv_1 _22766_ (.Y(_05159_),
    .A(_00102_));
 sg13g2_mux2_1 _22767_ (.A0(\cpu.dcache.r_data[5][27] ),
    .A1(\cpu.dcache.r_data[7][27] ),
    .S(_09104_),
    .X(_05160_));
 sg13g2_a22oi_1 _22768_ (.Y(_05161_),
    .B1(_05160_),
    .B2(net517),
    .A2(_09426_),
    .A1(\cpu.dcache.r_data[4][27] ));
 sg13g2_nor2_1 _22769_ (.A(net777),
    .B(_05161_),
    .Y(_05162_));
 sg13g2_a221oi_1 _22770_ (.B2(\cpu.dcache.r_data[6][27] ),
    .C1(_05162_),
    .B1(net489),
    .A1(_05159_),
    .Y(_05163_),
    .A2(net603));
 sg13g2_o21ai_1 _22771_ (.B1(_05163_),
    .Y(_05164_),
    .A1(_09305_),
    .A2(_05158_));
 sg13g2_inv_1 _22772_ (.Y(_05165_),
    .A(_00103_));
 sg13g2_a22oi_1 _22773_ (.Y(_05166_),
    .B1(net603),
    .B2(_05165_),
    .A2(net511),
    .A1(\cpu.dcache.r_data[3][11] ));
 sg13g2_a22oi_1 _22774_ (.Y(_05167_),
    .B1(_09779_),
    .B2(\cpu.dcache.r_data[7][11] ),
    .A2(net455),
    .A1(\cpu.dcache.r_data[1][11] ));
 sg13g2_a22oi_1 _22775_ (.Y(_05168_),
    .B1(_03080_),
    .B2(\cpu.dcache.r_data[5][11] ),
    .A2(net529),
    .A1(\cpu.dcache.r_data[4][11] ));
 sg13g2_a22oi_1 _22776_ (.Y(_05169_),
    .B1(net489),
    .B2(\cpu.dcache.r_data[6][11] ),
    .A2(_03072_),
    .A1(\cpu.dcache.r_data[2][11] ));
 sg13g2_nand4_1 _22777_ (.B(_05167_),
    .C(_05168_),
    .A(_05166_),
    .Y(_05170_),
    .D(_05169_));
 sg13g2_mux2_1 _22778_ (.A0(_05164_),
    .A1(_05170_),
    .S(net673),
    .X(_05171_));
 sg13g2_a22oi_1 _22779_ (.Y(_05172_),
    .B1(_05171_),
    .B2(net485),
    .A2(_05156_),
    .A1(_05022_));
 sg13g2_o21ai_1 _22780_ (.B1(_05141_),
    .Y(_05173_),
    .A1(net831),
    .A2(_05172_));
 sg13g2_nand2b_1 _22781_ (.Y(_05174_),
    .B(_05144_),
    .A_N(_10907_));
 sg13g2_o21ai_1 _22782_ (.B1(_05174_),
    .Y(_05175_),
    .A1(_05144_),
    .A2(_05173_));
 sg13g2_a221oi_1 _22783_ (.B2(_04243_),
    .C1(_05175_),
    .B1(_05150_),
    .A1(net94),
    .Y(_01007_),
    .A2(_05149_));
 sg13g2_a22oi_1 _22784_ (.Y(_05176_),
    .B1(net487),
    .B2(\cpu.intr.r_timer_count[12] ),
    .A2(net488),
    .A1(\cpu.intr.r_timer_reload[12] ));
 sg13g2_a22oi_1 _22785_ (.Y(_05177_),
    .B1(net444),
    .B2(\cpu.intr.r_clock_cmp[28] ),
    .A2(net462),
    .A1(_09998_));
 sg13g2_buf_2 _22786_ (.A(\cpu.intr.r_clock_count[28] ),
    .X(_05178_));
 sg13g2_a22oi_1 _22787_ (.Y(_05179_),
    .B1(net403),
    .B2(\cpu.intr.r_clock_cmp[12] ),
    .A2(_09966_),
    .A1(_05178_));
 sg13g2_nand3_1 _22788_ (.B(_05177_),
    .C(_05179_),
    .A(_05176_),
    .Y(_05180_));
 sg13g2_inv_1 _22789_ (.Y(_05181_),
    .A(_00112_));
 sg13g2_a22oi_1 _22790_ (.Y(_05182_),
    .B1(net603),
    .B2(_05181_),
    .A2(net582),
    .A1(\cpu.dcache.r_data[3][28] ));
 sg13g2_a22oi_1 _22791_ (.Y(_05183_),
    .B1(_09778_),
    .B2(\cpu.dcache.r_data[7][28] ),
    .A2(net513),
    .A1(\cpu.dcache.r_data[1][28] ));
 sg13g2_a22oi_1 _22792_ (.Y(_05184_),
    .B1(net510),
    .B2(\cpu.dcache.r_data[5][28] ),
    .A2(net529),
    .A1(\cpu.dcache.r_data[4][28] ));
 sg13g2_a22oi_1 _22793_ (.Y(_05185_),
    .B1(_03083_),
    .B2(\cpu.dcache.r_data[6][28] ),
    .A2(_03072_),
    .A1(\cpu.dcache.r_data[2][28] ));
 sg13g2_nand4_1 _22794_ (.B(_05183_),
    .C(_05184_),
    .A(_05182_),
    .Y(_05186_),
    .D(_05185_));
 sg13g2_buf_1 _22795_ (.A(_05186_),
    .X(_05187_));
 sg13g2_inv_1 _22796_ (.Y(_05188_),
    .A(_00113_));
 sg13g2_a22oi_1 _22797_ (.Y(_05189_),
    .B1(net486),
    .B2(_05188_),
    .A2(_09779_),
    .A1(\cpu.dcache.r_data[7][12] ));
 sg13g2_nand2_1 _22798_ (.Y(_05190_),
    .A(\cpu.dcache.r_data[6][12] ),
    .B(_04862_));
 sg13g2_a22oi_1 _22799_ (.Y(_05191_),
    .B1(_09915_),
    .B2(\cpu.dcache.r_data[4][12] ),
    .A2(net455),
    .A1(\cpu.dcache.r_data[1][12] ));
 sg13g2_mux2_1 _22800_ (.A0(\cpu.dcache.r_data[2][12] ),
    .A1(\cpu.dcache.r_data[3][12] ),
    .S(net517),
    .X(_05192_));
 sg13g2_a22oi_1 _22801_ (.Y(_05193_),
    .B1(_05192_),
    .B2(net890),
    .A2(net510),
    .A1(\cpu.dcache.r_data[5][12] ));
 sg13g2_nand4_1 _22802_ (.B(_05190_),
    .C(_05191_),
    .A(_05189_),
    .Y(_05194_),
    .D(_05193_));
 sg13g2_and2_1 _22803_ (.A(net754),
    .B(_05194_),
    .X(_05195_));
 sg13g2_a21o_1 _22804_ (.A2(_05187_),
    .A1(net637),
    .B1(_05195_),
    .X(_05196_));
 sg13g2_a22oi_1 _22805_ (.Y(_05197_),
    .B1(_05196_),
    .B2(net485),
    .A2(_05180_),
    .A1(_05022_));
 sg13g2_o21ai_1 _22806_ (.B1(_05141_),
    .Y(_05198_),
    .A1(net832),
    .A2(_05197_));
 sg13g2_mux2_1 _22807_ (.A0(_05198_),
    .A1(net589),
    .S(_05144_),
    .X(_05199_));
 sg13g2_o21ai_1 _22808_ (.B1(_05199_),
    .Y(_05200_),
    .A1(_08464_),
    .A2(_05017_));
 sg13g2_a21oi_1 _22809_ (.A1(net563),
    .A2(_04300_),
    .Y(_05201_),
    .B1(_05010_));
 sg13g2_o21ai_1 _22810_ (.B1(_05201_),
    .Y(_05202_),
    .A1(net563),
    .A2(_04298_));
 sg13g2_nor2b_1 _22811_ (.A(_05200_),
    .B_N(_05202_),
    .Y(_01008_));
 sg13g2_or2_1 _22812_ (.X(_05203_),
    .B(_04338_),
    .A(net630));
 sg13g2_a21o_1 _22813_ (.A2(_04002_),
    .A1(_11823_),
    .B1(_05203_),
    .X(_05204_));
 sg13g2_a21oi_1 _22814_ (.A1(net563),
    .A2(_04341_),
    .Y(_05205_),
    .B1(_05010_));
 sg13g2_a22oi_1 _22815_ (.Y(_05206_),
    .B1(net488),
    .B2(\cpu.intr.r_timer_reload[13] ),
    .A2(net462),
    .A1(_10002_));
 sg13g2_a22oi_1 _22816_ (.Y(_05207_),
    .B1(net403),
    .B2(\cpu.intr.r_clock_cmp[13] ),
    .A2(net487),
    .A1(\cpu.intr.r_timer_count[13] ));
 sg13g2_buf_2 _22817_ (.A(\cpu.intr.r_clock_count[29] ),
    .X(_05208_));
 sg13g2_a22oi_1 _22818_ (.Y(_05209_),
    .B1(net444),
    .B2(\cpu.intr.r_clock_cmp[29] ),
    .A2(net423),
    .A1(_05208_));
 sg13g2_nand3_1 _22819_ (.B(_05207_),
    .C(_05209_),
    .A(_05206_),
    .Y(_05210_));
 sg13g2_inv_1 _22820_ (.Y(_05211_),
    .A(_00118_));
 sg13g2_a22oi_1 _22821_ (.Y(_05212_),
    .B1(_05033_),
    .B2(_05211_),
    .A2(net511),
    .A1(\cpu.dcache.r_data[3][29] ));
 sg13g2_a22oi_1 _22822_ (.Y(_05213_),
    .B1(_09780_),
    .B2(\cpu.dcache.r_data[7][29] ),
    .A2(net413),
    .A1(\cpu.dcache.r_data[1][29] ));
 sg13g2_a22oi_1 _22823_ (.Y(_05214_),
    .B1(net453),
    .B2(\cpu.dcache.r_data[5][29] ),
    .A2(net463),
    .A1(\cpu.dcache.r_data[4][29] ));
 sg13g2_a22oi_1 _22824_ (.Y(_05215_),
    .B1(_03084_),
    .B2(\cpu.dcache.r_data[6][29] ),
    .A2(_03073_),
    .A1(\cpu.dcache.r_data[2][29] ));
 sg13g2_nand4_1 _22825_ (.B(_05213_),
    .C(_05214_),
    .A(_05212_),
    .Y(_05216_),
    .D(_05215_));
 sg13g2_mux2_1 _22826_ (.A0(\cpu.dcache.r_data[4][13] ),
    .A1(\cpu.dcache.r_data[6][13] ),
    .S(net532),
    .X(_05217_));
 sg13g2_a22oi_1 _22827_ (.Y(_05218_),
    .B1(_05217_),
    .B2(net644),
    .A2(_09379_),
    .A1(\cpu.dcache.r_data[7][13] ));
 sg13g2_a22oi_1 _22828_ (.Y(_05219_),
    .B1(net510),
    .B2(\cpu.dcache.r_data[5][13] ),
    .A2(net582),
    .A1(\cpu.dcache.r_data[3][13] ));
 sg13g2_o21ai_1 _22829_ (.B1(_05219_),
    .Y(_05220_),
    .A1(_00119_),
    .A2(net490));
 sg13g2_a221oi_1 _22830_ (.B2(\cpu.dcache.r_data[2][13] ),
    .C1(_05220_),
    .B1(net454),
    .A1(\cpu.dcache.r_data[1][13] ),
    .Y(_05221_),
    .A2(net455));
 sg13g2_o21ai_1 _22831_ (.B1(_05221_),
    .Y(_05222_),
    .A1(net645),
    .A2(_05218_));
 sg13g2_mux2_1 _22832_ (.A0(_05216_),
    .A1(_05222_),
    .S(net631),
    .X(_05223_));
 sg13g2_a22oi_1 _22833_ (.Y(_05224_),
    .B1(_05223_),
    .B2(net485),
    .A2(_05210_),
    .A1(_05022_));
 sg13g2_o21ai_1 _22834_ (.B1(_05141_),
    .Y(_05225_),
    .A1(net832),
    .A2(_05224_));
 sg13g2_mux2_1 _22835_ (.A0(_05225_),
    .A1(net601),
    .S(_05144_),
    .X(_05226_));
 sg13g2_o21ai_1 _22836_ (.B1(_05226_),
    .Y(_05227_),
    .A1(net616),
    .A2(_05017_));
 sg13g2_a21oi_1 _22837_ (.A1(_05204_),
    .A2(_05205_),
    .Y(_01009_),
    .B1(_05227_));
 sg13g2_buf_1 _22838_ (.A(net144),
    .X(_05228_));
 sg13g2_a22oi_1 _22839_ (.Y(_05229_),
    .B1(net403),
    .B2(\cpu.intr.r_clock_cmp[14] ),
    .A2(net488),
    .A1(\cpu.intr.r_timer_reload[14] ));
 sg13g2_a22oi_1 _22840_ (.Y(_05230_),
    .B1(net487),
    .B2(\cpu.intr.r_timer_count[14] ),
    .A2(net528),
    .A1(_10008_));
 sg13g2_buf_1 _22841_ (.A(\cpu.intr.r_clock_count[30] ),
    .X(_05231_));
 sg13g2_a22oi_1 _22842_ (.Y(_05232_),
    .B1(net444),
    .B2(\cpu.intr.r_clock_cmp[30] ),
    .A2(net423),
    .A1(_05231_));
 sg13g2_nand3_1 _22843_ (.B(_05230_),
    .C(_05232_),
    .A(_05229_),
    .Y(_05233_));
 sg13g2_mux2_1 _22844_ (.A0(\cpu.dcache.r_data[4][30] ),
    .A1(\cpu.dcache.r_data[6][30] ),
    .S(_09105_),
    .X(_05234_));
 sg13g2_a22oi_1 _22845_ (.Y(_05235_),
    .B1(_05234_),
    .B2(net768),
    .A2(_09379_),
    .A1(\cpu.dcache.r_data[7][30] ));
 sg13g2_a22oi_1 _22846_ (.Y(_05236_),
    .B1(_03079_),
    .B2(\cpu.dcache.r_data[5][30] ),
    .A2(_03075_),
    .A1(\cpu.dcache.r_data[3][30] ));
 sg13g2_o21ai_1 _22847_ (.B1(_05236_),
    .Y(_05237_),
    .A1(_00129_),
    .A2(_04855_));
 sg13g2_a221oi_1 _22848_ (.B2(\cpu.dcache.r_data[2][30] ),
    .C1(_05237_),
    .B1(net454),
    .A1(\cpu.dcache.r_data[1][30] ),
    .Y(_05238_),
    .A2(_03069_));
 sg13g2_o21ai_1 _22849_ (.B1(_05238_),
    .Y(_05239_),
    .A1(net645),
    .A2(_05235_));
 sg13g2_mux2_1 _22850_ (.A0(\cpu.dcache.r_data[1][14] ),
    .A1(\cpu.dcache.r_data[3][14] ),
    .S(net608),
    .X(_05240_));
 sg13g2_a22oi_1 _22851_ (.Y(_05241_),
    .B1(_05240_),
    .B2(net517),
    .A2(net680),
    .A1(\cpu.dcache.r_data[2][14] ));
 sg13g2_nand2b_1 _22852_ (.Y(_05242_),
    .B(net1028),
    .A_N(_05241_));
 sg13g2_mux2_1 _22853_ (.A0(\cpu.dcache.r_data[5][14] ),
    .A1(\cpu.dcache.r_data[7][14] ),
    .S(net608),
    .X(_05243_));
 sg13g2_a22oi_1 _22854_ (.Y(_05244_),
    .B1(_05243_),
    .B2(_12460_),
    .A2(_09426_),
    .A1(\cpu.dcache.r_data[4][14] ));
 sg13g2_nand2b_1 _22855_ (.Y(_05245_),
    .B(_11939_),
    .A_N(_05244_));
 sg13g2_inv_1 _22856_ (.Y(_05246_),
    .A(_00130_));
 sg13g2_a22oi_1 _22857_ (.Y(_05247_),
    .B1(net489),
    .B2(\cpu.dcache.r_data[6][14] ),
    .A2(net486),
    .A1(_05246_));
 sg13g2_nand3_1 _22858_ (.B(_05245_),
    .C(_05247_),
    .A(_05242_),
    .Y(_05248_));
 sg13g2_mux2_1 _22859_ (.A0(_05239_),
    .A1(_05248_),
    .S(net631),
    .X(_05249_));
 sg13g2_a22oi_1 _22860_ (.Y(_05250_),
    .B1(_05249_),
    .B2(net485),
    .A2(_05233_),
    .A1(_05022_));
 sg13g2_o21ai_1 _22861_ (.B1(_05141_),
    .Y(_05251_),
    .A1(net832),
    .A2(_05250_));
 sg13g2_mux2_1 _22862_ (.A0(_05251_),
    .A1(net732),
    .S(_05003_),
    .X(_05252_));
 sg13g2_nand2_1 _22863_ (.Y(_05253_),
    .A(net110),
    .B(_05252_));
 sg13g2_o21ai_1 _22864_ (.B1(net111),
    .Y(_05254_),
    .A1(net906),
    .A2(net214));
 sg13g2_nand3_1 _22865_ (.B(_04343_),
    .C(_04387_),
    .A(_11507_),
    .Y(_05255_));
 sg13g2_a21oi_1 _22866_ (.A1(net563),
    .A2(_04390_),
    .Y(_05256_),
    .B1(_05010_));
 sg13g2_a22oi_1 _22867_ (.Y(_01010_),
    .B1(_05255_),
    .B2(_05256_),
    .A2(_05254_),
    .A1(_05253_));
 sg13g2_nor2_1 _22868_ (.A(net649),
    .B(_04437_),
    .Y(_05257_));
 sg13g2_nor2_1 _22869_ (.A(net288),
    .B(net144),
    .Y(_05258_));
 sg13g2_buf_1 _22870_ (.A(_05258_),
    .X(_05259_));
 sg13g2_a22oi_1 _22871_ (.Y(_05260_),
    .B1(_05030_),
    .B2(\cpu.intr.r_timer_count[15] ),
    .A2(_05023_),
    .A1(\cpu.intr.r_timer_reload[15] ));
 sg13g2_a22oi_1 _22872_ (.Y(_05261_),
    .B1(_05027_),
    .B2(\cpu.intr.r_clock_cmp[31] ),
    .A2(net528),
    .A1(_10013_));
 sg13g2_buf_1 _22873_ (.A(\cpu.intr.r_clock_count[31] ),
    .X(_05262_));
 sg13g2_a22oi_1 _22874_ (.Y(_05263_),
    .B1(_04918_),
    .B2(\cpu.intr.r_clock_cmp[15] ),
    .A2(net461),
    .A1(_05262_));
 sg13g2_nand3_1 _22875_ (.B(_05261_),
    .C(_05263_),
    .A(_05260_),
    .Y(_05264_));
 sg13g2_mux2_1 _22876_ (.A0(_05056_),
    .A1(_05070_),
    .S(net631),
    .X(_05265_));
 sg13g2_a22oi_1 _22877_ (.Y(_05266_),
    .B1(_05265_),
    .B2(net564),
    .A2(_05264_),
    .A1(_05022_));
 sg13g2_o21ai_1 _22878_ (.B1(_05141_),
    .Y(_05267_),
    .A1(net1038),
    .A2(_05266_));
 sg13g2_mux2_1 _22879_ (.A0(_05267_),
    .A1(net731),
    .S(_05003_),
    .X(_05268_));
 sg13g2_nand3_1 _22880_ (.B(net288),
    .C(_11515_),
    .A(net790),
    .Y(_05269_));
 sg13g2_o21ai_1 _22881_ (.B1(_05269_),
    .Y(_05270_),
    .A1(net111),
    .A2(_05268_));
 sg13g2_a221oi_1 _22882_ (.B2(_05259_),
    .C1(_05270_),
    .B1(_05257_),
    .A1(_04435_),
    .Y(_01011_),
    .A2(_05150_));
 sg13g2_inv_1 _22883_ (.Y(_05271_),
    .A(_11562_));
 sg13g2_nand2b_1 _22884_ (.Y(_05272_),
    .B(_11538_),
    .A_N(_05008_));
 sg13g2_buf_8 _22885_ (.A(_05272_),
    .X(_05273_));
 sg13g2_nand2_1 _22886_ (.Y(_05274_),
    .A(_10326_),
    .B(net630));
 sg13g2_o21ai_1 _22887_ (.B1(_05274_),
    .Y(_05275_),
    .A1(net563),
    .A2(_04125_));
 sg13g2_o21ai_1 _22888_ (.B1(_05275_),
    .Y(_05276_),
    .A1(_05271_),
    .A2(_05273_));
 sg13g2_nand2_1 _22889_ (.Y(_05277_),
    .A(\cpu.dcache.r_data[0][1] ),
    .B(net486));
 sg13g2_a22oi_1 _22890_ (.Y(_05278_),
    .B1(net509),
    .B2(\cpu.dcache.r_data[6][1] ),
    .A2(_03076_),
    .A1(\cpu.dcache.r_data[3][1] ));
 sg13g2_a22oi_1 _22891_ (.Y(_05279_),
    .B1(net454),
    .B2(\cpu.dcache.r_data[2][1] ),
    .A2(net413),
    .A1(\cpu.dcache.r_data[1][1] ));
 sg13g2_mux2_1 _22892_ (.A0(\cpu.dcache.r_data[5][1] ),
    .A1(\cpu.dcache.r_data[7][1] ),
    .S(net532),
    .X(_05280_));
 sg13g2_a22oi_1 _22893_ (.Y(_05281_),
    .B1(_05280_),
    .B2(_12461_),
    .A2(_09426_),
    .A1(\cpu.dcache.r_data[4][1] ));
 sg13g2_nand2b_1 _22894_ (.Y(_05282_),
    .B(net646),
    .A_N(_05281_));
 sg13g2_nand4_1 _22895_ (.B(_05278_),
    .C(_05279_),
    .A(_05277_),
    .Y(_05283_),
    .D(_05282_));
 sg13g2_mux2_1 _22896_ (.A0(\cpu.dcache.r_data[4][17] ),
    .A1(\cpu.dcache.r_data[6][17] ),
    .S(net464),
    .X(_05284_));
 sg13g2_a22oi_1 _22897_ (.Y(_05285_),
    .B1(_05284_),
    .B2(net644),
    .A2(_09367_),
    .A1(\cpu.dcache.r_data[5][17] ));
 sg13g2_a22oi_1 _22898_ (.Y(_05286_),
    .B1(net511),
    .B2(\cpu.dcache.r_data[3][17] ),
    .A2(net599),
    .A1(\cpu.dcache.r_data[7][17] ));
 sg13g2_o21ai_1 _22899_ (.B1(_05286_),
    .Y(_05287_),
    .A1(_00282_),
    .A2(net490));
 sg13g2_a221oi_1 _22900_ (.B2(\cpu.dcache.r_data[2][17] ),
    .C1(_05287_),
    .B1(net454),
    .A1(\cpu.dcache.r_data[1][17] ),
    .Y(_05288_),
    .A2(net413));
 sg13g2_o21ai_1 _22901_ (.B1(_05288_),
    .Y(_05289_),
    .A1(net645),
    .A2(_05285_));
 sg13g2_mux2_1 _22902_ (.A0(_05283_),
    .A1(_05289_),
    .S(net637),
    .X(_05290_));
 sg13g2_nor2_1 _22903_ (.A(net754),
    .B(_11984_),
    .Y(_05291_));
 sg13g2_a221oi_1 _22904_ (.B2(_05291_),
    .C1(_05050_),
    .B1(_05289_),
    .A1(net993),
    .Y(_05292_),
    .A2(_05283_));
 sg13g2_inv_1 _22905_ (.Y(_05293_),
    .A(_00284_));
 sg13g2_a22oi_1 _22906_ (.Y(_05294_),
    .B1(_05033_),
    .B2(_05293_),
    .A2(net511),
    .A1(\cpu.dcache.r_data[3][9] ));
 sg13g2_a22oi_1 _22907_ (.Y(_05295_),
    .B1(_09780_),
    .B2(\cpu.dcache.r_data[7][9] ),
    .A2(net455),
    .A1(\cpu.dcache.r_data[1][9] ));
 sg13g2_a22oi_1 _22908_ (.Y(_05296_),
    .B1(net453),
    .B2(\cpu.dcache.r_data[5][9] ),
    .A2(net463),
    .A1(\cpu.dcache.r_data[4][9] ));
 sg13g2_a22oi_1 _22909_ (.Y(_05297_),
    .B1(_04862_),
    .B2(\cpu.dcache.r_data[6][9] ),
    .A2(net454),
    .A1(\cpu.dcache.r_data[2][9] ));
 sg13g2_nand4_1 _22910_ (.B(_05295_),
    .C(_05296_),
    .A(_05294_),
    .Y(_05298_),
    .D(_05297_));
 sg13g2_a22oi_1 _22911_ (.Y(_05299_),
    .B1(net580),
    .B2(\cpu.dcache.r_data[6][25] ),
    .A2(net602),
    .A1(\cpu.dcache.r_data[2][25] ));
 sg13g2_a22oi_1 _22912_ (.Y(_05300_),
    .B1(_03079_),
    .B2(\cpu.dcache.r_data[5][25] ),
    .A2(_09778_),
    .A1(\cpu.dcache.r_data[7][25] ));
 sg13g2_a22oi_1 _22913_ (.Y(_05301_),
    .B1(net604),
    .B2(\cpu.dcache.r_data[4][25] ),
    .A2(_03075_),
    .A1(\cpu.dcache.r_data[3][25] ));
 sg13g2_nand3_1 _22914_ (.B(_05300_),
    .C(_05301_),
    .A(_05299_),
    .Y(_05302_));
 sg13g2_nand2_1 _22915_ (.Y(_05303_),
    .A(_00283_),
    .B(_09462_));
 sg13g2_o21ai_1 _22916_ (.B1(_05303_),
    .Y(_05304_),
    .A1(_09462_),
    .A2(_05302_));
 sg13g2_nor3_1 _22917_ (.A(\cpu.dcache.r_data[1][25] ),
    .B(net531),
    .C(_05302_),
    .Y(_05305_));
 sg13g2_a21o_1 _22918_ (.A2(_05304_),
    .A1(net531),
    .B1(_05305_),
    .X(_05306_));
 sg13g2_inv_1 _22919_ (.Y(_05307_),
    .A(_05306_));
 sg13g2_a221oi_1 _22920_ (.B2(_04844_),
    .C1(_04847_),
    .B1(_05307_),
    .A1(_09874_),
    .Y(_05308_),
    .A2(_05298_));
 sg13g2_o21ai_1 _22921_ (.B1(_04880_),
    .Y(_05309_),
    .A1(_05292_),
    .A2(_05308_));
 sg13g2_o21ai_1 _22922_ (.B1(_05309_),
    .Y(_05310_),
    .A1(_04880_),
    .A2(_05290_));
 sg13g2_nor3_1 _22923_ (.A(net994),
    .B(_00290_),
    .C(_04908_),
    .Y(_05311_));
 sg13g2_nor2b_1 _22924_ (.A(_00291_),
    .B_N(_04966_),
    .Y(_05312_));
 sg13g2_nand4_1 _22925_ (.B(_09776_),
    .C(net883),
    .A(net456),
    .Y(_05313_),
    .D(_04887_));
 sg13g2_buf_1 _22926_ (.A(_05313_),
    .X(_05314_));
 sg13g2_buf_2 _22927_ (.A(\cpu.gpio.r_src_io[4][1] ),
    .X(_05315_));
 sg13g2_nand2_1 _22928_ (.Y(_05316_),
    .A(_05315_),
    .B(net354));
 sg13g2_o21ai_1 _22929_ (.B1(_05316_),
    .Y(_05317_),
    .A1(_00287_),
    .A2(_05314_));
 sg13g2_inv_1 _22930_ (.Y(_05318_),
    .A(_00289_));
 sg13g2_a22oi_1 _22931_ (.Y(_05319_),
    .B1(net883),
    .B2(_05318_),
    .A2(net848),
    .A1(_09004_));
 sg13g2_nand2b_1 _22932_ (.Y(_05320_),
    .B(net356),
    .A_N(_05319_));
 sg13g2_o21ai_1 _22933_ (.B1(_05320_),
    .Y(_05321_),
    .A1(_00288_),
    .A2(_04979_));
 sg13g2_nor4_1 _22934_ (.A(_05311_),
    .B(_05312_),
    .C(_05317_),
    .D(_05321_),
    .Y(_05322_));
 sg13g2_a21oi_1 _22935_ (.A1(_09004_),
    .A2(_04996_),
    .Y(_05323_),
    .B1(_05089_));
 sg13g2_nand2b_1 _22936_ (.Y(_05324_),
    .B(\cpu.gpio.r_enable_in[1] ),
    .A_N(_05323_));
 sg13g2_a21oi_1 _22937_ (.A1(_05322_),
    .A2(_05324_),
    .Y(_05325_),
    .B1(_04999_));
 sg13g2_nor2_1 _22938_ (.A(_00286_),
    .B(_04940_),
    .Y(_05326_));
 sg13g2_a221oi_1 _22939_ (.B2(_11928_),
    .C1(_05326_),
    .B1(_04948_),
    .A1(_11927_),
    .Y(_05327_),
    .A2(net405));
 sg13g2_buf_1 _22940_ (.A(\cpu.spi.r_clk_count[2][1] ),
    .X(_05328_));
 sg13g2_nand2_1 _22941_ (.Y(_05329_),
    .A(\cpu.spi.r_timeout[1] ),
    .B(_05127_));
 sg13g2_o21ai_1 _22942_ (.B1(_05329_),
    .Y(_05330_),
    .A1(_00285_),
    .A2(_04959_));
 sg13g2_a221oi_1 _22943_ (.B2(_05328_),
    .C1(_05330_),
    .B1(_04956_),
    .A1(_11933_),
    .Y(_05331_),
    .A2(_04953_));
 sg13g2_o21ai_1 _22944_ (.B1(_05331_),
    .Y(_05332_),
    .A1(net857),
    .A2(_05327_));
 sg13g2_a21oi_1 _22945_ (.A1(_09072_),
    .A2(_04943_),
    .Y(_05333_),
    .B1(_05332_));
 sg13g2_nor2_1 _22946_ (.A(_09030_),
    .B(_05333_),
    .Y(_05334_));
 sg13g2_inv_1 _22947_ (.Y(_05335_),
    .A(\cpu.intr.r_timer_reload[17] ));
 sg13g2_a22oi_1 _22948_ (.Y(_05336_),
    .B1(net509),
    .B2(_09791_),
    .A2(net453),
    .A1(\cpu.intr.r_clock_cmp[17] ));
 sg13g2_o21ai_1 _22949_ (.B1(_05336_),
    .Y(_05337_),
    .A1(_05335_),
    .A2(_09616_));
 sg13g2_nand2_1 _22950_ (.Y(_05338_),
    .A(_09931_),
    .B(net528));
 sg13g2_buf_1 _22951_ (.A(\cpu.intr.r_clock_count[17] ),
    .X(_05339_));
 sg13g2_buf_1 _22952_ (.A(_05094_),
    .X(_05340_));
 sg13g2_a22oi_1 _22953_ (.Y(_05341_),
    .B1(net402),
    .B2(_08968_),
    .A2(net461),
    .A1(_05339_));
 sg13g2_a22oi_1 _22954_ (.Y(_05342_),
    .B1(_04948_),
    .B2(_09796_),
    .A2(_04910_),
    .A1(\cpu.intr.r_timer_reload[1] ));
 sg13g2_nand3_1 _22955_ (.B(_05341_),
    .C(_05342_),
    .A(_05338_),
    .Y(_05343_));
 sg13g2_a221oi_1 _22956_ (.B2(net755),
    .C1(_05343_),
    .B1(_05337_),
    .A1(\cpu.intr.r_clock_cmp[1] ),
    .Y(_05344_),
    .A2(_04918_));
 sg13g2_a21oi_1 _22957_ (.A1(_08968_),
    .A2(_05020_),
    .Y(_05345_),
    .B1(net289));
 sg13g2_nand2b_1 _22958_ (.Y(_05346_),
    .B(\cpu.intr.r_enable[1] ),
    .A_N(_05345_));
 sg13g2_a21oi_1 _22959_ (.A1(_05344_),
    .A2(_05346_),
    .Y(_05347_),
    .B1(net674));
 sg13g2_a22oi_1 _22960_ (.Y(_05348_),
    .B1(_04901_),
    .B2(\cpu.uart.r_div_value[9] ),
    .A2(net405),
    .A1(\cpu.uart.r_div_value[1] ));
 sg13g2_a22oi_1 _22961_ (.Y(_05349_),
    .B1(_04898_),
    .B2(_08973_),
    .A2(net404),
    .A1(\cpu.uart.r_r_invert ));
 sg13g2_nand2_1 _22962_ (.Y(_05350_),
    .A(_05348_),
    .B(_05349_));
 sg13g2_a21oi_1 _22963_ (.A1(\cpu.uart.r_in[1] ),
    .A2(_04886_),
    .Y(_05351_),
    .B1(_05350_));
 sg13g2_o21ai_1 _22964_ (.B1(_08181_),
    .Y(_05352_),
    .A1(_04884_),
    .A2(_05351_));
 sg13g2_nor4_1 _22965_ (.A(_05325_),
    .B(_05334_),
    .C(_05347_),
    .D(_05352_),
    .Y(_05353_));
 sg13g2_a21oi_1 _22966_ (.A1(net896),
    .A2(_05310_),
    .Y(_05354_),
    .B1(_05353_));
 sg13g2_mux2_1 _22967_ (.A0(_05354_),
    .A1(_03651_),
    .S(_05003_),
    .X(_05355_));
 sg13g2_nand3_1 _22968_ (.B(net288),
    .C(net111),
    .A(net1044),
    .Y(_05356_));
 sg13g2_o21ai_1 _22969_ (.B1(_05356_),
    .Y(_05357_),
    .A1(net111),
    .A2(_05355_));
 sg13g2_a21oi_1 _22970_ (.A1(_05259_),
    .A2(_05276_),
    .Y(_01012_),
    .B1(_05357_));
 sg13g2_nand3_1 _22971_ (.B(net688),
    .C(net630),
    .A(_08302_),
    .Y(_05358_));
 sg13g2_o21ai_1 _22972_ (.B1(_05358_),
    .Y(_05359_),
    .A1(net563),
    .A2(_04482_));
 sg13g2_o21ai_1 _22973_ (.B1(_05359_),
    .Y(_05360_),
    .A1(_11579_),
    .A2(_05273_));
 sg13g2_nor2_1 _22974_ (.A(net688),
    .B(net649),
    .Y(_05361_));
 sg13g2_o21ai_1 _22975_ (.B1(net691),
    .Y(_05362_),
    .A1(net288),
    .A2(_05361_));
 sg13g2_nor2b_1 _22976_ (.A(net966),
    .B_N(_09028_),
    .Y(_05363_));
 sg13g2_inv_1 _22977_ (.Y(_05364_),
    .A(_00100_));
 sg13g2_nor2_2 _22978_ (.A(net994),
    .B(_04908_),
    .Y(_05365_));
 sg13g2_inv_1 _22979_ (.Y(_05366_),
    .A(_00099_));
 sg13g2_a22oi_1 _22980_ (.Y(_05367_),
    .B1(_05365_),
    .B2(_05366_),
    .A2(_04966_),
    .A1(_05364_));
 sg13g2_buf_1 _22981_ (.A(\cpu.gpio.r_src_io[4][2] ),
    .X(_05368_));
 sg13g2_buf_1 _22982_ (.A(net952),
    .X(_05369_));
 sg13g2_nand2_1 _22983_ (.Y(_05370_),
    .A(_09000_),
    .B(net848));
 sg13g2_o21ai_1 _22984_ (.B1(_05370_),
    .Y(_05371_),
    .A1(net830),
    .A2(_00098_));
 sg13g2_nand2b_1 _22985_ (.Y(_05372_),
    .B(_04974_),
    .A_N(_00096_));
 sg13g2_o21ai_1 _22986_ (.B1(_05372_),
    .Y(_05373_),
    .A1(_00097_),
    .A2(_04979_));
 sg13g2_a221oi_1 _22987_ (.B2(_04924_),
    .C1(_05373_),
    .B1(_05371_),
    .A1(_05368_),
    .Y(_05374_),
    .A2(net354));
 sg13g2_a21oi_1 _22988_ (.A1(_09000_),
    .A2(_04996_),
    .Y(_05375_),
    .B1(_05089_));
 sg13g2_nand2b_1 _22989_ (.Y(_05376_),
    .B(\cpu.gpio.r_enable_in[2] ),
    .A_N(_05375_));
 sg13g2_nand3_1 _22990_ (.B(_05374_),
    .C(_05376_),
    .A(_05367_),
    .Y(_05377_));
 sg13g2_nand2_1 _22991_ (.Y(_05378_),
    .A(_09076_),
    .B(_04943_));
 sg13g2_buf_1 _22992_ (.A(\cpu.spi.r_clk_count[2][2] ),
    .X(_05379_));
 sg13g2_a22oi_1 _22993_ (.Y(_05380_),
    .B1(_04956_),
    .B2(_05379_),
    .A2(_04953_),
    .A1(_11915_));
 sg13g2_nor2_1 _22994_ (.A(_00094_),
    .B(_04959_),
    .Y(_05381_));
 sg13g2_a21oi_1 _22995_ (.A1(\cpu.spi.r_timeout[2] ),
    .A2(_05127_),
    .Y(_05382_),
    .B1(_05381_));
 sg13g2_inv_1 _22996_ (.Y(_05383_),
    .A(_00095_));
 sg13g2_a22oi_1 _22997_ (.Y(_05384_),
    .B1(_04901_),
    .B2(_05383_),
    .A2(net405),
    .A1(_11916_));
 sg13g2_o21ai_1 _22998_ (.B1(_05384_),
    .Y(_05385_),
    .A1(_00262_),
    .A2(_04908_));
 sg13g2_nand2_1 _22999_ (.Y(_05386_),
    .A(net848),
    .B(_05385_));
 sg13g2_nand4_1 _23000_ (.B(_05380_),
    .C(_05382_),
    .A(_05378_),
    .Y(_05387_),
    .D(_05386_));
 sg13g2_buf_1 _23001_ (.A(\cpu.intr.r_clock_count[18] ),
    .X(_05388_));
 sg13g2_nand2_1 _23002_ (.Y(_05389_),
    .A(_05388_),
    .B(net461));
 sg13g2_nand3_1 _23003_ (.B(\cpu.intr.r_timer_reload[18] ),
    .C(net530),
    .A(net881),
    .Y(_05390_));
 sg13g2_mux2_1 _23004_ (.A0(\cpu.intr.r_clock_cmp[2] ),
    .A1(\cpu.intr.r_clock_cmp[18] ),
    .S(net881),
    .X(_05391_));
 sg13g2_a22oi_1 _23005_ (.Y(_05392_),
    .B1(_05391_),
    .B2(net453),
    .A2(net402),
    .A1(_08969_));
 sg13g2_mux2_1 _23006_ (.A0(\cpu.intr.r_timer_count[2] ),
    .A1(_09790_),
    .S(net881),
    .X(_05393_));
 sg13g2_a22oi_1 _23007_ (.Y(_05394_),
    .B1(_05393_),
    .B2(net509),
    .A2(net356),
    .A1(_08970_));
 sg13g2_nand4_1 _23008_ (.B(_05390_),
    .C(_05392_),
    .A(_05389_),
    .Y(_05395_),
    .D(_05394_));
 sg13g2_a22oi_1 _23009_ (.Y(_05396_),
    .B1(net463),
    .B2(_09938_),
    .A2(net530),
    .A1(\cpu.intr.r_timer_reload[2] ));
 sg13g2_nand3_1 _23010_ (.B(_08970_),
    .C(_05020_),
    .A(_08969_),
    .Y(_05397_));
 sg13g2_o21ai_1 _23011_ (.B1(_05397_),
    .Y(_05398_),
    .A1(net755),
    .A2(_05396_));
 sg13g2_and2_1 _23012_ (.A(net966),
    .B(_09782_),
    .X(_05399_));
 sg13g2_buf_1 _23013_ (.A(_05399_),
    .X(_05400_));
 sg13g2_o21ai_1 _23014_ (.B1(_05400_),
    .Y(_05401_),
    .A1(_05395_),
    .A2(_05398_));
 sg13g2_nand2_1 _23015_ (.Y(_05402_),
    .A(\cpu.uart.r_div_value[2] ),
    .B(net357));
 sg13g2_a22oi_1 _23016_ (.Y(_05403_),
    .B1(_04886_),
    .B2(\cpu.uart.r_in[2] ),
    .A2(_04902_),
    .A1(_09766_));
 sg13g2_a21o_1 _23017_ (.A2(_05403_),
    .A1(_05402_),
    .B1(_04884_),
    .X(_05404_));
 sg13g2_nand3_1 _23018_ (.B(_05401_),
    .C(_05404_),
    .A(_08181_),
    .Y(_05405_));
 sg13g2_a221oi_1 _23019_ (.B2(_05133_),
    .C1(_05405_),
    .B1(_05387_),
    .A1(_05363_),
    .Y(_05406_),
    .A2(_05377_));
 sg13g2_mux2_1 _23020_ (.A0(\cpu.dcache.r_data[4][18] ),
    .A1(\cpu.dcache.r_data[6][18] ),
    .S(net532),
    .X(_05407_));
 sg13g2_a22oi_1 _23021_ (.Y(_05408_),
    .B1(_05407_),
    .B2(net768),
    .A2(_09367_),
    .A1(\cpu.dcache.r_data[5][18] ));
 sg13g2_a22oi_1 _23022_ (.Y(_05409_),
    .B1(net582),
    .B2(\cpu.dcache.r_data[3][18] ),
    .A2(net675),
    .A1(\cpu.dcache.r_data[7][18] ));
 sg13g2_o21ai_1 _23023_ (.B1(_05409_),
    .Y(_05410_),
    .A1(_00091_),
    .A2(net490));
 sg13g2_a221oi_1 _23024_ (.B2(\cpu.dcache.r_data[2][18] ),
    .C1(_05410_),
    .B1(net454),
    .A1(\cpu.dcache.r_data[1][18] ),
    .Y(_05411_),
    .A2(net455));
 sg13g2_o21ai_1 _23025_ (.B1(_05411_),
    .Y(_05412_),
    .A1(net645),
    .A2(_05408_));
 sg13g2_a22oi_1 _23026_ (.Y(_05413_),
    .B1(_05412_),
    .B2(_05063_),
    .A2(_05039_),
    .A1(_05050_));
 sg13g2_mux2_1 _23027_ (.A0(\cpu.dcache.r_data[4][2] ),
    .A1(\cpu.dcache.r_data[6][2] ),
    .S(_09104_),
    .X(_05414_));
 sg13g2_a22oi_1 _23028_ (.Y(_05415_),
    .B1(_05414_),
    .B2(net768),
    .A2(_09367_),
    .A1(\cpu.dcache.r_data[5][2] ));
 sg13g2_mux2_1 _23029_ (.A0(\cpu.dcache.r_data[2][2] ),
    .A1(\cpu.dcache.r_data[3][2] ),
    .S(net517),
    .X(_05416_));
 sg13g2_a22oi_1 _23030_ (.Y(_05417_),
    .B1(net890),
    .B2(_05416_),
    .A2(net675),
    .A1(\cpu.dcache.r_data[7][2] ));
 sg13g2_o21ai_1 _23031_ (.B1(_05417_),
    .Y(_05418_),
    .A1(net777),
    .A2(_05415_));
 sg13g2_mux2_1 _23032_ (.A0(\cpu.dcache.r_data[0][2] ),
    .A1(_05418_),
    .S(_09582_),
    .X(_05419_));
 sg13g2_or3_1 _23033_ (.A(\cpu.dcache.r_data[1][2] ),
    .B(net531),
    .C(_05418_),
    .X(_05420_));
 sg13g2_o21ai_1 _23034_ (.B1(_05420_),
    .Y(_05421_),
    .A1(_03070_),
    .A2(_05419_));
 sg13g2_inv_1 _23035_ (.Y(_05422_),
    .A(_04875_));
 sg13g2_nand2b_1 _23036_ (.Y(_05423_),
    .B(_05422_),
    .A_N(_05421_));
 sg13g2_o21ai_1 _23037_ (.B1(_05423_),
    .Y(_05424_),
    .A1(net993),
    .A2(_05413_));
 sg13g2_a21oi_1 _23038_ (.A1(_05071_),
    .A2(_05046_),
    .Y(_05425_),
    .B1(_05424_));
 sg13g2_and2_1 _23039_ (.A(net755),
    .B(_05412_),
    .X(_05426_));
 sg13g2_nor2_1 _23040_ (.A(_09777_),
    .B(_05421_),
    .Y(_05427_));
 sg13g2_nor3_1 _23041_ (.A(_04880_),
    .B(_05426_),
    .C(_05427_),
    .Y(_05428_));
 sg13g2_a21oi_1 _23042_ (.A1(_04880_),
    .A2(_05425_),
    .Y(_05429_),
    .B1(_05428_));
 sg13g2_nor2_1 _23043_ (.A(net967),
    .B(_05429_),
    .Y(_05430_));
 sg13g2_nor3_1 _23044_ (.A(_05003_),
    .B(_05406_),
    .C(_05430_),
    .Y(_05431_));
 sg13g2_a21oi_1 _23045_ (.A1(net410),
    .A2(net68),
    .Y(_05432_),
    .B1(_05431_));
 sg13g2_mux2_1 _23046_ (.A0(_05362_),
    .A1(_05432_),
    .S(_11518_),
    .X(_05433_));
 sg13g2_o21ai_1 _23047_ (.B1(_05433_),
    .Y(_01013_),
    .A1(_05010_),
    .A2(_05360_));
 sg13g2_buf_1 _23048_ (.A(\cpu.intr.r_clock_count[19] ),
    .X(_05434_));
 sg13g2_nand2_1 _23049_ (.Y(_05435_),
    .A(_05434_),
    .B(_09966_));
 sg13g2_mux2_1 _23050_ (.A0(\cpu.intr.r_timer_reload[3] ),
    .A1(\cpu.intr.r_timer_reload[19] ),
    .S(net755),
    .X(_05436_));
 sg13g2_a22oi_1 _23051_ (.Y(_05437_),
    .B1(_05436_),
    .B2(net530),
    .A2(net402),
    .A1(_08975_));
 sg13g2_a22oi_1 _23052_ (.Y(_05438_),
    .B1(net487),
    .B2(\cpu.intr.r_timer_count[3] ),
    .A2(net462),
    .A1(_09943_));
 sg13g2_a22oi_1 _23053_ (.Y(_05439_),
    .B1(net509),
    .B2(_09789_),
    .A2(net453),
    .A1(\cpu.intr.r_clock_cmp[19] ));
 sg13g2_inv_1 _23054_ (.Y(_05440_),
    .A(_05439_));
 sg13g2_a22oi_1 _23055_ (.Y(_05441_),
    .B1(_05440_),
    .B2(net637),
    .A2(_05024_),
    .A1(\cpu.intr.r_clock_cmp[3] ));
 sg13g2_nand4_1 _23056_ (.B(_05437_),
    .C(_05438_),
    .A(_05435_),
    .Y(_05442_),
    .D(_05441_));
 sg13g2_a21oi_1 _23057_ (.A1(_08975_),
    .A2(_05020_),
    .Y(_05443_),
    .B1(net289));
 sg13g2_nor2b_1 _23058_ (.A(_05443_),
    .B_N(\cpu.intr.r_enable[3] ),
    .Y(_05444_));
 sg13g2_o21ai_1 _23059_ (.B1(_05400_),
    .Y(_05445_),
    .A1(_05442_),
    .A2(_05444_));
 sg13g2_inv_1 _23060_ (.Y(_05446_),
    .A(_00107_));
 sg13g2_nand2_1 _23061_ (.Y(_05447_),
    .A(_08980_),
    .B(net848));
 sg13g2_o21ai_1 _23062_ (.B1(_05447_),
    .Y(_05448_),
    .A1(net830),
    .A2(_00108_));
 sg13g2_a22oi_1 _23063_ (.Y(_05449_),
    .B1(_05448_),
    .B2(net289),
    .A2(_04980_),
    .A1(_05446_));
 sg13g2_inv_1 _23064_ (.Y(_05450_),
    .A(_00109_));
 sg13g2_a22oi_1 _23065_ (.Y(_05451_),
    .B1(_05027_),
    .B2(_05450_),
    .A2(_09922_),
    .A1(\cpu.gpio.genblk1[3].srcs_o[0] ));
 sg13g2_nand2b_1 _23066_ (.Y(_05452_),
    .B(net830),
    .A_N(_05451_));
 sg13g2_buf_1 _23067_ (.A(\cpu.gpio.r_src_io[4][3] ),
    .X(_05453_));
 sg13g2_nor2_1 _23068_ (.A(_00106_),
    .B(_05314_),
    .Y(_05454_));
 sg13g2_a221oi_1 _23069_ (.B2(\cpu.gpio.r_enable_in[3] ),
    .C1(_05454_),
    .B1(_05089_),
    .A1(_05453_),
    .Y(_05455_),
    .A2(net354));
 sg13g2_nand2b_1 _23070_ (.Y(_05456_),
    .B(_04996_),
    .A_N(_08981_));
 sg13g2_nand4_1 _23071_ (.B(_05452_),
    .C(_05455_),
    .A(_05449_),
    .Y(_05457_),
    .D(_05456_));
 sg13g2_buf_1 _23072_ (.A(\cpu.spi.r_clk_count[2][3] ),
    .X(_05458_));
 sg13g2_buf_1 _23073_ (.A(_05110_),
    .X(_05459_));
 sg13g2_inv_1 _23074_ (.Y(_05460_),
    .A(_00105_));
 sg13g2_a22oi_1 _23075_ (.Y(_05461_),
    .B1(net287),
    .B2(_05460_),
    .A2(_04956_),
    .A1(_05458_));
 sg13g2_nor2_1 _23076_ (.A(_00104_),
    .B(_04959_),
    .Y(_05462_));
 sg13g2_a21oi_1 _23077_ (.A1(\cpu.spi.r_timeout[3] ),
    .A2(_05127_),
    .Y(_05463_),
    .B1(_05462_));
 sg13g2_nand2_1 _23078_ (.Y(_05464_),
    .A(_09070_),
    .B(_04943_));
 sg13g2_nand3_1 _23079_ (.B(_05463_),
    .C(_05464_),
    .A(_05461_),
    .Y(_05465_));
 sg13g2_and2_1 _23080_ (.A(\cpu.uart.r_div_value[11] ),
    .B(_04902_),
    .X(_05466_));
 sg13g2_a221oi_1 _23081_ (.B2(\cpu.uart.r_in[3] ),
    .C1(_05466_),
    .B1(_04886_),
    .A1(\cpu.uart.r_div_value[3] ),
    .Y(_05467_),
    .A2(net357));
 sg13g2_o21ai_1 _23082_ (.B1(net967),
    .Y(_05468_),
    .A1(_04884_),
    .A2(_05467_));
 sg13g2_a221oi_1 _23083_ (.B2(_05133_),
    .C1(_05468_),
    .B1(_05465_),
    .A1(_05363_),
    .Y(_05469_),
    .A2(_05457_));
 sg13g2_inv_1 _23084_ (.Y(_05470_),
    .A(_00101_));
 sg13g2_a22oi_1 _23085_ (.Y(_05471_),
    .B1(net486),
    .B2(_05470_),
    .A2(net463),
    .A1(\cpu.dcache.r_data[4][19] ));
 sg13g2_a22oi_1 _23086_ (.Y(_05472_),
    .B1(net489),
    .B2(\cpu.dcache.r_data[6][19] ),
    .A2(net455),
    .A1(\cpu.dcache.r_data[1][19] ));
 sg13g2_a22oi_1 _23087_ (.Y(_05473_),
    .B1(net511),
    .B2(\cpu.dcache.r_data[3][19] ),
    .A2(net599),
    .A1(\cpu.dcache.r_data[7][19] ));
 sg13g2_a22oi_1 _23088_ (.Y(_05474_),
    .B1(net453),
    .B2(\cpu.dcache.r_data[5][19] ),
    .A2(net454),
    .A1(\cpu.dcache.r_data[2][19] ));
 sg13g2_nand4_1 _23089_ (.B(_05472_),
    .C(_05473_),
    .A(_05471_),
    .Y(_05475_),
    .D(_05474_));
 sg13g2_buf_1 _23090_ (.A(_05475_),
    .X(_05476_));
 sg13g2_a22oi_1 _23091_ (.Y(_05477_),
    .B1(_05476_),
    .B2(_05063_),
    .A2(_05164_),
    .A1(_05050_));
 sg13g2_nand2_1 _23092_ (.Y(_05478_),
    .A(\cpu.dcache.r_data[2][3] ),
    .B(net512));
 sg13g2_a22oi_1 _23093_ (.Y(_05479_),
    .B1(net580),
    .B2(\cpu.dcache.r_data[6][3] ),
    .A2(net675),
    .A1(\cpu.dcache.r_data[7][3] ));
 sg13g2_a22oi_1 _23094_ (.Y(_05480_),
    .B1(net581),
    .B2(\cpu.dcache.r_data[5][3] ),
    .A2(net513),
    .A1(\cpu.dcache.r_data[1][3] ));
 sg13g2_a22oi_1 _23095_ (.Y(_05481_),
    .B1(net529),
    .B2(\cpu.dcache.r_data[4][3] ),
    .A2(net582),
    .A1(\cpu.dcache.r_data[3][3] ));
 sg13g2_nand4_1 _23096_ (.B(_05479_),
    .C(_05480_),
    .A(_05478_),
    .Y(_05482_),
    .D(_05481_));
 sg13g2_mux2_1 _23097_ (.A0(\cpu.dcache.r_data[0][3] ),
    .A1(_05482_),
    .S(_04855_),
    .X(_05483_));
 sg13g2_buf_1 _23098_ (.A(_05483_),
    .X(_05484_));
 sg13g2_a22oi_1 _23099_ (.Y(_05485_),
    .B1(_05484_),
    .B2(_05422_),
    .A2(_05170_),
    .A1(_05071_));
 sg13g2_o21ai_1 _23100_ (.B1(_05485_),
    .Y(_05486_),
    .A1(net993),
    .A2(_05477_));
 sg13g2_and2_1 _23101_ (.A(net637),
    .B(_05476_),
    .X(_05487_));
 sg13g2_a21oi_1 _23102_ (.A1(_04852_),
    .A2(_05484_),
    .Y(_05488_),
    .B1(_05487_));
 sg13g2_nand2_1 _23103_ (.Y(_05489_),
    .A(_04849_),
    .B(_05488_));
 sg13g2_o21ai_1 _23104_ (.B1(_05489_),
    .Y(_05490_),
    .A1(_05048_),
    .A2(_05486_));
 sg13g2_a221oi_1 _23105_ (.B2(net896),
    .C1(_05003_),
    .B1(_05490_),
    .A1(_05445_),
    .Y(_05491_),
    .A2(_05469_));
 sg13g2_a21oi_1 _23106_ (.A1(net464),
    .A2(net68),
    .Y(_05492_),
    .B1(_05491_));
 sg13g2_mux2_1 _23107_ (.A0(_04556_),
    .A1(_04521_),
    .S(net649),
    .X(_05493_));
 sg13g2_o21ai_1 _23108_ (.B1(_05493_),
    .Y(_05494_),
    .A1(_11606_),
    .A2(_05273_));
 sg13g2_a21oi_1 _23109_ (.A1(net563),
    .A2(_04488_),
    .Y(_05495_),
    .B1(net288));
 sg13g2_nor3_1 _23110_ (.A(net692),
    .B(net144),
    .C(_05495_),
    .Y(_05496_));
 sg13g2_a221oi_1 _23111_ (.B2(_05259_),
    .C1(_05496_),
    .B1(_05494_),
    .A1(net110),
    .Y(_01014_),
    .A2(_05492_));
 sg13g2_a21oi_1 _23112_ (.A1(_04811_),
    .A2(_04556_),
    .Y(_05497_),
    .B1(net373));
 sg13g2_nand4_1 _23113_ (.B(_04005_),
    .C(net630),
    .A(net1046),
    .Y(_05498_),
    .D(_04247_));
 sg13g2_o21ai_1 _23114_ (.B1(_05498_),
    .Y(_05499_),
    .A1(net1046),
    .A2(_05497_));
 sg13g2_or2_1 _23115_ (.X(_05500_),
    .B(_05499_),
    .A(net144));
 sg13g2_a21oi_1 _23116_ (.A1(_04844_),
    .A2(_05187_),
    .Y(_05501_),
    .B1(_05195_));
 sg13g2_mux2_1 _23117_ (.A0(\cpu.dcache.r_data[4][4] ),
    .A1(\cpu.dcache.r_data[6][4] ),
    .S(net532),
    .X(_05502_));
 sg13g2_a22oi_1 _23118_ (.Y(_05503_),
    .B1(_05502_),
    .B2(net644),
    .A2(_09379_),
    .A1(\cpu.dcache.r_data[7][4] ));
 sg13g2_a22oi_1 _23119_ (.Y(_05504_),
    .B1(net510),
    .B2(\cpu.dcache.r_data[5][4] ),
    .A2(net582),
    .A1(\cpu.dcache.r_data[3][4] ));
 sg13g2_o21ai_1 _23120_ (.B1(_05504_),
    .Y(_05505_),
    .A1(_00110_),
    .A2(net490));
 sg13g2_a221oi_1 _23121_ (.B2(\cpu.dcache.r_data[2][4] ),
    .C1(_05505_),
    .B1(net454),
    .A1(\cpu.dcache.r_data[1][4] ),
    .Y(_05506_),
    .A2(net413));
 sg13g2_o21ai_1 _23122_ (.B1(_05506_),
    .Y(_05507_),
    .A1(_11942_),
    .A2(_05503_));
 sg13g2_inv_1 _23123_ (.Y(_05508_),
    .A(_00111_));
 sg13g2_a22oi_1 _23124_ (.Y(_05509_),
    .B1(net486),
    .B2(_05508_),
    .A2(net530),
    .A1(\cpu.dcache.r_data[7][20] ));
 sg13g2_nand2_1 _23125_ (.Y(_05510_),
    .A(\cpu.dcache.r_data[5][20] ),
    .B(_03081_));
 sg13g2_a22oi_1 _23126_ (.Y(_05511_),
    .B1(net509),
    .B2(\cpu.dcache.r_data[6][20] ),
    .A2(net413),
    .A1(\cpu.dcache.r_data[1][20] ));
 sg13g2_mux2_1 _23127_ (.A0(\cpu.dcache.r_data[2][20] ),
    .A1(\cpu.dcache.r_data[3][20] ),
    .S(net456),
    .X(_05512_));
 sg13g2_a22oi_1 _23128_ (.Y(_05513_),
    .B1(_05512_),
    .B2(net890),
    .A2(net463),
    .A1(\cpu.dcache.r_data[4][20] ));
 sg13g2_nand4_1 _23129_ (.B(_05510_),
    .C(_05511_),
    .A(_05509_),
    .Y(_05514_),
    .D(_05513_));
 sg13g2_a221oi_1 _23130_ (.B2(_05291_),
    .C1(_05050_),
    .B1(_05514_),
    .A1(net993),
    .Y(_05515_),
    .A2(_05507_));
 sg13g2_a21o_1 _23131_ (.A2(_05501_),
    .A1(_05050_),
    .B1(_05515_),
    .X(_05516_));
 sg13g2_mux2_1 _23132_ (.A0(_05507_),
    .A1(_05514_),
    .S(_03650_),
    .X(_05517_));
 sg13g2_nand2_1 _23133_ (.Y(_05518_),
    .A(net564),
    .B(_05517_));
 sg13g2_o21ai_1 _23134_ (.B1(_05518_),
    .Y(_05519_),
    .A1(_05048_),
    .A2(_05516_));
 sg13g2_a22oi_1 _23135_ (.Y(_05520_),
    .B1(_04886_),
    .B2(\cpu.uart.r_in[4] ),
    .A2(net357),
    .A1(\cpu.uart.r_div_value[4] ));
 sg13g2_nor2_1 _23136_ (.A(_04884_),
    .B(_05520_),
    .Y(_05521_));
 sg13g2_buf_1 _23137_ (.A(\cpu.spi.r_clk_count[2][4] ),
    .X(_05522_));
 sg13g2_inv_1 _23138_ (.Y(_05523_),
    .A(_00115_));
 sg13g2_nand2_1 _23139_ (.Y(_05524_),
    .A(\cpu.spi.r_timeout[4] ),
    .B(_05127_));
 sg13g2_o21ai_1 _23140_ (.B1(_05524_),
    .Y(_05525_),
    .A1(_00114_),
    .A2(_04959_));
 sg13g2_a221oi_1 _23141_ (.B2(_05523_),
    .C1(_05525_),
    .B1(net287),
    .A1(_05522_),
    .Y(_05526_),
    .A2(_04956_));
 sg13g2_nand2_1 _23142_ (.Y(_05527_),
    .A(_09078_),
    .B(_04943_));
 sg13g2_a21oi_1 _23143_ (.A1(_05526_),
    .A2(_05527_),
    .Y(_05528_),
    .B1(_09030_));
 sg13g2_a22oi_1 _23144_ (.Y(_05529_),
    .B1(net356),
    .B2(_08996_),
    .A2(net405),
    .A1(_08995_));
 sg13g2_buf_2 _23145_ (.A(\cpu.gpio.r_src_o[7][0] ),
    .X(_05530_));
 sg13g2_buf_2 _23146_ (.A(\cpu.gpio.r_src_o[3][0] ),
    .X(_05531_));
 sg13g2_a221oi_1 _23147_ (.B2(_05531_),
    .C1(_03087_),
    .B1(net402),
    .A1(_05530_),
    .Y(_05532_),
    .A2(net404));
 sg13g2_a21oi_1 _23148_ (.A1(_03087_),
    .A2(_05529_),
    .Y(_05533_),
    .B1(_05532_));
 sg13g2_nand3_1 _23149_ (.B(\cpu.gpio.genblk2[4].srcs_io[0] ),
    .C(net461),
    .A(net830),
    .Y(_05534_));
 sg13g2_buf_2 _23150_ (.A(\cpu.gpio.r_src_io[5][0] ),
    .X(_05535_));
 sg13g2_nand2_1 _23151_ (.Y(_05536_),
    .A(_05535_),
    .B(net354));
 sg13g2_buf_2 _23152_ (.A(\cpu.gpio.r_src_io[7][0] ),
    .X(_05537_));
 sg13g2_buf_2 _23153_ (.A(\cpu.gpio.r_src_o[5][0] ),
    .X(_05538_));
 sg13g2_a22oi_1 _23154_ (.Y(_05539_),
    .B1(_04981_),
    .B2(_05538_),
    .A2(_04974_),
    .A1(_05537_));
 sg13g2_nand3_1 _23155_ (.B(_05536_),
    .C(_05539_),
    .A(_05534_),
    .Y(_05540_));
 sg13g2_buf_2 _23156_ (.A(\cpu.gpio.r_spi_miso_src[1][0] ),
    .X(_05541_));
 sg13g2_and2_1 _23157_ (.A(_09775_),
    .B(_05541_),
    .X(_05542_));
 sg13g2_a21oi_1 _23158_ (.A1(net879),
    .A2(net7),
    .Y(_05543_),
    .B1(_05542_));
 sg13g2_nor2_1 _23159_ (.A(_02697_),
    .B(_05543_),
    .Y(_05544_));
 sg13g2_a221oi_1 _23160_ (.B2(_08982_),
    .C1(_05544_),
    .B1(_04893_),
    .A1(\cpu.gpio.genblk1[4].srcs_o[0] ),
    .Y(_05545_),
    .A2(net528));
 sg13g2_and3_1 _23161_ (.X(_05546_),
    .A(_08982_),
    .B(net952),
    .C(_05094_));
 sg13g2_o21ai_1 _23162_ (.B1(\cpu.gpio.r_enable_io[4] ),
    .Y(_05547_),
    .A1(_05110_),
    .A2(_05546_));
 sg13g2_o21ai_1 _23163_ (.B1(_05547_),
    .Y(_05548_),
    .A1(net883),
    .A2(_05545_));
 sg13g2_nor3_1 _23164_ (.A(_05533_),
    .B(_05540_),
    .C(_05548_),
    .Y(_05549_));
 sg13g2_nand3_1 _23165_ (.B(_08996_),
    .C(_04996_),
    .A(_08995_),
    .Y(_05550_));
 sg13g2_a21oi_1 _23166_ (.A1(_05549_),
    .A2(_05550_),
    .Y(_05551_),
    .B1(_04999_));
 sg13g2_a21oi_1 _23167_ (.A1(\cpu.intr.r_clock_cmp[20] ),
    .A2(_05026_),
    .Y(_05552_),
    .B1(_05020_));
 sg13g2_mux2_1 _23168_ (.A0(\cpu.intr.r_timer_count[4] ),
    .A1(_09814_),
    .S(net881),
    .X(_05553_));
 sg13g2_a22oi_1 _23169_ (.Y(_05554_),
    .B1(_05553_),
    .B2(net509),
    .A2(net356),
    .A1(_09008_));
 sg13g2_buf_1 _23170_ (.A(\cpu.intr.r_clock_count[20] ),
    .X(_05555_));
 sg13g2_mux2_1 _23171_ (.A0(\cpu.intr.r_timer_reload[4] ),
    .A1(\cpu.intr.r_timer_reload[20] ),
    .S(net1025),
    .X(_05556_));
 sg13g2_a22oi_1 _23172_ (.Y(_05557_),
    .B1(_05556_),
    .B2(net599),
    .A2(_09964_),
    .A1(_05555_));
 sg13g2_a22oi_1 _23173_ (.Y(_05558_),
    .B1(_04918_),
    .B2(\cpu.intr.r_clock_cmp[4] ),
    .A2(_09921_),
    .A1(_09948_));
 sg13g2_and3_1 _23174_ (.X(_05559_),
    .A(_05554_),
    .B(_05557_),
    .C(_05558_));
 sg13g2_nand2_1 _23175_ (.Y(_05560_),
    .A(_05552_),
    .B(_05559_));
 sg13g2_nor2_1 _23176_ (.A(net402),
    .B(_05560_),
    .Y(_05561_));
 sg13g2_nor3_1 _23177_ (.A(_09008_),
    .B(net646),
    .C(_04926_),
    .Y(_05562_));
 sg13g2_a21oi_1 _23178_ (.A1(_05552_),
    .A2(_05559_),
    .Y(_05563_),
    .B1(_05020_));
 sg13g2_nor3_1 _23179_ (.A(_10105_),
    .B(_10106_),
    .C(_05563_),
    .Y(_05564_));
 sg13g2_nor4_1 _23180_ (.A(net674),
    .B(_05561_),
    .C(_05562_),
    .D(_05564_),
    .Y(_05565_));
 sg13g2_nor4_1 _23181_ (.A(_05521_),
    .B(_05528_),
    .C(_05551_),
    .D(_05565_),
    .Y(_05566_));
 sg13g2_nand2_1 _23182_ (.Y(_05567_),
    .A(net967),
    .B(_05566_));
 sg13g2_o21ai_1 _23183_ (.B1(_05567_),
    .Y(_05568_),
    .A1(net967),
    .A2(_05519_));
 sg13g2_nand2_1 _23184_ (.Y(_05569_),
    .A(net448),
    .B(_05003_));
 sg13g2_o21ai_1 _23185_ (.B1(_05569_),
    .Y(_05570_),
    .A1(net68),
    .A2(_05568_));
 sg13g2_nand2_1 _23186_ (.Y(_05571_),
    .A(_05228_),
    .B(_05570_));
 sg13g2_a22oi_1 _23187_ (.Y(_01015_),
    .B1(_05500_),
    .B2(_05571_),
    .A2(_05150_),
    .A1(_04555_));
 sg13g2_nand2_1 _23188_ (.Y(_05572_),
    .A(net630),
    .B(_04563_));
 sg13g2_o21ai_1 _23189_ (.B1(_05572_),
    .Y(_05573_),
    .A1(net630),
    .A2(_04592_));
 sg13g2_o21ai_1 _23190_ (.B1(_05573_),
    .Y(_05574_),
    .A1(_11639_),
    .A2(_05273_));
 sg13g2_a22oi_1 _23191_ (.Y(_05575_),
    .B1(net580),
    .B2(\cpu.dcache.r_data[6][21] ),
    .A2(net582),
    .A1(\cpu.dcache.r_data[3][21] ));
 sg13g2_a22oi_1 _23192_ (.Y(_05576_),
    .B1(net581),
    .B2(\cpu.dcache.r_data[5][21] ),
    .A2(net675),
    .A1(\cpu.dcache.r_data[7][21] ));
 sg13g2_a22oi_1 _23193_ (.Y(_05577_),
    .B1(net529),
    .B2(\cpu.dcache.r_data[4][21] ),
    .A2(net602),
    .A1(\cpu.dcache.r_data[2][21] ));
 sg13g2_nand3_1 _23194_ (.B(_05576_),
    .C(_05577_),
    .A(_05575_),
    .Y(_05578_));
 sg13g2_nand2_1 _23195_ (.Y(_05579_),
    .A(_00117_),
    .B(net758));
 sg13g2_o21ai_1 _23196_ (.B1(_05579_),
    .Y(_05580_),
    .A1(net758),
    .A2(_05578_));
 sg13g2_o21ai_1 _23197_ (.B1(net413),
    .Y(_05581_),
    .A1(\cpu.dcache.r_data[1][21] ),
    .A2(_05578_));
 sg13g2_o21ai_1 _23198_ (.B1(_05581_),
    .Y(_05582_),
    .A1(net413),
    .A2(_05580_));
 sg13g2_and2_1 _23199_ (.A(_09777_),
    .B(_05582_),
    .X(_05583_));
 sg13g2_mux2_1 _23200_ (.A0(\cpu.dcache.r_data[5][5] ),
    .A1(\cpu.dcache.r_data[7][5] ),
    .S(_09105_),
    .X(_05584_));
 sg13g2_a22oi_1 _23201_ (.Y(_05585_),
    .B1(_05584_),
    .B2(_12461_),
    .A2(net680),
    .A1(\cpu.dcache.r_data[6][5] ));
 sg13g2_inv_1 _23202_ (.Y(_05586_),
    .A(_00116_));
 sg13g2_mux2_1 _23203_ (.A0(\cpu.dcache.r_data[1][5] ),
    .A1(\cpu.dcache.r_data[3][5] ),
    .S(net532),
    .X(_05587_));
 sg13g2_a22oi_1 _23204_ (.Y(_05588_),
    .B1(_05587_),
    .B2(net517),
    .A2(net680),
    .A1(\cpu.dcache.r_data[2][5] ));
 sg13g2_nor2_1 _23205_ (.A(_09305_),
    .B(_05588_),
    .Y(_05589_));
 sg13g2_a221oi_1 _23206_ (.B2(_05586_),
    .C1(_05589_),
    .B1(net486),
    .A1(\cpu.dcache.r_data[4][5] ),
    .Y(_05590_),
    .A2(_09916_));
 sg13g2_o21ai_1 _23207_ (.B1(_05590_),
    .Y(_05591_),
    .A1(_11942_),
    .A2(_05585_));
 sg13g2_and2_1 _23208_ (.A(net993),
    .B(_05591_),
    .X(_05592_));
 sg13g2_a21oi_1 _23209_ (.A1(_04844_),
    .A2(_05583_),
    .Y(_05593_),
    .B1(_05592_));
 sg13g2_a221oi_1 _23210_ (.B2(_09874_),
    .C1(_04847_),
    .B1(_05222_),
    .A1(_04844_),
    .Y(_05594_),
    .A2(_05216_));
 sg13g2_a21oi_1 _23211_ (.A1(_04847_),
    .A2(_05593_),
    .Y(_05595_),
    .B1(_05594_));
 sg13g2_a21oi_1 _23212_ (.A1(net631),
    .A2(_05591_),
    .Y(_05596_),
    .B1(_05583_));
 sg13g2_nand2_1 _23213_ (.Y(_05597_),
    .A(net564),
    .B(_05596_));
 sg13g2_o21ai_1 _23214_ (.B1(_05597_),
    .Y(_05598_),
    .A1(net485),
    .A2(_05595_));
 sg13g2_nand3_1 _23215_ (.B(_09002_),
    .C(_04996_),
    .A(_09001_),
    .Y(_05599_));
 sg13g2_nor3_1 _23216_ (.A(net754),
    .B(_00126_),
    .C(_02697_),
    .Y(_05600_));
 sg13g2_a22oi_1 _23217_ (.Y(_05601_),
    .B1(net453),
    .B2(net8),
    .A2(net463),
    .A1(\cpu.gpio.genblk1[5].srcs_o[0] ));
 sg13g2_a21oi_1 _23218_ (.A1(_08984_),
    .A2(_05094_),
    .Y(_05602_),
    .B1(net404));
 sg13g2_nand2b_1 _23219_ (.Y(_05603_),
    .B(_08985_),
    .A_N(_05602_));
 sg13g2_o21ai_1 _23220_ (.B1(_05603_),
    .Y(_05604_),
    .A1(net755),
    .A2(_05601_));
 sg13g2_or2_1 _23221_ (.X(_05605_),
    .B(_05604_),
    .A(_05600_));
 sg13g2_nand2_1 _23222_ (.Y(_05606_),
    .A(_11937_),
    .B(_05094_));
 sg13g2_buf_2 _23223_ (.A(\cpu.gpio.r_src_io[5][1] ),
    .X(_05607_));
 sg13g2_nand2_1 _23224_ (.Y(_05608_),
    .A(_05607_),
    .B(net354));
 sg13g2_o21ai_1 _23225_ (.B1(_05608_),
    .Y(_05609_),
    .A1(_00123_),
    .A2(_04979_));
 sg13g2_nand3_1 _23226_ (.B(\cpu.gpio.genblk2[5].srcs_io[0] ),
    .C(_09965_),
    .A(net830),
    .Y(_05610_));
 sg13g2_o21ai_1 _23227_ (.B1(_05610_),
    .Y(_05611_),
    .A1(_00122_),
    .A2(_05314_));
 sg13g2_a22oi_1 _23228_ (.Y(_05612_),
    .B1(_04901_),
    .B2(_08984_),
    .A2(net356),
    .A1(_09002_));
 sg13g2_inv_1 _23229_ (.Y(_05613_),
    .A(_00124_));
 sg13g2_a22oi_1 _23230_ (.Y(_05614_),
    .B1(_05089_),
    .B2(_09001_),
    .A2(_04981_),
    .A1(_05613_));
 sg13g2_o21ai_1 _23231_ (.B1(_05614_),
    .Y(_05615_),
    .A1(_11937_),
    .A2(_05612_));
 sg13g2_nor3_1 _23232_ (.A(_05609_),
    .B(_05611_),
    .C(_05615_),
    .Y(_05616_));
 sg13g2_o21ai_1 _23233_ (.B1(_05616_),
    .Y(_05617_),
    .A1(_00125_),
    .A2(_05606_));
 sg13g2_a21oi_1 _23234_ (.A1(_05369_),
    .A2(_05605_),
    .Y(_05618_),
    .B1(_05617_));
 sg13g2_a21o_1 _23235_ (.A2(_05618_),
    .A1(_05599_),
    .B1(_04999_),
    .X(_05619_));
 sg13g2_buf_1 _23236_ (.A(\cpu.spi.r_clk_count[2][5] ),
    .X(_05620_));
 sg13g2_inv_1 _23237_ (.Y(_05621_),
    .A(_00121_));
 sg13g2_a22oi_1 _23238_ (.Y(_05622_),
    .B1(net287),
    .B2(_05621_),
    .A2(_04956_),
    .A1(_05620_));
 sg13g2_nor2_1 _23239_ (.A(_00120_),
    .B(_04959_),
    .Y(_05623_));
 sg13g2_a21oi_1 _23240_ (.A1(\cpu.spi.r_timeout[5] ),
    .A2(_05127_),
    .Y(_05624_),
    .B1(_05623_));
 sg13g2_nand2_1 _23241_ (.Y(_05625_),
    .A(_09077_),
    .B(_04943_));
 sg13g2_nand3_1 _23242_ (.B(_05624_),
    .C(_05625_),
    .A(_05622_),
    .Y(_05626_));
 sg13g2_and2_1 _23243_ (.A(net881),
    .B(\cpu.intr.r_clock_cmp[21] ),
    .X(_05627_));
 sg13g2_a21oi_1 _23244_ (.A1(net879),
    .A2(\cpu.intr.r_clock_cmp[5] ),
    .Y(_05628_),
    .B1(_05627_));
 sg13g2_buf_1 _23245_ (.A(\cpu.intr.r_clock_count[21] ),
    .X(_05629_));
 sg13g2_a22oi_1 _23246_ (.Y(_05630_),
    .B1(net402),
    .B2(_08976_),
    .A2(net461),
    .A1(_05629_));
 sg13g2_o21ai_1 _23247_ (.B1(_05630_),
    .Y(_05631_),
    .A1(_02697_),
    .A2(_05628_));
 sg13g2_a221oi_1 _23248_ (.B2(\cpu.intr.r_timer_count[5] ),
    .C1(_05631_),
    .B1(_05030_),
    .A1(_09953_),
    .Y(_05632_),
    .A2(net462));
 sg13g2_a22oi_1 _23249_ (.Y(_05633_),
    .B1(net509),
    .B2(_09813_),
    .A2(net530),
    .A1(\cpu.intr.r_timer_reload[21] ));
 sg13g2_inv_1 _23250_ (.Y(_05634_),
    .A(_05633_));
 sg13g2_a22oi_1 _23251_ (.Y(_05635_),
    .B1(_05634_),
    .B2(net637),
    .A2(_05023_),
    .A1(\cpu.intr.r_timer_reload[5] ));
 sg13g2_a21oi_1 _23252_ (.A1(_08976_),
    .A2(_05020_),
    .Y(_05636_),
    .B1(net289));
 sg13g2_nand2b_1 _23253_ (.Y(_05637_),
    .B(\cpu.intr.r_enable[5] ),
    .A_N(_05636_));
 sg13g2_nand3_1 _23254_ (.B(_05635_),
    .C(_05637_),
    .A(_05632_),
    .Y(_05638_));
 sg13g2_a22oi_1 _23255_ (.Y(_05639_),
    .B1(_04886_),
    .B2(\cpu.uart.r_in[5] ),
    .A2(net357),
    .A1(\cpu.uart.r_div_value[5] ));
 sg13g2_o21ai_1 _23256_ (.B1(net967),
    .Y(_05640_),
    .A1(_04884_),
    .A2(_05639_));
 sg13g2_a221oi_1 _23257_ (.B2(_05400_),
    .C1(_05640_),
    .B1(_05638_),
    .A1(_05133_),
    .Y(_05641_),
    .A2(_05626_));
 sg13g2_a221oi_1 _23258_ (.B2(_05641_),
    .C1(_05003_),
    .B1(_05619_),
    .A1(net896),
    .Y(_05642_),
    .A2(_05598_));
 sg13g2_a21oi_1 _23259_ (.A1(net640),
    .A2(_05004_),
    .Y(_05643_),
    .B1(_05642_));
 sg13g2_nor3_1 _23260_ (.A(net957),
    .B(net214),
    .C(_11518_),
    .Y(_05644_));
 sg13g2_a221oi_1 _23261_ (.B2(net110),
    .C1(_05644_),
    .B1(_05643_),
    .A1(_05259_),
    .Y(_01016_),
    .A2(_05574_));
 sg13g2_inv_1 _23262_ (.Y(_05645_),
    .A(_00128_));
 sg13g2_a22oi_1 _23263_ (.Y(_05646_),
    .B1(net486),
    .B2(_05645_),
    .A2(net511),
    .A1(\cpu.dcache.r_data[3][22] ));
 sg13g2_a22oi_1 _23264_ (.Y(_05647_),
    .B1(net599),
    .B2(\cpu.dcache.r_data[7][22] ),
    .A2(net513),
    .A1(\cpu.dcache.r_data[1][22] ));
 sg13g2_a22oi_1 _23265_ (.Y(_05648_),
    .B1(net489),
    .B2(\cpu.dcache.r_data[6][22] ),
    .A2(net529),
    .A1(\cpu.dcache.r_data[4][22] ));
 sg13g2_a22oi_1 _23266_ (.Y(_05649_),
    .B1(net510),
    .B2(\cpu.dcache.r_data[5][22] ),
    .A2(net512),
    .A1(\cpu.dcache.r_data[2][22] ));
 sg13g2_nand4_1 _23267_ (.B(_05647_),
    .C(_05648_),
    .A(_05646_),
    .Y(_05650_),
    .D(_05649_));
 sg13g2_buf_1 _23268_ (.A(_05650_),
    .X(_05651_));
 sg13g2_inv_1 _23269_ (.Y(_05652_),
    .A(_00127_));
 sg13g2_a22oi_1 _23270_ (.Y(_05653_),
    .B1(net603),
    .B2(_05652_),
    .A2(net529),
    .A1(\cpu.dcache.r_data[4][6] ));
 sg13g2_a22oi_1 _23271_ (.Y(_05654_),
    .B1(net489),
    .B2(\cpu.dcache.r_data[6][6] ),
    .A2(net513),
    .A1(\cpu.dcache.r_data[1][6] ));
 sg13g2_a22oi_1 _23272_ (.Y(_05655_),
    .B1(net511),
    .B2(\cpu.dcache.r_data[3][6] ),
    .A2(net599),
    .A1(\cpu.dcache.r_data[7][6] ));
 sg13g2_a22oi_1 _23273_ (.Y(_05656_),
    .B1(net510),
    .B2(\cpu.dcache.r_data[5][6] ),
    .A2(net512),
    .A1(\cpu.dcache.r_data[2][6] ));
 sg13g2_and4_1 _23274_ (.A(_05653_),
    .B(_05654_),
    .C(_05655_),
    .D(_05656_),
    .X(_05657_));
 sg13g2_buf_1 _23275_ (.A(_05657_),
    .X(_05658_));
 sg13g2_nand2_1 _23276_ (.Y(_05659_),
    .A(net631),
    .B(_05658_));
 sg13g2_o21ai_1 _23277_ (.B1(_05659_),
    .Y(_05660_),
    .A1(net631),
    .A2(_05651_));
 sg13g2_a22oi_1 _23278_ (.Y(_05661_),
    .B1(_05651_),
    .B2(_05063_),
    .A2(_05239_),
    .A1(_05050_));
 sg13g2_nor2_1 _23279_ (.A(_04875_),
    .B(_05658_),
    .Y(_05662_));
 sg13g2_a21oi_1 _23280_ (.A1(_05071_),
    .A2(_05248_),
    .Y(_05663_),
    .B1(_05662_));
 sg13g2_o21ai_1 _23281_ (.B1(_05663_),
    .Y(_05664_),
    .A1(net993),
    .A2(_05661_));
 sg13g2_nor2_1 _23282_ (.A(net564),
    .B(_05664_),
    .Y(_05665_));
 sg13g2_a21oi_1 _23283_ (.A1(net564),
    .A2(_05660_),
    .Y(_05666_),
    .B1(_05665_));
 sg13g2_a22oi_1 _23284_ (.Y(_05667_),
    .B1(_04886_),
    .B2(\cpu.uart.r_in[6] ),
    .A2(net357),
    .A1(\cpu.uart.r_div_value[6] ));
 sg13g2_buf_2 _23285_ (.A(\cpu.intr.r_clock_count[22] ),
    .X(_05668_));
 sg13g2_mux2_1 _23286_ (.A0(\cpu.intr.r_clock_cmp[6] ),
    .A1(\cpu.intr.r_clock_cmp[22] ),
    .S(net881),
    .X(_05669_));
 sg13g2_a22oi_1 _23287_ (.Y(_05670_),
    .B1(_05669_),
    .B2(net453),
    .A2(net461),
    .A1(_05668_));
 sg13g2_nand2_1 _23288_ (.Y(_05671_),
    .A(_09959_),
    .B(net528));
 sg13g2_nand2_1 _23289_ (.Y(_05672_),
    .A(_05670_),
    .B(_05671_));
 sg13g2_a22oi_1 _23290_ (.Y(_05673_),
    .B1(net509),
    .B2(_09816_),
    .A2(net530),
    .A1(\cpu.intr.r_timer_reload[22] ));
 sg13g2_a22oi_1 _23291_ (.Y(_05674_),
    .B1(_04948_),
    .B2(\cpu.intr.r_timer_count[6] ),
    .A2(_04910_),
    .A1(\cpu.intr.r_timer_reload[6] ));
 sg13g2_o21ai_1 _23292_ (.B1(_05674_),
    .Y(_05675_),
    .A1(net754),
    .A2(_05673_));
 sg13g2_o21ai_1 _23293_ (.B1(_05114_),
    .Y(_05676_),
    .A1(_05672_),
    .A2(_05675_));
 sg13g2_o21ai_1 _23294_ (.B1(_05676_),
    .Y(_05677_),
    .A1(_04884_),
    .A2(_05667_));
 sg13g2_buf_1 _23295_ (.A(\cpu.spi.r_clk_count[2][6] ),
    .X(_05678_));
 sg13g2_inv_1 _23296_ (.Y(_05679_),
    .A(_00132_));
 sg13g2_nand2_1 _23297_ (.Y(_05680_),
    .A(\cpu.spi.r_timeout[6] ),
    .B(_05127_));
 sg13g2_o21ai_1 _23298_ (.B1(_05680_),
    .Y(_05681_),
    .A1(_00131_),
    .A2(_04959_));
 sg13g2_a221oi_1 _23299_ (.B2(_05679_),
    .C1(_05681_),
    .B1(net287),
    .A1(_05678_),
    .Y(_05682_),
    .A2(_04956_));
 sg13g2_nand2_1 _23300_ (.Y(_05683_),
    .A(_09071_),
    .B(_04943_));
 sg13g2_a21oi_1 _23301_ (.A1(_05682_),
    .A2(_05683_),
    .Y(_05684_),
    .B1(_09030_));
 sg13g2_nand3_1 _23302_ (.B(net952),
    .C(net402),
    .A(_09005_),
    .Y(_05685_));
 sg13g2_nand2b_1 _23303_ (.Y(_05686_),
    .B(_05685_),
    .A_N(net287));
 sg13g2_nand2b_1 _23304_ (.Y(_05687_),
    .B(_05026_),
    .A_N(_00137_));
 sg13g2_a22oi_1 _23305_ (.Y(_05688_),
    .B1(_04893_),
    .B2(_09005_),
    .A2(_09965_),
    .A1(\cpu.gpio.genblk2[6].srcs_io[0] ));
 sg13g2_a22oi_1 _23306_ (.Y(_05689_),
    .B1(_04918_),
    .B2(net9),
    .A2(_09922_),
    .A1(\cpu.gpio.genblk1[6].srcs_o[0] ));
 sg13g2_nand3_1 _23307_ (.B(_05688_),
    .C(_05689_),
    .A(_05687_),
    .Y(_05690_));
 sg13g2_nand2b_1 _23308_ (.Y(_05691_),
    .B(_04974_),
    .A_N(_00133_));
 sg13g2_or2_1 _23309_ (.X(_05692_),
    .B(_05606_),
    .A(_00136_));
 sg13g2_buf_1 _23310_ (.A(\cpu.gpio.r_src_io[5][2] ),
    .X(_05693_));
 sg13g2_a22oi_1 _23311_ (.Y(_05694_),
    .B1(_05089_),
    .B2(_08997_),
    .A2(_04973_),
    .A1(_05693_));
 sg13g2_inv_1 _23312_ (.Y(_05695_),
    .A(_00134_));
 sg13g2_nand2_1 _23313_ (.Y(_05696_),
    .A(_08998_),
    .B(_10473_));
 sg13g2_o21ai_1 _23314_ (.B1(_05696_),
    .Y(_05697_),
    .A1(net952),
    .A2(_00135_));
 sg13g2_a22oi_1 _23315_ (.Y(_05698_),
    .B1(_05697_),
    .B2(net356),
    .A2(_04980_),
    .A1(_05695_));
 sg13g2_nand4_1 _23316_ (.B(_05692_),
    .C(_05694_),
    .A(_05691_),
    .Y(_05699_),
    .D(_05698_));
 sg13g2_a221oi_1 _23317_ (.B2(net830),
    .C1(_05699_),
    .B1(_05690_),
    .A1(\cpu.gpio.r_enable_io[6] ),
    .Y(_05700_),
    .A2(_05686_));
 sg13g2_nand3_1 _23318_ (.B(_08998_),
    .C(_04996_),
    .A(_08997_),
    .Y(_05701_));
 sg13g2_a21oi_1 _23319_ (.A1(_05700_),
    .A2(_05701_),
    .Y(_05702_),
    .B1(_04999_));
 sg13g2_or4_1 _23320_ (.A(net896),
    .B(_05677_),
    .C(_05684_),
    .D(_05702_),
    .X(_05703_));
 sg13g2_o21ai_1 _23321_ (.B1(_05703_),
    .Y(_05704_),
    .A1(net967),
    .A2(_05666_));
 sg13g2_nor2_1 _23322_ (.A(net68),
    .B(_05704_),
    .Y(_05705_));
 sg13g2_a21oi_1 _23323_ (.A1(net966),
    .A2(net68),
    .Y(_05706_),
    .B1(_05705_));
 sg13g2_mux2_1 _23324_ (.A0(_04595_),
    .A1(_04624_),
    .S(net649),
    .X(_05707_));
 sg13g2_o21ai_1 _23325_ (.B1(_05707_),
    .Y(_05708_),
    .A1(_11663_),
    .A2(_05273_));
 sg13g2_nor3_1 _23326_ (.A(\cpu.ex.pc[6] ),
    .B(net214),
    .C(net144),
    .Y(_05709_));
 sg13g2_a221oi_1 _23327_ (.B2(_05259_),
    .C1(_05709_),
    .B1(_05708_),
    .A1(_05228_),
    .Y(_01017_),
    .A2(_05706_));
 sg13g2_nand2_1 _23328_ (.Y(_05710_),
    .A(_05013_),
    .B(_04657_));
 sg13g2_o21ai_1 _23329_ (.B1(_05710_),
    .Y(_05711_),
    .A1(_05013_),
    .A2(_04654_));
 sg13g2_o21ai_1 _23330_ (.B1(_05711_),
    .Y(_05712_),
    .A1(_04627_),
    .A2(_05273_));
 sg13g2_nor2_1 _23331_ (.A(net956),
    .B(net214),
    .Y(_05713_));
 sg13g2_nor2b_1 _23332_ (.A(net68),
    .B_N(_05139_),
    .Y(_05714_));
 sg13g2_a221oi_1 _23333_ (.B2(net965),
    .C1(_05714_),
    .B1(_05004_),
    .A1(net783),
    .Y(_05715_),
    .A2(_11513_));
 sg13g2_a221oi_1 _23334_ (.B2(_05147_),
    .C1(_05715_),
    .B1(_05713_),
    .A1(_05259_),
    .Y(_01018_),
    .A2(_05712_));
 sg13g2_or3_1 _23335_ (.A(net288),
    .B(_11507_),
    .C(_04695_),
    .X(_05716_));
 sg13g2_o21ai_1 _23336_ (.B1(_05716_),
    .Y(_05717_),
    .A1(net955),
    .A2(_04005_));
 sg13g2_a22oi_1 _23337_ (.Y(_05718_),
    .B1(net444),
    .B2(\cpu.intr.r_clock_cmp[24] ),
    .A2(net488),
    .A1(\cpu.intr.r_timer_reload[8] ));
 sg13g2_a22oi_1 _23338_ (.Y(_05719_),
    .B1(net487),
    .B2(\cpu.intr.r_timer_count[8] ),
    .A2(net462),
    .A1(_09976_));
 sg13g2_buf_1 _23339_ (.A(\cpu.intr.r_clock_count[24] ),
    .X(_05720_));
 sg13g2_a22oi_1 _23340_ (.Y(_05721_),
    .B1(net403),
    .B2(\cpu.intr.r_clock_cmp[8] ),
    .A2(net423),
    .A1(_05720_));
 sg13g2_nand3_1 _23341_ (.B(_05719_),
    .C(_05721_),
    .A(_05718_),
    .Y(_05722_));
 sg13g2_mux2_1 _23342_ (.A0(_04859_),
    .A1(_04866_),
    .S(_03650_),
    .X(_05723_));
 sg13g2_a22oi_1 _23343_ (.Y(_05724_),
    .B1(_05723_),
    .B2(net485),
    .A2(_05722_),
    .A1(_05022_));
 sg13g2_o21ai_1 _23344_ (.B1(_05141_),
    .Y(_05725_),
    .A1(net832),
    .A2(_05724_));
 sg13g2_nand2b_1 _23345_ (.Y(_05726_),
    .B(_05144_),
    .A_N(net1037));
 sg13g2_o21ai_1 _23346_ (.B1(_05726_),
    .Y(_05727_),
    .A1(_05144_),
    .A2(_05725_));
 sg13g2_a221oi_1 _23347_ (.B2(_05147_),
    .C1(_05727_),
    .B1(_05717_),
    .A1(_04692_),
    .Y(_01019_),
    .A2(_05150_));
 sg13g2_a21o_1 _23348_ (.A2(_04729_),
    .A1(_04706_),
    .B1(net630),
    .X(_05728_));
 sg13g2_nand2b_1 _23349_ (.Y(_05729_),
    .B(_05014_),
    .A_N(_04732_));
 sg13g2_o21ai_1 _23350_ (.B1(_05729_),
    .Y(_05730_),
    .A1(_04730_),
    .A2(_05728_));
 sg13g2_a22oi_1 _23351_ (.Y(_05731_),
    .B1(net444),
    .B2(\cpu.intr.r_clock_cmp[25] ),
    .A2(net488),
    .A1(\cpu.intr.r_timer_reload[9] ));
 sg13g2_a22oi_1 _23352_ (.Y(_05732_),
    .B1(net487),
    .B2(\cpu.intr.r_timer_count[9] ),
    .A2(net528),
    .A1(_09982_));
 sg13g2_buf_2 _23353_ (.A(\cpu.intr.r_clock_count[25] ),
    .X(_05733_));
 sg13g2_a22oi_1 _23354_ (.Y(_05734_),
    .B1(net403),
    .B2(\cpu.intr.r_clock_cmp[9] ),
    .A2(net423),
    .A1(_05733_));
 sg13g2_nand3_1 _23355_ (.B(_05732_),
    .C(_05734_),
    .A(_05731_),
    .Y(_05735_));
 sg13g2_nand2_1 _23356_ (.Y(_05736_),
    .A(net631),
    .B(_05298_));
 sg13g2_o21ai_1 _23357_ (.B1(_05736_),
    .Y(_05737_),
    .A1(net673),
    .A2(_05306_));
 sg13g2_a22oi_1 _23358_ (.Y(_05738_),
    .B1(_05737_),
    .B2(net485),
    .A2(_05735_),
    .A1(_05022_));
 sg13g2_o21ai_1 _23359_ (.B1(_05141_),
    .Y(_05739_),
    .A1(net832),
    .A2(_05738_));
 sg13g2_mux2_1 _23360_ (.A0(_05739_),
    .A1(_10831_),
    .S(_05144_),
    .X(_05740_));
 sg13g2_o21ai_1 _23361_ (.B1(_05740_),
    .Y(_05741_),
    .A1(_08656_),
    .A2(_05017_));
 sg13g2_a21oi_1 _23362_ (.A1(_05259_),
    .A2(_05730_),
    .Y(_01020_),
    .B1(_05741_));
 sg13g2_buf_1 _23363_ (.A(net111),
    .X(_05742_));
 sg13g2_inv_1 _23364_ (.Y(_05743_),
    .A(_03590_));
 sg13g2_a21oi_1 _23365_ (.A1(_05743_),
    .A2(\cpu.dec.r_rd[0] ),
    .Y(_05744_),
    .B1(_05016_));
 sg13g2_buf_1 _23366_ (.A(_11515_),
    .X(_05745_));
 sg13g2_nor2_1 _23367_ (.A(_10025_),
    .B(_05745_),
    .Y(_05746_));
 sg13g2_a21oi_1 _23368_ (.A1(net93),
    .A2(_05744_),
    .Y(_01021_),
    .B1(_05746_));
 sg13g2_a21oi_1 _23369_ (.A1(_05743_),
    .A2(\cpu.dec.r_rd[1] ),
    .Y(_05747_),
    .B1(_05016_));
 sg13g2_nor2_1 _23370_ (.A(_10023_),
    .B(_05745_),
    .Y(_05748_));
 sg13g2_a21oi_1 _23371_ (.A1(net93),
    .A2(_05747_),
    .Y(_01022_),
    .B1(_05748_));
 sg13g2_nor3_1 _23372_ (.A(_03590_),
    .B(_09123_),
    .C(net288),
    .Y(_05749_));
 sg13g2_nand3_1 _23373_ (.B(_04810_),
    .C(_05749_),
    .A(\cpu.dec.r_rd[2] ),
    .Y(_05750_));
 sg13g2_o21ai_1 _23374_ (.B1(_05750_),
    .Y(_01023_),
    .A1(_03636_),
    .A2(_05742_));
 sg13g2_nand3_1 _23375_ (.B(_04810_),
    .C(_05749_),
    .A(\cpu.dec.r_rd[3] ),
    .Y(_05751_));
 sg13g2_o21ai_1 _23376_ (.B1(_05751_),
    .Y(_01024_),
    .A1(_10020_),
    .A2(_05742_));
 sg13g2_mux2_1 _23377_ (.A0(\cpu.dec.r_swapsp ),
    .A1(\cpu.ex.r_wb_swapsp ),
    .S(net110),
    .X(_01025_));
 sg13g2_nand2_1 _23378_ (.Y(_05752_),
    .A(net960),
    .B(_11043_));
 sg13g2_o21ai_1 _23379_ (.B1(_05752_),
    .Y(_05753_),
    .A1(_10344_),
    .A2(_10196_));
 sg13g2_mux2_1 _23380_ (.A0(_09861_),
    .A1(_05753_),
    .S(net94),
    .X(_01026_));
 sg13g2_a21oi_2 _23381_ (.B1(_10457_),
    .Y(_05754_),
    .A2(_11587_),
    .A1(net525));
 sg13g2_a221oi_1 _23382_ (.B2(_10991_),
    .C1(net832),
    .B1(net525),
    .A1(net1095),
    .Y(_05755_),
    .A2(net459));
 sg13g2_a21o_1 _23383_ (.A2(_05754_),
    .A1(net831),
    .B1(_05755_),
    .X(_05756_));
 sg13g2_nand2_1 _23384_ (.Y(_05757_),
    .A(_09986_),
    .B(net110));
 sg13g2_o21ai_1 _23385_ (.B1(_05757_),
    .Y(_01027_),
    .A1(net110),
    .A2(_05756_));
 sg13g2_and2_1 _23386_ (.A(net525),
    .B(_10423_),
    .X(_05758_));
 sg13g2_a21o_1 _23387_ (.A2(net459),
    .A1(_09106_),
    .B1(_05758_),
    .X(_05759_));
 sg13g2_a21oi_1 _23388_ (.A1(_10906_),
    .A2(_10908_),
    .Y(_05760_),
    .B1(net831));
 sg13g2_a21oi_1 _23389_ (.A1(net831),
    .A2(_05759_),
    .Y(_05761_),
    .B1(_05760_));
 sg13g2_nand2_1 _23390_ (.Y(_05762_),
    .A(_09991_),
    .B(net110));
 sg13g2_o21ai_1 _23391_ (.B1(_05762_),
    .Y(_01028_),
    .A1(net110),
    .A2(_05761_));
 sg13g2_nand2_1 _23392_ (.Y(_05763_),
    .A(_10550_),
    .B(_10570_));
 sg13g2_a22oi_1 _23393_ (.Y(_05764_),
    .B1(net525),
    .B2(_05763_),
    .A2(net459),
    .A1(_03656_));
 sg13g2_nand2_1 _23394_ (.Y(_05765_),
    .A(_11505_),
    .B(_11173_));
 sg13g2_o21ai_1 _23395_ (.B1(_05765_),
    .Y(_05766_),
    .A1(_11505_),
    .A2(_05764_));
 sg13g2_nand2_1 _23396_ (.Y(_05767_),
    .A(net109),
    .B(_05766_));
 sg13g2_o21ai_1 _23397_ (.B1(_05767_),
    .Y(_01029_),
    .A1(_12060_),
    .A2(net93));
 sg13g2_nand2_1 _23398_ (.Y(_05768_),
    .A(net831),
    .B(_10536_));
 sg13g2_inv_1 _23399_ (.Y(_05769_),
    .A(_11148_));
 sg13g2_o21ai_1 _23400_ (.B1(_11505_),
    .Y(_05770_),
    .A1(_11147_),
    .A2(_05769_));
 sg13g2_a21o_1 _23401_ (.A2(_05770_),
    .A1(_05768_),
    .B1(net144),
    .X(_05771_));
 sg13g2_o21ai_1 _23402_ (.B1(_05771_),
    .Y(_01030_),
    .A1(_12070_),
    .A2(net93));
 sg13g2_nand2_1 _23403_ (.Y(_05772_),
    .A(_05018_),
    .B(_10708_));
 sg13g2_o21ai_1 _23404_ (.B1(_05772_),
    .Y(_05773_),
    .A1(net831),
    .A2(_11067_));
 sg13g2_nand2_1 _23405_ (.Y(_05774_),
    .A(net109),
    .B(_05773_));
 sg13g2_o21ai_1 _23406_ (.B1(_05774_),
    .Y(_01031_),
    .A1(_12077_),
    .A2(net93));
 sg13g2_nand2_1 _23407_ (.Y(_05775_),
    .A(net965),
    .B(net459));
 sg13g2_nand2_1 _23408_ (.Y(_05776_),
    .A(_10793_),
    .B(_05775_));
 sg13g2_nand2_1 _23409_ (.Y(_05777_),
    .A(net832),
    .B(_05776_));
 sg13g2_o21ai_1 _23410_ (.B1(_05777_),
    .Y(_05778_),
    .A1(net831),
    .A2(_11208_));
 sg13g2_nand2_1 _23411_ (.Y(_05779_),
    .A(net109),
    .B(_05778_));
 sg13g2_o21ai_1 _23412_ (.B1(_05779_),
    .Y(_01032_),
    .A1(_12084_),
    .A2(net93));
 sg13g2_buf_1 _23413_ (.A(net1023),
    .X(_05780_));
 sg13g2_nand2_1 _23414_ (.Y(_05781_),
    .A(_03651_),
    .B(_11043_));
 sg13g2_o21ai_1 _23415_ (.B1(_05781_),
    .Y(_05782_),
    .A1(_10344_),
    .A2(_10325_));
 sg13g2_mux2_1 _23416_ (.A0(_05780_),
    .A1(_05782_),
    .S(net94),
    .X(_01033_));
 sg13g2_nor2_1 _23417_ (.A(net876),
    .B(net109),
    .Y(_05783_));
 sg13g2_a21oi_1 _23418_ (.A1(_05754_),
    .A2(net93),
    .Y(_01034_),
    .B1(_05783_));
 sg13g2_nand2_1 _23419_ (.Y(_05784_),
    .A(net109),
    .B(_05759_));
 sg13g2_o21ai_1 _23420_ (.B1(_05784_),
    .Y(_01035_),
    .A1(net721),
    .A2(net94));
 sg13g2_nor2_1 _23421_ (.A(net1105),
    .B(net109),
    .Y(_05785_));
 sg13g2_a21oi_1 _23422_ (.A1(net93),
    .A2(_05764_),
    .Y(_01036_),
    .B1(_05785_));
 sg13g2_mux2_1 _23423_ (.A0(_12522_),
    .A1(_10536_),
    .S(net94),
    .X(_01037_));
 sg13g2_mux2_1 _23424_ (.A0(_09957_),
    .A1(_10708_),
    .S(net94),
    .X(_01038_));
 sg13g2_nand2_1 _23425_ (.Y(_05786_),
    .A(_05776_),
    .B(net111));
 sg13g2_o21ai_1 _23426_ (.B1(_05786_),
    .Y(_01039_),
    .A1(_02766_),
    .A2(net94));
 sg13g2_a22oi_1 _23427_ (.Y(_05787_),
    .B1(net525),
    .B2(_10639_),
    .A2(net459),
    .A1(net1037));
 sg13g2_nand2_1 _23428_ (.Y(_05788_),
    .A(_05151_),
    .B(_05753_));
 sg13g2_o21ai_1 _23429_ (.B1(_05788_),
    .Y(_05789_),
    .A1(_05151_),
    .A2(_05787_));
 sg13g2_mux2_1 _23430_ (.A0(_09975_),
    .A1(_05789_),
    .S(net109),
    .X(_01040_));
 sg13g2_nand2_1 _23431_ (.Y(_05790_),
    .A(_05018_),
    .B(_05782_));
 sg13g2_o21ai_1 _23432_ (.B1(_05790_),
    .Y(_05791_),
    .A1(net831),
    .A2(_10873_));
 sg13g2_nand2_1 _23433_ (.Y(_05792_),
    .A(net109),
    .B(_05791_));
 sg13g2_o21ai_1 _23434_ (.B1(_05792_),
    .Y(_01041_),
    .A1(_12157_),
    .A2(net94));
 sg13g2_inv_1 _23435_ (.Y(_05793_),
    .A(_11010_));
 sg13g2_or3_1 _23436_ (.A(_10205_),
    .B(_10458_),
    .C(_10427_),
    .X(_05794_));
 sg13g2_buf_1 _23437_ (.A(_05794_),
    .X(_05795_));
 sg13g2_o21ai_1 _23438_ (.B1(_03465_),
    .Y(_05796_),
    .A1(_10327_),
    .A2(_05795_));
 sg13g2_buf_2 _23439_ (.A(_05796_),
    .X(_05797_));
 sg13g2_nor4_2 _23440_ (.A(_08132_),
    .B(_04765_),
    .C(_10022_),
    .Y(_05798_),
    .D(_03671_));
 sg13g2_and2_1 _23441_ (.A(_05797_),
    .B(_05798_),
    .X(_05799_));
 sg13g2_buf_1 _23442_ (.A(_05799_),
    .X(_05800_));
 sg13g2_o21ai_1 _23443_ (.B1(_08963_),
    .Y(_05801_),
    .A1(_11496_),
    .A2(_05800_));
 sg13g2_buf_1 _23444_ (.A(_05801_),
    .X(_05802_));
 sg13g2_buf_1 _23445_ (.A(_00267_),
    .X(_05803_));
 sg13g2_nand2b_1 _23446_ (.Y(_05804_),
    .B(net960),
    .A_N(_05803_));
 sg13g2_o21ai_1 _23447_ (.B1(_05804_),
    .Y(_05805_),
    .A1(net960),
    .A2(_11023_));
 sg13g2_nand3_1 _23448_ (.B(_05800_),
    .C(_05805_),
    .A(net290),
    .Y(_05806_));
 sg13g2_nand2_1 _23449_ (.Y(_05807_),
    .A(net589),
    .B(_08256_));
 sg13g2_o21ai_1 _23450_ (.B1(_05807_),
    .Y(_05808_),
    .A1(_08229_),
    .A2(_08256_));
 sg13g2_or2_1 _23451_ (.X(_05809_),
    .B(_05808_),
    .A(net387));
 sg13g2_a21oi_1 _23452_ (.A1(_05806_),
    .A2(_05809_),
    .Y(_05810_),
    .B1(net684));
 sg13g2_a21oi_1 _23453_ (.A1(_05793_),
    .A2(_05802_),
    .Y(_01044_),
    .B1(_05810_));
 sg13g2_buf_1 _23454_ (.A(_11115_),
    .X(_05811_));
 sg13g2_mux2_1 _23455_ (.A0(_08339_),
    .A1(_09483_),
    .S(_08256_),
    .X(_05812_));
 sg13g2_nand2_1 _23456_ (.Y(_05813_),
    .A(_05797_),
    .B(_05798_));
 sg13g2_and2_1 _23457_ (.A(_11010_),
    .B(_11115_),
    .X(_05814_));
 sg13g2_buf_1 _23458_ (.A(_05814_),
    .X(_05815_));
 sg13g2_buf_1 _23459_ (.A(_11010_),
    .X(_05816_));
 sg13g2_nor2_1 _23460_ (.A(net950),
    .B(net951),
    .Y(_05817_));
 sg13g2_o21ai_1 _23461_ (.B1(net960),
    .Y(_05818_),
    .A1(_05815_),
    .A2(_05817_));
 sg13g2_o21ai_1 _23462_ (.B1(_05818_),
    .Y(_05819_),
    .A1(net960),
    .A2(net601));
 sg13g2_nor2_1 _23463_ (.A(_05813_),
    .B(_05819_),
    .Y(_05820_));
 sg13g2_mux2_1 _23464_ (.A0(_05812_),
    .A1(_05820_),
    .S(net387),
    .X(_05821_));
 sg13g2_a22oi_1 _23465_ (.Y(_05822_),
    .B1(_05821_),
    .B2(_09118_),
    .A2(_05802_),
    .A1(_05811_));
 sg13g2_inv_1 _23466_ (.Y(_01045_),
    .A(_05822_));
 sg13g2_inv_2 _23467_ (.Y(_05823_),
    .A(_11062_));
 sg13g2_buf_1 _23468_ (.A(_11062_),
    .X(_05824_));
 sg13g2_nand2_1 _23469_ (.Y(_05825_),
    .A(_11010_),
    .B(_11115_));
 sg13g2_buf_1 _23470_ (.A(_05825_),
    .X(_05826_));
 sg13g2_nor2_1 _23471_ (.A(_05824_),
    .B(net828),
    .Y(_05827_));
 sg13g2_buf_1 _23472_ (.A(net949),
    .X(_05828_));
 sg13g2_nand2_1 _23473_ (.Y(_05829_),
    .A(net827),
    .B(_05826_));
 sg13g2_nand3b_1 _23474_ (.B(_05829_),
    .C(_03632_),
    .Y(_05830_),
    .A_N(_05827_));
 sg13g2_o21ai_1 _23475_ (.B1(_05830_),
    .Y(_05831_),
    .A1(net960),
    .A2(net732));
 sg13g2_nand3_1 _23476_ (.B(_05800_),
    .C(_05831_),
    .A(net290),
    .Y(_05832_));
 sg13g2_nand2b_1 _23477_ (.Y(_05833_),
    .B(_08438_),
    .A_N(_08256_));
 sg13g2_nand2_1 _23478_ (.Y(_05834_),
    .A(_11042_),
    .B(_08256_));
 sg13g2_nand3_1 _23479_ (.B(_05833_),
    .C(_05834_),
    .A(_11496_),
    .Y(_05835_));
 sg13g2_a21oi_1 _23480_ (.A1(_05832_),
    .A2(_05835_),
    .Y(_05836_),
    .B1(_09124_));
 sg13g2_a21oi_1 _23481_ (.A1(_05823_),
    .A2(_05802_),
    .Y(_01046_),
    .B1(_05836_));
 sg13g2_inv_2 _23482_ (.Y(_05837_),
    .A(_11188_));
 sg13g2_nand2_1 _23483_ (.Y(_05838_),
    .A(net949),
    .B(_05815_));
 sg13g2_buf_2 _23484_ (.A(_05838_),
    .X(_05839_));
 sg13g2_xnor2_1 _23485_ (.Y(_05840_),
    .A(_05837_),
    .B(_05839_));
 sg13g2_nand2_1 _23486_ (.Y(_05841_),
    .A(_03632_),
    .B(_05840_));
 sg13g2_o21ai_1 _23487_ (.B1(_05841_),
    .Y(_05842_),
    .A1(net960),
    .A2(net731));
 sg13g2_nand3_1 _23488_ (.B(_05800_),
    .C(_05842_),
    .A(net290),
    .Y(_05843_));
 sg13g2_nand2_1 _23489_ (.Y(_05844_),
    .A(_11186_),
    .B(_08256_));
 sg13g2_o21ai_1 _23490_ (.B1(_05844_),
    .Y(_05845_),
    .A1(_08389_),
    .A2(_08256_));
 sg13g2_or2_1 _23491_ (.X(_05846_),
    .B(_05845_),
    .A(_08259_));
 sg13g2_a21oi_1 _23492_ (.A1(_05843_),
    .A2(_05846_),
    .Y(_05847_),
    .B1(_09129_));
 sg13g2_a21oi_1 _23493_ (.A1(_05837_),
    .A2(_05802_),
    .Y(_01047_),
    .B1(_05847_));
 sg13g2_buf_1 _23494_ (.A(net448),
    .X(_05848_));
 sg13g2_buf_2 _23495_ (.A(_00172_),
    .X(_05849_));
 sg13g2_nor2_1 _23496_ (.A(_10079_),
    .B(_11188_),
    .Y(_05850_));
 sg13g2_buf_1 _23497_ (.A(_05850_),
    .X(_05851_));
 sg13g2_nand2_1 _23498_ (.Y(_05852_),
    .A(_05849_),
    .B(_05851_));
 sg13g2_nand3b_1 _23499_ (.B(_05798_),
    .C(net1118),
    .Y(_05853_),
    .A_N(_10382_));
 sg13g2_buf_1 _23500_ (.A(_05853_),
    .X(_05854_));
 sg13g2_or3_1 _23501_ (.A(net950),
    .B(net951),
    .C(_05854_),
    .X(_05855_));
 sg13g2_buf_1 _23502_ (.A(_05855_),
    .X(_05856_));
 sg13g2_nor2_1 _23503_ (.A(_05852_),
    .B(_05856_),
    .Y(_05857_));
 sg13g2_buf_1 _23504_ (.A(_05857_),
    .X(_05858_));
 sg13g2_buf_1 _23505_ (.A(_05858_),
    .X(_05859_));
 sg13g2_mux2_1 _23506_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][0] ),
    .A1(net401),
    .S(net286),
    .X(_01115_));
 sg13g2_mux2_1 _23507_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][10] ),
    .A1(net565),
    .S(net286),
    .X(_01116_));
 sg13g2_mux2_1 _23508_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][11] ),
    .A1(net635),
    .S(_05859_),
    .X(_01117_));
 sg13g2_mux2_1 _23509_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][1] ),
    .A1(net570),
    .S(net286),
    .X(_01118_));
 sg13g2_mux2_1 _23510_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][2] ),
    .A1(_03133_),
    .S(net286),
    .X(_01119_));
 sg13g2_buf_1 _23511_ (.A(net965),
    .X(_05860_));
 sg13g2_mux2_1 _23512_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][3] ),
    .A1(_05860_),
    .S(net286),
    .X(_01120_));
 sg13g2_mux2_1 _23513_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][4] ),
    .A1(net833),
    .S(net286),
    .X(_01121_));
 sg13g2_mux2_1 _23514_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][5] ),
    .A1(net953),
    .S(net286),
    .X(_01122_));
 sg13g2_buf_1 _23515_ (.A(net963),
    .X(_05861_));
 sg13g2_mux2_1 _23516_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][6] ),
    .A1(net825),
    .S(_05859_),
    .X(_01123_));
 sg13g2_buf_1 _23517_ (.A(net962),
    .X(_05862_));
 sg13g2_mux2_1 _23518_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][7] ),
    .A1(_05862_),
    .S(net286),
    .X(_01124_));
 sg13g2_mux2_1 _23519_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][8] ),
    .A1(net496),
    .S(_05858_),
    .X(_01125_));
 sg13g2_mux2_1 _23520_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][9] ),
    .A1(net447),
    .S(_05858_),
    .X(_01126_));
 sg13g2_buf_1 _23521_ (.A(_05854_),
    .X(_05863_));
 sg13g2_nand2_1 _23522_ (.Y(_05864_),
    .A(_05793_),
    .B(net951));
 sg13g2_buf_1 _23523_ (.A(_05864_),
    .X(_05865_));
 sg13g2_nand2_1 _23524_ (.Y(_05866_),
    .A(_10080_),
    .B(_11188_));
 sg13g2_buf_1 _23525_ (.A(_05866_),
    .X(_05867_));
 sg13g2_nor3_2 _23526_ (.A(net949),
    .B(net708),
    .C(_05867_),
    .Y(_05868_));
 sg13g2_nor2b_1 _23527_ (.A(net484),
    .B_N(_05868_),
    .Y(_05869_));
 sg13g2_buf_1 _23528_ (.A(_05869_),
    .X(_05870_));
 sg13g2_buf_1 _23529_ (.A(_05870_),
    .X(_05871_));
 sg13g2_mux2_1 _23530_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][0] ),
    .A1(net401),
    .S(net353),
    .X(_01127_));
 sg13g2_mux2_1 _23531_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][10] ),
    .A1(net565),
    .S(net353),
    .X(_01128_));
 sg13g2_mux2_1 _23532_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][11] ),
    .A1(net635),
    .S(net353),
    .X(_01129_));
 sg13g2_mux2_1 _23533_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][1] ),
    .A1(net570),
    .S(net353),
    .X(_01130_));
 sg13g2_mux2_1 _23534_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][2] ),
    .A1(_03133_),
    .S(net353),
    .X(_01131_));
 sg13g2_mux2_1 _23535_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][3] ),
    .A1(net826),
    .S(net353),
    .X(_01132_));
 sg13g2_mux2_1 _23536_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][4] ),
    .A1(_04770_),
    .S(net353),
    .X(_01133_));
 sg13g2_mux2_1 _23537_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][5] ),
    .A1(net953),
    .S(_05871_),
    .X(_01134_));
 sg13g2_mux2_1 _23538_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][6] ),
    .A1(net825),
    .S(_05871_),
    .X(_01135_));
 sg13g2_mux2_1 _23539_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][7] ),
    .A1(net824),
    .S(net353),
    .X(_01136_));
 sg13g2_mux2_1 _23540_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][8] ),
    .A1(net496),
    .S(_05870_),
    .X(_01137_));
 sg13g2_mux2_1 _23541_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][9] ),
    .A1(net447),
    .S(_05870_),
    .X(_01138_));
 sg13g2_nor3_1 _23542_ (.A(net949),
    .B(_05826_),
    .C(_05867_),
    .Y(_05872_));
 sg13g2_buf_2 _23543_ (.A(_05872_),
    .X(_05873_));
 sg13g2_nor2b_1 _23544_ (.A(net484),
    .B_N(_05873_),
    .Y(_05874_));
 sg13g2_buf_1 _23545_ (.A(_05874_),
    .X(_05875_));
 sg13g2_buf_1 _23546_ (.A(_05875_),
    .X(_05876_));
 sg13g2_mux2_1 _23547_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][0] ),
    .A1(net401),
    .S(net352),
    .X(_01139_));
 sg13g2_mux2_1 _23548_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][10] ),
    .A1(net565),
    .S(net352),
    .X(_01140_));
 sg13g2_mux2_1 _23549_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][11] ),
    .A1(net635),
    .S(net352),
    .X(_01141_));
 sg13g2_mux2_1 _23550_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][1] ),
    .A1(net570),
    .S(net352),
    .X(_01142_));
 sg13g2_buf_1 _23551_ (.A(net966),
    .X(_05877_));
 sg13g2_mux2_1 _23552_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][2] ),
    .A1(_05877_),
    .S(net352),
    .X(_01143_));
 sg13g2_mux2_1 _23553_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][3] ),
    .A1(net826),
    .S(net352),
    .X(_01144_));
 sg13g2_mux2_1 _23554_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][4] ),
    .A1(net833),
    .S(_05876_),
    .X(_01145_));
 sg13g2_mux2_1 _23555_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][5] ),
    .A1(net953),
    .S(_05876_),
    .X(_01146_));
 sg13g2_mux2_1 _23556_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][6] ),
    .A1(net825),
    .S(net352),
    .X(_01147_));
 sg13g2_mux2_1 _23557_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][7] ),
    .A1(_05862_),
    .S(net352),
    .X(_01148_));
 sg13g2_mux2_1 _23558_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][8] ),
    .A1(net496),
    .S(_05875_),
    .X(_01149_));
 sg13g2_mux2_1 _23559_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][9] ),
    .A1(net447),
    .S(_05875_),
    .X(_01150_));
 sg13g2_nor2_1 _23560_ (.A(_10079_),
    .B(_05837_),
    .Y(_05878_));
 sg13g2_nand2b_1 _23561_ (.Y(_05879_),
    .B(_05878_),
    .A_N(_05849_));
 sg13g2_buf_1 _23562_ (.A(_05879_),
    .X(_05880_));
 sg13g2_nor2_1 _23563_ (.A(_05856_),
    .B(_05880_),
    .Y(_05881_));
 sg13g2_buf_1 _23564_ (.A(_05881_),
    .X(_05882_));
 sg13g2_buf_1 _23565_ (.A(_05882_),
    .X(_05883_));
 sg13g2_mux2_1 _23566_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][0] ),
    .A1(net401),
    .S(net285),
    .X(_01151_));
 sg13g2_mux2_1 _23567_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][10] ),
    .A1(net565),
    .S(net285),
    .X(_01152_));
 sg13g2_mux2_1 _23568_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][11] ),
    .A1(net635),
    .S(_05883_),
    .X(_01153_));
 sg13g2_mux2_1 _23569_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][1] ),
    .A1(_03688_),
    .S(net285),
    .X(_01154_));
 sg13g2_mux2_1 _23570_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][2] ),
    .A1(_05877_),
    .S(_05883_),
    .X(_01155_));
 sg13g2_mux2_1 _23571_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][3] ),
    .A1(net826),
    .S(net285),
    .X(_01156_));
 sg13g2_mux2_1 _23572_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][4] ),
    .A1(net833),
    .S(net285),
    .X(_01157_));
 sg13g2_mux2_1 _23573_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][5] ),
    .A1(net953),
    .S(net285),
    .X(_01158_));
 sg13g2_mux2_1 _23574_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][6] ),
    .A1(net825),
    .S(net285),
    .X(_01159_));
 sg13g2_mux2_1 _23575_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][7] ),
    .A1(net824),
    .S(net285),
    .X(_01160_));
 sg13g2_mux2_1 _23576_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][8] ),
    .A1(net496),
    .S(_05882_),
    .X(_01161_));
 sg13g2_mux2_1 _23577_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][9] ),
    .A1(net447),
    .S(_05882_),
    .X(_01162_));
 sg13g2_nand2b_1 _23578_ (.Y(_05884_),
    .B(_11010_),
    .A_N(net951));
 sg13g2_buf_2 _23579_ (.A(_05884_),
    .X(_05885_));
 sg13g2_or2_1 _23580_ (.X(_05886_),
    .B(_05854_),
    .A(_05885_));
 sg13g2_buf_2 _23581_ (.A(_05886_),
    .X(_05887_));
 sg13g2_nor2_1 _23582_ (.A(_05880_),
    .B(_05887_),
    .Y(_05888_));
 sg13g2_buf_1 _23583_ (.A(_05888_),
    .X(_05889_));
 sg13g2_buf_1 _23584_ (.A(_05889_),
    .X(_05890_));
 sg13g2_mux2_1 _23585_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][0] ),
    .A1(net401),
    .S(net284),
    .X(_01163_));
 sg13g2_mux2_1 _23586_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][10] ),
    .A1(_04769_),
    .S(net284),
    .X(_01164_));
 sg13g2_mux2_1 _23587_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][11] ),
    .A1(net635),
    .S(net284),
    .X(_01165_));
 sg13g2_mux2_1 _23588_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][1] ),
    .A1(_03688_),
    .S(net284),
    .X(_01166_));
 sg13g2_mux2_1 _23589_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][2] ),
    .A1(net823),
    .S(_05890_),
    .X(_01167_));
 sg13g2_mux2_1 _23590_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][3] ),
    .A1(net826),
    .S(net284),
    .X(_01168_));
 sg13g2_mux2_1 _23591_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][4] ),
    .A1(net833),
    .S(net284),
    .X(_01169_));
 sg13g2_mux2_1 _23592_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][5] ),
    .A1(net953),
    .S(net284),
    .X(_01170_));
 sg13g2_mux2_1 _23593_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][6] ),
    .A1(_05861_),
    .S(_05890_),
    .X(_01171_));
 sg13g2_mux2_1 _23594_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][7] ),
    .A1(net824),
    .S(net284),
    .X(_01172_));
 sg13g2_mux2_1 _23595_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][8] ),
    .A1(net496),
    .S(_05889_),
    .X(_01173_));
 sg13g2_mux2_1 _23596_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][9] ),
    .A1(net447),
    .S(_05889_),
    .X(_01174_));
 sg13g2_buf_1 _23597_ (.A(_05854_),
    .X(_05891_));
 sg13g2_nor3_1 _23598_ (.A(net708),
    .B(_05891_),
    .C(_05880_),
    .Y(_05892_));
 sg13g2_buf_1 _23599_ (.A(_05892_),
    .X(_05893_));
 sg13g2_buf_1 _23600_ (.A(_05893_),
    .X(_05894_));
 sg13g2_mux2_1 _23601_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][0] ),
    .A1(_05848_),
    .S(net351),
    .X(_01175_));
 sg13g2_mux2_1 _23602_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][10] ),
    .A1(net565),
    .S(net351),
    .X(_01176_));
 sg13g2_mux2_1 _23603_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][11] ),
    .A1(net635),
    .S(net351),
    .X(_01177_));
 sg13g2_buf_1 _23604_ (.A(net640),
    .X(_05895_));
 sg13g2_mux2_1 _23605_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][1] ),
    .A1(_05895_),
    .S(net351),
    .X(_01178_));
 sg13g2_mux2_1 _23606_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][2] ),
    .A1(net823),
    .S(_05894_),
    .X(_01179_));
 sg13g2_mux2_1 _23607_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][3] ),
    .A1(net826),
    .S(net351),
    .X(_01180_));
 sg13g2_mux2_1 _23608_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][4] ),
    .A1(net833),
    .S(net351),
    .X(_01181_));
 sg13g2_mux2_1 _23609_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][5] ),
    .A1(net953),
    .S(net351),
    .X(_01182_));
 sg13g2_mux2_1 _23610_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][6] ),
    .A1(_05861_),
    .S(_05894_),
    .X(_01183_));
 sg13g2_mux2_1 _23611_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][7] ),
    .A1(net824),
    .S(net351),
    .X(_01184_));
 sg13g2_mux2_1 _23612_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][8] ),
    .A1(_03696_),
    .S(_05893_),
    .X(_01185_));
 sg13g2_mux2_1 _23613_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][9] ),
    .A1(_03697_),
    .S(_05893_),
    .X(_01186_));
 sg13g2_nor3_1 _23614_ (.A(net828),
    .B(net483),
    .C(_05880_),
    .Y(_05896_));
 sg13g2_buf_1 _23615_ (.A(_05896_),
    .X(_05897_));
 sg13g2_buf_1 _23616_ (.A(_05897_),
    .X(_05898_));
 sg13g2_mux2_1 _23617_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][0] ),
    .A1(_05848_),
    .S(net350),
    .X(_01187_));
 sg13g2_mux2_1 _23618_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][10] ),
    .A1(net565),
    .S(net350),
    .X(_01188_));
 sg13g2_mux2_1 _23619_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][11] ),
    .A1(_03705_),
    .S(_05898_),
    .X(_01189_));
 sg13g2_mux2_1 _23620_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][1] ),
    .A1(net562),
    .S(net350),
    .X(_01190_));
 sg13g2_mux2_1 _23621_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][2] ),
    .A1(net823),
    .S(_05898_),
    .X(_01191_));
 sg13g2_mux2_1 _23622_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][3] ),
    .A1(net826),
    .S(net350),
    .X(_01192_));
 sg13g2_mux2_1 _23623_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][4] ),
    .A1(net833),
    .S(net350),
    .X(_01193_));
 sg13g2_mux2_1 _23624_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][5] ),
    .A1(_04771_),
    .S(net350),
    .X(_01194_));
 sg13g2_mux2_1 _23625_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][6] ),
    .A1(net825),
    .S(net350),
    .X(_01195_));
 sg13g2_mux2_1 _23626_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][7] ),
    .A1(net824),
    .S(net350),
    .X(_01196_));
 sg13g2_mux2_1 _23627_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][8] ),
    .A1(_03696_),
    .S(_05897_),
    .X(_01197_));
 sg13g2_mux2_1 _23628_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][9] ),
    .A1(_03697_),
    .S(_05897_),
    .X(_01198_));
 sg13g2_nand2_1 _23629_ (.Y(_05899_),
    .A(_10079_),
    .B(_05837_));
 sg13g2_buf_2 _23630_ (.A(_05899_),
    .X(_05900_));
 sg13g2_nor2_1 _23631_ (.A(_11115_),
    .B(_11062_),
    .Y(_05901_));
 sg13g2_buf_1 _23632_ (.A(_05901_),
    .X(_05902_));
 sg13g2_nand2_1 _23633_ (.Y(_05903_),
    .A(_05793_),
    .B(_05902_));
 sg13g2_nor3_1 _23634_ (.A(net483),
    .B(_05900_),
    .C(_05903_),
    .Y(_05904_));
 sg13g2_buf_1 _23635_ (.A(_05904_),
    .X(_05905_));
 sg13g2_buf_1 _23636_ (.A(_05905_),
    .X(_05906_));
 sg13g2_mux2_1 _23637_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][0] ),
    .A1(net401),
    .S(net349),
    .X(_01199_));
 sg13g2_mux2_1 _23638_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][10] ),
    .A1(net565),
    .S(net349),
    .X(_01200_));
 sg13g2_mux2_1 _23639_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][11] ),
    .A1(_03705_),
    .S(_05906_),
    .X(_01201_));
 sg13g2_mux2_1 _23640_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][1] ),
    .A1(net562),
    .S(net349),
    .X(_01202_));
 sg13g2_mux2_1 _23641_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][2] ),
    .A1(net823),
    .S(net349),
    .X(_01203_));
 sg13g2_mux2_1 _23642_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][3] ),
    .A1(net826),
    .S(net349),
    .X(_01204_));
 sg13g2_mux2_1 _23643_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][4] ),
    .A1(net833),
    .S(net349),
    .X(_01205_));
 sg13g2_mux2_1 _23644_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][5] ),
    .A1(net953),
    .S(net349),
    .X(_01206_));
 sg13g2_mux2_1 _23645_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][6] ),
    .A1(net825),
    .S(_05906_),
    .X(_01207_));
 sg13g2_mux2_1 _23646_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][7] ),
    .A1(net824),
    .S(net349),
    .X(_01208_));
 sg13g2_buf_1 _23647_ (.A(_11023_),
    .X(_05907_));
 sg13g2_mux2_1 _23648_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][8] ),
    .A1(net482),
    .S(_05905_),
    .X(_01209_));
 sg13g2_buf_1 _23649_ (.A(net601),
    .X(_05908_));
 sg13g2_mux2_1 _23650_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][9] ),
    .A1(net481),
    .S(_05905_),
    .X(_01210_));
 sg13g2_nor3_1 _23651_ (.A(net827),
    .B(_05887_),
    .C(_05900_),
    .Y(_05909_));
 sg13g2_buf_1 _23652_ (.A(_05909_),
    .X(_05910_));
 sg13g2_buf_1 _23653_ (.A(_05910_),
    .X(_05911_));
 sg13g2_mux2_1 _23654_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][0] ),
    .A1(net401),
    .S(net283),
    .X(_01211_));
 sg13g2_mux2_1 _23655_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][10] ),
    .A1(net565),
    .S(net283),
    .X(_01212_));
 sg13g2_buf_1 _23656_ (.A(net731),
    .X(_05912_));
 sg13g2_mux2_1 _23657_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][11] ),
    .A1(net629),
    .S(net283),
    .X(_01213_));
 sg13g2_mux2_1 _23658_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][1] ),
    .A1(net562),
    .S(net283),
    .X(_01214_));
 sg13g2_mux2_1 _23659_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][2] ),
    .A1(net823),
    .S(net283),
    .X(_01215_));
 sg13g2_mux2_1 _23660_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][3] ),
    .A1(net826),
    .S(net283),
    .X(_01216_));
 sg13g2_mux2_1 _23661_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][4] ),
    .A1(net833),
    .S(net283),
    .X(_01217_));
 sg13g2_mux2_1 _23662_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][5] ),
    .A1(net953),
    .S(_05911_),
    .X(_01218_));
 sg13g2_mux2_1 _23663_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][6] ),
    .A1(net825),
    .S(_05911_),
    .X(_01219_));
 sg13g2_mux2_1 _23664_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][7] ),
    .A1(net824),
    .S(net283),
    .X(_01220_));
 sg13g2_mux2_1 _23665_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][8] ),
    .A1(net482),
    .S(_05910_),
    .X(_01221_));
 sg13g2_mux2_1 _23666_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][9] ),
    .A1(_05908_),
    .S(_05910_),
    .X(_01222_));
 sg13g2_buf_1 _23667_ (.A(_11188_),
    .X(_05913_));
 sg13g2_nor2_1 _23668_ (.A(_10080_),
    .B(net950),
    .Y(_05914_));
 sg13g2_nand3_1 _23669_ (.B(_05823_),
    .C(_05914_),
    .A(net951),
    .Y(_05915_));
 sg13g2_nor2_2 _23670_ (.A(net948),
    .B(_05915_),
    .Y(_05916_));
 sg13g2_nor2b_1 _23671_ (.A(net484),
    .B_N(_05916_),
    .Y(_05917_));
 sg13g2_buf_1 _23672_ (.A(_05917_),
    .X(_05918_));
 sg13g2_buf_1 _23673_ (.A(_05918_),
    .X(_05919_));
 sg13g2_mux2_1 _23674_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][0] ),
    .A1(net401),
    .S(net348),
    .X(_01223_));
 sg13g2_buf_1 _23675_ (.A(net732),
    .X(_05920_));
 sg13g2_mux2_1 _23676_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][10] ),
    .A1(_05920_),
    .S(net348),
    .X(_01224_));
 sg13g2_mux2_1 _23677_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][11] ),
    .A1(net629),
    .S(net348),
    .X(_01225_));
 sg13g2_mux2_1 _23678_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][1] ),
    .A1(net562),
    .S(net348),
    .X(_01226_));
 sg13g2_mux2_1 _23679_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][2] ),
    .A1(net823),
    .S(net348),
    .X(_01227_));
 sg13g2_mux2_1 _23680_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][3] ),
    .A1(_05860_),
    .S(net348),
    .X(_01228_));
 sg13g2_buf_1 _23681_ (.A(_09025_),
    .X(_05921_));
 sg13g2_mux2_1 _23682_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][4] ),
    .A1(_05921_),
    .S(net348),
    .X(_01229_));
 sg13g2_buf_1 _23683_ (.A(_10831_),
    .X(_05922_));
 sg13g2_mux2_1 _23684_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][5] ),
    .A1(_05922_),
    .S(_05919_),
    .X(_01230_));
 sg13g2_mux2_1 _23685_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][6] ),
    .A1(net825),
    .S(_05919_),
    .X(_01231_));
 sg13g2_mux2_1 _23686_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][7] ),
    .A1(net824),
    .S(net348),
    .X(_01232_));
 sg13g2_mux2_1 _23687_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][8] ),
    .A1(_05907_),
    .S(_05918_),
    .X(_01233_));
 sg13g2_mux2_1 _23688_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][9] ),
    .A1(net481),
    .S(_05918_),
    .X(_01234_));
 sg13g2_buf_1 _23689_ (.A(net448),
    .X(_05923_));
 sg13g2_nor3_1 _23690_ (.A(net949),
    .B(net828),
    .C(_05900_),
    .Y(_05924_));
 sg13g2_buf_1 _23691_ (.A(_05924_),
    .X(_05925_));
 sg13g2_nor2b_1 _23692_ (.A(net484),
    .B_N(_05925_),
    .Y(_05926_));
 sg13g2_buf_1 _23693_ (.A(_05926_),
    .X(_05927_));
 sg13g2_buf_1 _23694_ (.A(_05927_),
    .X(_05928_));
 sg13g2_mux2_1 _23695_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][0] ),
    .A1(_05923_),
    .S(net347),
    .X(_01235_));
 sg13g2_mux2_1 _23696_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][10] ),
    .A1(net628),
    .S(net347),
    .X(_01236_));
 sg13g2_mux2_1 _23697_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][11] ),
    .A1(_05912_),
    .S(net347),
    .X(_01237_));
 sg13g2_mux2_1 _23698_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][1] ),
    .A1(net562),
    .S(net347),
    .X(_01238_));
 sg13g2_mux2_1 _23699_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][2] ),
    .A1(net823),
    .S(net347),
    .X(_01239_));
 sg13g2_buf_1 _23700_ (.A(_03096_),
    .X(_05929_));
 sg13g2_mux2_1 _23701_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][3] ),
    .A1(_05929_),
    .S(net347),
    .X(_01240_));
 sg13g2_mux2_1 _23702_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][4] ),
    .A1(net822),
    .S(net347),
    .X(_01241_));
 sg13g2_mux2_1 _23703_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][5] ),
    .A1(net947),
    .S(_05928_),
    .X(_01242_));
 sg13g2_buf_1 _23704_ (.A(net1095),
    .X(_05930_));
 sg13g2_mux2_1 _23705_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][6] ),
    .A1(_05930_),
    .S(_05928_),
    .X(_01243_));
 sg13g2_buf_1 _23706_ (.A(_10907_),
    .X(_05931_));
 sg13g2_mux2_1 _23707_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][7] ),
    .A1(_05931_),
    .S(net347),
    .X(_01244_));
 sg13g2_mux2_1 _23708_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][8] ),
    .A1(_05907_),
    .S(_05927_),
    .X(_01245_));
 sg13g2_mux2_1 _23709_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][9] ),
    .A1(net481),
    .S(_05927_),
    .X(_01246_));
 sg13g2_nor2_1 _23710_ (.A(_05852_),
    .B(_05887_),
    .Y(_05932_));
 sg13g2_buf_1 _23711_ (.A(_05932_),
    .X(_05933_));
 sg13g2_buf_1 _23712_ (.A(_05933_),
    .X(_05934_));
 sg13g2_mux2_1 _23713_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][0] ),
    .A1(_05923_),
    .S(net282),
    .X(_01247_));
 sg13g2_mux2_1 _23714_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][10] ),
    .A1(_05920_),
    .S(net282),
    .X(_01248_));
 sg13g2_mux2_1 _23715_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][11] ),
    .A1(_05912_),
    .S(net282),
    .X(_01249_));
 sg13g2_mux2_1 _23716_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][1] ),
    .A1(_05895_),
    .S(net282),
    .X(_01250_));
 sg13g2_mux2_1 _23717_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][2] ),
    .A1(net823),
    .S(net282),
    .X(_01251_));
 sg13g2_mux2_1 _23718_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][3] ),
    .A1(_05929_),
    .S(net282),
    .X(_01252_));
 sg13g2_mux2_1 _23719_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][4] ),
    .A1(_05921_),
    .S(net282),
    .X(_01253_));
 sg13g2_mux2_1 _23720_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][5] ),
    .A1(_05922_),
    .S(_05934_),
    .X(_01254_));
 sg13g2_mux2_1 _23721_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][6] ),
    .A1(_05930_),
    .S(_05934_),
    .X(_01255_));
 sg13g2_mux2_1 _23722_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][7] ),
    .A1(_05931_),
    .S(net282),
    .X(_01256_));
 sg13g2_mux2_1 _23723_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][8] ),
    .A1(net482),
    .S(_05933_),
    .X(_01257_));
 sg13g2_mux2_1 _23724_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][9] ),
    .A1(_05908_),
    .S(_05933_),
    .X(_01258_));
 sg13g2_or2_1 _23725_ (.X(_05935_),
    .B(_05900_),
    .A(_05849_));
 sg13g2_buf_1 _23726_ (.A(_05935_),
    .X(_05936_));
 sg13g2_nor2_1 _23727_ (.A(_05856_),
    .B(_05936_),
    .Y(_05937_));
 sg13g2_buf_1 _23728_ (.A(_05937_),
    .X(_05938_));
 sg13g2_buf_1 _23729_ (.A(_05938_),
    .X(_05939_));
 sg13g2_mux2_1 _23730_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][0] ),
    .A1(net400),
    .S(net281),
    .X(_01259_));
 sg13g2_mux2_1 _23731_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][10] ),
    .A1(net628),
    .S(net281),
    .X(_01260_));
 sg13g2_mux2_1 _23732_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][11] ),
    .A1(net629),
    .S(net281),
    .X(_01261_));
 sg13g2_mux2_1 _23733_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][1] ),
    .A1(net562),
    .S(net281),
    .X(_01262_));
 sg13g2_buf_1 _23734_ (.A(net966),
    .X(_05940_));
 sg13g2_mux2_1 _23735_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][2] ),
    .A1(_05940_),
    .S(_05939_),
    .X(_01263_));
 sg13g2_mux2_1 _23736_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][3] ),
    .A1(net821),
    .S(net281),
    .X(_01264_));
 sg13g2_mux2_1 _23737_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][4] ),
    .A1(net822),
    .S(net281),
    .X(_01265_));
 sg13g2_mux2_1 _23738_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][5] ),
    .A1(net947),
    .S(_05939_),
    .X(_01266_));
 sg13g2_mux2_1 _23739_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][6] ),
    .A1(net946),
    .S(net281),
    .X(_01267_));
 sg13g2_mux2_1 _23740_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][7] ),
    .A1(net945),
    .S(net281),
    .X(_01268_));
 sg13g2_mux2_1 _23741_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][8] ),
    .A1(net482),
    .S(_05938_),
    .X(_01269_));
 sg13g2_mux2_1 _23742_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][9] ),
    .A1(net481),
    .S(_05938_),
    .X(_01270_));
 sg13g2_nor2_1 _23743_ (.A(_05887_),
    .B(_05936_),
    .Y(_05941_));
 sg13g2_buf_1 _23744_ (.A(_05941_),
    .X(_05942_));
 sg13g2_buf_1 _23745_ (.A(_05942_),
    .X(_05943_));
 sg13g2_mux2_1 _23746_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][0] ),
    .A1(net400),
    .S(net280),
    .X(_01271_));
 sg13g2_mux2_1 _23747_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][10] ),
    .A1(net628),
    .S(net280),
    .X(_01272_));
 sg13g2_mux2_1 _23748_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][11] ),
    .A1(net629),
    .S(net280),
    .X(_01273_));
 sg13g2_mux2_1 _23749_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][1] ),
    .A1(net562),
    .S(net280),
    .X(_01274_));
 sg13g2_mux2_1 _23750_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][2] ),
    .A1(net820),
    .S(_05943_),
    .X(_01275_));
 sg13g2_mux2_1 _23751_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][3] ),
    .A1(net821),
    .S(net280),
    .X(_01276_));
 sg13g2_mux2_1 _23752_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][4] ),
    .A1(net822),
    .S(net280),
    .X(_01277_));
 sg13g2_mux2_1 _23753_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][5] ),
    .A1(net947),
    .S(_05943_),
    .X(_01278_));
 sg13g2_mux2_1 _23754_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][6] ),
    .A1(net946),
    .S(net280),
    .X(_01279_));
 sg13g2_mux2_1 _23755_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][7] ),
    .A1(net945),
    .S(net280),
    .X(_01280_));
 sg13g2_mux2_1 _23756_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][8] ),
    .A1(net482),
    .S(_05942_),
    .X(_01281_));
 sg13g2_mux2_1 _23757_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][9] ),
    .A1(net481),
    .S(_05942_),
    .X(_01282_));
 sg13g2_nor3_1 _23758_ (.A(net708),
    .B(net483),
    .C(_05936_),
    .Y(_05944_));
 sg13g2_buf_1 _23759_ (.A(_05944_),
    .X(_05945_));
 sg13g2_buf_1 _23760_ (.A(_05945_),
    .X(_05946_));
 sg13g2_mux2_1 _23761_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][0] ),
    .A1(net400),
    .S(net346),
    .X(_01283_));
 sg13g2_mux2_1 _23762_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][10] ),
    .A1(net628),
    .S(net346),
    .X(_01284_));
 sg13g2_mux2_1 _23763_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][11] ),
    .A1(net629),
    .S(net346),
    .X(_01285_));
 sg13g2_mux2_1 _23764_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][1] ),
    .A1(net562),
    .S(net346),
    .X(_01286_));
 sg13g2_mux2_1 _23765_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][2] ),
    .A1(net820),
    .S(_05946_),
    .X(_01287_));
 sg13g2_mux2_1 _23766_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][3] ),
    .A1(net821),
    .S(net346),
    .X(_01288_));
 sg13g2_mux2_1 _23767_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][4] ),
    .A1(net822),
    .S(net346),
    .X(_01289_));
 sg13g2_mux2_1 _23768_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][5] ),
    .A1(net947),
    .S(_05946_),
    .X(_01290_));
 sg13g2_mux2_1 _23769_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][6] ),
    .A1(net946),
    .S(net346),
    .X(_01291_));
 sg13g2_mux2_1 _23770_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][7] ),
    .A1(net945),
    .S(net346),
    .X(_01292_));
 sg13g2_mux2_1 _23771_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][8] ),
    .A1(net482),
    .S(_05945_),
    .X(_01293_));
 sg13g2_mux2_1 _23772_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][9] ),
    .A1(net481),
    .S(_05945_),
    .X(_01294_));
 sg13g2_nor3_1 _23773_ (.A(net828),
    .B(net483),
    .C(_05936_),
    .Y(_05947_));
 sg13g2_buf_1 _23774_ (.A(_05947_),
    .X(_05948_));
 sg13g2_buf_1 _23775_ (.A(_05948_),
    .X(_05949_));
 sg13g2_mux2_1 _23776_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][0] ),
    .A1(net400),
    .S(net345),
    .X(_01295_));
 sg13g2_mux2_1 _23777_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][10] ),
    .A1(net628),
    .S(net345),
    .X(_01296_));
 sg13g2_mux2_1 _23778_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][11] ),
    .A1(net629),
    .S(net345),
    .X(_01297_));
 sg13g2_buf_1 _23779_ (.A(_03107_),
    .X(_05950_));
 sg13g2_mux2_1 _23780_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][1] ),
    .A1(net561),
    .S(net345),
    .X(_01298_));
 sg13g2_mux2_1 _23781_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][2] ),
    .A1(_05940_),
    .S(_05949_),
    .X(_01299_));
 sg13g2_mux2_1 _23782_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][3] ),
    .A1(net821),
    .S(net345),
    .X(_01300_));
 sg13g2_mux2_1 _23783_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][4] ),
    .A1(net822),
    .S(net345),
    .X(_01301_));
 sg13g2_mux2_1 _23784_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][5] ),
    .A1(net947),
    .S(net345),
    .X(_01302_));
 sg13g2_mux2_1 _23785_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][6] ),
    .A1(net946),
    .S(_05949_),
    .X(_01303_));
 sg13g2_mux2_1 _23786_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][7] ),
    .A1(net945),
    .S(net345),
    .X(_01304_));
 sg13g2_mux2_1 _23787_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][8] ),
    .A1(net482),
    .S(_05948_),
    .X(_01305_));
 sg13g2_mux2_1 _23788_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][9] ),
    .A1(net481),
    .S(_05948_),
    .X(_01306_));
 sg13g2_buf_1 _23789_ (.A(_10079_),
    .X(_05951_));
 sg13g2_nand2_2 _23790_ (.Y(_05952_),
    .A(net944),
    .B(net948));
 sg13g2_nor3_1 _23791_ (.A(net483),
    .B(_05903_),
    .C(_05952_),
    .Y(_05953_));
 sg13g2_buf_1 _23792_ (.A(_05953_),
    .X(_05954_));
 sg13g2_buf_1 _23793_ (.A(_05954_),
    .X(_05955_));
 sg13g2_mux2_1 _23794_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][0] ),
    .A1(net400),
    .S(net344),
    .X(_01307_));
 sg13g2_mux2_1 _23795_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][10] ),
    .A1(net628),
    .S(net344),
    .X(_01308_));
 sg13g2_mux2_1 _23796_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][11] ),
    .A1(net629),
    .S(net344),
    .X(_01309_));
 sg13g2_mux2_1 _23797_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][1] ),
    .A1(net561),
    .S(net344),
    .X(_01310_));
 sg13g2_mux2_1 _23798_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][2] ),
    .A1(net820),
    .S(_05955_),
    .X(_01311_));
 sg13g2_mux2_1 _23799_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][3] ),
    .A1(net821),
    .S(net344),
    .X(_01312_));
 sg13g2_mux2_1 _23800_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][4] ),
    .A1(net822),
    .S(net344),
    .X(_01313_));
 sg13g2_mux2_1 _23801_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][5] ),
    .A1(net947),
    .S(_05955_),
    .X(_01314_));
 sg13g2_mux2_1 _23802_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][6] ),
    .A1(net946),
    .S(net344),
    .X(_01315_));
 sg13g2_mux2_1 _23803_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][7] ),
    .A1(net945),
    .S(net344),
    .X(_01316_));
 sg13g2_mux2_1 _23804_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][8] ),
    .A1(net482),
    .S(_05954_),
    .X(_01317_));
 sg13g2_mux2_1 _23805_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][9] ),
    .A1(net481),
    .S(_05954_),
    .X(_01318_));
 sg13g2_nor3_1 _23806_ (.A(net827),
    .B(_05887_),
    .C(_05952_),
    .Y(_05956_));
 sg13g2_buf_1 _23807_ (.A(_05956_),
    .X(_05957_));
 sg13g2_buf_1 _23808_ (.A(_05957_),
    .X(_05958_));
 sg13g2_mux2_1 _23809_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][0] ),
    .A1(net400),
    .S(net279),
    .X(_01319_));
 sg13g2_mux2_1 _23810_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][10] ),
    .A1(net628),
    .S(net279),
    .X(_01320_));
 sg13g2_mux2_1 _23811_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][11] ),
    .A1(net629),
    .S(net279),
    .X(_01321_));
 sg13g2_mux2_1 _23812_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][1] ),
    .A1(net561),
    .S(net279),
    .X(_01322_));
 sg13g2_mux2_1 _23813_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][2] ),
    .A1(net820),
    .S(net279),
    .X(_01323_));
 sg13g2_mux2_1 _23814_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][3] ),
    .A1(net821),
    .S(net279),
    .X(_01324_));
 sg13g2_mux2_1 _23815_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][4] ),
    .A1(net822),
    .S(net279),
    .X(_01325_));
 sg13g2_mux2_1 _23816_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][5] ),
    .A1(net947),
    .S(_05958_),
    .X(_01326_));
 sg13g2_mux2_1 _23817_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][6] ),
    .A1(net946),
    .S(_05958_),
    .X(_01327_));
 sg13g2_mux2_1 _23818_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][7] ),
    .A1(net945),
    .S(net279),
    .X(_01328_));
 sg13g2_buf_1 _23819_ (.A(net589),
    .X(_05959_));
 sg13g2_mux2_1 _23820_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][8] ),
    .A1(net480),
    .S(_05957_),
    .X(_01329_));
 sg13g2_buf_1 _23821_ (.A(net601),
    .X(_05960_));
 sg13g2_mux2_1 _23822_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][9] ),
    .A1(net479),
    .S(_05957_),
    .X(_01330_));
 sg13g2_nor2_2 _23823_ (.A(_05837_),
    .B(_05915_),
    .Y(_05961_));
 sg13g2_nor2b_1 _23824_ (.A(net484),
    .B_N(_05961_),
    .Y(_05962_));
 sg13g2_buf_1 _23825_ (.A(_05962_),
    .X(_05963_));
 sg13g2_buf_1 _23826_ (.A(_05963_),
    .X(_05964_));
 sg13g2_mux2_1 _23827_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][0] ),
    .A1(net400),
    .S(net343),
    .X(_01331_));
 sg13g2_mux2_1 _23828_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][10] ),
    .A1(net628),
    .S(net343),
    .X(_01332_));
 sg13g2_buf_1 _23829_ (.A(_11186_),
    .X(_05965_));
 sg13g2_mux2_1 _23830_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][11] ),
    .A1(net627),
    .S(net343),
    .X(_01333_));
 sg13g2_mux2_1 _23831_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][1] ),
    .A1(net561),
    .S(net343),
    .X(_01334_));
 sg13g2_mux2_1 _23832_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][2] ),
    .A1(net820),
    .S(net343),
    .X(_01335_));
 sg13g2_mux2_1 _23833_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][3] ),
    .A1(net821),
    .S(net343),
    .X(_01336_));
 sg13g2_mux2_1 _23834_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][4] ),
    .A1(net822),
    .S(net343),
    .X(_01337_));
 sg13g2_mux2_1 _23835_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][5] ),
    .A1(net947),
    .S(_05964_),
    .X(_01338_));
 sg13g2_mux2_1 _23836_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][6] ),
    .A1(net946),
    .S(_05964_),
    .X(_01339_));
 sg13g2_mux2_1 _23837_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][7] ),
    .A1(net945),
    .S(net343),
    .X(_01340_));
 sg13g2_mux2_1 _23838_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][8] ),
    .A1(net480),
    .S(_05963_),
    .X(_01341_));
 sg13g2_mux2_1 _23839_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][9] ),
    .A1(net479),
    .S(_05963_),
    .X(_01342_));
 sg13g2_nor3_1 _23840_ (.A(net949),
    .B(net828),
    .C(_05952_),
    .Y(_05966_));
 sg13g2_buf_2 _23841_ (.A(_05966_),
    .X(_05967_));
 sg13g2_nor2b_1 _23842_ (.A(net484),
    .B_N(_05967_),
    .Y(_05968_));
 sg13g2_buf_1 _23843_ (.A(_05968_),
    .X(_05969_));
 sg13g2_buf_1 _23844_ (.A(_05969_),
    .X(_05970_));
 sg13g2_mux2_1 _23845_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][0] ),
    .A1(net400),
    .S(net342),
    .X(_01343_));
 sg13g2_buf_1 _23846_ (.A(net732),
    .X(_05971_));
 sg13g2_mux2_1 _23847_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][10] ),
    .A1(net626),
    .S(net342),
    .X(_01344_));
 sg13g2_mux2_1 _23848_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][11] ),
    .A1(net627),
    .S(net342),
    .X(_01345_));
 sg13g2_mux2_1 _23849_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][1] ),
    .A1(net561),
    .S(net342),
    .X(_01346_));
 sg13g2_mux2_1 _23850_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][2] ),
    .A1(net820),
    .S(net342),
    .X(_01347_));
 sg13g2_mux2_1 _23851_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][3] ),
    .A1(net821),
    .S(net342),
    .X(_01348_));
 sg13g2_buf_1 _23852_ (.A(_09025_),
    .X(_05972_));
 sg13g2_mux2_1 _23853_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][4] ),
    .A1(net819),
    .S(net342),
    .X(_01349_));
 sg13g2_buf_1 _23854_ (.A(_10831_),
    .X(_05973_));
 sg13g2_mux2_1 _23855_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][5] ),
    .A1(net943),
    .S(_05970_),
    .X(_01350_));
 sg13g2_mux2_1 _23856_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][6] ),
    .A1(net946),
    .S(_05970_),
    .X(_01351_));
 sg13g2_mux2_1 _23857_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][7] ),
    .A1(net945),
    .S(net342),
    .X(_01352_));
 sg13g2_mux2_1 _23858_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][8] ),
    .A1(net480),
    .S(_05969_),
    .X(_01353_));
 sg13g2_mux2_1 _23859_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][9] ),
    .A1(net479),
    .S(_05969_),
    .X(_01354_));
 sg13g2_buf_1 _23860_ (.A(net448),
    .X(_05974_));
 sg13g2_or2_1 _23861_ (.X(_05975_),
    .B(_05952_),
    .A(_05849_));
 sg13g2_buf_1 _23862_ (.A(_05975_),
    .X(_05976_));
 sg13g2_nor2_1 _23863_ (.A(_05856_),
    .B(_05976_),
    .Y(_05977_));
 sg13g2_buf_1 _23864_ (.A(_05977_),
    .X(_05978_));
 sg13g2_buf_1 _23865_ (.A(_05978_),
    .X(_05979_));
 sg13g2_mux2_1 _23866_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][0] ),
    .A1(net399),
    .S(net278),
    .X(_01355_));
 sg13g2_mux2_1 _23867_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][10] ),
    .A1(net626),
    .S(net278),
    .X(_01356_));
 sg13g2_mux2_1 _23868_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][11] ),
    .A1(net627),
    .S(net278),
    .X(_01357_));
 sg13g2_mux2_1 _23869_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][1] ),
    .A1(net561),
    .S(net278),
    .X(_01358_));
 sg13g2_mux2_1 _23870_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][2] ),
    .A1(net820),
    .S(net278),
    .X(_01359_));
 sg13g2_buf_1 _23871_ (.A(_03096_),
    .X(_05980_));
 sg13g2_mux2_1 _23872_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][3] ),
    .A1(net818),
    .S(net278),
    .X(_01360_));
 sg13g2_mux2_1 _23873_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][4] ),
    .A1(net819),
    .S(net278),
    .X(_01361_));
 sg13g2_mux2_1 _23874_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][5] ),
    .A1(net943),
    .S(_05979_),
    .X(_01362_));
 sg13g2_buf_1 _23875_ (.A(_10963_),
    .X(_05981_));
 sg13g2_mux2_1 _23876_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][6] ),
    .A1(net942),
    .S(_05979_),
    .X(_01363_));
 sg13g2_buf_1 _23877_ (.A(_10907_),
    .X(_05982_));
 sg13g2_mux2_1 _23878_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][7] ),
    .A1(net941),
    .S(net278),
    .X(_01364_));
 sg13g2_mux2_1 _23879_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][8] ),
    .A1(net480),
    .S(_05978_),
    .X(_01365_));
 sg13g2_mux2_1 _23880_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][9] ),
    .A1(net479),
    .S(_05978_),
    .X(_01366_));
 sg13g2_nor2_1 _23881_ (.A(_05887_),
    .B(_05976_),
    .Y(_05983_));
 sg13g2_buf_1 _23882_ (.A(_05983_),
    .X(_05984_));
 sg13g2_buf_1 _23883_ (.A(_05984_),
    .X(_05985_));
 sg13g2_mux2_1 _23884_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][0] ),
    .A1(net399),
    .S(net277),
    .X(_01367_));
 sg13g2_mux2_1 _23885_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][10] ),
    .A1(net626),
    .S(net277),
    .X(_01368_));
 sg13g2_mux2_1 _23886_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][11] ),
    .A1(net627),
    .S(net277),
    .X(_01369_));
 sg13g2_mux2_1 _23887_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][1] ),
    .A1(net561),
    .S(net277),
    .X(_01370_));
 sg13g2_mux2_1 _23888_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][2] ),
    .A1(net820),
    .S(net277),
    .X(_01371_));
 sg13g2_mux2_1 _23889_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][3] ),
    .A1(net818),
    .S(net277),
    .X(_01372_));
 sg13g2_mux2_1 _23890_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][4] ),
    .A1(net819),
    .S(net277),
    .X(_01373_));
 sg13g2_mux2_1 _23891_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][5] ),
    .A1(net943),
    .S(_05985_),
    .X(_01374_));
 sg13g2_mux2_1 _23892_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][6] ),
    .A1(net942),
    .S(_05985_),
    .X(_01375_));
 sg13g2_mux2_1 _23893_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][7] ),
    .A1(net941),
    .S(net277),
    .X(_01376_));
 sg13g2_mux2_1 _23894_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][8] ),
    .A1(net480),
    .S(_05984_),
    .X(_01377_));
 sg13g2_mux2_1 _23895_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][9] ),
    .A1(net479),
    .S(_05984_),
    .X(_01378_));
 sg13g2_nor3_1 _23896_ (.A(net708),
    .B(_05852_),
    .C(_05863_),
    .Y(_05986_));
 sg13g2_buf_1 _23897_ (.A(_05986_),
    .X(_05987_));
 sg13g2_buf_1 _23898_ (.A(_05987_),
    .X(_05988_));
 sg13g2_mux2_1 _23899_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][0] ),
    .A1(net399),
    .S(net341),
    .X(_01379_));
 sg13g2_mux2_1 _23900_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][10] ),
    .A1(net626),
    .S(net341),
    .X(_01380_));
 sg13g2_mux2_1 _23901_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][11] ),
    .A1(net627),
    .S(net341),
    .X(_01381_));
 sg13g2_mux2_1 _23902_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][1] ),
    .A1(_05950_),
    .S(net341),
    .X(_01382_));
 sg13g2_buf_1 _23903_ (.A(_03093_),
    .X(_05989_));
 sg13g2_mux2_1 _23904_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][2] ),
    .A1(_05989_),
    .S(net341),
    .X(_01383_));
 sg13g2_mux2_1 _23905_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][3] ),
    .A1(net818),
    .S(net341),
    .X(_01384_));
 sg13g2_mux2_1 _23906_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][4] ),
    .A1(net819),
    .S(net341),
    .X(_01385_));
 sg13g2_mux2_1 _23907_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][5] ),
    .A1(net943),
    .S(_05988_),
    .X(_01386_));
 sg13g2_mux2_1 _23908_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][6] ),
    .A1(net942),
    .S(_05988_),
    .X(_01387_));
 sg13g2_mux2_1 _23909_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][7] ),
    .A1(net941),
    .S(net341),
    .X(_01388_));
 sg13g2_mux2_1 _23910_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][8] ),
    .A1(_05959_),
    .S(_05987_),
    .X(_01389_));
 sg13g2_mux2_1 _23911_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][9] ),
    .A1(_05960_),
    .S(_05987_),
    .X(_01390_));
 sg13g2_nor3_1 _23912_ (.A(net708),
    .B(net483),
    .C(_05976_),
    .Y(_05990_));
 sg13g2_buf_1 _23913_ (.A(_05990_),
    .X(_05991_));
 sg13g2_buf_1 _23914_ (.A(_05991_),
    .X(_05992_));
 sg13g2_mux2_1 _23915_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][0] ),
    .A1(net399),
    .S(net340),
    .X(_01391_));
 sg13g2_mux2_1 _23916_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][10] ),
    .A1(net626),
    .S(net340),
    .X(_01392_));
 sg13g2_mux2_1 _23917_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][11] ),
    .A1(net627),
    .S(net340),
    .X(_01393_));
 sg13g2_mux2_1 _23918_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][1] ),
    .A1(_05950_),
    .S(net340),
    .X(_01394_));
 sg13g2_mux2_1 _23919_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][2] ),
    .A1(net817),
    .S(net340),
    .X(_01395_));
 sg13g2_mux2_1 _23920_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][3] ),
    .A1(net818),
    .S(net340),
    .X(_01396_));
 sg13g2_mux2_1 _23921_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][4] ),
    .A1(net819),
    .S(net340),
    .X(_01397_));
 sg13g2_mux2_1 _23922_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][5] ),
    .A1(net943),
    .S(_05992_),
    .X(_01398_));
 sg13g2_mux2_1 _23923_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][6] ),
    .A1(_05981_),
    .S(_05992_),
    .X(_01399_));
 sg13g2_mux2_1 _23924_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][7] ),
    .A1(net941),
    .S(net340),
    .X(_01400_));
 sg13g2_mux2_1 _23925_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][8] ),
    .A1(net480),
    .S(_05991_),
    .X(_01401_));
 sg13g2_mux2_1 _23926_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][9] ),
    .A1(net479),
    .S(_05991_),
    .X(_01402_));
 sg13g2_nor3_1 _23927_ (.A(net828),
    .B(net483),
    .C(_05976_),
    .Y(_05993_));
 sg13g2_buf_1 _23928_ (.A(_05993_),
    .X(_05994_));
 sg13g2_buf_1 _23929_ (.A(_05994_),
    .X(_05995_));
 sg13g2_mux2_1 _23930_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][0] ),
    .A1(net399),
    .S(net339),
    .X(_01403_));
 sg13g2_mux2_1 _23931_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][10] ),
    .A1(net626),
    .S(net339),
    .X(_01404_));
 sg13g2_mux2_1 _23932_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][11] ),
    .A1(net627),
    .S(net339),
    .X(_01405_));
 sg13g2_mux2_1 _23933_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][1] ),
    .A1(net561),
    .S(net339),
    .X(_01406_));
 sg13g2_mux2_1 _23934_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][2] ),
    .A1(net817),
    .S(net339),
    .X(_01407_));
 sg13g2_mux2_1 _23935_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][3] ),
    .A1(net818),
    .S(net339),
    .X(_01408_));
 sg13g2_mux2_1 _23936_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][4] ),
    .A1(net819),
    .S(net339),
    .X(_01409_));
 sg13g2_mux2_1 _23937_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][5] ),
    .A1(net943),
    .S(_05995_),
    .X(_01410_));
 sg13g2_mux2_1 _23938_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][6] ),
    .A1(_05981_),
    .S(_05995_),
    .X(_01411_));
 sg13g2_mux2_1 _23939_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][7] ),
    .A1(net941),
    .S(net339),
    .X(_01412_));
 sg13g2_mux2_1 _23940_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][8] ),
    .A1(net480),
    .S(_05994_),
    .X(_01413_));
 sg13g2_mux2_1 _23941_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][9] ),
    .A1(net479),
    .S(_05994_),
    .X(_01414_));
 sg13g2_nor3_1 _23942_ (.A(net828),
    .B(_05852_),
    .C(net483),
    .Y(_05996_));
 sg13g2_buf_1 _23943_ (.A(_05996_),
    .X(_05997_));
 sg13g2_buf_1 _23944_ (.A(_05997_),
    .X(_05998_));
 sg13g2_mux2_1 _23945_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][0] ),
    .A1(_05974_),
    .S(net338),
    .X(_01415_));
 sg13g2_mux2_1 _23946_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][10] ),
    .A1(net626),
    .S(net338),
    .X(_01416_));
 sg13g2_mux2_1 _23947_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][11] ),
    .A1(net627),
    .S(net338),
    .X(_01417_));
 sg13g2_mux2_1 _23948_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][1] ),
    .A1(net579),
    .S(net338),
    .X(_01418_));
 sg13g2_mux2_1 _23949_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][2] ),
    .A1(_05989_),
    .S(net338),
    .X(_01419_));
 sg13g2_mux2_1 _23950_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][3] ),
    .A1(net818),
    .S(net338),
    .X(_01420_));
 sg13g2_mux2_1 _23951_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][4] ),
    .A1(net819),
    .S(net338),
    .X(_01421_));
 sg13g2_mux2_1 _23952_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][5] ),
    .A1(net943),
    .S(_05998_),
    .X(_01422_));
 sg13g2_mux2_1 _23953_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][6] ),
    .A1(net942),
    .S(_05998_),
    .X(_01423_));
 sg13g2_mux2_1 _23954_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][7] ),
    .A1(_05982_),
    .S(net338),
    .X(_01424_));
 sg13g2_mux2_1 _23955_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][8] ),
    .A1(net480),
    .S(_05997_),
    .X(_01425_));
 sg13g2_mux2_1 _23956_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][9] ),
    .A1(net479),
    .S(_05997_),
    .X(_01426_));
 sg13g2_nand2_1 _23957_ (.Y(_05999_),
    .A(_11062_),
    .B(_05851_));
 sg13g2_nor2_1 _23958_ (.A(_05856_),
    .B(_05999_),
    .Y(_06000_));
 sg13g2_buf_1 _23959_ (.A(_06000_),
    .X(_06001_));
 sg13g2_buf_1 _23960_ (.A(_06001_),
    .X(_06002_));
 sg13g2_mux2_1 _23961_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][0] ),
    .A1(_05974_),
    .S(net276),
    .X(_01427_));
 sg13g2_mux2_1 _23962_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][10] ),
    .A1(net626),
    .S(net276),
    .X(_01428_));
 sg13g2_mux2_1 _23963_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][11] ),
    .A1(_05965_),
    .S(_06002_),
    .X(_01429_));
 sg13g2_mux2_1 _23964_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][1] ),
    .A1(net579),
    .S(net276),
    .X(_01430_));
 sg13g2_mux2_1 _23965_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][2] ),
    .A1(net817),
    .S(_06002_),
    .X(_01431_));
 sg13g2_mux2_1 _23966_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][3] ),
    .A1(_05980_),
    .S(net276),
    .X(_01432_));
 sg13g2_mux2_1 _23967_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][4] ),
    .A1(net819),
    .S(net276),
    .X(_01433_));
 sg13g2_mux2_1 _23968_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][5] ),
    .A1(net943),
    .S(net276),
    .X(_01434_));
 sg13g2_mux2_1 _23969_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][6] ),
    .A1(net942),
    .S(net276),
    .X(_01435_));
 sg13g2_mux2_1 _23970_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][7] ),
    .A1(net941),
    .S(net276),
    .X(_01436_));
 sg13g2_mux2_1 _23971_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][8] ),
    .A1(_05959_),
    .S(_06001_),
    .X(_01437_));
 sg13g2_mux2_1 _23972_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][9] ),
    .A1(_05960_),
    .S(_06001_),
    .X(_01438_));
 sg13g2_nor2_1 _23973_ (.A(_05885_),
    .B(_05999_),
    .Y(_06003_));
 sg13g2_buf_2 _23974_ (.A(_06003_),
    .X(_06004_));
 sg13g2_nor2b_1 _23975_ (.A(net484),
    .B_N(_06004_),
    .Y(_06005_));
 sg13g2_buf_1 _23976_ (.A(_06005_),
    .X(_06006_));
 sg13g2_buf_1 _23977_ (.A(_06006_),
    .X(_06007_));
 sg13g2_mux2_1 _23978_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][0] ),
    .A1(net399),
    .S(net337),
    .X(_01439_));
 sg13g2_mux2_1 _23979_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][10] ),
    .A1(_05971_),
    .S(net337),
    .X(_01440_));
 sg13g2_mux2_1 _23980_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][11] ),
    .A1(_05965_),
    .S(_06007_),
    .X(_01441_));
 sg13g2_mux2_1 _23981_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][1] ),
    .A1(net579),
    .S(net337),
    .X(_01442_));
 sg13g2_mux2_1 _23982_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][2] ),
    .A1(net817),
    .S(net337),
    .X(_01443_));
 sg13g2_mux2_1 _23983_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][3] ),
    .A1(_05980_),
    .S(net337),
    .X(_01444_));
 sg13g2_mux2_1 _23984_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][4] ),
    .A1(_05972_),
    .S(net337),
    .X(_01445_));
 sg13g2_mux2_1 _23985_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][5] ),
    .A1(_05973_),
    .S(net337),
    .X(_01446_));
 sg13g2_mux2_1 _23986_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][6] ),
    .A1(net942),
    .S(_06007_),
    .X(_01447_));
 sg13g2_mux2_1 _23987_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][7] ),
    .A1(net941),
    .S(net337),
    .X(_01448_));
 sg13g2_mux2_1 _23988_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][8] ),
    .A1(net504),
    .S(_06006_),
    .X(_01449_));
 sg13g2_mux2_1 _23989_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][9] ),
    .A1(net503),
    .S(_06006_),
    .X(_01450_));
 sg13g2_nor2b_1 _23990_ (.A(_11010_),
    .B_N(net951),
    .Y(_06008_));
 sg13g2_buf_1 _23991_ (.A(_06008_),
    .X(_06009_));
 sg13g2_nand2_2 _23992_ (.Y(_06010_),
    .A(net949),
    .B(_06009_));
 sg13g2_nor3_2 _23993_ (.A(net944),
    .B(net948),
    .C(_06010_),
    .Y(_06011_));
 sg13g2_nor2b_1 _23994_ (.A(net484),
    .B_N(_06011_),
    .Y(_06012_));
 sg13g2_buf_1 _23995_ (.A(_06012_),
    .X(_06013_));
 sg13g2_buf_1 _23996_ (.A(_06013_),
    .X(_06014_));
 sg13g2_mux2_1 _23997_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][0] ),
    .A1(net399),
    .S(net336),
    .X(_01451_));
 sg13g2_mux2_1 _23998_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][10] ),
    .A1(_05971_),
    .S(net336),
    .X(_01452_));
 sg13g2_mux2_1 _23999_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][11] ),
    .A1(net638),
    .S(net336),
    .X(_01453_));
 sg13g2_mux2_1 _24000_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][1] ),
    .A1(net579),
    .S(net336),
    .X(_01454_));
 sg13g2_mux2_1 _24001_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][2] ),
    .A1(net817),
    .S(net336),
    .X(_01455_));
 sg13g2_mux2_1 _24002_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][3] ),
    .A1(net818),
    .S(net336),
    .X(_01456_));
 sg13g2_mux2_1 _24003_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][4] ),
    .A1(_05972_),
    .S(net336),
    .X(_01457_));
 sg13g2_mux2_1 _24004_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][5] ),
    .A1(_05973_),
    .S(_06014_),
    .X(_01458_));
 sg13g2_mux2_1 _24005_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][6] ),
    .A1(net942),
    .S(_06014_),
    .X(_01459_));
 sg13g2_mux2_1 _24006_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][7] ),
    .A1(net941),
    .S(net336),
    .X(_01460_));
 sg13g2_mux2_1 _24007_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][8] ),
    .A1(net504),
    .S(_06013_),
    .X(_01461_));
 sg13g2_mux2_1 _24008_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][9] ),
    .A1(net503),
    .S(_06013_),
    .X(_01462_));
 sg13g2_nor2_1 _24009_ (.A(net828),
    .B(_05999_),
    .Y(_06015_));
 sg13g2_buf_2 _24010_ (.A(_06015_),
    .X(_06016_));
 sg13g2_nor2b_1 _24011_ (.A(_05863_),
    .B_N(_06016_),
    .Y(_06017_));
 sg13g2_buf_1 _24012_ (.A(_06017_),
    .X(_06018_));
 sg13g2_buf_1 _24013_ (.A(_06018_),
    .X(_06019_));
 sg13g2_mux2_1 _24014_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][0] ),
    .A1(net399),
    .S(net335),
    .X(_01463_));
 sg13g2_mux2_1 _24015_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][10] ),
    .A1(net639),
    .S(net335),
    .X(_01464_));
 sg13g2_mux2_1 _24016_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][11] ),
    .A1(net638),
    .S(net335),
    .X(_01465_));
 sg13g2_mux2_1 _24017_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][1] ),
    .A1(net579),
    .S(net335),
    .X(_01466_));
 sg13g2_mux2_1 _24018_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][2] ),
    .A1(net817),
    .S(_06019_),
    .X(_01467_));
 sg13g2_mux2_1 _24019_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][3] ),
    .A1(net818),
    .S(net335),
    .X(_01468_));
 sg13g2_mux2_1 _24020_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][4] ),
    .A1(net845),
    .S(net335),
    .X(_01469_));
 sg13g2_mux2_1 _24021_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][5] ),
    .A1(net964),
    .S(_06019_),
    .X(_01470_));
 sg13g2_mux2_1 _24022_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][6] ),
    .A1(net942),
    .S(net335),
    .X(_01471_));
 sg13g2_mux2_1 _24023_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][7] ),
    .A1(_05982_),
    .S(net335),
    .X(_01472_));
 sg13g2_mux2_1 _24024_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][8] ),
    .A1(net504),
    .S(_06018_),
    .X(_01473_));
 sg13g2_mux2_1 _24025_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][9] ),
    .A1(net503),
    .S(_06018_),
    .X(_01474_));
 sg13g2_nor3_1 _24026_ (.A(_05891_),
    .B(_05867_),
    .C(_05903_),
    .Y(_06020_));
 sg13g2_buf_1 _24027_ (.A(_06020_),
    .X(_06021_));
 sg13g2_buf_1 _24028_ (.A(_06021_),
    .X(_06022_));
 sg13g2_mux2_1 _24029_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][0] ),
    .A1(_03657_),
    .S(net334),
    .X(_01475_));
 sg13g2_mux2_1 _24030_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][10] ),
    .A1(_03646_),
    .S(net334),
    .X(_01476_));
 sg13g2_mux2_1 _24031_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][11] ),
    .A1(_03648_),
    .S(net334),
    .X(_01477_));
 sg13g2_mux2_1 _24032_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][1] ),
    .A1(_03108_),
    .S(net334),
    .X(_01478_));
 sg13g2_mux2_1 _24033_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][2] ),
    .A1(net817),
    .S(net334),
    .X(_01479_));
 sg13g2_mux2_1 _24034_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][3] ),
    .A1(net846),
    .S(net334),
    .X(_01480_));
 sg13g2_mux2_1 _24035_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][4] ),
    .A1(net845),
    .S(net334),
    .X(_01481_));
 sg13g2_mux2_1 _24036_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][5] ),
    .A1(net964),
    .S(_06022_),
    .X(_01482_));
 sg13g2_mux2_1 _24037_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][6] ),
    .A1(net963),
    .S(_06022_),
    .X(_01483_));
 sg13g2_mux2_1 _24038_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][7] ),
    .A1(net962),
    .S(net334),
    .X(_01484_));
 sg13g2_mux2_1 _24039_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][8] ),
    .A1(net504),
    .S(_06021_),
    .X(_01485_));
 sg13g2_mux2_1 _24040_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][9] ),
    .A1(_03644_),
    .S(_06021_),
    .X(_01486_));
 sg13g2_nor3_1 _24041_ (.A(net827),
    .B(_05867_),
    .C(_05887_),
    .Y(_06023_));
 sg13g2_buf_1 _24042_ (.A(_06023_),
    .X(_06024_));
 sg13g2_buf_1 _24043_ (.A(_06024_),
    .X(_06025_));
 sg13g2_mux2_1 _24044_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][0] ),
    .A1(net448),
    .S(net275),
    .X(_01487_));
 sg13g2_mux2_1 _24045_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][10] ),
    .A1(_03646_),
    .S(net275),
    .X(_01488_));
 sg13g2_mux2_1 _24046_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][11] ),
    .A1(_03648_),
    .S(net275),
    .X(_01489_));
 sg13g2_mux2_1 _24047_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][1] ),
    .A1(_03108_),
    .S(net275),
    .X(_01490_));
 sg13g2_mux2_1 _24048_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][2] ),
    .A1(net817),
    .S(net275),
    .X(_01491_));
 sg13g2_mux2_1 _24049_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][3] ),
    .A1(_03097_),
    .S(net275),
    .X(_01492_));
 sg13g2_mux2_1 _24050_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][4] ),
    .A1(_03099_),
    .S(net275),
    .X(_01493_));
 sg13g2_mux2_1 _24051_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][5] ),
    .A1(_03101_),
    .S(_06025_),
    .X(_01494_));
 sg13g2_mux2_1 _24052_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][6] ),
    .A1(_03103_),
    .S(_06025_),
    .X(_01495_));
 sg13g2_mux2_1 _24053_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][7] ),
    .A1(_03105_),
    .S(net275),
    .X(_01496_));
 sg13g2_mux2_1 _24054_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][8] ),
    .A1(net504),
    .S(_06024_),
    .X(_01497_));
 sg13g2_mux2_1 _24055_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][9] ),
    .A1(_03644_),
    .S(_06024_),
    .X(_01498_));
 sg13g2_and2_1 _24056_ (.A(_05849_),
    .B(_05851_),
    .X(_06026_));
 sg13g2_buf_1 _24057_ (.A(_06026_),
    .X(_06027_));
 sg13g2_and3_1 _24058_ (.X(_06028_),
    .A(net1118),
    .B(_10382_),
    .C(_05798_));
 sg13g2_buf_1 _24059_ (.A(_06028_),
    .X(_06029_));
 sg13g2_and2_1 _24060_ (.A(_05817_),
    .B(_06029_),
    .X(_06030_));
 sg13g2_buf_1 _24061_ (.A(_06030_),
    .X(_06031_));
 sg13g2_nand2_1 _24062_ (.Y(_06032_),
    .A(_06027_),
    .B(_06031_));
 sg13g2_buf_2 _24063_ (.A(_06032_),
    .X(_06033_));
 sg13g2_buf_1 _24064_ (.A(_06033_),
    .X(_06034_));
 sg13g2_nand2_1 _24065_ (.Y(_06035_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][0] ),
    .B(_06033_));
 sg13g2_o21ai_1 _24066_ (.B1(_06035_),
    .Y(_01499_),
    .A1(net495),
    .A2(net274));
 sg13g2_mux2_1 _24067_ (.A0(net568),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][10] ),
    .S(net274),
    .X(_01500_));
 sg13g2_mux2_1 _24068_ (.A0(net567),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][11] ),
    .S(_06034_),
    .X(_01501_));
 sg13g2_nand2_1 _24069_ (.Y(_06036_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][1] ),
    .B(_06033_));
 sg13g2_o21ai_1 _24070_ (.B1(_06036_),
    .Y(_01502_),
    .A1(net641),
    .A2(_06034_));
 sg13g2_mux2_1 _24071_ (.A0(net717),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][2] ),
    .S(net274),
    .X(_01503_));
 sg13g2_mux2_1 _24072_ (.A0(net716),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][3] ),
    .S(net274),
    .X(_01504_));
 sg13g2_mux2_1 _24073_ (.A0(net715),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][4] ),
    .S(net274),
    .X(_01505_));
 sg13g2_mux2_1 _24074_ (.A0(net844),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][5] ),
    .S(net274),
    .X(_01506_));
 sg13g2_mux2_1 _24075_ (.A0(net843),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][6] ),
    .S(net274),
    .X(_01507_));
 sg13g2_mux2_1 _24076_ (.A0(net842),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][7] ),
    .S(net274),
    .X(_01508_));
 sg13g2_mux2_1 _24077_ (.A0(net446),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][8] ),
    .S(_06033_),
    .X(_01509_));
 sg13g2_mux2_1 _24078_ (.A0(net445),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][9] ),
    .S(_06033_),
    .X(_01510_));
 sg13g2_buf_1 _24079_ (.A(_06029_),
    .X(_06037_));
 sg13g2_nand2_1 _24080_ (.Y(_06038_),
    .A(_05868_),
    .B(net478));
 sg13g2_buf_2 _24081_ (.A(_06038_),
    .X(_06039_));
 sg13g2_buf_1 _24082_ (.A(_06039_),
    .X(_06040_));
 sg13g2_nand2_1 _24083_ (.Y(_06041_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][0] ),
    .B(_06039_));
 sg13g2_o21ai_1 _24084_ (.B1(_06041_),
    .Y(_01511_),
    .A1(net495),
    .A2(_06040_));
 sg13g2_mux2_1 _24085_ (.A0(net568),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][10] ),
    .S(net333),
    .X(_01512_));
 sg13g2_mux2_1 _24086_ (.A0(net567),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][11] ),
    .S(_06040_),
    .X(_01513_));
 sg13g2_nand2_1 _24087_ (.Y(_06042_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][1] ),
    .B(_06039_));
 sg13g2_o21ai_1 _24088_ (.B1(_06042_),
    .Y(_01514_),
    .A1(net641),
    .A2(net333));
 sg13g2_mux2_1 _24089_ (.A0(_03095_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][2] ),
    .S(net333),
    .X(_01515_));
 sg13g2_mux2_1 _24090_ (.A0(net716),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][3] ),
    .S(net333),
    .X(_01516_));
 sg13g2_mux2_1 _24091_ (.A0(net715),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][4] ),
    .S(net333),
    .X(_01517_));
 sg13g2_mux2_1 _24092_ (.A0(net844),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][5] ),
    .S(net333),
    .X(_01518_));
 sg13g2_mux2_1 _24093_ (.A0(net843),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][6] ),
    .S(net333),
    .X(_01519_));
 sg13g2_mux2_1 _24094_ (.A0(_03106_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][7] ),
    .S(net333),
    .X(_01520_));
 sg13g2_mux2_1 _24095_ (.A0(net446),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][8] ),
    .S(_06039_),
    .X(_01521_));
 sg13g2_mux2_1 _24096_ (.A0(_03712_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][9] ),
    .S(_06039_),
    .X(_01522_));
 sg13g2_nand2_1 _24097_ (.Y(_06043_),
    .A(_05873_),
    .B(net478));
 sg13g2_buf_2 _24098_ (.A(_06043_),
    .X(_06044_));
 sg13g2_buf_1 _24099_ (.A(_06044_),
    .X(_06045_));
 sg13g2_nand2_1 _24100_ (.Y(_06046_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][0] ),
    .B(_06044_));
 sg13g2_o21ai_1 _24101_ (.B1(_06046_),
    .Y(_01523_),
    .A1(_03718_),
    .A2(_06045_));
 sg13g2_mux2_1 _24102_ (.A0(_03713_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][10] ),
    .S(net332),
    .X(_01524_));
 sg13g2_mux2_1 _24103_ (.A0(net567),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][11] ),
    .S(_06045_),
    .X(_01525_));
 sg13g2_nand2_1 _24104_ (.Y(_06047_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][1] ),
    .B(_06044_));
 sg13g2_o21ai_1 _24105_ (.B1(_06047_),
    .Y(_01526_),
    .A1(net641),
    .A2(net332));
 sg13g2_mux2_1 _24106_ (.A0(net717),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][2] ),
    .S(net332),
    .X(_01527_));
 sg13g2_mux2_1 _24107_ (.A0(net716),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][3] ),
    .S(net332),
    .X(_01528_));
 sg13g2_mux2_1 _24108_ (.A0(net715),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][4] ),
    .S(net332),
    .X(_01529_));
 sg13g2_mux2_1 _24109_ (.A0(net844),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][5] ),
    .S(net332),
    .X(_01530_));
 sg13g2_mux2_1 _24110_ (.A0(net843),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][6] ),
    .S(net332),
    .X(_01531_));
 sg13g2_mux2_1 _24111_ (.A0(_03106_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][7] ),
    .S(net332),
    .X(_01532_));
 sg13g2_mux2_1 _24112_ (.A0(net446),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][8] ),
    .S(_06044_),
    .X(_01533_));
 sg13g2_mux2_1 _24113_ (.A0(net445),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][9] ),
    .S(_06044_),
    .X(_01534_));
 sg13g2_nor2_1 _24114_ (.A(_05849_),
    .B(_05867_),
    .Y(_06048_));
 sg13g2_nand2_1 _24115_ (.Y(_06049_),
    .A(_06048_),
    .B(_06031_));
 sg13g2_buf_2 _24116_ (.A(_06049_),
    .X(_06050_));
 sg13g2_buf_1 _24117_ (.A(_06050_),
    .X(_06051_));
 sg13g2_nand2_1 _24118_ (.Y(_06052_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][0] ),
    .B(_06050_));
 sg13g2_o21ai_1 _24119_ (.B1(_06052_),
    .Y(_01535_),
    .A1(net495),
    .A2(_06051_));
 sg13g2_mux2_1 _24120_ (.A0(net568),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][10] ),
    .S(net273),
    .X(_01536_));
 sg13g2_mux2_1 _24121_ (.A0(net567),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][11] ),
    .S(_06051_),
    .X(_01537_));
 sg13g2_nand2_1 _24122_ (.Y(_06053_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][1] ),
    .B(_06050_));
 sg13g2_o21ai_1 _24123_ (.B1(_06053_),
    .Y(_01538_),
    .A1(net641),
    .A2(net273));
 sg13g2_mux2_1 _24124_ (.A0(net717),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][2] ),
    .S(net273),
    .X(_01539_));
 sg13g2_mux2_1 _24125_ (.A0(net716),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][3] ),
    .S(net273),
    .X(_01540_));
 sg13g2_mux2_1 _24126_ (.A0(net715),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][4] ),
    .S(net273),
    .X(_01541_));
 sg13g2_mux2_1 _24127_ (.A0(net844),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][5] ),
    .S(net273),
    .X(_01542_));
 sg13g2_mux2_1 _24128_ (.A0(net843),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][6] ),
    .S(net273),
    .X(_01543_));
 sg13g2_mux2_1 _24129_ (.A0(net842),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][7] ),
    .S(net273),
    .X(_01544_));
 sg13g2_mux2_1 _24130_ (.A0(net446),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][8] ),
    .S(_06050_),
    .X(_01545_));
 sg13g2_mux2_1 _24131_ (.A0(net445),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][9] ),
    .S(_06050_),
    .X(_01546_));
 sg13g2_nor2b_1 _24132_ (.A(_05885_),
    .B_N(_06029_),
    .Y(_06054_));
 sg13g2_buf_2 _24133_ (.A(_06054_),
    .X(_06055_));
 sg13g2_nand2_1 _24134_ (.Y(_06056_),
    .A(_06048_),
    .B(_06055_));
 sg13g2_buf_2 _24135_ (.A(_06056_),
    .X(_06057_));
 sg13g2_buf_1 _24136_ (.A(_06057_),
    .X(_06058_));
 sg13g2_nand2_1 _24137_ (.Y(_06059_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][0] ),
    .B(_06057_));
 sg13g2_o21ai_1 _24138_ (.B1(_06059_),
    .Y(_01547_),
    .A1(net495),
    .A2(_06058_));
 sg13g2_mux2_1 _24139_ (.A0(net568),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][10] ),
    .S(net272),
    .X(_01548_));
 sg13g2_mux2_1 _24140_ (.A0(net567),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][11] ),
    .S(_06058_),
    .X(_01549_));
 sg13g2_nand2_1 _24141_ (.Y(_06060_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][1] ),
    .B(_06057_));
 sg13g2_o21ai_1 _24142_ (.B1(_06060_),
    .Y(_01550_),
    .A1(net641),
    .A2(net272));
 sg13g2_mux2_1 _24143_ (.A0(net717),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][2] ),
    .S(net272),
    .X(_01551_));
 sg13g2_mux2_1 _24144_ (.A0(net716),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][3] ),
    .S(net272),
    .X(_01552_));
 sg13g2_mux2_1 _24145_ (.A0(net715),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][4] ),
    .S(net272),
    .X(_01553_));
 sg13g2_mux2_1 _24146_ (.A0(net844),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][5] ),
    .S(net272),
    .X(_01554_));
 sg13g2_mux2_1 _24147_ (.A0(net843),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][6] ),
    .S(net272),
    .X(_01555_));
 sg13g2_mux2_1 _24148_ (.A0(net842),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][7] ),
    .S(net272),
    .X(_01556_));
 sg13g2_mux2_1 _24149_ (.A0(net446),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][8] ),
    .S(_06057_),
    .X(_01557_));
 sg13g2_mux2_1 _24150_ (.A0(net445),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][9] ),
    .S(_06057_),
    .X(_01558_));
 sg13g2_nand3_1 _24151_ (.B(_06048_),
    .C(net478),
    .A(_06009_),
    .Y(_06061_));
 sg13g2_buf_2 _24152_ (.A(_06061_),
    .X(_06062_));
 sg13g2_buf_1 _24153_ (.A(_06062_),
    .X(_06063_));
 sg13g2_nand2_1 _24154_ (.Y(_06064_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][0] ),
    .B(_06062_));
 sg13g2_o21ai_1 _24155_ (.B1(_06064_),
    .Y(_01559_),
    .A1(net495),
    .A2(_06063_));
 sg13g2_mux2_1 _24156_ (.A0(net568),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][10] ),
    .S(net331),
    .X(_01560_));
 sg13g2_mux2_1 _24157_ (.A0(_03714_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][11] ),
    .S(_06063_),
    .X(_01561_));
 sg13g2_nand2_1 _24158_ (.Y(_06065_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][1] ),
    .B(_06062_));
 sg13g2_o21ai_1 _24159_ (.B1(_06065_),
    .Y(_01562_),
    .A1(net641),
    .A2(net331));
 sg13g2_mux2_1 _24160_ (.A0(net717),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][2] ),
    .S(net331),
    .X(_01563_));
 sg13g2_mux2_1 _24161_ (.A0(_03098_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][3] ),
    .S(net331),
    .X(_01564_));
 sg13g2_mux2_1 _24162_ (.A0(_03100_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][4] ),
    .S(net331),
    .X(_01565_));
 sg13g2_mux2_1 _24163_ (.A0(net844),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][5] ),
    .S(net331),
    .X(_01566_));
 sg13g2_mux2_1 _24164_ (.A0(_03104_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][6] ),
    .S(net331),
    .X(_01567_));
 sg13g2_mux2_1 _24165_ (.A0(net842),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][7] ),
    .S(net331),
    .X(_01568_));
 sg13g2_mux2_1 _24166_ (.A0(_03711_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][8] ),
    .S(_06062_),
    .X(_01569_));
 sg13g2_mux2_1 _24167_ (.A0(net445),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][9] ),
    .S(_06062_),
    .X(_01570_));
 sg13g2_buf_1 _24168_ (.A(_06029_),
    .X(_06066_));
 sg13g2_nand3_1 _24169_ (.B(_06048_),
    .C(_06066_),
    .A(_05815_),
    .Y(_06067_));
 sg13g2_buf_2 _24170_ (.A(_06067_),
    .X(_06068_));
 sg13g2_buf_1 _24171_ (.A(_06068_),
    .X(_06069_));
 sg13g2_nand2_1 _24172_ (.Y(_06070_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][0] ),
    .B(_06068_));
 sg13g2_o21ai_1 _24173_ (.B1(_06070_),
    .Y(_01571_),
    .A1(net495),
    .A2(_06069_));
 sg13g2_mux2_1 _24174_ (.A0(net568),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][10] ),
    .S(net330),
    .X(_01572_));
 sg13g2_mux2_1 _24175_ (.A0(_03714_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][11] ),
    .S(_06069_),
    .X(_01573_));
 sg13g2_nand2_1 _24176_ (.Y(_06071_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][1] ),
    .B(_06068_));
 sg13g2_o21ai_1 _24177_ (.B1(_06071_),
    .Y(_01574_),
    .A1(net641),
    .A2(net330));
 sg13g2_mux2_1 _24178_ (.A0(net717),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][2] ),
    .S(net330),
    .X(_01575_));
 sg13g2_mux2_1 _24179_ (.A0(_03098_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][3] ),
    .S(net330),
    .X(_01576_));
 sg13g2_mux2_1 _24180_ (.A0(_03100_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][4] ),
    .S(net330),
    .X(_01577_));
 sg13g2_mux2_1 _24181_ (.A0(net844),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][5] ),
    .S(net330),
    .X(_01578_));
 sg13g2_mux2_1 _24182_ (.A0(_03104_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][6] ),
    .S(net330),
    .X(_01579_));
 sg13g2_mux2_1 _24183_ (.A0(net842),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][7] ),
    .S(net330),
    .X(_01580_));
 sg13g2_mux2_1 _24184_ (.A0(_03711_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][8] ),
    .S(_06068_),
    .X(_01581_));
 sg13g2_mux2_1 _24185_ (.A0(net445),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][9] ),
    .S(_06068_),
    .X(_01582_));
 sg13g2_nor3_2 _24186_ (.A(net950),
    .B(net951),
    .C(net949),
    .Y(_06072_));
 sg13g2_nand4_1 _24187_ (.B(_05837_),
    .C(_06072_),
    .A(net944),
    .Y(_06073_),
    .D(net477));
 sg13g2_buf_2 _24188_ (.A(_06073_),
    .X(_06074_));
 sg13g2_buf_1 _24189_ (.A(_06074_),
    .X(_06075_));
 sg13g2_nand2_1 _24190_ (.Y(_06076_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][0] ),
    .B(_06074_));
 sg13g2_o21ai_1 _24191_ (.B1(_06076_),
    .Y(_01583_),
    .A1(net495),
    .A2(_06075_));
 sg13g2_mux2_1 _24192_ (.A0(net568),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][10] ),
    .S(net329),
    .X(_01584_));
 sg13g2_mux2_1 _24193_ (.A0(net567),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][11] ),
    .S(net329),
    .X(_01585_));
 sg13g2_buf_1 _24194_ (.A(_03088_),
    .X(_06077_));
 sg13g2_nand2_1 _24195_ (.Y(_06078_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][1] ),
    .B(_06074_));
 sg13g2_o21ai_1 _24196_ (.B1(_06078_),
    .Y(_01586_),
    .A1(_06077_),
    .A2(_06075_));
 sg13g2_buf_1 _24197_ (.A(net847),
    .X(_06079_));
 sg13g2_mux2_1 _24198_ (.A0(net707),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][2] ),
    .S(net329),
    .X(_01587_));
 sg13g2_buf_1 _24199_ (.A(net846),
    .X(_06080_));
 sg13g2_mux2_1 _24200_ (.A0(net706),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][3] ),
    .S(net329),
    .X(_01588_));
 sg13g2_buf_1 _24201_ (.A(net845),
    .X(_06081_));
 sg13g2_mux2_1 _24202_ (.A0(net705),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][4] ),
    .S(net329),
    .X(_01589_));
 sg13g2_buf_1 _24203_ (.A(net964),
    .X(_06082_));
 sg13g2_mux2_1 _24204_ (.A0(net816),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][5] ),
    .S(net329),
    .X(_01590_));
 sg13g2_buf_1 _24205_ (.A(net963),
    .X(_06083_));
 sg13g2_mux2_1 _24206_ (.A0(net815),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][6] ),
    .S(net329),
    .X(_01591_));
 sg13g2_buf_1 _24207_ (.A(net962),
    .X(_06084_));
 sg13g2_mux2_1 _24208_ (.A0(net814),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][7] ),
    .S(net329),
    .X(_01592_));
 sg13g2_mux2_1 _24209_ (.A0(net446),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][8] ),
    .S(_06074_),
    .X(_01593_));
 sg13g2_mux2_1 _24210_ (.A0(net445),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][9] ),
    .S(_06074_),
    .X(_01594_));
 sg13g2_nand4_1 _24211_ (.B(_05823_),
    .C(_05837_),
    .A(net944),
    .Y(_06085_),
    .D(_06055_));
 sg13g2_buf_2 _24212_ (.A(_06085_),
    .X(_06086_));
 sg13g2_buf_1 _24213_ (.A(_06086_),
    .X(_06087_));
 sg13g2_nand2_1 _24214_ (.Y(_06088_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][0] ),
    .B(_06086_));
 sg13g2_o21ai_1 _24215_ (.B1(_06088_),
    .Y(_01595_),
    .A1(net495),
    .A2(_06087_));
 sg13g2_mux2_1 _24216_ (.A0(net568),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][10] ),
    .S(net271),
    .X(_01596_));
 sg13g2_mux2_1 _24217_ (.A0(net567),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][11] ),
    .S(net271),
    .X(_01597_));
 sg13g2_nand2_1 _24218_ (.Y(_06089_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][1] ),
    .B(_06086_));
 sg13g2_o21ai_1 _24219_ (.B1(_06089_),
    .Y(_01598_),
    .A1(_06077_),
    .A2(_06087_));
 sg13g2_mux2_1 _24220_ (.A0(net707),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][2] ),
    .S(net271),
    .X(_01599_));
 sg13g2_mux2_1 _24221_ (.A0(net706),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][3] ),
    .S(net271),
    .X(_01600_));
 sg13g2_mux2_1 _24222_ (.A0(net705),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][4] ),
    .S(net271),
    .X(_01601_));
 sg13g2_mux2_1 _24223_ (.A0(_06082_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][5] ),
    .S(net271),
    .X(_01602_));
 sg13g2_mux2_1 _24224_ (.A0(net815),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][6] ),
    .S(net271),
    .X(_01603_));
 sg13g2_mux2_1 _24225_ (.A0(net814),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][7] ),
    .S(net271),
    .X(_01604_));
 sg13g2_mux2_1 _24226_ (.A0(net446),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][8] ),
    .S(_06086_),
    .X(_01605_));
 sg13g2_mux2_1 _24227_ (.A0(net445),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][9] ),
    .S(_06086_),
    .X(_01606_));
 sg13g2_buf_1 _24228_ (.A(net566),
    .X(_06090_));
 sg13g2_nand2_1 _24229_ (.Y(_06091_),
    .A(_05916_),
    .B(net478));
 sg13g2_buf_2 _24230_ (.A(_06091_),
    .X(_06092_));
 sg13g2_buf_1 _24231_ (.A(_06092_),
    .X(_06093_));
 sg13g2_nand2_1 _24232_ (.Y(_06094_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][0] ),
    .B(_06092_));
 sg13g2_o21ai_1 _24233_ (.B1(_06094_),
    .Y(_01607_),
    .A1(net476),
    .A2(_06093_));
 sg13g2_buf_1 _24234_ (.A(net639),
    .X(_06095_));
 sg13g2_mux2_1 _24235_ (.A0(net560),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][10] ),
    .S(net328),
    .X(_01608_));
 sg13g2_buf_1 _24236_ (.A(net638),
    .X(_06096_));
 sg13g2_mux2_1 _24237_ (.A0(net559),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][11] ),
    .S(net328),
    .X(_01609_));
 sg13g2_nand2_1 _24238_ (.Y(_06097_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][1] ),
    .B(_06092_));
 sg13g2_o21ai_1 _24239_ (.B1(_06097_),
    .Y(_01610_),
    .A1(net625),
    .A2(_06093_));
 sg13g2_mux2_1 _24240_ (.A0(net707),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][2] ),
    .S(net328),
    .X(_01611_));
 sg13g2_mux2_1 _24241_ (.A0(net706),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][3] ),
    .S(net328),
    .X(_01612_));
 sg13g2_mux2_1 _24242_ (.A0(net705),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][4] ),
    .S(net328),
    .X(_01613_));
 sg13g2_mux2_1 _24243_ (.A0(net816),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][5] ),
    .S(net328),
    .X(_01614_));
 sg13g2_mux2_1 _24244_ (.A0(net815),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][6] ),
    .S(net328),
    .X(_01615_));
 sg13g2_mux2_1 _24245_ (.A0(net814),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][7] ),
    .S(net328),
    .X(_01616_));
 sg13g2_buf_1 _24246_ (.A(net504),
    .X(_06098_));
 sg13g2_mux2_1 _24247_ (.A0(net443),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][8] ),
    .S(_06092_),
    .X(_01617_));
 sg13g2_buf_1 _24248_ (.A(net503),
    .X(_06099_));
 sg13g2_mux2_1 _24249_ (.A0(net442),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][9] ),
    .S(_06092_),
    .X(_01618_));
 sg13g2_nand2_1 _24250_ (.Y(_06100_),
    .A(_05925_),
    .B(net478));
 sg13g2_buf_2 _24251_ (.A(_06100_),
    .X(_06101_));
 sg13g2_buf_1 _24252_ (.A(_06101_),
    .X(_06102_));
 sg13g2_nand2_1 _24253_ (.Y(_06103_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][0] ),
    .B(_06101_));
 sg13g2_o21ai_1 _24254_ (.B1(_06103_),
    .Y(_01619_),
    .A1(_06090_),
    .A2(_06102_));
 sg13g2_mux2_1 _24255_ (.A0(net560),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][10] ),
    .S(net327),
    .X(_01620_));
 sg13g2_mux2_1 _24256_ (.A0(net559),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][11] ),
    .S(net327),
    .X(_01621_));
 sg13g2_nand2_1 _24257_ (.Y(_06104_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][1] ),
    .B(_06101_));
 sg13g2_o21ai_1 _24258_ (.B1(_06104_),
    .Y(_01622_),
    .A1(net625),
    .A2(_06102_));
 sg13g2_mux2_1 _24259_ (.A0(_06079_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][2] ),
    .S(net327),
    .X(_01623_));
 sg13g2_mux2_1 _24260_ (.A0(net706),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][3] ),
    .S(net327),
    .X(_01624_));
 sg13g2_mux2_1 _24261_ (.A0(net705),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][4] ),
    .S(net327),
    .X(_01625_));
 sg13g2_mux2_1 _24262_ (.A0(net816),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][5] ),
    .S(net327),
    .X(_01626_));
 sg13g2_mux2_1 _24263_ (.A0(net815),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][6] ),
    .S(net327),
    .X(_01627_));
 sg13g2_mux2_1 _24264_ (.A0(net814),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][7] ),
    .S(net327),
    .X(_01628_));
 sg13g2_mux2_1 _24265_ (.A0(net443),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][8] ),
    .S(_06101_),
    .X(_01629_));
 sg13g2_mux2_1 _24266_ (.A0(net442),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][9] ),
    .S(_06101_),
    .X(_01630_));
 sg13g2_nand2_1 _24267_ (.Y(_06105_),
    .A(_06027_),
    .B(_06055_));
 sg13g2_buf_2 _24268_ (.A(_06105_),
    .X(_06106_));
 sg13g2_buf_1 _24269_ (.A(_06106_),
    .X(_06107_));
 sg13g2_nand2_1 _24270_ (.Y(_06108_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][0] ),
    .B(_06106_));
 sg13g2_o21ai_1 _24271_ (.B1(_06108_),
    .Y(_01631_),
    .A1(net476),
    .A2(_06107_));
 sg13g2_mux2_1 _24272_ (.A0(_06095_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][10] ),
    .S(net270),
    .X(_01632_));
 sg13g2_mux2_1 _24273_ (.A0(net559),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][11] ),
    .S(net270),
    .X(_01633_));
 sg13g2_nand2_1 _24274_ (.Y(_06109_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][1] ),
    .B(_06106_));
 sg13g2_o21ai_1 _24275_ (.B1(_06109_),
    .Y(_01634_),
    .A1(net625),
    .A2(_06107_));
 sg13g2_mux2_1 _24276_ (.A0(_06079_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][2] ),
    .S(net270),
    .X(_01635_));
 sg13g2_mux2_1 _24277_ (.A0(_06080_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][3] ),
    .S(net270),
    .X(_01636_));
 sg13g2_mux2_1 _24278_ (.A0(_06081_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][4] ),
    .S(net270),
    .X(_01637_));
 sg13g2_mux2_1 _24279_ (.A0(_06082_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][5] ),
    .S(net270),
    .X(_01638_));
 sg13g2_mux2_1 _24280_ (.A0(_06083_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][6] ),
    .S(net270),
    .X(_01639_));
 sg13g2_mux2_1 _24281_ (.A0(net814),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][7] ),
    .S(net270),
    .X(_01640_));
 sg13g2_mux2_1 _24282_ (.A0(net443),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][8] ),
    .S(_06106_),
    .X(_01641_));
 sg13g2_mux2_1 _24283_ (.A0(net442),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][9] ),
    .S(_06106_),
    .X(_01642_));
 sg13g2_nor2_1 _24284_ (.A(_05849_),
    .B(_05900_),
    .Y(_06110_));
 sg13g2_nand2_1 _24285_ (.Y(_06111_),
    .A(_06110_),
    .B(_06031_));
 sg13g2_buf_2 _24286_ (.A(_06111_),
    .X(_06112_));
 sg13g2_buf_1 _24287_ (.A(_06112_),
    .X(_06113_));
 sg13g2_nand2_1 _24288_ (.Y(_06114_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][0] ),
    .B(_06112_));
 sg13g2_o21ai_1 _24289_ (.B1(_06114_),
    .Y(_01643_),
    .A1(net476),
    .A2(_06113_));
 sg13g2_mux2_1 _24290_ (.A0(net560),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][10] ),
    .S(net269),
    .X(_01644_));
 sg13g2_mux2_1 _24291_ (.A0(net559),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][11] ),
    .S(net269),
    .X(_01645_));
 sg13g2_nand2_1 _24292_ (.Y(_06115_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][1] ),
    .B(_06112_));
 sg13g2_o21ai_1 _24293_ (.B1(_06115_),
    .Y(_01646_),
    .A1(net625),
    .A2(_06113_));
 sg13g2_mux2_1 _24294_ (.A0(net707),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][2] ),
    .S(net269),
    .X(_01647_));
 sg13g2_mux2_1 _24295_ (.A0(net706),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][3] ),
    .S(net269),
    .X(_01648_));
 sg13g2_mux2_1 _24296_ (.A0(net705),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][4] ),
    .S(net269),
    .X(_01649_));
 sg13g2_mux2_1 _24297_ (.A0(net816),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][5] ),
    .S(net269),
    .X(_01650_));
 sg13g2_mux2_1 _24298_ (.A0(net815),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][6] ),
    .S(net269),
    .X(_01651_));
 sg13g2_mux2_1 _24299_ (.A0(net814),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][7] ),
    .S(net269),
    .X(_01652_));
 sg13g2_mux2_1 _24300_ (.A0(net443),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][8] ),
    .S(_06112_),
    .X(_01653_));
 sg13g2_mux2_1 _24301_ (.A0(_06099_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][9] ),
    .S(_06112_),
    .X(_01654_));
 sg13g2_nand2_1 _24302_ (.Y(_06116_),
    .A(_06110_),
    .B(_06055_));
 sg13g2_buf_2 _24303_ (.A(_06116_),
    .X(_06117_));
 sg13g2_buf_1 _24304_ (.A(_06117_),
    .X(_06118_));
 sg13g2_nand2_1 _24305_ (.Y(_06119_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][0] ),
    .B(_06117_));
 sg13g2_o21ai_1 _24306_ (.B1(_06119_),
    .Y(_01655_),
    .A1(net476),
    .A2(_06118_));
 sg13g2_mux2_1 _24307_ (.A0(net560),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][10] ),
    .S(net268),
    .X(_01656_));
 sg13g2_mux2_1 _24308_ (.A0(net559),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][11] ),
    .S(net268),
    .X(_01657_));
 sg13g2_nand2_1 _24309_ (.Y(_06120_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][1] ),
    .B(_06117_));
 sg13g2_o21ai_1 _24310_ (.B1(_06120_),
    .Y(_01658_),
    .A1(net625),
    .A2(_06118_));
 sg13g2_mux2_1 _24311_ (.A0(net707),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][2] ),
    .S(net268),
    .X(_01659_));
 sg13g2_mux2_1 _24312_ (.A0(net706),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][3] ),
    .S(net268),
    .X(_01660_));
 sg13g2_mux2_1 _24313_ (.A0(net705),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][4] ),
    .S(net268),
    .X(_01661_));
 sg13g2_mux2_1 _24314_ (.A0(net816),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][5] ),
    .S(net268),
    .X(_01662_));
 sg13g2_mux2_1 _24315_ (.A0(net815),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][6] ),
    .S(net268),
    .X(_01663_));
 sg13g2_mux2_1 _24316_ (.A0(net814),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][7] ),
    .S(net268),
    .X(_01664_));
 sg13g2_mux2_1 _24317_ (.A0(net443),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][8] ),
    .S(_06117_),
    .X(_01665_));
 sg13g2_mux2_1 _24318_ (.A0(net442),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][9] ),
    .S(_06117_),
    .X(_01666_));
 sg13g2_nand3_1 _24319_ (.B(_06110_),
    .C(net477),
    .A(_06009_),
    .Y(_06121_));
 sg13g2_buf_2 _24320_ (.A(_06121_),
    .X(_06122_));
 sg13g2_buf_1 _24321_ (.A(_06122_),
    .X(_06123_));
 sg13g2_nand2_1 _24322_ (.Y(_06124_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][0] ),
    .B(_06122_));
 sg13g2_o21ai_1 _24323_ (.B1(_06124_),
    .Y(_01667_),
    .A1(net476),
    .A2(_06123_));
 sg13g2_mux2_1 _24324_ (.A0(net560),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][10] ),
    .S(net326),
    .X(_01668_));
 sg13g2_mux2_1 _24325_ (.A0(_06096_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][11] ),
    .S(net326),
    .X(_01669_));
 sg13g2_nand2_1 _24326_ (.Y(_06125_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][1] ),
    .B(_06122_));
 sg13g2_o21ai_1 _24327_ (.B1(_06125_),
    .Y(_01670_),
    .A1(net625),
    .A2(_06123_));
 sg13g2_mux2_1 _24328_ (.A0(net707),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][2] ),
    .S(net326),
    .X(_01671_));
 sg13g2_mux2_1 _24329_ (.A0(net706),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][3] ),
    .S(net326),
    .X(_01672_));
 sg13g2_mux2_1 _24330_ (.A0(net705),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][4] ),
    .S(net326),
    .X(_01673_));
 sg13g2_mux2_1 _24331_ (.A0(net816),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][5] ),
    .S(net326),
    .X(_01674_));
 sg13g2_mux2_1 _24332_ (.A0(net815),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][6] ),
    .S(net326),
    .X(_01675_));
 sg13g2_mux2_1 _24333_ (.A0(_06084_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][7] ),
    .S(net326),
    .X(_01676_));
 sg13g2_mux2_1 _24334_ (.A0(net443),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][8] ),
    .S(_06122_),
    .X(_01677_));
 sg13g2_mux2_1 _24335_ (.A0(_06099_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][9] ),
    .S(_06122_),
    .X(_01678_));
 sg13g2_nand3_1 _24336_ (.B(_06110_),
    .C(net477),
    .A(_05815_),
    .Y(_06126_));
 sg13g2_buf_2 _24337_ (.A(_06126_),
    .X(_06127_));
 sg13g2_buf_1 _24338_ (.A(_06127_),
    .X(_06128_));
 sg13g2_nand2_1 _24339_ (.Y(_06129_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][0] ),
    .B(_06127_));
 sg13g2_o21ai_1 _24340_ (.B1(_06129_),
    .Y(_01679_),
    .A1(_06090_),
    .A2(_06128_));
 sg13g2_mux2_1 _24341_ (.A0(net560),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][10] ),
    .S(net325),
    .X(_01680_));
 sg13g2_mux2_1 _24342_ (.A0(_06096_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][11] ),
    .S(net325),
    .X(_01681_));
 sg13g2_nand2_1 _24343_ (.Y(_06130_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][1] ),
    .B(_06127_));
 sg13g2_o21ai_1 _24344_ (.B1(_06130_),
    .Y(_01682_),
    .A1(net625),
    .A2(_06128_));
 sg13g2_mux2_1 _24345_ (.A0(net707),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][2] ),
    .S(net325),
    .X(_01683_));
 sg13g2_mux2_1 _24346_ (.A0(net706),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][3] ),
    .S(net325),
    .X(_01684_));
 sg13g2_mux2_1 _24347_ (.A0(net705),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][4] ),
    .S(net325),
    .X(_01685_));
 sg13g2_mux2_1 _24348_ (.A0(net816),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][5] ),
    .S(net325),
    .X(_01686_));
 sg13g2_mux2_1 _24349_ (.A0(_06083_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][6] ),
    .S(net325),
    .X(_01687_));
 sg13g2_mux2_1 _24350_ (.A0(_06084_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][7] ),
    .S(net325),
    .X(_01688_));
 sg13g2_mux2_1 _24351_ (.A0(net443),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][8] ),
    .S(_06127_),
    .X(_01689_));
 sg13g2_mux2_1 _24352_ (.A0(net442),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][9] ),
    .S(_06127_),
    .X(_01690_));
 sg13g2_nand4_1 _24353_ (.B(net948),
    .C(_06072_),
    .A(net944),
    .Y(_06131_),
    .D(net477));
 sg13g2_buf_2 _24354_ (.A(_06131_),
    .X(_06132_));
 sg13g2_buf_1 _24355_ (.A(_06132_),
    .X(_06133_));
 sg13g2_nand2_1 _24356_ (.Y(_06134_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][0] ),
    .B(_06132_));
 sg13g2_o21ai_1 _24357_ (.B1(_06134_),
    .Y(_01691_),
    .A1(net476),
    .A2(_06133_));
 sg13g2_mux2_1 _24358_ (.A0(net560),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][10] ),
    .S(net324),
    .X(_01692_));
 sg13g2_mux2_1 _24359_ (.A0(net559),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][11] ),
    .S(net324),
    .X(_01693_));
 sg13g2_nand2_1 _24360_ (.Y(_06135_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][1] ),
    .B(_06132_));
 sg13g2_o21ai_1 _24361_ (.B1(_06135_),
    .Y(_01694_),
    .A1(net625),
    .A2(_06133_));
 sg13g2_mux2_1 _24362_ (.A0(net707),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][2] ),
    .S(net324),
    .X(_01695_));
 sg13g2_mux2_1 _24363_ (.A0(_06080_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][3] ),
    .S(net324),
    .X(_01696_));
 sg13g2_mux2_1 _24364_ (.A0(_06081_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][4] ),
    .S(net324),
    .X(_01697_));
 sg13g2_mux2_1 _24365_ (.A0(net816),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][5] ),
    .S(net324),
    .X(_01698_));
 sg13g2_mux2_1 _24366_ (.A0(net815),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][6] ),
    .S(net324),
    .X(_01699_));
 sg13g2_mux2_1 _24367_ (.A0(net814),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][7] ),
    .S(net324),
    .X(_01700_));
 sg13g2_mux2_1 _24368_ (.A0(net443),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][8] ),
    .S(_06132_),
    .X(_01701_));
 sg13g2_mux2_1 _24369_ (.A0(net442),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][9] ),
    .S(_06132_),
    .X(_01702_));
 sg13g2_nand4_1 _24370_ (.B(_05823_),
    .C(net948),
    .A(net944),
    .Y(_06136_),
    .D(_06055_));
 sg13g2_buf_2 _24371_ (.A(_06136_),
    .X(_06137_));
 sg13g2_buf_1 _24372_ (.A(_06137_),
    .X(_06138_));
 sg13g2_nand2_1 _24373_ (.Y(_06139_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][0] ),
    .B(_06137_));
 sg13g2_o21ai_1 _24374_ (.B1(_06139_),
    .Y(_01703_),
    .A1(net476),
    .A2(_06138_));
 sg13g2_mux2_1 _24375_ (.A0(_06095_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][10] ),
    .S(net267),
    .X(_01704_));
 sg13g2_mux2_1 _24376_ (.A0(net559),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][11] ),
    .S(net267),
    .X(_01705_));
 sg13g2_buf_1 _24377_ (.A(net718),
    .X(_06140_));
 sg13g2_nand2_1 _24378_ (.Y(_06141_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][1] ),
    .B(_06137_));
 sg13g2_o21ai_1 _24379_ (.B1(_06141_),
    .Y(_01706_),
    .A1(net624),
    .A2(_06138_));
 sg13g2_buf_1 _24380_ (.A(net847),
    .X(_06142_));
 sg13g2_mux2_1 _24381_ (.A0(net704),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][2] ),
    .S(net267),
    .X(_01707_));
 sg13g2_buf_1 _24382_ (.A(net846),
    .X(_06143_));
 sg13g2_mux2_1 _24383_ (.A0(net703),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][3] ),
    .S(net267),
    .X(_01708_));
 sg13g2_buf_1 _24384_ (.A(net845),
    .X(_06144_));
 sg13g2_mux2_1 _24385_ (.A0(net702),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][4] ),
    .S(net267),
    .X(_01709_));
 sg13g2_buf_1 _24386_ (.A(net964),
    .X(_06145_));
 sg13g2_mux2_1 _24387_ (.A0(net813),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][5] ),
    .S(net267),
    .X(_01710_));
 sg13g2_buf_1 _24388_ (.A(net963),
    .X(_06146_));
 sg13g2_mux2_1 _24389_ (.A0(net812),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][6] ),
    .S(net267),
    .X(_01711_));
 sg13g2_buf_1 _24390_ (.A(net962),
    .X(_06147_));
 sg13g2_mux2_1 _24391_ (.A0(net811),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][7] ),
    .S(net267),
    .X(_01712_));
 sg13g2_mux2_1 _24392_ (.A0(_06098_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][8] ),
    .S(_06137_),
    .X(_01713_));
 sg13g2_mux2_1 _24393_ (.A0(net442),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][9] ),
    .S(_06137_),
    .X(_01714_));
 sg13g2_nand2_1 _24394_ (.Y(_06148_),
    .A(_05961_),
    .B(net478));
 sg13g2_buf_2 _24395_ (.A(_06148_),
    .X(_06149_));
 sg13g2_buf_1 _24396_ (.A(_06149_),
    .X(_06150_));
 sg13g2_nand2_1 _24397_ (.Y(_06151_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][0] ),
    .B(_06149_));
 sg13g2_o21ai_1 _24398_ (.B1(_06151_),
    .Y(_01715_),
    .A1(net476),
    .A2(_06150_));
 sg13g2_mux2_1 _24399_ (.A0(net560),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][10] ),
    .S(net323),
    .X(_01716_));
 sg13g2_mux2_1 _24400_ (.A0(net559),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][11] ),
    .S(net323),
    .X(_01717_));
 sg13g2_nand2_1 _24401_ (.Y(_06152_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][1] ),
    .B(_06149_));
 sg13g2_o21ai_1 _24402_ (.B1(_06152_),
    .Y(_01718_),
    .A1(net624),
    .A2(_06150_));
 sg13g2_mux2_1 _24403_ (.A0(net704),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][2] ),
    .S(net323),
    .X(_01719_));
 sg13g2_mux2_1 _24404_ (.A0(net703),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][3] ),
    .S(net323),
    .X(_01720_));
 sg13g2_mux2_1 _24405_ (.A0(net702),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][4] ),
    .S(net323),
    .X(_01721_));
 sg13g2_mux2_1 _24406_ (.A0(net813),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][5] ),
    .S(net323),
    .X(_01722_));
 sg13g2_mux2_1 _24407_ (.A0(net812),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][6] ),
    .S(net323),
    .X(_01723_));
 sg13g2_mux2_1 _24408_ (.A0(net811),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][7] ),
    .S(net323),
    .X(_01724_));
 sg13g2_mux2_1 _24409_ (.A0(_06098_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][8] ),
    .S(_06149_),
    .X(_01725_));
 sg13g2_mux2_1 _24410_ (.A0(net442),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][9] ),
    .S(_06149_),
    .X(_01726_));
 sg13g2_buf_1 _24411_ (.A(net566),
    .X(_06153_));
 sg13g2_nand2_1 _24412_ (.Y(_06154_),
    .A(_05967_),
    .B(net478));
 sg13g2_buf_2 _24413_ (.A(_06154_),
    .X(_06155_));
 sg13g2_buf_1 _24414_ (.A(_06155_),
    .X(_06156_));
 sg13g2_nand2_1 _24415_ (.Y(_06157_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][0] ),
    .B(_06155_));
 sg13g2_o21ai_1 _24416_ (.B1(_06157_),
    .Y(_01727_),
    .A1(net475),
    .A2(_06156_));
 sg13g2_buf_1 _24417_ (.A(net639),
    .X(_06158_));
 sg13g2_mux2_1 _24418_ (.A0(net558),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][10] ),
    .S(net322),
    .X(_01728_));
 sg13g2_buf_1 _24419_ (.A(net638),
    .X(_06159_));
 sg13g2_mux2_1 _24420_ (.A0(net557),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][11] ),
    .S(net322),
    .X(_01729_));
 sg13g2_nand2_1 _24421_ (.Y(_06160_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][1] ),
    .B(_06155_));
 sg13g2_o21ai_1 _24422_ (.B1(_06160_),
    .Y(_01730_),
    .A1(net624),
    .A2(_06156_));
 sg13g2_mux2_1 _24423_ (.A0(net704),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][2] ),
    .S(net322),
    .X(_01731_));
 sg13g2_mux2_1 _24424_ (.A0(net703),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][3] ),
    .S(net322),
    .X(_01732_));
 sg13g2_mux2_1 _24425_ (.A0(net702),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][4] ),
    .S(net322),
    .X(_01733_));
 sg13g2_mux2_1 _24426_ (.A0(net813),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][5] ),
    .S(net322),
    .X(_01734_));
 sg13g2_mux2_1 _24427_ (.A0(net812),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][6] ),
    .S(net322),
    .X(_01735_));
 sg13g2_mux2_1 _24428_ (.A0(net811),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][7] ),
    .S(net322),
    .X(_01736_));
 sg13g2_buf_1 _24429_ (.A(_03642_),
    .X(_06161_));
 sg13g2_mux2_1 _24430_ (.A0(net441),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][8] ),
    .S(_06155_),
    .X(_01737_));
 sg13g2_buf_1 _24431_ (.A(net503),
    .X(_06162_));
 sg13g2_mux2_1 _24432_ (.A0(_06162_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][9] ),
    .S(_06155_),
    .X(_01738_));
 sg13g2_nor2_1 _24433_ (.A(_05849_),
    .B(_05952_),
    .Y(_06163_));
 sg13g2_nand2_1 _24434_ (.Y(_06164_),
    .A(_06163_),
    .B(_06031_));
 sg13g2_buf_2 _24435_ (.A(_06164_),
    .X(_06165_));
 sg13g2_buf_1 _24436_ (.A(_06165_),
    .X(_06166_));
 sg13g2_nand2_1 _24437_ (.Y(_06167_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][0] ),
    .B(_06165_));
 sg13g2_o21ai_1 _24438_ (.B1(_06167_),
    .Y(_01739_),
    .A1(net475),
    .A2(net266));
 sg13g2_mux2_1 _24439_ (.A0(net558),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][10] ),
    .S(net266),
    .X(_01740_));
 sg13g2_mux2_1 _24440_ (.A0(net557),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][11] ),
    .S(_06166_),
    .X(_01741_));
 sg13g2_nand2_1 _24441_ (.Y(_06168_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][1] ),
    .B(_06165_));
 sg13g2_o21ai_1 _24442_ (.B1(_06168_),
    .Y(_01742_),
    .A1(net624),
    .A2(_06166_));
 sg13g2_mux2_1 _24443_ (.A0(net704),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][2] ),
    .S(net266),
    .X(_01743_));
 sg13g2_mux2_1 _24444_ (.A0(net703),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][3] ),
    .S(net266),
    .X(_01744_));
 sg13g2_mux2_1 _24445_ (.A0(net702),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][4] ),
    .S(net266),
    .X(_01745_));
 sg13g2_mux2_1 _24446_ (.A0(net813),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][5] ),
    .S(net266),
    .X(_01746_));
 sg13g2_mux2_1 _24447_ (.A0(net812),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][6] ),
    .S(net266),
    .X(_01747_));
 sg13g2_mux2_1 _24448_ (.A0(net811),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][7] ),
    .S(net266),
    .X(_01748_));
 sg13g2_mux2_1 _24449_ (.A0(net441),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][8] ),
    .S(_06165_),
    .X(_01749_));
 sg13g2_mux2_1 _24450_ (.A0(net440),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][9] ),
    .S(_06165_),
    .X(_01750_));
 sg13g2_nand2_1 _24451_ (.Y(_06169_),
    .A(_06163_),
    .B(_06055_));
 sg13g2_buf_2 _24452_ (.A(_06169_),
    .X(_06170_));
 sg13g2_buf_1 _24453_ (.A(_06170_),
    .X(_06171_));
 sg13g2_nand2_1 _24454_ (.Y(_06172_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][0] ),
    .B(_06170_));
 sg13g2_o21ai_1 _24455_ (.B1(_06172_),
    .Y(_01751_),
    .A1(net475),
    .A2(net265));
 sg13g2_mux2_1 _24456_ (.A0(net558),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][10] ),
    .S(net265),
    .X(_01752_));
 sg13g2_mux2_1 _24457_ (.A0(net557),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][11] ),
    .S(_06171_),
    .X(_01753_));
 sg13g2_nand2_1 _24458_ (.Y(_06173_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][1] ),
    .B(_06170_));
 sg13g2_o21ai_1 _24459_ (.B1(_06173_),
    .Y(_01754_),
    .A1(net624),
    .A2(_06171_));
 sg13g2_mux2_1 _24460_ (.A0(net704),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][2] ),
    .S(net265),
    .X(_01755_));
 sg13g2_mux2_1 _24461_ (.A0(net703),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][3] ),
    .S(net265),
    .X(_01756_));
 sg13g2_mux2_1 _24462_ (.A0(net702),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][4] ),
    .S(net265),
    .X(_01757_));
 sg13g2_mux2_1 _24463_ (.A0(net813),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][5] ),
    .S(net265),
    .X(_01758_));
 sg13g2_mux2_1 _24464_ (.A0(net812),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][6] ),
    .S(net265),
    .X(_01759_));
 sg13g2_mux2_1 _24465_ (.A0(net811),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][7] ),
    .S(net265),
    .X(_01760_));
 sg13g2_mux2_1 _24466_ (.A0(net441),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][8] ),
    .S(_06170_),
    .X(_01761_));
 sg13g2_mux2_1 _24467_ (.A0(net440),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][9] ),
    .S(_06170_),
    .X(_01762_));
 sg13g2_nand3_1 _24468_ (.B(_06027_),
    .C(net477),
    .A(_06009_),
    .Y(_06174_));
 sg13g2_buf_2 _24469_ (.A(_06174_),
    .X(_06175_));
 sg13g2_buf_1 _24470_ (.A(_06175_),
    .X(_06176_));
 sg13g2_nand2_1 _24471_ (.Y(_06177_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][0] ),
    .B(_06175_));
 sg13g2_o21ai_1 _24472_ (.B1(_06177_),
    .Y(_01763_),
    .A1(net475),
    .A2(net321));
 sg13g2_mux2_1 _24473_ (.A0(net558),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][10] ),
    .S(_06176_),
    .X(_01764_));
 sg13g2_mux2_1 _24474_ (.A0(net557),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][11] ),
    .S(_06176_),
    .X(_01765_));
 sg13g2_nand2_1 _24475_ (.Y(_06178_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][1] ),
    .B(_06175_));
 sg13g2_o21ai_1 _24476_ (.B1(_06178_),
    .Y(_01766_),
    .A1(_06140_),
    .A2(net321));
 sg13g2_mux2_1 _24477_ (.A0(net704),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][2] ),
    .S(net321),
    .X(_01767_));
 sg13g2_mux2_1 _24478_ (.A0(net703),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][3] ),
    .S(net321),
    .X(_01768_));
 sg13g2_mux2_1 _24479_ (.A0(net702),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][4] ),
    .S(net321),
    .X(_01769_));
 sg13g2_mux2_1 _24480_ (.A0(net813),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][5] ),
    .S(net321),
    .X(_01770_));
 sg13g2_mux2_1 _24481_ (.A0(_06146_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][6] ),
    .S(net321),
    .X(_01771_));
 sg13g2_mux2_1 _24482_ (.A0(net811),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][7] ),
    .S(net321),
    .X(_01772_));
 sg13g2_mux2_1 _24483_ (.A0(_06161_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][8] ),
    .S(_06175_),
    .X(_01773_));
 sg13g2_mux2_1 _24484_ (.A0(net440),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][9] ),
    .S(_06175_),
    .X(_01774_));
 sg13g2_nand3_1 _24485_ (.B(_06163_),
    .C(net477),
    .A(_06009_),
    .Y(_06179_));
 sg13g2_buf_2 _24486_ (.A(_06179_),
    .X(_06180_));
 sg13g2_buf_1 _24487_ (.A(_06180_),
    .X(_06181_));
 sg13g2_nand2_1 _24488_ (.Y(_06182_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][0] ),
    .B(_06180_));
 sg13g2_o21ai_1 _24489_ (.B1(_06182_),
    .Y(_01775_),
    .A1(net475),
    .A2(net320));
 sg13g2_mux2_1 _24490_ (.A0(net558),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][10] ),
    .S(net320),
    .X(_01776_));
 sg13g2_mux2_1 _24491_ (.A0(net557),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][11] ),
    .S(_06181_),
    .X(_01777_));
 sg13g2_nand2_1 _24492_ (.Y(_06183_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][1] ),
    .B(_06180_));
 sg13g2_o21ai_1 _24493_ (.B1(_06183_),
    .Y(_01778_),
    .A1(net624),
    .A2(net320));
 sg13g2_mux2_1 _24494_ (.A0(net704),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][2] ),
    .S(_06181_),
    .X(_01779_));
 sg13g2_mux2_1 _24495_ (.A0(net703),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][3] ),
    .S(net320),
    .X(_01780_));
 sg13g2_mux2_1 _24496_ (.A0(net702),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][4] ),
    .S(net320),
    .X(_01781_));
 sg13g2_mux2_1 _24497_ (.A0(net813),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][5] ),
    .S(net320),
    .X(_01782_));
 sg13g2_mux2_1 _24498_ (.A0(net812),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][6] ),
    .S(net320),
    .X(_01783_));
 sg13g2_mux2_1 _24499_ (.A0(net811),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][7] ),
    .S(net320),
    .X(_01784_));
 sg13g2_mux2_1 _24500_ (.A0(net441),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][8] ),
    .S(_06180_),
    .X(_01785_));
 sg13g2_mux2_1 _24501_ (.A0(net440),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][9] ),
    .S(_06180_),
    .X(_01786_));
 sg13g2_nand3_1 _24502_ (.B(_06163_),
    .C(net477),
    .A(_05815_),
    .Y(_06184_));
 sg13g2_buf_2 _24503_ (.A(_06184_),
    .X(_06185_));
 sg13g2_buf_1 _24504_ (.A(_06185_),
    .X(_06186_));
 sg13g2_nand2_1 _24505_ (.Y(_06187_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][0] ),
    .B(_06185_));
 sg13g2_o21ai_1 _24506_ (.B1(_06187_),
    .Y(_01787_),
    .A1(net475),
    .A2(net319));
 sg13g2_mux2_1 _24507_ (.A0(net558),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][10] ),
    .S(net319),
    .X(_01788_));
 sg13g2_mux2_1 _24508_ (.A0(net557),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][11] ),
    .S(_06186_),
    .X(_01789_));
 sg13g2_nand2_1 _24509_ (.Y(_06188_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][1] ),
    .B(_06185_));
 sg13g2_o21ai_1 _24510_ (.B1(_06188_),
    .Y(_01790_),
    .A1(net624),
    .A2(net319));
 sg13g2_mux2_1 _24511_ (.A0(net704),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][2] ),
    .S(_06186_),
    .X(_01791_));
 sg13g2_mux2_1 _24512_ (.A0(net703),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][3] ),
    .S(net319),
    .X(_01792_));
 sg13g2_mux2_1 _24513_ (.A0(net702),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][4] ),
    .S(net319),
    .X(_01793_));
 sg13g2_mux2_1 _24514_ (.A0(net813),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][5] ),
    .S(net319),
    .X(_01794_));
 sg13g2_mux2_1 _24515_ (.A0(net812),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][6] ),
    .S(net319),
    .X(_01795_));
 sg13g2_mux2_1 _24516_ (.A0(net811),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][7] ),
    .S(net319),
    .X(_01796_));
 sg13g2_mux2_1 _24517_ (.A0(net441),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][8] ),
    .S(_06185_),
    .X(_01797_));
 sg13g2_mux2_1 _24518_ (.A0(net440),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][9] ),
    .S(_06185_),
    .X(_01798_));
 sg13g2_nand3_1 _24519_ (.B(_06027_),
    .C(net477),
    .A(_05815_),
    .Y(_06189_));
 sg13g2_buf_2 _24520_ (.A(_06189_),
    .X(_06190_));
 sg13g2_buf_1 _24521_ (.A(_06190_),
    .X(_06191_));
 sg13g2_nand2_1 _24522_ (.Y(_06192_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][0] ),
    .B(_06190_));
 sg13g2_o21ai_1 _24523_ (.B1(_06192_),
    .Y(_01799_),
    .A1(net475),
    .A2(net318));
 sg13g2_mux2_1 _24524_ (.A0(net558),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][10] ),
    .S(net318),
    .X(_01800_));
 sg13g2_mux2_1 _24525_ (.A0(net557),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][11] ),
    .S(_06191_),
    .X(_01801_));
 sg13g2_nand2_1 _24526_ (.Y(_06193_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][1] ),
    .B(_06190_));
 sg13g2_o21ai_1 _24527_ (.B1(_06193_),
    .Y(_01802_),
    .A1(_06140_),
    .A2(_06191_));
 sg13g2_mux2_1 _24528_ (.A0(_06142_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][2] ),
    .S(net318),
    .X(_01803_));
 sg13g2_mux2_1 _24529_ (.A0(_06143_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][3] ),
    .S(net318),
    .X(_01804_));
 sg13g2_mux2_1 _24530_ (.A0(_06144_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][4] ),
    .S(net318),
    .X(_01805_));
 sg13g2_mux2_1 _24531_ (.A0(_06145_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][5] ),
    .S(net318),
    .X(_01806_));
 sg13g2_mux2_1 _24532_ (.A0(_06146_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][6] ),
    .S(net318),
    .X(_01807_));
 sg13g2_mux2_1 _24533_ (.A0(_06147_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][7] ),
    .S(net318),
    .X(_01808_));
 sg13g2_mux2_1 _24534_ (.A0(net441),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][8] ),
    .S(_06190_),
    .X(_01809_));
 sg13g2_mux2_1 _24535_ (.A0(_06162_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][9] ),
    .S(_06190_),
    .X(_01810_));
 sg13g2_nand2b_1 _24536_ (.Y(_06194_),
    .B(_06031_),
    .A_N(_05999_));
 sg13g2_buf_2 _24537_ (.A(_06194_),
    .X(_06195_));
 sg13g2_buf_1 _24538_ (.A(_06195_),
    .X(_06196_));
 sg13g2_nand2_1 _24539_ (.Y(_06197_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][0] ),
    .B(_06195_));
 sg13g2_o21ai_1 _24540_ (.B1(_06197_),
    .Y(_01811_),
    .A1(net475),
    .A2(_06196_));
 sg13g2_mux2_1 _24541_ (.A0(net558),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][10] ),
    .S(net264),
    .X(_01812_));
 sg13g2_mux2_1 _24542_ (.A0(_06159_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][11] ),
    .S(_06196_),
    .X(_01813_));
 sg13g2_nand2_1 _24543_ (.Y(_06198_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][1] ),
    .B(_06195_));
 sg13g2_o21ai_1 _24544_ (.B1(_06198_),
    .Y(_01814_),
    .A1(net624),
    .A2(net264));
 sg13g2_mux2_1 _24545_ (.A0(_06142_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][2] ),
    .S(net264),
    .X(_01815_));
 sg13g2_mux2_1 _24546_ (.A0(_06143_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][3] ),
    .S(net264),
    .X(_01816_));
 sg13g2_mux2_1 _24547_ (.A0(_06144_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][4] ),
    .S(net264),
    .X(_01817_));
 sg13g2_mux2_1 _24548_ (.A0(_06145_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][5] ),
    .S(net264),
    .X(_01818_));
 sg13g2_mux2_1 _24549_ (.A0(net812),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][6] ),
    .S(net264),
    .X(_01819_));
 sg13g2_mux2_1 _24550_ (.A0(_06147_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][7] ),
    .S(net264),
    .X(_01820_));
 sg13g2_mux2_1 _24551_ (.A0(net441),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][8] ),
    .S(_06195_),
    .X(_01821_));
 sg13g2_mux2_1 _24552_ (.A0(net440),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][9] ),
    .S(_06195_),
    .X(_01822_));
 sg13g2_nand2_1 _24553_ (.Y(_06199_),
    .A(_06004_),
    .B(net478));
 sg13g2_buf_2 _24554_ (.A(_06199_),
    .X(_06200_));
 sg13g2_buf_1 _24555_ (.A(_06200_),
    .X(_06201_));
 sg13g2_nand2_1 _24556_ (.Y(_06202_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][0] ),
    .B(_06200_));
 sg13g2_o21ai_1 _24557_ (.B1(_06202_),
    .Y(_01823_),
    .A1(_06153_),
    .A2(_06201_));
 sg13g2_mux2_1 _24558_ (.A0(_06158_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][10] ),
    .S(net317),
    .X(_01824_));
 sg13g2_mux2_1 _24559_ (.A0(_06159_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][11] ),
    .S(_06201_),
    .X(_01825_));
 sg13g2_nand2_1 _24560_ (.Y(_06203_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][1] ),
    .B(_06200_));
 sg13g2_o21ai_1 _24561_ (.B1(_06203_),
    .Y(_01826_),
    .A1(net718),
    .A2(net317));
 sg13g2_mux2_1 _24562_ (.A0(net714),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][2] ),
    .S(net317),
    .X(_01827_));
 sg13g2_mux2_1 _24563_ (.A0(net713),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][3] ),
    .S(net317),
    .X(_01828_));
 sg13g2_mux2_1 _24564_ (.A0(net712),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][4] ),
    .S(net317),
    .X(_01829_));
 sg13g2_mux2_1 _24565_ (.A0(net841),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][5] ),
    .S(net317),
    .X(_01830_));
 sg13g2_mux2_1 _24566_ (.A0(net840),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][6] ),
    .S(net317),
    .X(_01831_));
 sg13g2_mux2_1 _24567_ (.A0(net839),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][7] ),
    .S(net317),
    .X(_01832_));
 sg13g2_mux2_1 _24568_ (.A0(net441),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][8] ),
    .S(_06200_),
    .X(_01833_));
 sg13g2_mux2_1 _24569_ (.A0(net440),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][9] ),
    .S(_06200_),
    .X(_01834_));
 sg13g2_nand2_1 _24570_ (.Y(_06204_),
    .A(_06011_),
    .B(_06037_));
 sg13g2_buf_2 _24571_ (.A(_06204_),
    .X(_06205_));
 sg13g2_buf_1 _24572_ (.A(_06205_),
    .X(_06206_));
 sg13g2_nand2_1 _24573_ (.Y(_06207_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][0] ),
    .B(_06205_));
 sg13g2_o21ai_1 _24574_ (.B1(_06207_),
    .Y(_01835_),
    .A1(_06153_),
    .A2(_06206_));
 sg13g2_mux2_1 _24575_ (.A0(_06158_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][10] ),
    .S(net316),
    .X(_01836_));
 sg13g2_mux2_1 _24576_ (.A0(net557),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][11] ),
    .S(_06206_),
    .X(_01837_));
 sg13g2_nand2_1 _24577_ (.Y(_06208_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][1] ),
    .B(_06205_));
 sg13g2_o21ai_1 _24578_ (.B1(_06208_),
    .Y(_01838_),
    .A1(net718),
    .A2(net316));
 sg13g2_mux2_1 _24579_ (.A0(net714),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][2] ),
    .S(net316),
    .X(_01839_));
 sg13g2_mux2_1 _24580_ (.A0(net713),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][3] ),
    .S(net316),
    .X(_01840_));
 sg13g2_mux2_1 _24581_ (.A0(net712),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][4] ),
    .S(net316),
    .X(_01841_));
 sg13g2_mux2_1 _24582_ (.A0(net841),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][5] ),
    .S(net316),
    .X(_01842_));
 sg13g2_mux2_1 _24583_ (.A0(net840),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][6] ),
    .S(net316),
    .X(_01843_));
 sg13g2_mux2_1 _24584_ (.A0(net839),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][7] ),
    .S(net316),
    .X(_01844_));
 sg13g2_mux2_1 _24585_ (.A0(_06161_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][8] ),
    .S(_06205_),
    .X(_01845_));
 sg13g2_mux2_1 _24586_ (.A0(net440),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][9] ),
    .S(_06205_),
    .X(_01846_));
 sg13g2_nand2_1 _24587_ (.Y(_06209_),
    .A(_06016_),
    .B(_06037_));
 sg13g2_buf_2 _24588_ (.A(_06209_),
    .X(_06210_));
 sg13g2_buf_1 _24589_ (.A(_06210_),
    .X(_06211_));
 sg13g2_nand2_1 _24590_ (.Y(_06212_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][0] ),
    .B(_06210_));
 sg13g2_o21ai_1 _24591_ (.B1(_06212_),
    .Y(_01847_),
    .A1(net566),
    .A2(net315));
 sg13g2_mux2_1 _24592_ (.A0(net577),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][10] ),
    .S(net315),
    .X(_01848_));
 sg13g2_mux2_1 _24593_ (.A0(net576),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][11] ),
    .S(_06211_),
    .X(_01849_));
 sg13g2_nand2_1 _24594_ (.Y(_06213_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][1] ),
    .B(_06210_));
 sg13g2_o21ai_1 _24595_ (.B1(_06213_),
    .Y(_01850_),
    .A1(net718),
    .A2(_06211_));
 sg13g2_mux2_1 _24596_ (.A0(net714),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][2] ),
    .S(net315),
    .X(_01851_));
 sg13g2_mux2_1 _24597_ (.A0(net713),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][3] ),
    .S(net315),
    .X(_01852_));
 sg13g2_mux2_1 _24598_ (.A0(net712),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][4] ),
    .S(net315),
    .X(_01853_));
 sg13g2_mux2_1 _24599_ (.A0(net841),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][5] ),
    .S(net315),
    .X(_01854_));
 sg13g2_mux2_1 _24600_ (.A0(net840),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][6] ),
    .S(net315),
    .X(_01855_));
 sg13g2_mux2_1 _24601_ (.A0(net839),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][7] ),
    .S(net315),
    .X(_01856_));
 sg13g2_mux2_1 _24602_ (.A0(_03643_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][8] ),
    .S(_06210_),
    .X(_01857_));
 sg13g2_mux2_1 _24603_ (.A0(_03645_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][9] ),
    .S(_06210_),
    .X(_01858_));
 sg13g2_nand3_1 _24604_ (.B(_06072_),
    .C(_06066_),
    .A(_05878_),
    .Y(_06214_));
 sg13g2_buf_2 _24605_ (.A(_06214_),
    .X(_06215_));
 sg13g2_buf_1 _24606_ (.A(_06215_),
    .X(_06216_));
 sg13g2_nand2_1 _24607_ (.Y(_06217_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][0] ),
    .B(_06215_));
 sg13g2_o21ai_1 _24608_ (.B1(_06217_),
    .Y(_01859_),
    .A1(net566),
    .A2(net314));
 sg13g2_mux2_1 _24609_ (.A0(net577),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][10] ),
    .S(_06216_),
    .X(_01860_));
 sg13g2_mux2_1 _24610_ (.A0(net576),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][11] ),
    .S(net314),
    .X(_01861_));
 sg13g2_nand2_1 _24611_ (.Y(_06218_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][1] ),
    .B(_06215_));
 sg13g2_o21ai_1 _24612_ (.B1(_06218_),
    .Y(_01862_),
    .A1(net718),
    .A2(_06216_));
 sg13g2_mux2_1 _24613_ (.A0(net714),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][2] ),
    .S(net314),
    .X(_01863_));
 sg13g2_mux2_1 _24614_ (.A0(net713),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][3] ),
    .S(net314),
    .X(_01864_));
 sg13g2_mux2_1 _24615_ (.A0(net712),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][4] ),
    .S(net314),
    .X(_01865_));
 sg13g2_mux2_1 _24616_ (.A0(net841),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][5] ),
    .S(net314),
    .X(_01866_));
 sg13g2_mux2_1 _24617_ (.A0(net840),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][6] ),
    .S(net314),
    .X(_01867_));
 sg13g2_mux2_1 _24618_ (.A0(_03117_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][7] ),
    .S(net314),
    .X(_01868_));
 sg13g2_mux2_1 _24619_ (.A0(net450),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][8] ),
    .S(_06215_),
    .X(_01869_));
 sg13g2_mux2_1 _24620_ (.A0(net449),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][9] ),
    .S(_06215_),
    .X(_01870_));
 sg13g2_nand3_1 _24621_ (.B(_05878_),
    .C(_06055_),
    .A(_05823_),
    .Y(_06219_));
 sg13g2_buf_2 _24622_ (.A(_06219_),
    .X(_06220_));
 sg13g2_buf_1 _24623_ (.A(_06220_),
    .X(_06221_));
 sg13g2_nand2_1 _24624_ (.Y(_06222_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][0] ),
    .B(_06220_));
 sg13g2_o21ai_1 _24625_ (.B1(_06222_),
    .Y(_01871_),
    .A1(_03717_),
    .A2(net263));
 sg13g2_mux2_1 _24626_ (.A0(net577),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][10] ),
    .S(_06221_),
    .X(_01872_));
 sg13g2_mux2_1 _24627_ (.A0(net576),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][11] ),
    .S(_06221_),
    .X(_01873_));
 sg13g2_nand2_1 _24628_ (.Y(_06223_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][1] ),
    .B(_06220_));
 sg13g2_o21ai_1 _24629_ (.B1(_06223_),
    .Y(_01874_),
    .A1(net718),
    .A2(net263));
 sg13g2_mux2_1 _24630_ (.A0(net714),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][2] ),
    .S(net263),
    .X(_01875_));
 sg13g2_mux2_1 _24631_ (.A0(net713),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][3] ),
    .S(net263),
    .X(_01876_));
 sg13g2_mux2_1 _24632_ (.A0(net712),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][4] ),
    .S(net263),
    .X(_01877_));
 sg13g2_mux2_1 _24633_ (.A0(net841),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][5] ),
    .S(net263),
    .X(_01878_));
 sg13g2_mux2_1 _24634_ (.A0(net840),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][6] ),
    .S(net263),
    .X(_01879_));
 sg13g2_mux2_1 _24635_ (.A0(_03117_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][7] ),
    .S(net263),
    .X(_01880_));
 sg13g2_mux2_1 _24636_ (.A0(_03643_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][8] ),
    .S(_06220_),
    .X(_01881_));
 sg13g2_mux2_1 _24637_ (.A0(_03645_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][9] ),
    .S(_06220_),
    .X(_01882_));
 sg13g2_mux2_1 _24638_ (.A0(\cpu.genblk1.mmu.r_writeable_d[0] ),
    .A1(_03663_),
    .S(_05858_),
    .X(_01883_));
 sg13g2_buf_1 _24639_ (.A(net410),
    .X(_06224_));
 sg13g2_mux2_1 _24640_ (.A0(\cpu.genblk1.mmu.r_writeable_d[10] ),
    .A1(net313),
    .S(_05870_),
    .X(_01884_));
 sg13g2_mux2_1 _24641_ (.A0(\cpu.genblk1.mmu.r_writeable_d[11] ),
    .A1(net313),
    .S(_05875_),
    .X(_01885_));
 sg13g2_mux2_1 _24642_ (.A0(\cpu.genblk1.mmu.r_writeable_d[12] ),
    .A1(net313),
    .S(_05882_),
    .X(_01886_));
 sg13g2_mux2_1 _24643_ (.A0(\cpu.genblk1.mmu.r_writeable_d[13] ),
    .A1(net313),
    .S(_05889_),
    .X(_01887_));
 sg13g2_mux2_1 _24644_ (.A0(\cpu.genblk1.mmu.r_writeable_d[14] ),
    .A1(_06224_),
    .S(_05893_),
    .X(_01888_));
 sg13g2_mux2_1 _24645_ (.A0(\cpu.genblk1.mmu.r_writeable_d[15] ),
    .A1(_06224_),
    .S(_05897_),
    .X(_01889_));
 sg13g2_mux2_1 _24646_ (.A0(\cpu.genblk1.mmu.r_writeable_d[16] ),
    .A1(net313),
    .S(_05905_),
    .X(_01890_));
 sg13g2_mux2_1 _24647_ (.A0(\cpu.genblk1.mmu.r_writeable_d[17] ),
    .A1(net313),
    .S(_05910_),
    .X(_01891_));
 sg13g2_mux2_1 _24648_ (.A0(\cpu.genblk1.mmu.r_writeable_d[18] ),
    .A1(net313),
    .S(_05918_),
    .X(_01892_));
 sg13g2_mux2_1 _24649_ (.A0(\cpu.genblk1.mmu.r_writeable_d[19] ),
    .A1(net313),
    .S(_05927_),
    .X(_01893_));
 sg13g2_buf_1 _24650_ (.A(net410),
    .X(_06225_));
 sg13g2_mux2_1 _24651_ (.A0(\cpu.genblk1.mmu.r_writeable_d[1] ),
    .A1(_06225_),
    .S(_05933_),
    .X(_01894_));
 sg13g2_mux2_1 _24652_ (.A0(\cpu.genblk1.mmu.r_writeable_d[20] ),
    .A1(net312),
    .S(_05938_),
    .X(_01895_));
 sg13g2_mux2_1 _24653_ (.A0(\cpu.genblk1.mmu.r_writeable_d[21] ),
    .A1(net312),
    .S(_05942_),
    .X(_01896_));
 sg13g2_mux2_1 _24654_ (.A0(\cpu.genblk1.mmu.r_writeable_d[22] ),
    .A1(_06225_),
    .S(_05945_),
    .X(_01897_));
 sg13g2_mux2_1 _24655_ (.A0(\cpu.genblk1.mmu.r_writeable_d[23] ),
    .A1(net312),
    .S(_05948_),
    .X(_01898_));
 sg13g2_mux2_1 _24656_ (.A0(\cpu.genblk1.mmu.r_writeable_d[24] ),
    .A1(net312),
    .S(_05954_),
    .X(_01899_));
 sg13g2_mux2_1 _24657_ (.A0(\cpu.genblk1.mmu.r_writeable_d[25] ),
    .A1(net312),
    .S(_05957_),
    .X(_01900_));
 sg13g2_mux2_1 _24658_ (.A0(\cpu.genblk1.mmu.r_writeable_d[26] ),
    .A1(net312),
    .S(_05963_),
    .X(_01901_));
 sg13g2_mux2_1 _24659_ (.A0(\cpu.genblk1.mmu.r_writeable_d[27] ),
    .A1(net312),
    .S(_05969_),
    .X(_01902_));
 sg13g2_mux2_1 _24660_ (.A0(\cpu.genblk1.mmu.r_writeable_d[28] ),
    .A1(net312),
    .S(_05978_),
    .X(_01903_));
 sg13g2_buf_1 _24661_ (.A(_03653_),
    .X(_06226_));
 sg13g2_mux2_1 _24662_ (.A0(\cpu.genblk1.mmu.r_writeable_d[29] ),
    .A1(net311),
    .S(_05984_),
    .X(_01904_));
 sg13g2_mux2_1 _24663_ (.A0(\cpu.genblk1.mmu.r_writeable_d[2] ),
    .A1(net311),
    .S(_05987_),
    .X(_01905_));
 sg13g2_mux2_1 _24664_ (.A0(\cpu.genblk1.mmu.r_writeable_d[30] ),
    .A1(net311),
    .S(_05991_),
    .X(_01906_));
 sg13g2_mux2_1 _24665_ (.A0(\cpu.genblk1.mmu.r_writeable_d[31] ),
    .A1(net311),
    .S(_05994_),
    .X(_01907_));
 sg13g2_mux2_1 _24666_ (.A0(\cpu.genblk1.mmu.r_writeable_d[3] ),
    .A1(net311),
    .S(_05997_),
    .X(_01908_));
 sg13g2_mux2_1 _24667_ (.A0(\cpu.genblk1.mmu.r_writeable_d[4] ),
    .A1(net311),
    .S(_06001_),
    .X(_01909_));
 sg13g2_mux2_1 _24668_ (.A0(\cpu.genblk1.mmu.r_writeable_d[5] ),
    .A1(_06226_),
    .S(_06006_),
    .X(_01910_));
 sg13g2_mux2_1 _24669_ (.A0(\cpu.genblk1.mmu.r_writeable_d[6] ),
    .A1(net311),
    .S(_06013_),
    .X(_01911_));
 sg13g2_mux2_1 _24670_ (.A0(\cpu.genblk1.mmu.r_writeable_d[7] ),
    .A1(_06226_),
    .S(_06018_),
    .X(_01912_));
 sg13g2_mux2_1 _24671_ (.A0(\cpu.genblk1.mmu.r_writeable_d[8] ),
    .A1(net311),
    .S(_06021_),
    .X(_01913_));
 sg13g2_mux2_1 _24672_ (.A0(\cpu.genblk1.mmu.r_writeable_d[9] ),
    .A1(_03653_),
    .S(_06024_),
    .X(_01914_));
 sg13g2_nor2_2 _24673_ (.A(_09023_),
    .B(_09046_),
    .Y(_06227_));
 sg13g2_and3_1 _24674_ (.X(_06228_),
    .A(net965),
    .B(_00213_),
    .C(_06227_));
 sg13g2_buf_2 _24675_ (.A(_06228_),
    .X(_06229_));
 sg13g2_nand2_2 _24676_ (.Y(_06230_),
    .A(net1039),
    .B(_06229_));
 sg13g2_nor4_2 _24677_ (.A(net883),
    .B(_09335_),
    .C(net598),
    .Y(_06231_),
    .D(_06230_));
 sg13g2_mux2_1 _24678_ (.A0(\cpu.gpio.genblk2[4].srcs_io[0] ),
    .A1(net1022),
    .S(_06231_),
    .X(_01931_));
 sg13g2_mux2_1 _24679_ (.A0(\cpu.gpio.genblk2[5].srcs_io[0] ),
    .A1(net986),
    .S(_06231_),
    .X(_01932_));
 sg13g2_mux2_1 _24680_ (.A0(\cpu.gpio.genblk2[6].srcs_io[0] ),
    .A1(net974),
    .S(_06231_),
    .X(_01933_));
 sg13g2_mux2_1 _24681_ (.A0(\cpu.gpio.genblk2[7].srcs_io[0] ),
    .A1(net1019),
    .S(_06231_),
    .X(_01934_));
 sg13g2_and2_1 _24682_ (.A(net1039),
    .B(_06229_),
    .X(_06232_));
 sg13g2_buf_1 _24683_ (.A(_06232_),
    .X(_06233_));
 sg13g2_nand3_1 _24684_ (.B(_09923_),
    .C(_06233_),
    .A(net830),
    .Y(_06234_));
 sg13g2_buf_2 _24685_ (.A(_06234_),
    .X(_06235_));
 sg13g2_nand2_1 _24686_ (.Y(_06236_),
    .A(\cpu.gpio.genblk1[3].srcs_o[0] ),
    .B(_06235_));
 sg13g2_o21ai_1 _24687_ (.B1(_06236_),
    .Y(_01935_),
    .A1(_02749_),
    .A2(_06235_));
 sg13g2_nand2_1 _24688_ (.Y(_06237_),
    .A(\cpu.gpio.genblk1[4].srcs_o[0] ),
    .B(_06235_));
 sg13g2_o21ai_1 _24689_ (.B1(_06237_),
    .Y(_01936_),
    .A1(net720),
    .A2(_06235_));
 sg13g2_mux2_1 _24690_ (.A0(net849),
    .A1(\cpu.gpio.genblk1[5].srcs_o[0] ),
    .S(_06235_),
    .X(_01937_));
 sg13g2_mux2_1 _24691_ (.A0(_09957_),
    .A1(\cpu.gpio.genblk1[6].srcs_o[0] ),
    .S(_06235_),
    .X(_01938_));
 sg13g2_nand2_1 _24692_ (.Y(_06238_),
    .A(\cpu.gpio.genblk1[7].srcs_o[0] ),
    .B(_06235_));
 sg13g2_o21ai_1 _24693_ (.B1(_06238_),
    .Y(_01939_),
    .A1(net719),
    .A2(_06235_));
 sg13g2_and2_1 _24694_ (.A(_04966_),
    .B(_06233_),
    .X(_06239_));
 sg13g2_buf_1 _24695_ (.A(_06239_),
    .X(_06240_));
 sg13g2_mux2_1 _24696_ (.A0(_04965_),
    .A1(net880),
    .S(net76),
    .X(_01940_));
 sg13g2_buf_1 _24697_ (.A(\cpu.gpio.r_spi_miso_src[0][1] ),
    .X(_06241_));
 sg13g2_mux2_1 _24698_ (.A0(_06241_),
    .A1(net829),
    .S(net76),
    .X(_01941_));
 sg13g2_mux2_1 _24699_ (.A0(\cpu.gpio.r_spi_miso_src[0][2] ),
    .A1(_09937_),
    .S(net76),
    .X(_01942_));
 sg13g2_buf_1 _24700_ (.A(\cpu.gpio.r_spi_miso_src[0][3] ),
    .X(_06242_));
 sg13g2_mux2_1 _24701_ (.A0(_06242_),
    .A1(net1016),
    .S(net76),
    .X(_01943_));
 sg13g2_mux2_1 _24702_ (.A0(_05541_),
    .A1(net1022),
    .S(net76),
    .X(_01944_));
 sg13g2_inv_1 _24703_ (.Y(_06243_),
    .A(\cpu.gpio.r_spi_miso_src[1][1] ));
 sg13g2_nand2_1 _24704_ (.Y(_06244_),
    .A(net1021),
    .B(net76));
 sg13g2_o21ai_1 _24705_ (.B1(_06244_),
    .Y(_01945_),
    .A1(_06243_),
    .A2(_06240_));
 sg13g2_mux2_1 _24706_ (.A0(\cpu.gpio.r_spi_miso_src[1][2] ),
    .A1(net974),
    .S(net76),
    .X(_01946_));
 sg13g2_buf_1 _24707_ (.A(\cpu.gpio.r_spi_miso_src[1][3] ),
    .X(_06245_));
 sg13g2_mux2_1 _24708_ (.A0(_06245_),
    .A1(_09911_),
    .S(net76),
    .X(_01947_));
 sg13g2_and2_1 _24709_ (.A(net354),
    .B(_06233_),
    .X(_06246_));
 sg13g2_buf_4 _24710_ (.X(_06247_),
    .A(_06246_));
 sg13g2_mux2_1 _24711_ (.A0(_04971_),
    .A1(net877),
    .S(_06247_),
    .X(_01948_));
 sg13g2_mux2_1 _24712_ (.A0(_05315_),
    .A1(net829),
    .S(_06247_),
    .X(_01949_));
 sg13g2_mux2_1 _24713_ (.A0(_05368_),
    .A1(net876),
    .S(_06247_),
    .X(_01950_));
 sg13g2_mux2_1 _24714_ (.A0(_05453_),
    .A1(net1016),
    .S(_06247_),
    .X(_01951_));
 sg13g2_mux2_1 _24715_ (.A0(_05535_),
    .A1(net1022),
    .S(_06247_),
    .X(_01952_));
 sg13g2_mux2_1 _24716_ (.A0(_05607_),
    .A1(net986),
    .S(_06247_),
    .X(_01953_));
 sg13g2_mux2_1 _24717_ (.A0(_05693_),
    .A1(net974),
    .S(_06247_),
    .X(_01954_));
 sg13g2_mux2_1 _24718_ (.A0(_05105_),
    .A1(net1019),
    .S(_06247_),
    .X(_01955_));
 sg13g2_nor2_1 _24719_ (.A(_05314_),
    .B(_06230_),
    .Y(_06248_));
 sg13g2_buf_4 _24720_ (.X(_06249_),
    .A(_06248_));
 sg13g2_mux2_1 _24721_ (.A0(_04975_),
    .A1(net877),
    .S(_06249_),
    .X(_01956_));
 sg13g2_buf_1 _24722_ (.A(\cpu.gpio.r_src_io[6][1] ),
    .X(_06250_));
 sg13g2_mux2_1 _24723_ (.A0(_06250_),
    .A1(_12104_),
    .S(_06249_),
    .X(_01957_));
 sg13g2_mux2_1 _24724_ (.A0(\cpu.gpio.r_src_io[6][2] ),
    .A1(net876),
    .S(_06249_),
    .X(_01958_));
 sg13g2_mux2_1 _24725_ (.A0(\cpu.gpio.r_src_io[6][3] ),
    .A1(net1016),
    .S(_06249_),
    .X(_01959_));
 sg13g2_mux2_1 _24726_ (.A0(_05537_),
    .A1(net1022),
    .S(_06249_),
    .X(_01960_));
 sg13g2_buf_1 _24727_ (.A(\cpu.gpio.r_src_io[7][1] ),
    .X(_06251_));
 sg13g2_mux2_1 _24728_ (.A0(_06251_),
    .A1(net986),
    .S(_06249_),
    .X(_01961_));
 sg13g2_mux2_1 _24729_ (.A0(\cpu.gpio.r_src_io[7][2] ),
    .A1(net974),
    .S(_06249_),
    .X(_01962_));
 sg13g2_mux2_1 _24730_ (.A0(\cpu.gpio.r_src_io[7][3] ),
    .A1(net1019),
    .S(_06249_),
    .X(_01963_));
 sg13g2_nor2_2 _24731_ (.A(_05606_),
    .B(_06230_),
    .Y(_06252_));
 sg13g2_mux2_1 _24732_ (.A0(_05531_),
    .A1(_09896_),
    .S(_06252_),
    .X(_01964_));
 sg13g2_buf_1 _24733_ (.A(\cpu.gpio.r_src_o[3][1] ),
    .X(_06253_));
 sg13g2_mux2_1 _24734_ (.A0(_06253_),
    .A1(net986),
    .S(_06252_),
    .X(_01965_));
 sg13g2_mux2_1 _24735_ (.A0(\cpu.gpio.r_src_o[3][2] ),
    .A1(_12569_),
    .S(_06252_),
    .X(_01966_));
 sg13g2_mux2_1 _24736_ (.A0(\cpu.gpio.r_src_o[3][3] ),
    .A1(net1019),
    .S(_06252_),
    .X(_01967_));
 sg13g2_nand2_1 _24737_ (.Y(_06254_),
    .A(_04981_),
    .B(_06233_));
 sg13g2_buf_1 _24738_ (.A(_06254_),
    .X(_06255_));
 sg13g2_mux2_1 _24739_ (.A0(_09861_),
    .A1(_04982_),
    .S(net75),
    .X(_01968_));
 sg13g2_buf_1 _24740_ (.A(\cpu.gpio.r_src_o[4][1] ),
    .X(_06256_));
 sg13g2_mux2_1 _24741_ (.A0(_05780_),
    .A1(_06256_),
    .S(net75),
    .X(_01969_));
 sg13g2_nand2_1 _24742_ (.Y(_06257_),
    .A(\cpu.gpio.r_src_o[4][2] ),
    .B(_06255_));
 sg13g2_o21ai_1 _24743_ (.B1(_06257_),
    .Y(_01970_),
    .A1(_09884_),
    .A2(_06255_));
 sg13g2_nand2_1 _24744_ (.Y(_06258_),
    .A(\cpu.gpio.r_src_o[4][3] ),
    .B(net75));
 sg13g2_o21ai_1 _24745_ (.B1(_06258_),
    .Y(_01971_),
    .A1(_02749_),
    .A2(net75));
 sg13g2_nand2_1 _24746_ (.Y(_06259_),
    .A(_05538_),
    .B(_06254_));
 sg13g2_o21ai_1 _24747_ (.B1(_06259_),
    .Y(_01972_),
    .A1(net720),
    .A2(net75));
 sg13g2_buf_1 _24748_ (.A(\cpu.gpio.r_src_o[5][1] ),
    .X(_06260_));
 sg13g2_mux2_1 _24749_ (.A0(_12522_),
    .A1(_06260_),
    .S(net75),
    .X(_01973_));
 sg13g2_mux2_1 _24750_ (.A0(net875),
    .A1(\cpu.gpio.r_src_o[5][2] ),
    .S(net75),
    .X(_01974_));
 sg13g2_nand2_1 _24751_ (.Y(_06261_),
    .A(\cpu.gpio.r_src_o[5][3] ),
    .B(_06254_));
 sg13g2_o21ai_1 _24752_ (.B1(_06261_),
    .Y(_01975_),
    .A1(net719),
    .A2(net75));
 sg13g2_nor2_2 _24753_ (.A(_04979_),
    .B(_06230_),
    .Y(_06262_));
 sg13g2_mux2_1 _24754_ (.A0(_05530_),
    .A1(_09896_),
    .S(_06262_),
    .X(_01980_));
 sg13g2_buf_1 _24755_ (.A(\cpu.gpio.r_src_o[7][1] ),
    .X(_06263_));
 sg13g2_mux2_1 _24756_ (.A0(_06263_),
    .A1(net986),
    .S(_06262_),
    .X(_01981_));
 sg13g2_mux2_1 _24757_ (.A0(\cpu.gpio.r_src_o[7][2] ),
    .A1(_12569_),
    .S(_06262_),
    .X(_01982_));
 sg13g2_mux2_1 _24758_ (.A0(\cpu.gpio.r_src_o[7][3] ),
    .A1(_09911_),
    .S(_06262_),
    .X(_01983_));
 sg13g2_buf_1 _24759_ (.A(_12143_),
    .X(_06264_));
 sg13g2_and2_1 _24760_ (.A(net689),
    .B(_08742_),
    .X(_06265_));
 sg13g2_buf_4 _24761_ (.X(_06266_),
    .A(_06265_));
 sg13g2_nor2_1 _24762_ (.A(\cpu.icache.r_offset[2] ),
    .B(_00231_),
    .Y(_06267_));
 sg13g2_buf_2 _24763_ (.A(_06267_),
    .X(_06268_));
 sg13g2_buf_1 _24764_ (.A(\cpu.icache.r_offset[1] ),
    .X(_06269_));
 sg13g2_buf_1 _24765_ (.A(\cpu.icache.r_offset[0] ),
    .X(_06270_));
 sg13g2_nor2b_1 _24766_ (.A(_06269_),
    .B_N(_06270_),
    .Y(_06271_));
 sg13g2_buf_1 _24767_ (.A(_06271_),
    .X(_06272_));
 sg13g2_and2_1 _24768_ (.A(_06268_),
    .B(_06272_),
    .X(_06273_));
 sg13g2_buf_2 _24769_ (.A(_06273_),
    .X(_06274_));
 sg13g2_nand2_2 _24770_ (.Y(_06275_),
    .A(_06266_),
    .B(_06274_));
 sg13g2_mux2_1 _24771_ (.A0(net940),
    .A1(\cpu.icache.r_data[0][0] ),
    .S(_06275_),
    .X(_01987_));
 sg13g2_buf_1 _24772_ (.A(net969),
    .X(_06276_));
 sg13g2_inv_1 _24773_ (.Y(_06277_),
    .A(_00231_));
 sg13g2_buf_1 _24774_ (.A(_00232_),
    .X(_06278_));
 sg13g2_nand4_1 _24775_ (.B(_06270_),
    .C(_06277_),
    .A(_06269_),
    .Y(_06279_),
    .D(_06278_));
 sg13g2_buf_2 _24776_ (.A(_06279_),
    .X(_06280_));
 sg13g2_inv_1 _24777_ (.Y(_06281_),
    .A(_06280_));
 sg13g2_nand2_2 _24778_ (.Y(_06282_),
    .A(_06266_),
    .B(_06281_));
 sg13g2_mux2_1 _24779_ (.A0(net810),
    .A1(\cpu.icache.r_data[0][10] ),
    .S(_06282_),
    .X(_01988_));
 sg13g2_buf_1 _24780_ (.A(net968),
    .X(_06283_));
 sg13g2_mux2_1 _24781_ (.A0(net809),
    .A1(\cpu.icache.r_data[0][11] ),
    .S(_06282_),
    .X(_01989_));
 sg13g2_nor2b_1 _24782_ (.A(_06270_),
    .B_N(_06269_),
    .Y(_06284_));
 sg13g2_buf_1 _24783_ (.A(_06284_),
    .X(_06285_));
 sg13g2_and2_1 _24784_ (.A(_06268_),
    .B(_06285_),
    .X(_06286_));
 sg13g2_buf_2 _24785_ (.A(_06286_),
    .X(_06287_));
 sg13g2_nand2_2 _24786_ (.Y(_06288_),
    .A(_06266_),
    .B(_06287_));
 sg13g2_mux2_1 _24787_ (.A0(_06264_),
    .A1(\cpu.icache.r_data[0][12] ),
    .S(_06288_),
    .X(_01990_));
 sg13g2_buf_1 _24788_ (.A(_03029_),
    .X(_06289_));
 sg13g2_mux2_1 _24789_ (.A0(net939),
    .A1(\cpu.icache.r_data[0][13] ),
    .S(_06288_),
    .X(_01991_));
 sg13g2_mux2_1 _24790_ (.A0(net810),
    .A1(\cpu.icache.r_data[0][14] ),
    .S(_06288_),
    .X(_01992_));
 sg13g2_mux2_1 _24791_ (.A0(net809),
    .A1(\cpu.icache.r_data[0][15] ),
    .S(_06288_),
    .X(_01993_));
 sg13g2_nor2_1 _24792_ (.A(_00231_),
    .B(_06278_),
    .Y(_06290_));
 sg13g2_buf_2 _24793_ (.A(_06290_),
    .X(_06291_));
 sg13g2_and2_1 _24794_ (.A(_06272_),
    .B(_06291_),
    .X(_06292_));
 sg13g2_buf_2 _24795_ (.A(_06292_),
    .X(_06293_));
 sg13g2_nand2_2 _24796_ (.Y(_06294_),
    .A(_06266_),
    .B(_06293_));
 sg13g2_mux2_1 _24797_ (.A0(net940),
    .A1(\cpu.icache.r_data[0][16] ),
    .S(_06294_),
    .X(_01994_));
 sg13g2_mux2_1 _24798_ (.A0(net939),
    .A1(\cpu.icache.r_data[0][17] ),
    .S(_06294_),
    .X(_01995_));
 sg13g2_mux2_1 _24799_ (.A0(_06276_),
    .A1(\cpu.icache.r_data[0][18] ),
    .S(_06294_),
    .X(_01996_));
 sg13g2_mux2_1 _24800_ (.A0(net809),
    .A1(\cpu.icache.r_data[0][19] ),
    .S(_06294_),
    .X(_01997_));
 sg13g2_mux2_1 _24801_ (.A0(net939),
    .A1(\cpu.icache.r_data[0][1] ),
    .S(_06275_),
    .X(_01998_));
 sg13g2_nor2_2 _24802_ (.A(_06269_),
    .B(_06270_),
    .Y(_06295_));
 sg13g2_and2_1 _24803_ (.A(_06291_),
    .B(_06295_),
    .X(_06296_));
 sg13g2_buf_2 _24804_ (.A(_06296_),
    .X(_06297_));
 sg13g2_nand2_2 _24805_ (.Y(_06298_),
    .A(_06266_),
    .B(_06297_));
 sg13g2_mux2_1 _24806_ (.A0(net940),
    .A1(\cpu.icache.r_data[0][20] ),
    .S(_06298_),
    .X(_01999_));
 sg13g2_mux2_1 _24807_ (.A0(net939),
    .A1(\cpu.icache.r_data[0][21] ),
    .S(_06298_),
    .X(_02000_));
 sg13g2_mux2_1 _24808_ (.A0(net810),
    .A1(\cpu.icache.r_data[0][22] ),
    .S(_06298_),
    .X(_02001_));
 sg13g2_mux2_1 _24809_ (.A0(net809),
    .A1(\cpu.icache.r_data[0][23] ),
    .S(_06298_),
    .X(_02002_));
 sg13g2_inv_1 _24810_ (.Y(_06299_),
    .A(\cpu.i_wstrobe_d ));
 sg13g2_nand2_2 _24811_ (.Y(_06300_),
    .A(_06269_),
    .B(_06270_));
 sg13g2_nor3_2 _24812_ (.A(_06278_),
    .B(_06299_),
    .C(_06300_),
    .Y(_06301_));
 sg13g2_nand2_1 _24813_ (.Y(_06302_),
    .A(_06266_),
    .B(_06301_));
 sg13g2_buf_1 _24814_ (.A(_06302_),
    .X(_06303_));
 sg13g2_buf_1 _24815_ (.A(net398),
    .X(_06304_));
 sg13g2_mux2_1 _24816_ (.A0(net940),
    .A1(\cpu.icache.r_data[0][24] ),
    .S(net310),
    .X(_02003_));
 sg13g2_mux2_1 _24817_ (.A0(net939),
    .A1(\cpu.icache.r_data[0][25] ),
    .S(net310),
    .X(_02004_));
 sg13g2_mux2_1 _24818_ (.A0(net810),
    .A1(\cpu.icache.r_data[0][26] ),
    .S(_06304_),
    .X(_02005_));
 sg13g2_mux2_1 _24819_ (.A0(net809),
    .A1(\cpu.icache.r_data[0][27] ),
    .S(_06304_),
    .X(_02006_));
 sg13g2_and2_1 _24820_ (.A(_06285_),
    .B(_06291_),
    .X(_06305_));
 sg13g2_buf_2 _24821_ (.A(_06305_),
    .X(_06306_));
 sg13g2_nand2_2 _24822_ (.Y(_06307_),
    .A(_06266_),
    .B(_06306_));
 sg13g2_mux2_1 _24823_ (.A0(net940),
    .A1(\cpu.icache.r_data[0][28] ),
    .S(_06307_),
    .X(_02007_));
 sg13g2_mux2_1 _24824_ (.A0(net939),
    .A1(\cpu.icache.r_data[0][29] ),
    .S(_06307_),
    .X(_02008_));
 sg13g2_mux2_1 _24825_ (.A0(net810),
    .A1(\cpu.icache.r_data[0][2] ),
    .S(_06275_),
    .X(_02009_));
 sg13g2_mux2_1 _24826_ (.A0(net810),
    .A1(\cpu.icache.r_data[0][30] ),
    .S(_06307_),
    .X(_02010_));
 sg13g2_mux2_1 _24827_ (.A0(net809),
    .A1(\cpu.icache.r_data[0][31] ),
    .S(_06307_),
    .X(_02011_));
 sg13g2_mux2_1 _24828_ (.A0(_06283_),
    .A1(\cpu.icache.r_data[0][3] ),
    .S(_06275_),
    .X(_02012_));
 sg13g2_and2_1 _24829_ (.A(_06268_),
    .B(_06295_),
    .X(_06308_));
 sg13g2_buf_2 _24830_ (.A(_06308_),
    .X(_06309_));
 sg13g2_nand2_2 _24831_ (.Y(_06310_),
    .A(_06266_),
    .B(_06309_));
 sg13g2_mux2_1 _24832_ (.A0(net940),
    .A1(\cpu.icache.r_data[0][4] ),
    .S(_06310_),
    .X(_02013_));
 sg13g2_mux2_1 _24833_ (.A0(net939),
    .A1(\cpu.icache.r_data[0][5] ),
    .S(_06310_),
    .X(_02014_));
 sg13g2_mux2_1 _24834_ (.A0(net810),
    .A1(\cpu.icache.r_data[0][6] ),
    .S(_06310_),
    .X(_02015_));
 sg13g2_mux2_1 _24835_ (.A0(net809),
    .A1(\cpu.icache.r_data[0][7] ),
    .S(_06310_),
    .X(_02016_));
 sg13g2_mux2_1 _24836_ (.A0(_06264_),
    .A1(\cpu.icache.r_data[0][8] ),
    .S(_06282_),
    .X(_02017_));
 sg13g2_mux2_1 _24837_ (.A0(_06289_),
    .A1(\cpu.icache.r_data[0][9] ),
    .S(_06282_),
    .X(_02018_));
 sg13g2_buf_1 _24838_ (.A(_12143_),
    .X(_06311_));
 sg13g2_nand2b_1 _24839_ (.Y(_06312_),
    .B(_08752_),
    .A_N(_08667_));
 sg13g2_buf_4 _24840_ (.X(_06313_),
    .A(_06312_));
 sg13g2_nand2_2 _24841_ (.Y(_06314_),
    .A(_06268_),
    .B(_06272_));
 sg13g2_nor2_2 _24842_ (.A(_06313_),
    .B(_06314_),
    .Y(_06315_));
 sg13g2_mux2_1 _24843_ (.A0(\cpu.icache.r_data[1][0] ),
    .A1(net938),
    .S(_06315_),
    .X(_02019_));
 sg13g2_buf_1 _24844_ (.A(net969),
    .X(_06316_));
 sg13g2_nor2_2 _24845_ (.A(_06313_),
    .B(_06280_),
    .Y(_06317_));
 sg13g2_mux2_1 _24846_ (.A0(\cpu.icache.r_data[1][10] ),
    .A1(net808),
    .S(_06317_),
    .X(_02020_));
 sg13g2_buf_1 _24847_ (.A(net968),
    .X(_06318_));
 sg13g2_mux2_1 _24848_ (.A0(\cpu.icache.r_data[1][11] ),
    .A1(_06318_),
    .S(_06317_),
    .X(_02021_));
 sg13g2_buf_1 _24849_ (.A(_12143_),
    .X(_06319_));
 sg13g2_nand2_2 _24850_ (.Y(_06320_),
    .A(_06268_),
    .B(_06285_));
 sg13g2_nor2_2 _24851_ (.A(_06313_),
    .B(_06320_),
    .Y(_06321_));
 sg13g2_mux2_1 _24852_ (.A0(\cpu.icache.r_data[1][12] ),
    .A1(net937),
    .S(_06321_),
    .X(_02022_));
 sg13g2_buf_1 _24853_ (.A(_03029_),
    .X(_06322_));
 sg13g2_mux2_1 _24854_ (.A0(\cpu.icache.r_data[1][13] ),
    .A1(net936),
    .S(_06321_),
    .X(_02023_));
 sg13g2_buf_1 _24855_ (.A(_02918_),
    .X(_06323_));
 sg13g2_mux2_1 _24856_ (.A0(\cpu.icache.r_data[1][14] ),
    .A1(net806),
    .S(_06321_),
    .X(_02024_));
 sg13g2_buf_1 _24857_ (.A(net968),
    .X(_06324_));
 sg13g2_mux2_1 _24858_ (.A0(\cpu.icache.r_data[1][15] ),
    .A1(net805),
    .S(_06321_),
    .X(_02025_));
 sg13g2_nand2_2 _24859_ (.Y(_06325_),
    .A(_06272_),
    .B(_06291_));
 sg13g2_nor2_2 _24860_ (.A(_06313_),
    .B(_06325_),
    .Y(_06326_));
 sg13g2_mux2_1 _24861_ (.A0(\cpu.icache.r_data[1][16] ),
    .A1(net937),
    .S(_06326_),
    .X(_02026_));
 sg13g2_buf_1 _24862_ (.A(_03029_),
    .X(_06327_));
 sg13g2_mux2_1 _24863_ (.A0(\cpu.icache.r_data[1][17] ),
    .A1(net935),
    .S(_06326_),
    .X(_02027_));
 sg13g2_mux2_1 _24864_ (.A0(\cpu.icache.r_data[1][18] ),
    .A1(net806),
    .S(_06326_),
    .X(_02028_));
 sg13g2_mux2_1 _24865_ (.A0(\cpu.icache.r_data[1][19] ),
    .A1(net805),
    .S(_06326_),
    .X(_02029_));
 sg13g2_mux2_1 _24866_ (.A0(\cpu.icache.r_data[1][1] ),
    .A1(net935),
    .S(_06315_),
    .X(_02030_));
 sg13g2_nand2_2 _24867_ (.Y(_06328_),
    .A(_06291_),
    .B(_06295_));
 sg13g2_nor2_2 _24868_ (.A(_06313_),
    .B(_06328_),
    .Y(_06329_));
 sg13g2_mux2_1 _24869_ (.A0(\cpu.icache.r_data[1][20] ),
    .A1(net937),
    .S(_06329_),
    .X(_02031_));
 sg13g2_mux2_1 _24870_ (.A0(\cpu.icache.r_data[1][21] ),
    .A1(net935),
    .S(_06329_),
    .X(_02032_));
 sg13g2_mux2_1 _24871_ (.A0(\cpu.icache.r_data[1][22] ),
    .A1(net806),
    .S(_06329_),
    .X(_02033_));
 sg13g2_mux2_1 _24872_ (.A0(\cpu.icache.r_data[1][23] ),
    .A1(net805),
    .S(_06329_),
    .X(_02034_));
 sg13g2_or3_1 _24873_ (.A(_06278_),
    .B(_06299_),
    .C(_06300_),
    .X(_06330_));
 sg13g2_buf_1 _24874_ (.A(_06330_),
    .X(_06331_));
 sg13g2_nor2_1 _24875_ (.A(_06313_),
    .B(_06331_),
    .Y(_06332_));
 sg13g2_buf_2 _24876_ (.A(_06332_),
    .X(_06333_));
 sg13g2_mux2_1 _24877_ (.A0(\cpu.icache.r_data[1][24] ),
    .A1(net937),
    .S(_06333_),
    .X(_02035_));
 sg13g2_mux2_1 _24878_ (.A0(\cpu.icache.r_data[1][25] ),
    .A1(net935),
    .S(_06333_),
    .X(_02036_));
 sg13g2_mux2_1 _24879_ (.A0(\cpu.icache.r_data[1][26] ),
    .A1(_06323_),
    .S(_06333_),
    .X(_02037_));
 sg13g2_mux2_1 _24880_ (.A0(\cpu.icache.r_data[1][27] ),
    .A1(_06324_),
    .S(_06333_),
    .X(_02038_));
 sg13g2_nand2_2 _24881_ (.Y(_06334_),
    .A(_06285_),
    .B(_06291_));
 sg13g2_nor2_2 _24882_ (.A(_06313_),
    .B(_06334_),
    .Y(_06335_));
 sg13g2_mux2_1 _24883_ (.A0(\cpu.icache.r_data[1][28] ),
    .A1(net937),
    .S(_06335_),
    .X(_02039_));
 sg13g2_mux2_1 _24884_ (.A0(\cpu.icache.r_data[1][29] ),
    .A1(net935),
    .S(_06335_),
    .X(_02040_));
 sg13g2_mux2_1 _24885_ (.A0(\cpu.icache.r_data[1][2] ),
    .A1(net806),
    .S(_06315_),
    .X(_02041_));
 sg13g2_mux2_1 _24886_ (.A0(\cpu.icache.r_data[1][30] ),
    .A1(net806),
    .S(_06335_),
    .X(_02042_));
 sg13g2_mux2_1 _24887_ (.A0(\cpu.icache.r_data[1][31] ),
    .A1(net805),
    .S(_06335_),
    .X(_02043_));
 sg13g2_mux2_1 _24888_ (.A0(\cpu.icache.r_data[1][3] ),
    .A1(net805),
    .S(_06315_),
    .X(_02044_));
 sg13g2_nand2_2 _24889_ (.Y(_06336_),
    .A(_06268_),
    .B(_06295_));
 sg13g2_nor2_2 _24890_ (.A(_06313_),
    .B(_06336_),
    .Y(_06337_));
 sg13g2_mux2_1 _24891_ (.A0(\cpu.icache.r_data[1][4] ),
    .A1(net937),
    .S(_06337_),
    .X(_02045_));
 sg13g2_mux2_1 _24892_ (.A0(\cpu.icache.r_data[1][5] ),
    .A1(net935),
    .S(_06337_),
    .X(_02046_));
 sg13g2_mux2_1 _24893_ (.A0(\cpu.icache.r_data[1][6] ),
    .A1(net806),
    .S(_06337_),
    .X(_02047_));
 sg13g2_mux2_1 _24894_ (.A0(\cpu.icache.r_data[1][7] ),
    .A1(net805),
    .S(_06337_),
    .X(_02048_));
 sg13g2_mux2_1 _24895_ (.A0(\cpu.icache.r_data[1][8] ),
    .A1(net937),
    .S(_06317_),
    .X(_02049_));
 sg13g2_mux2_1 _24896_ (.A0(\cpu.icache.r_data[1][9] ),
    .A1(net935),
    .S(_06317_),
    .X(_02050_));
 sg13g2_nand2_1 _24897_ (.Y(_06338_),
    .A(net915),
    .B(_08291_));
 sg13g2_buf_4 _24898_ (.X(_06339_),
    .A(_06338_));
 sg13g2_nor2_2 _24899_ (.A(_06339_),
    .B(_06314_),
    .Y(_06340_));
 sg13g2_mux2_1 _24900_ (.A0(\cpu.icache.r_data[2][0] ),
    .A1(_06319_),
    .S(_06340_),
    .X(_02051_));
 sg13g2_nor2_2 _24901_ (.A(_06339_),
    .B(_06280_),
    .Y(_06341_));
 sg13g2_mux2_1 _24902_ (.A0(\cpu.icache.r_data[2][10] ),
    .A1(_06323_),
    .S(_06341_),
    .X(_02052_));
 sg13g2_mux2_1 _24903_ (.A0(\cpu.icache.r_data[2][11] ),
    .A1(net805),
    .S(_06341_),
    .X(_02053_));
 sg13g2_nor2_2 _24904_ (.A(_06339_),
    .B(_06320_),
    .Y(_06342_));
 sg13g2_mux2_1 _24905_ (.A0(\cpu.icache.r_data[2][12] ),
    .A1(net937),
    .S(_06342_),
    .X(_02054_));
 sg13g2_mux2_1 _24906_ (.A0(\cpu.icache.r_data[2][13] ),
    .A1(net935),
    .S(_06342_),
    .X(_02055_));
 sg13g2_mux2_1 _24907_ (.A0(\cpu.icache.r_data[2][14] ),
    .A1(net806),
    .S(_06342_),
    .X(_02056_));
 sg13g2_mux2_1 _24908_ (.A0(\cpu.icache.r_data[2][15] ),
    .A1(net805),
    .S(_06342_),
    .X(_02057_));
 sg13g2_nor2_2 _24909_ (.A(_06339_),
    .B(_06325_),
    .Y(_06343_));
 sg13g2_mux2_1 _24910_ (.A0(\cpu.icache.r_data[2][16] ),
    .A1(_06319_),
    .S(_06343_),
    .X(_02058_));
 sg13g2_mux2_1 _24911_ (.A0(\cpu.icache.r_data[2][17] ),
    .A1(_06327_),
    .S(_06343_),
    .X(_02059_));
 sg13g2_mux2_1 _24912_ (.A0(\cpu.icache.r_data[2][18] ),
    .A1(net806),
    .S(_06343_),
    .X(_02060_));
 sg13g2_mux2_1 _24913_ (.A0(\cpu.icache.r_data[2][19] ),
    .A1(_06324_),
    .S(_06343_),
    .X(_02061_));
 sg13g2_mux2_1 _24914_ (.A0(\cpu.icache.r_data[2][1] ),
    .A1(_06327_),
    .S(_06340_),
    .X(_02062_));
 sg13g2_buf_1 _24915_ (.A(_12143_),
    .X(_06344_));
 sg13g2_nor2_2 _24916_ (.A(_06339_),
    .B(_06328_),
    .Y(_06345_));
 sg13g2_mux2_1 _24917_ (.A0(\cpu.icache.r_data[2][20] ),
    .A1(net934),
    .S(_06345_),
    .X(_02063_));
 sg13g2_buf_1 _24918_ (.A(_03029_),
    .X(_06346_));
 sg13g2_mux2_1 _24919_ (.A0(\cpu.icache.r_data[2][21] ),
    .A1(net933),
    .S(_06345_),
    .X(_02064_));
 sg13g2_buf_1 _24920_ (.A(_12107_),
    .X(_06347_));
 sg13g2_mux2_1 _24921_ (.A0(\cpu.icache.r_data[2][22] ),
    .A1(net932),
    .S(_06345_),
    .X(_02065_));
 sg13g2_buf_1 _24922_ (.A(net968),
    .X(_06348_));
 sg13g2_mux2_1 _24923_ (.A0(\cpu.icache.r_data[2][23] ),
    .A1(net804),
    .S(_06345_),
    .X(_02066_));
 sg13g2_nor2_1 _24924_ (.A(_06339_),
    .B(_06331_),
    .Y(_06349_));
 sg13g2_buf_2 _24925_ (.A(_06349_),
    .X(_06350_));
 sg13g2_mux2_1 _24926_ (.A0(\cpu.icache.r_data[2][24] ),
    .A1(net934),
    .S(_06350_),
    .X(_02067_));
 sg13g2_mux2_1 _24927_ (.A0(\cpu.icache.r_data[2][25] ),
    .A1(net933),
    .S(_06350_),
    .X(_02068_));
 sg13g2_mux2_1 _24928_ (.A0(\cpu.icache.r_data[2][26] ),
    .A1(_06347_),
    .S(_06350_),
    .X(_02069_));
 sg13g2_mux2_1 _24929_ (.A0(\cpu.icache.r_data[2][27] ),
    .A1(net804),
    .S(_06350_),
    .X(_02070_));
 sg13g2_nor2_2 _24930_ (.A(_06339_),
    .B(_06334_),
    .Y(_06351_));
 sg13g2_mux2_1 _24931_ (.A0(\cpu.icache.r_data[2][28] ),
    .A1(net934),
    .S(_06351_),
    .X(_02071_));
 sg13g2_mux2_1 _24932_ (.A0(\cpu.icache.r_data[2][29] ),
    .A1(net933),
    .S(_06351_),
    .X(_02072_));
 sg13g2_mux2_1 _24933_ (.A0(\cpu.icache.r_data[2][2] ),
    .A1(net932),
    .S(_06340_),
    .X(_02073_));
 sg13g2_mux2_1 _24934_ (.A0(\cpu.icache.r_data[2][30] ),
    .A1(net932),
    .S(_06351_),
    .X(_02074_));
 sg13g2_mux2_1 _24935_ (.A0(\cpu.icache.r_data[2][31] ),
    .A1(net804),
    .S(_06351_),
    .X(_02075_));
 sg13g2_mux2_1 _24936_ (.A0(\cpu.icache.r_data[2][3] ),
    .A1(net804),
    .S(_06340_),
    .X(_02076_));
 sg13g2_nor2_2 _24937_ (.A(_06339_),
    .B(_06336_),
    .Y(_06352_));
 sg13g2_mux2_1 _24938_ (.A0(\cpu.icache.r_data[2][4] ),
    .A1(net934),
    .S(_06352_),
    .X(_02077_));
 sg13g2_mux2_1 _24939_ (.A0(\cpu.icache.r_data[2][5] ),
    .A1(net933),
    .S(_06352_),
    .X(_02078_));
 sg13g2_mux2_1 _24940_ (.A0(\cpu.icache.r_data[2][6] ),
    .A1(net932),
    .S(_06352_),
    .X(_02079_));
 sg13g2_mux2_1 _24941_ (.A0(\cpu.icache.r_data[2][7] ),
    .A1(net804),
    .S(_06352_),
    .X(_02080_));
 sg13g2_mux2_1 _24942_ (.A0(\cpu.icache.r_data[2][8] ),
    .A1(net934),
    .S(_06341_),
    .X(_02081_));
 sg13g2_mux2_1 _24943_ (.A0(\cpu.icache.r_data[2][9] ),
    .A1(net933),
    .S(_06341_),
    .X(_02082_));
 sg13g2_nand2_2 _24944_ (.Y(_06353_),
    .A(_08889_),
    .B(_06274_));
 sg13g2_mux2_1 _24945_ (.A0(net940),
    .A1(\cpu.icache.r_data[3][0] ),
    .S(_06353_),
    .X(_02083_));
 sg13g2_and2_1 _24946_ (.A(net433),
    .B(_06281_),
    .X(_06354_));
 sg13g2_buf_1 _24947_ (.A(_06354_),
    .X(_06355_));
 sg13g2_mux2_1 _24948_ (.A0(\cpu.icache.r_data[3][10] ),
    .A1(net932),
    .S(_06355_),
    .X(_02084_));
 sg13g2_mux2_1 _24949_ (.A0(\cpu.icache.r_data[3][11] ),
    .A1(net804),
    .S(_06355_),
    .X(_02085_));
 sg13g2_nand2_2 _24950_ (.Y(_06356_),
    .A(net433),
    .B(_06287_));
 sg13g2_mux2_1 _24951_ (.A0(net940),
    .A1(\cpu.icache.r_data[3][12] ),
    .S(_06356_),
    .X(_02086_));
 sg13g2_mux2_1 _24952_ (.A0(net939),
    .A1(\cpu.icache.r_data[3][13] ),
    .S(_06356_),
    .X(_02087_));
 sg13g2_mux2_1 _24953_ (.A0(net810),
    .A1(\cpu.icache.r_data[3][14] ),
    .S(_06356_),
    .X(_02088_));
 sg13g2_mux2_1 _24954_ (.A0(_06283_),
    .A1(\cpu.icache.r_data[3][15] ),
    .S(_06356_),
    .X(_02089_));
 sg13g2_buf_1 _24955_ (.A(_12143_),
    .X(_06357_));
 sg13g2_nand2_2 _24956_ (.Y(_06358_),
    .A(net433),
    .B(_06293_));
 sg13g2_mux2_1 _24957_ (.A0(net931),
    .A1(\cpu.icache.r_data[3][16] ),
    .S(_06358_),
    .X(_02090_));
 sg13g2_mux2_1 _24958_ (.A0(_06289_),
    .A1(\cpu.icache.r_data[3][17] ),
    .S(_06358_),
    .X(_02091_));
 sg13g2_mux2_1 _24959_ (.A0(_06276_),
    .A1(\cpu.icache.r_data[3][18] ),
    .S(_06358_),
    .X(_02092_));
 sg13g2_mux2_1 _24960_ (.A0(net809),
    .A1(\cpu.icache.r_data[3][19] ),
    .S(_06358_),
    .X(_02093_));
 sg13g2_buf_1 _24961_ (.A(_03029_),
    .X(_06359_));
 sg13g2_mux2_1 _24962_ (.A0(net930),
    .A1(\cpu.icache.r_data[3][1] ),
    .S(_06353_),
    .X(_02094_));
 sg13g2_nand2_2 _24963_ (.Y(_06360_),
    .A(net433),
    .B(_06297_));
 sg13g2_mux2_1 _24964_ (.A0(net931),
    .A1(\cpu.icache.r_data[3][20] ),
    .S(_06360_),
    .X(_02095_));
 sg13g2_mux2_1 _24965_ (.A0(net930),
    .A1(\cpu.icache.r_data[3][21] ),
    .S(_06360_),
    .X(_02096_));
 sg13g2_buf_1 _24966_ (.A(_02918_),
    .X(_06361_));
 sg13g2_mux2_1 _24967_ (.A0(net803),
    .A1(\cpu.icache.r_data[3][22] ),
    .S(_06360_),
    .X(_02097_));
 sg13g2_buf_1 _24968_ (.A(_02963_),
    .X(_06362_));
 sg13g2_mux2_1 _24969_ (.A0(net802),
    .A1(\cpu.icache.r_data[3][23] ),
    .S(_06360_),
    .X(_02098_));
 sg13g2_nand2_1 _24970_ (.Y(_06363_),
    .A(net433),
    .B(_06301_));
 sg13g2_buf_1 _24971_ (.A(_06363_),
    .X(_06364_));
 sg13g2_buf_1 _24972_ (.A(net262),
    .X(_06365_));
 sg13g2_mux2_1 _24973_ (.A0(_06357_),
    .A1(\cpu.icache.r_data[3][24] ),
    .S(net236),
    .X(_02099_));
 sg13g2_mux2_1 _24974_ (.A0(net930),
    .A1(\cpu.icache.r_data[3][25] ),
    .S(net236),
    .X(_02100_));
 sg13g2_mux2_1 _24975_ (.A0(net803),
    .A1(\cpu.icache.r_data[3][26] ),
    .S(_06365_),
    .X(_02101_));
 sg13g2_mux2_1 _24976_ (.A0(_06362_),
    .A1(\cpu.icache.r_data[3][27] ),
    .S(_06365_),
    .X(_02102_));
 sg13g2_nand2_2 _24977_ (.Y(_06366_),
    .A(net433),
    .B(_06306_));
 sg13g2_mux2_1 _24978_ (.A0(net931),
    .A1(\cpu.icache.r_data[3][28] ),
    .S(_06366_),
    .X(_02103_));
 sg13g2_mux2_1 _24979_ (.A0(net930),
    .A1(\cpu.icache.r_data[3][29] ),
    .S(_06366_),
    .X(_02104_));
 sg13g2_mux2_1 _24980_ (.A0(_06361_),
    .A1(\cpu.icache.r_data[3][2] ),
    .S(_06353_),
    .X(_02105_));
 sg13g2_mux2_1 _24981_ (.A0(net803),
    .A1(\cpu.icache.r_data[3][30] ),
    .S(_06366_),
    .X(_02106_));
 sg13g2_mux2_1 _24982_ (.A0(net802),
    .A1(\cpu.icache.r_data[3][31] ),
    .S(_06366_),
    .X(_02107_));
 sg13g2_mux2_1 _24983_ (.A0(net802),
    .A1(\cpu.icache.r_data[3][3] ),
    .S(_06353_),
    .X(_02108_));
 sg13g2_nand2_2 _24984_ (.Y(_06367_),
    .A(net433),
    .B(_06309_));
 sg13g2_mux2_1 _24985_ (.A0(net931),
    .A1(\cpu.icache.r_data[3][4] ),
    .S(_06367_),
    .X(_02109_));
 sg13g2_mux2_1 _24986_ (.A0(net930),
    .A1(\cpu.icache.r_data[3][5] ),
    .S(_06367_),
    .X(_02110_));
 sg13g2_mux2_1 _24987_ (.A0(net803),
    .A1(\cpu.icache.r_data[3][6] ),
    .S(_06367_),
    .X(_02111_));
 sg13g2_mux2_1 _24988_ (.A0(net802),
    .A1(\cpu.icache.r_data[3][7] ),
    .S(_06367_),
    .X(_02112_));
 sg13g2_mux2_1 _24989_ (.A0(\cpu.icache.r_data[3][8] ),
    .A1(_06344_),
    .S(_06355_),
    .X(_02113_));
 sg13g2_mux2_1 _24990_ (.A0(\cpu.icache.r_data[3][9] ),
    .A1(net933),
    .S(_06355_),
    .X(_02114_));
 sg13g2_nand2_2 _24991_ (.Y(_06368_),
    .A(net610),
    .B(_06274_));
 sg13g2_mux2_1 _24992_ (.A0(net931),
    .A1(\cpu.icache.r_data[4][0] ),
    .S(_06368_),
    .X(_02115_));
 sg13g2_and2_1 _24993_ (.A(net610),
    .B(_06281_),
    .X(_06369_));
 sg13g2_buf_1 _24994_ (.A(_06369_),
    .X(_06370_));
 sg13g2_mux2_1 _24995_ (.A0(\cpu.icache.r_data[4][10] ),
    .A1(net932),
    .S(_06370_),
    .X(_02116_));
 sg13g2_mux2_1 _24996_ (.A0(\cpu.icache.r_data[4][11] ),
    .A1(_06348_),
    .S(_06370_),
    .X(_02117_));
 sg13g2_nand2_2 _24997_ (.Y(_06371_),
    .A(_08888_),
    .B(_06287_));
 sg13g2_mux2_1 _24998_ (.A0(net931),
    .A1(\cpu.icache.r_data[4][12] ),
    .S(_06371_),
    .X(_02118_));
 sg13g2_mux2_1 _24999_ (.A0(net930),
    .A1(\cpu.icache.r_data[4][13] ),
    .S(_06371_),
    .X(_02119_));
 sg13g2_mux2_1 _25000_ (.A0(net803),
    .A1(\cpu.icache.r_data[4][14] ),
    .S(_06371_),
    .X(_02120_));
 sg13g2_mux2_1 _25001_ (.A0(net802),
    .A1(\cpu.icache.r_data[4][15] ),
    .S(_06371_),
    .X(_02121_));
 sg13g2_nand2_2 _25002_ (.Y(_06372_),
    .A(_08888_),
    .B(_06293_));
 sg13g2_mux2_1 _25003_ (.A0(_06357_),
    .A1(\cpu.icache.r_data[4][16] ),
    .S(_06372_),
    .X(_02122_));
 sg13g2_mux2_1 _25004_ (.A0(_06359_),
    .A1(\cpu.icache.r_data[4][17] ),
    .S(_06372_),
    .X(_02123_));
 sg13g2_mux2_1 _25005_ (.A0(net803),
    .A1(\cpu.icache.r_data[4][18] ),
    .S(_06372_),
    .X(_02124_));
 sg13g2_mux2_1 _25006_ (.A0(_06362_),
    .A1(\cpu.icache.r_data[4][19] ),
    .S(_06372_),
    .X(_02125_));
 sg13g2_mux2_1 _25007_ (.A0(_06359_),
    .A1(\cpu.icache.r_data[4][1] ),
    .S(_06368_),
    .X(_02126_));
 sg13g2_nand2_2 _25008_ (.Y(_06373_),
    .A(net610),
    .B(_06297_));
 sg13g2_mux2_1 _25009_ (.A0(net931),
    .A1(\cpu.icache.r_data[4][20] ),
    .S(_06373_),
    .X(_02127_));
 sg13g2_mux2_1 _25010_ (.A0(net930),
    .A1(\cpu.icache.r_data[4][21] ),
    .S(_06373_),
    .X(_02128_));
 sg13g2_mux2_1 _25011_ (.A0(net803),
    .A1(\cpu.icache.r_data[4][22] ),
    .S(_06373_),
    .X(_02129_));
 sg13g2_mux2_1 _25012_ (.A0(net802),
    .A1(\cpu.icache.r_data[4][23] ),
    .S(_06373_),
    .X(_02130_));
 sg13g2_and2_1 _25013_ (.A(net610),
    .B(_06301_),
    .X(_06374_));
 sg13g2_buf_2 _25014_ (.A(_06374_),
    .X(_06375_));
 sg13g2_mux2_1 _25015_ (.A0(\cpu.icache.r_data[4][24] ),
    .A1(net934),
    .S(_06375_),
    .X(_02131_));
 sg13g2_mux2_1 _25016_ (.A0(\cpu.icache.r_data[4][25] ),
    .A1(net933),
    .S(_06375_),
    .X(_02132_));
 sg13g2_mux2_1 _25017_ (.A0(\cpu.icache.r_data[4][26] ),
    .A1(net932),
    .S(_06375_),
    .X(_02133_));
 sg13g2_mux2_1 _25018_ (.A0(\cpu.icache.r_data[4][27] ),
    .A1(net804),
    .S(_06375_),
    .X(_02134_));
 sg13g2_nand2_2 _25019_ (.Y(_06376_),
    .A(net610),
    .B(_06306_));
 sg13g2_mux2_1 _25020_ (.A0(net931),
    .A1(\cpu.icache.r_data[4][28] ),
    .S(_06376_),
    .X(_02135_));
 sg13g2_mux2_1 _25021_ (.A0(net930),
    .A1(\cpu.icache.r_data[4][29] ),
    .S(_06376_),
    .X(_02136_));
 sg13g2_mux2_1 _25022_ (.A0(_06361_),
    .A1(\cpu.icache.r_data[4][2] ),
    .S(_06368_),
    .X(_02137_));
 sg13g2_mux2_1 _25023_ (.A0(net803),
    .A1(\cpu.icache.r_data[4][30] ),
    .S(_06376_),
    .X(_02138_));
 sg13g2_mux2_1 _25024_ (.A0(net802),
    .A1(\cpu.icache.r_data[4][31] ),
    .S(_06376_),
    .X(_02139_));
 sg13g2_mux2_1 _25025_ (.A0(net802),
    .A1(\cpu.icache.r_data[4][3] ),
    .S(_06368_),
    .X(_02140_));
 sg13g2_nand2_2 _25026_ (.Y(_06377_),
    .A(net610),
    .B(_06309_));
 sg13g2_mux2_1 _25027_ (.A0(net938),
    .A1(\cpu.icache.r_data[4][4] ),
    .S(_06377_),
    .X(_02141_));
 sg13g2_mux2_1 _25028_ (.A0(net936),
    .A1(\cpu.icache.r_data[4][5] ),
    .S(_06377_),
    .X(_02142_));
 sg13g2_mux2_1 _25029_ (.A0(net808),
    .A1(\cpu.icache.r_data[4][6] ),
    .S(_06377_),
    .X(_02143_));
 sg13g2_mux2_1 _25030_ (.A0(net807),
    .A1(\cpu.icache.r_data[4][7] ),
    .S(_06377_),
    .X(_02144_));
 sg13g2_mux2_1 _25031_ (.A0(\cpu.icache.r_data[4][8] ),
    .A1(_06344_),
    .S(_06370_),
    .X(_02145_));
 sg13g2_mux2_1 _25032_ (.A0(\cpu.icache.r_data[4][9] ),
    .A1(_06346_),
    .S(_06370_),
    .X(_02146_));
 sg13g2_nand2_1 _25033_ (.Y(_06378_),
    .A(net1050),
    .B(_08752_));
 sg13g2_buf_4 _25034_ (.X(_06379_),
    .A(_06378_));
 sg13g2_nor2_2 _25035_ (.A(_06379_),
    .B(_06314_),
    .Y(_06380_));
 sg13g2_mux2_1 _25036_ (.A0(\cpu.icache.r_data[5][0] ),
    .A1(net934),
    .S(_06380_),
    .X(_02147_));
 sg13g2_nor2_2 _25037_ (.A(_06379_),
    .B(_06280_),
    .Y(_06381_));
 sg13g2_mux2_1 _25038_ (.A0(\cpu.icache.r_data[5][10] ),
    .A1(_06347_),
    .S(_06381_),
    .X(_02148_));
 sg13g2_mux2_1 _25039_ (.A0(\cpu.icache.r_data[5][11] ),
    .A1(_06348_),
    .S(_06381_),
    .X(_02149_));
 sg13g2_nor2_2 _25040_ (.A(_06379_),
    .B(_06320_),
    .Y(_06382_));
 sg13g2_mux2_1 _25041_ (.A0(\cpu.icache.r_data[5][12] ),
    .A1(net934),
    .S(_06382_),
    .X(_02150_));
 sg13g2_mux2_1 _25042_ (.A0(\cpu.icache.r_data[5][13] ),
    .A1(net933),
    .S(_06382_),
    .X(_02151_));
 sg13g2_mux2_1 _25043_ (.A0(\cpu.icache.r_data[5][14] ),
    .A1(net932),
    .S(_06382_),
    .X(_02152_));
 sg13g2_mux2_1 _25044_ (.A0(\cpu.icache.r_data[5][15] ),
    .A1(net804),
    .S(_06382_),
    .X(_02153_));
 sg13g2_buf_1 _25045_ (.A(_12143_),
    .X(_06383_));
 sg13g2_nor2_2 _25046_ (.A(_06379_),
    .B(_06325_),
    .Y(_06384_));
 sg13g2_mux2_1 _25047_ (.A0(\cpu.icache.r_data[5][16] ),
    .A1(net929),
    .S(_06384_),
    .X(_02154_));
 sg13g2_mux2_1 _25048_ (.A0(\cpu.icache.r_data[5][17] ),
    .A1(_06346_),
    .S(_06384_),
    .X(_02155_));
 sg13g2_buf_1 _25049_ (.A(_12107_),
    .X(_06385_));
 sg13g2_mux2_1 _25050_ (.A0(\cpu.icache.r_data[5][18] ),
    .A1(net928),
    .S(_06384_),
    .X(_02156_));
 sg13g2_buf_2 _25051_ (.A(_12113_),
    .X(_06386_));
 sg13g2_mux2_1 _25052_ (.A0(\cpu.icache.r_data[5][19] ),
    .A1(_06386_),
    .S(_06384_),
    .X(_02157_));
 sg13g2_buf_1 _25053_ (.A(_03029_),
    .X(_06387_));
 sg13g2_mux2_1 _25054_ (.A0(\cpu.icache.r_data[5][1] ),
    .A1(_06387_),
    .S(_06380_),
    .X(_02158_));
 sg13g2_nor2_2 _25055_ (.A(_06379_),
    .B(_06328_),
    .Y(_06388_));
 sg13g2_mux2_1 _25056_ (.A0(\cpu.icache.r_data[5][20] ),
    .A1(net929),
    .S(_06388_),
    .X(_02159_));
 sg13g2_mux2_1 _25057_ (.A0(\cpu.icache.r_data[5][21] ),
    .A1(net926),
    .S(_06388_),
    .X(_02160_));
 sg13g2_mux2_1 _25058_ (.A0(\cpu.icache.r_data[5][22] ),
    .A1(net928),
    .S(_06388_),
    .X(_02161_));
 sg13g2_mux2_1 _25059_ (.A0(\cpu.icache.r_data[5][23] ),
    .A1(net927),
    .S(_06388_),
    .X(_02162_));
 sg13g2_nor2_1 _25060_ (.A(_06379_),
    .B(_06331_),
    .Y(_06389_));
 sg13g2_buf_2 _25061_ (.A(_06389_),
    .X(_06390_));
 sg13g2_mux2_1 _25062_ (.A0(\cpu.icache.r_data[5][24] ),
    .A1(net929),
    .S(_06390_),
    .X(_02163_));
 sg13g2_mux2_1 _25063_ (.A0(\cpu.icache.r_data[5][25] ),
    .A1(net926),
    .S(_06390_),
    .X(_02164_));
 sg13g2_mux2_1 _25064_ (.A0(\cpu.icache.r_data[5][26] ),
    .A1(net928),
    .S(_06390_),
    .X(_02165_));
 sg13g2_mux2_1 _25065_ (.A0(\cpu.icache.r_data[5][27] ),
    .A1(net927),
    .S(_06390_),
    .X(_02166_));
 sg13g2_nor2_2 _25066_ (.A(_06379_),
    .B(_06334_),
    .Y(_06391_));
 sg13g2_mux2_1 _25067_ (.A0(\cpu.icache.r_data[5][28] ),
    .A1(net929),
    .S(_06391_),
    .X(_02167_));
 sg13g2_mux2_1 _25068_ (.A0(\cpu.icache.r_data[5][29] ),
    .A1(net926),
    .S(_06391_),
    .X(_02168_));
 sg13g2_mux2_1 _25069_ (.A0(\cpu.icache.r_data[5][2] ),
    .A1(_06385_),
    .S(_06380_),
    .X(_02169_));
 sg13g2_mux2_1 _25070_ (.A0(\cpu.icache.r_data[5][30] ),
    .A1(net928),
    .S(_06391_),
    .X(_02170_));
 sg13g2_mux2_1 _25071_ (.A0(\cpu.icache.r_data[5][31] ),
    .A1(net927),
    .S(_06391_),
    .X(_02171_));
 sg13g2_mux2_1 _25072_ (.A0(\cpu.icache.r_data[5][3] ),
    .A1(net927),
    .S(_06380_),
    .X(_02172_));
 sg13g2_nor2_2 _25073_ (.A(_06379_),
    .B(_06336_),
    .Y(_06392_));
 sg13g2_mux2_1 _25074_ (.A0(\cpu.icache.r_data[5][4] ),
    .A1(net929),
    .S(_06392_),
    .X(_02173_));
 sg13g2_mux2_1 _25075_ (.A0(\cpu.icache.r_data[5][5] ),
    .A1(net926),
    .S(_06392_),
    .X(_02174_));
 sg13g2_mux2_1 _25076_ (.A0(\cpu.icache.r_data[5][6] ),
    .A1(net928),
    .S(_06392_),
    .X(_02175_));
 sg13g2_mux2_1 _25077_ (.A0(\cpu.icache.r_data[5][7] ),
    .A1(net927),
    .S(_06392_),
    .X(_02176_));
 sg13g2_mux2_1 _25078_ (.A0(\cpu.icache.r_data[5][8] ),
    .A1(net929),
    .S(_06381_),
    .X(_02177_));
 sg13g2_mux2_1 _25079_ (.A0(\cpu.icache.r_data[5][9] ),
    .A1(net926),
    .S(_06381_),
    .X(_02178_));
 sg13g2_nand2_2 _25080_ (.Y(_06393_),
    .A(net466),
    .B(_06274_));
 sg13g2_mux2_1 _25081_ (.A0(_06311_),
    .A1(\cpu.icache.r_data[6][0] ),
    .S(_06393_),
    .X(_02179_));
 sg13g2_nand2_2 _25082_ (.Y(_06394_),
    .A(net466),
    .B(_06281_));
 sg13g2_mux2_1 _25083_ (.A0(net808),
    .A1(\cpu.icache.r_data[6][10] ),
    .S(_06394_),
    .X(_02180_));
 sg13g2_mux2_1 _25084_ (.A0(net807),
    .A1(\cpu.icache.r_data[6][11] ),
    .S(_06394_),
    .X(_02181_));
 sg13g2_nand2_2 _25085_ (.Y(_06395_),
    .A(_08770_),
    .B(_06287_));
 sg13g2_mux2_1 _25086_ (.A0(net938),
    .A1(\cpu.icache.r_data[6][12] ),
    .S(_06395_),
    .X(_02182_));
 sg13g2_mux2_1 _25087_ (.A0(net936),
    .A1(\cpu.icache.r_data[6][13] ),
    .S(_06395_),
    .X(_02183_));
 sg13g2_mux2_1 _25088_ (.A0(net808),
    .A1(\cpu.icache.r_data[6][14] ),
    .S(_06395_),
    .X(_02184_));
 sg13g2_mux2_1 _25089_ (.A0(net807),
    .A1(\cpu.icache.r_data[6][15] ),
    .S(_06395_),
    .X(_02185_));
 sg13g2_nand2_2 _25090_ (.Y(_06396_),
    .A(_08770_),
    .B(_06293_));
 sg13g2_mux2_1 _25091_ (.A0(net938),
    .A1(\cpu.icache.r_data[6][16] ),
    .S(_06396_),
    .X(_02186_));
 sg13g2_mux2_1 _25092_ (.A0(net936),
    .A1(\cpu.icache.r_data[6][17] ),
    .S(_06396_),
    .X(_02187_));
 sg13g2_mux2_1 _25093_ (.A0(_06316_),
    .A1(\cpu.icache.r_data[6][18] ),
    .S(_06396_),
    .X(_02188_));
 sg13g2_mux2_1 _25094_ (.A0(_06318_),
    .A1(\cpu.icache.r_data[6][19] ),
    .S(_06396_),
    .X(_02189_));
 sg13g2_mux2_1 _25095_ (.A0(_06322_),
    .A1(\cpu.icache.r_data[6][1] ),
    .S(_06393_),
    .X(_02190_));
 sg13g2_nand2_2 _25096_ (.Y(_06397_),
    .A(net466),
    .B(_06297_));
 sg13g2_mux2_1 _25097_ (.A0(net938),
    .A1(\cpu.icache.r_data[6][20] ),
    .S(_06397_),
    .X(_02191_));
 sg13g2_mux2_1 _25098_ (.A0(net936),
    .A1(\cpu.icache.r_data[6][21] ),
    .S(_06397_),
    .X(_02192_));
 sg13g2_mux2_1 _25099_ (.A0(net808),
    .A1(\cpu.icache.r_data[6][22] ),
    .S(_06397_),
    .X(_02193_));
 sg13g2_mux2_1 _25100_ (.A0(net807),
    .A1(\cpu.icache.r_data[6][23] ),
    .S(_06397_),
    .X(_02194_));
 sg13g2_nand2_1 _25101_ (.Y(_06398_),
    .A(net466),
    .B(_06301_));
 sg13g2_buf_2 _25102_ (.A(_06398_),
    .X(_06399_));
 sg13g2_mux2_1 _25103_ (.A0(_06311_),
    .A1(\cpu.icache.r_data[6][24] ),
    .S(_06399_),
    .X(_02195_));
 sg13g2_mux2_1 _25104_ (.A0(net936),
    .A1(\cpu.icache.r_data[6][25] ),
    .S(_06399_),
    .X(_02196_));
 sg13g2_mux2_1 _25105_ (.A0(net808),
    .A1(\cpu.icache.r_data[6][26] ),
    .S(_06399_),
    .X(_02197_));
 sg13g2_mux2_1 _25106_ (.A0(net807),
    .A1(\cpu.icache.r_data[6][27] ),
    .S(_06399_),
    .X(_02198_));
 sg13g2_nand2_2 _25107_ (.Y(_06400_),
    .A(net466),
    .B(_06306_));
 sg13g2_mux2_1 _25108_ (.A0(net938),
    .A1(\cpu.icache.r_data[6][28] ),
    .S(_06400_),
    .X(_02199_));
 sg13g2_mux2_1 _25109_ (.A0(net936),
    .A1(\cpu.icache.r_data[6][29] ),
    .S(_06400_),
    .X(_02200_));
 sg13g2_mux2_1 _25110_ (.A0(_06316_),
    .A1(\cpu.icache.r_data[6][2] ),
    .S(_06393_),
    .X(_02201_));
 sg13g2_mux2_1 _25111_ (.A0(net808),
    .A1(\cpu.icache.r_data[6][30] ),
    .S(_06400_),
    .X(_02202_));
 sg13g2_mux2_1 _25112_ (.A0(net807),
    .A1(\cpu.icache.r_data[6][31] ),
    .S(_06400_),
    .X(_02203_));
 sg13g2_mux2_1 _25113_ (.A0(net807),
    .A1(\cpu.icache.r_data[6][3] ),
    .S(_06393_),
    .X(_02204_));
 sg13g2_nand2_2 _25114_ (.Y(_06401_),
    .A(net466),
    .B(_06309_));
 sg13g2_mux2_1 _25115_ (.A0(net938),
    .A1(\cpu.icache.r_data[6][4] ),
    .S(_06401_),
    .X(_02205_));
 sg13g2_mux2_1 _25116_ (.A0(net936),
    .A1(\cpu.icache.r_data[6][5] ),
    .S(_06401_),
    .X(_02206_));
 sg13g2_mux2_1 _25117_ (.A0(net808),
    .A1(\cpu.icache.r_data[6][6] ),
    .S(_06401_),
    .X(_02207_));
 sg13g2_mux2_1 _25118_ (.A0(net807),
    .A1(\cpu.icache.r_data[6][7] ),
    .S(_06401_),
    .X(_02208_));
 sg13g2_mux2_1 _25119_ (.A0(net938),
    .A1(\cpu.icache.r_data[6][8] ),
    .S(_06394_),
    .X(_02209_));
 sg13g2_mux2_1 _25120_ (.A0(_06322_),
    .A1(\cpu.icache.r_data[6][9] ),
    .S(_06394_),
    .X(_02210_));
 sg13g2_nand2_1 _25121_ (.Y(_06402_),
    .A(net1050),
    .B(_08424_));
 sg13g2_buf_4 _25122_ (.X(_06403_),
    .A(_06402_));
 sg13g2_nor2_2 _25123_ (.A(_06403_),
    .B(_06314_),
    .Y(_06404_));
 sg13g2_mux2_1 _25124_ (.A0(\cpu.icache.r_data[7][0] ),
    .A1(_06383_),
    .S(_06404_),
    .X(_02211_));
 sg13g2_nor2_2 _25125_ (.A(_06403_),
    .B(_06280_),
    .Y(_06405_));
 sg13g2_mux2_1 _25126_ (.A0(\cpu.icache.r_data[7][10] ),
    .A1(net928),
    .S(_06405_),
    .X(_02212_));
 sg13g2_mux2_1 _25127_ (.A0(\cpu.icache.r_data[7][11] ),
    .A1(net927),
    .S(_06405_),
    .X(_02213_));
 sg13g2_nor2_2 _25128_ (.A(_06403_),
    .B(_06320_),
    .Y(_06406_));
 sg13g2_mux2_1 _25129_ (.A0(\cpu.icache.r_data[7][12] ),
    .A1(net929),
    .S(_06406_),
    .X(_02214_));
 sg13g2_mux2_1 _25130_ (.A0(\cpu.icache.r_data[7][13] ),
    .A1(net926),
    .S(_06406_),
    .X(_02215_));
 sg13g2_mux2_1 _25131_ (.A0(\cpu.icache.r_data[7][14] ),
    .A1(net928),
    .S(_06406_),
    .X(_02216_));
 sg13g2_mux2_1 _25132_ (.A0(\cpu.icache.r_data[7][15] ),
    .A1(net927),
    .S(_06406_),
    .X(_02217_));
 sg13g2_nor2_2 _25133_ (.A(_06403_),
    .B(_06325_),
    .Y(_06407_));
 sg13g2_mux2_1 _25134_ (.A0(\cpu.icache.r_data[7][16] ),
    .A1(_06383_),
    .S(_06407_),
    .X(_02218_));
 sg13g2_mux2_1 _25135_ (.A0(\cpu.icache.r_data[7][17] ),
    .A1(net926),
    .S(_06407_),
    .X(_02219_));
 sg13g2_mux2_1 _25136_ (.A0(\cpu.icache.r_data[7][18] ),
    .A1(_06385_),
    .S(_06407_),
    .X(_02220_));
 sg13g2_mux2_1 _25137_ (.A0(\cpu.icache.r_data[7][19] ),
    .A1(_06386_),
    .S(_06407_),
    .X(_02221_));
 sg13g2_mux2_1 _25138_ (.A0(\cpu.icache.r_data[7][1] ),
    .A1(_06387_),
    .S(_06404_),
    .X(_02222_));
 sg13g2_nor2_2 _25139_ (.A(_06403_),
    .B(_06328_),
    .Y(_06408_));
 sg13g2_mux2_1 _25140_ (.A0(\cpu.icache.r_data[7][20] ),
    .A1(net929),
    .S(_06408_),
    .X(_02223_));
 sg13g2_mux2_1 _25141_ (.A0(\cpu.icache.r_data[7][21] ),
    .A1(net926),
    .S(_06408_),
    .X(_02224_));
 sg13g2_mux2_1 _25142_ (.A0(\cpu.icache.r_data[7][22] ),
    .A1(net928),
    .S(_06408_),
    .X(_02225_));
 sg13g2_mux2_1 _25143_ (.A0(\cpu.icache.r_data[7][23] ),
    .A1(net927),
    .S(_06408_),
    .X(_02226_));
 sg13g2_nor2_1 _25144_ (.A(_06403_),
    .B(_06331_),
    .Y(_06409_));
 sg13g2_buf_2 _25145_ (.A(_06409_),
    .X(_06410_));
 sg13g2_mux2_1 _25146_ (.A0(\cpu.icache.r_data[7][24] ),
    .A1(net992),
    .S(_06410_),
    .X(_02227_));
 sg13g2_mux2_1 _25147_ (.A0(\cpu.icache.r_data[7][25] ),
    .A1(net988),
    .S(_06410_),
    .X(_02228_));
 sg13g2_mux2_1 _25148_ (.A0(\cpu.icache.r_data[7][26] ),
    .A1(net990),
    .S(_06410_),
    .X(_02229_));
 sg13g2_mux2_1 _25149_ (.A0(\cpu.icache.r_data[7][27] ),
    .A1(net989),
    .S(_06410_),
    .X(_02230_));
 sg13g2_nor2_2 _25150_ (.A(_06403_),
    .B(_06334_),
    .Y(_06411_));
 sg13g2_mux2_1 _25151_ (.A0(\cpu.icache.r_data[7][28] ),
    .A1(net992),
    .S(_06411_),
    .X(_02231_));
 sg13g2_mux2_1 _25152_ (.A0(\cpu.icache.r_data[7][29] ),
    .A1(net988),
    .S(_06411_),
    .X(_02232_));
 sg13g2_mux2_1 _25153_ (.A0(\cpu.icache.r_data[7][2] ),
    .A1(net990),
    .S(_06404_),
    .X(_02233_));
 sg13g2_mux2_1 _25154_ (.A0(\cpu.icache.r_data[7][30] ),
    .A1(_12031_),
    .S(_06411_),
    .X(_02234_));
 sg13g2_mux2_1 _25155_ (.A0(\cpu.icache.r_data[7][31] ),
    .A1(net989),
    .S(_06411_),
    .X(_02235_));
 sg13g2_mux2_1 _25156_ (.A0(\cpu.icache.r_data[7][3] ),
    .A1(_12047_),
    .S(_06404_),
    .X(_02236_));
 sg13g2_nor2_2 _25157_ (.A(_06403_),
    .B(_06336_),
    .Y(_06412_));
 sg13g2_mux2_1 _25158_ (.A0(\cpu.icache.r_data[7][4] ),
    .A1(_12007_),
    .S(_06412_),
    .X(_02237_));
 sg13g2_mux2_1 _25159_ (.A0(\cpu.icache.r_data[7][5] ),
    .A1(_12067_),
    .S(_06412_),
    .X(_02238_));
 sg13g2_mux2_1 _25160_ (.A0(\cpu.icache.r_data[7][6] ),
    .A1(_12031_),
    .S(_06412_),
    .X(_02239_));
 sg13g2_mux2_1 _25161_ (.A0(\cpu.icache.r_data[7][7] ),
    .A1(_12047_),
    .S(_06412_),
    .X(_02240_));
 sg13g2_mux2_1 _25162_ (.A0(\cpu.icache.r_data[7][8] ),
    .A1(_12007_),
    .S(_06405_),
    .X(_02241_));
 sg13g2_mux2_1 _25163_ (.A0(\cpu.icache.r_data[7][9] ),
    .A1(_12067_),
    .S(_06405_),
    .X(_02242_));
 sg13g2_mux2_1 _25164_ (.A0(net957),
    .A1(\cpu.icache.r_tag[0][5] ),
    .S(net310),
    .X(_02246_));
 sg13g2_buf_1 _25165_ (.A(net398),
    .X(_06413_));
 sg13g2_buf_1 _25166_ (.A(_06302_),
    .X(_06414_));
 sg13g2_nand2_1 _25167_ (.Y(_06415_),
    .A(\cpu.icache.r_tag[0][15] ),
    .B(_06414_));
 sg13g2_o21ai_1 _25168_ (.B1(_06415_),
    .Y(_02247_),
    .A1(net380),
    .A2(net309));
 sg13g2_nand2_1 _25169_ (.Y(_06416_),
    .A(\cpu.icache.r_tag[0][16] ),
    .B(net397));
 sg13g2_o21ai_1 _25170_ (.B1(_06416_),
    .Y(_02248_),
    .A1(net383),
    .A2(net309));
 sg13g2_nand2_1 _25171_ (.Y(_06417_),
    .A(\cpu.icache.r_tag[0][17] ),
    .B(net397));
 sg13g2_o21ai_1 _25172_ (.B1(_06417_),
    .Y(_02249_),
    .A1(net437),
    .A2(net309));
 sg13g2_nand2_1 _25173_ (.Y(_06418_),
    .A(\cpu.icache.r_tag[0][18] ),
    .B(net397));
 sg13g2_o21ai_1 _25174_ (.B1(_06418_),
    .Y(_02250_),
    .A1(net436),
    .A2(net309));
 sg13g2_nand2_1 _25175_ (.Y(_06419_),
    .A(\cpu.icache.r_tag[0][19] ),
    .B(_06414_));
 sg13g2_o21ai_1 _25176_ (.B1(_06419_),
    .Y(_02251_),
    .A1(_08494_),
    .A2(_06413_));
 sg13g2_nand2_1 _25177_ (.Y(_06420_),
    .A(\cpu.icache.r_tag[0][20] ),
    .B(net397));
 sg13g2_o21ai_1 _25178_ (.B1(_06420_),
    .Y(_02252_),
    .A1(_08400_),
    .A2(net309));
 sg13g2_nand2_1 _25179_ (.Y(_06421_),
    .A(\cpu.icache.r_tag[0][21] ),
    .B(_06303_));
 sg13g2_o21ai_1 _25180_ (.B1(_06421_),
    .Y(_02253_),
    .A1(_08422_),
    .A2(_06413_));
 sg13g2_nand2_1 _25181_ (.Y(_06422_),
    .A(\cpu.icache.r_tag[0][22] ),
    .B(net398));
 sg13g2_o21ai_1 _25182_ (.B1(_06422_),
    .Y(_02254_),
    .A1(_08601_),
    .A2(net309));
 sg13g2_nand2_1 _25183_ (.Y(_06423_),
    .A(\cpu.icache.r_tag[0][23] ),
    .B(net398));
 sg13g2_o21ai_1 _25184_ (.B1(_06423_),
    .Y(_02255_),
    .A1(_08535_),
    .A2(net309));
 sg13g2_nand2_1 _25185_ (.Y(_06424_),
    .A(\cpu.icache.r_tag[0][6] ),
    .B(net398));
 sg13g2_o21ai_1 _25186_ (.B1(_06424_),
    .Y(_02256_),
    .A1(net1047),
    .A2(net310));
 sg13g2_mux2_1 _25187_ (.A0(net956),
    .A1(\cpu.icache.r_tag[0][7] ),
    .S(net397),
    .X(_02257_));
 sg13g2_mux2_1 _25188_ (.A0(net955),
    .A1(\cpu.icache.r_tag[0][8] ),
    .S(net397),
    .X(_02258_));
 sg13g2_nand2_1 _25189_ (.Y(_06425_),
    .A(\cpu.icache.r_tag[0][9] ),
    .B(net398));
 sg13g2_o21ai_1 _25190_ (.B1(_06425_),
    .Y(_02259_),
    .A1(net958),
    .A2(net310));
 sg13g2_mux2_1 _25191_ (.A0(net954),
    .A1(\cpu.icache.r_tag[0][10] ),
    .S(net397),
    .X(_02260_));
 sg13g2_mux2_1 _25192_ (.A0(net959),
    .A1(\cpu.icache.r_tag[0][11] ),
    .S(net397),
    .X(_02261_));
 sg13g2_nand2_1 _25193_ (.Y(_06426_),
    .A(\cpu.icache.r_tag[0][12] ),
    .B(net398));
 sg13g2_o21ai_1 _25194_ (.B1(_06426_),
    .Y(_02262_),
    .A1(_08285_),
    .A2(net310));
 sg13g2_nand2_1 _25195_ (.Y(_06427_),
    .A(\cpu.icache.r_tag[0][13] ),
    .B(net398));
 sg13g2_o21ai_1 _25196_ (.B1(_06427_),
    .Y(_02263_),
    .A1(net386),
    .A2(net310));
 sg13g2_nand2_1 _25197_ (.Y(_06428_),
    .A(\cpu.icache.r_tag[0][14] ),
    .B(_06303_));
 sg13g2_o21ai_1 _25198_ (.B1(_06428_),
    .Y(_02264_),
    .A1(net382),
    .A2(net310));
 sg13g2_nor2b_1 _25199_ (.A(_06300_),
    .B_N(_06291_),
    .Y(_06429_));
 sg13g2_buf_1 _25200_ (.A(_06429_),
    .X(_06430_));
 sg13g2_nand2_1 _25201_ (.Y(_06431_),
    .A(net535),
    .B(_06430_));
 sg13g2_buf_1 _25202_ (.A(_06431_),
    .X(_06432_));
 sg13g2_buf_1 _25203_ (.A(_06432_),
    .X(_06433_));
 sg13g2_mux2_1 _25204_ (.A0(net957),
    .A1(\cpu.icache.r_tag[1][5] ),
    .S(_06433_),
    .X(_02265_));
 sg13g2_buf_1 _25205_ (.A(_06432_),
    .X(_06434_));
 sg13g2_nand2_1 _25206_ (.Y(_06435_),
    .A(\cpu.icache.r_tag[1][15] ),
    .B(net308));
 sg13g2_o21ai_1 _25207_ (.B1(_06435_),
    .Y(_02266_),
    .A1(net380),
    .A2(net307));
 sg13g2_buf_1 _25208_ (.A(_06432_),
    .X(_06436_));
 sg13g2_nand2_1 _25209_ (.Y(_06437_),
    .A(\cpu.icache.r_tag[1][16] ),
    .B(_06436_));
 sg13g2_o21ai_1 _25210_ (.B1(_06437_),
    .Y(_02267_),
    .A1(net383),
    .A2(net307));
 sg13g2_nand2_1 _25211_ (.Y(_06438_),
    .A(\cpu.icache.r_tag[1][17] ),
    .B(net306));
 sg13g2_o21ai_1 _25212_ (.B1(_06438_),
    .Y(_02268_),
    .A1(net437),
    .A2(_06434_));
 sg13g2_nand2_1 _25213_ (.Y(_06439_),
    .A(\cpu.icache.r_tag[1][18] ),
    .B(net306));
 sg13g2_o21ai_1 _25214_ (.B1(_06439_),
    .Y(_02269_),
    .A1(net436),
    .A2(net307));
 sg13g2_nand2_1 _25215_ (.Y(_06440_),
    .A(\cpu.icache.r_tag[1][19] ),
    .B(net306));
 sg13g2_o21ai_1 _25216_ (.B1(_06440_),
    .Y(_02270_),
    .A1(net381),
    .A2(net307));
 sg13g2_nand2_1 _25217_ (.Y(_06441_),
    .A(\cpu.icache.r_tag[1][20] ),
    .B(net306));
 sg13g2_o21ai_1 _25218_ (.B1(_06441_),
    .Y(_02271_),
    .A1(net385),
    .A2(net307));
 sg13g2_nand2_1 _25219_ (.Y(_06442_),
    .A(\cpu.icache.r_tag[1][21] ),
    .B(_06436_));
 sg13g2_o21ai_1 _25220_ (.B1(_06442_),
    .Y(_02272_),
    .A1(net384),
    .A2(net307));
 sg13g2_nand2_1 _25221_ (.Y(_06443_),
    .A(\cpu.icache.r_tag[1][22] ),
    .B(net306));
 sg13g2_o21ai_1 _25222_ (.B1(_06443_),
    .Y(_02273_),
    .A1(net435),
    .A2(net307));
 sg13g2_nand2_1 _25223_ (.Y(_06444_),
    .A(\cpu.icache.r_tag[1][23] ),
    .B(net306));
 sg13g2_o21ai_1 _25224_ (.B1(_06444_),
    .Y(_02274_),
    .A1(net469),
    .A2(net307));
 sg13g2_nand2_1 _25225_ (.Y(_06445_),
    .A(\cpu.icache.r_tag[1][6] ),
    .B(net306));
 sg13g2_o21ai_1 _25226_ (.B1(_06445_),
    .Y(_02275_),
    .A1(net1047),
    .A2(_06434_));
 sg13g2_mux2_1 _25227_ (.A0(net956),
    .A1(\cpu.icache.r_tag[1][7] ),
    .S(net308),
    .X(_02276_));
 sg13g2_mux2_1 _25228_ (.A0(net955),
    .A1(\cpu.icache.r_tag[1][8] ),
    .S(net308),
    .X(_02277_));
 sg13g2_nand2_1 _25229_ (.Y(_06446_),
    .A(\cpu.icache.r_tag[1][9] ),
    .B(net306));
 sg13g2_o21ai_1 _25230_ (.B1(_06446_),
    .Y(_02278_),
    .A1(net958),
    .A2(_06433_));
 sg13g2_mux2_1 _25231_ (.A0(net954),
    .A1(\cpu.icache.r_tag[1][10] ),
    .S(net308),
    .X(_02279_));
 sg13g2_mux2_1 _25232_ (.A0(net959),
    .A1(\cpu.icache.r_tag[1][11] ),
    .S(net308),
    .X(_02280_));
 sg13g2_nand2_1 _25233_ (.Y(_06447_),
    .A(\cpu.icache.r_tag[1][12] ),
    .B(_06432_));
 sg13g2_o21ai_1 _25234_ (.B1(_06447_),
    .Y(_02281_),
    .A1(net438),
    .A2(net308));
 sg13g2_nand2_1 _25235_ (.Y(_06448_),
    .A(\cpu.icache.r_tag[1][13] ),
    .B(_06432_));
 sg13g2_o21ai_1 _25236_ (.B1(_06448_),
    .Y(_02282_),
    .A1(net386),
    .A2(net308));
 sg13g2_nand2_1 _25237_ (.Y(_06449_),
    .A(\cpu.icache.r_tag[1][14] ),
    .B(_06432_));
 sg13g2_o21ai_1 _25238_ (.B1(_06449_),
    .Y(_02283_),
    .A1(net382),
    .A2(net308));
 sg13g2_nand2_1 _25239_ (.Y(_06450_),
    .A(net468),
    .B(_06430_));
 sg13g2_buf_1 _25240_ (.A(_06450_),
    .X(_06451_));
 sg13g2_buf_1 _25241_ (.A(_06451_),
    .X(_06452_));
 sg13g2_mux2_1 _25242_ (.A0(net957),
    .A1(\cpu.icache.r_tag[2][5] ),
    .S(net261),
    .X(_02284_));
 sg13g2_buf_1 _25243_ (.A(_06451_),
    .X(_06453_));
 sg13g2_nand2_1 _25244_ (.Y(_06454_),
    .A(\cpu.icache.r_tag[2][15] ),
    .B(_06452_));
 sg13g2_o21ai_1 _25245_ (.B1(_06454_),
    .Y(_02285_),
    .A1(_08515_),
    .A2(_06453_));
 sg13g2_buf_1 _25246_ (.A(_06451_),
    .X(_06455_));
 sg13g2_nand2_1 _25247_ (.Y(_06456_),
    .A(\cpu.icache.r_tag[2][16] ),
    .B(_06455_));
 sg13g2_o21ai_1 _25248_ (.B1(_06456_),
    .Y(_02286_),
    .A1(net383),
    .A2(_06453_));
 sg13g2_nand2_1 _25249_ (.Y(_06457_),
    .A(\cpu.icache.r_tag[2][17] ),
    .B(net259));
 sg13g2_o21ai_1 _25250_ (.B1(_06457_),
    .Y(_02287_),
    .A1(net437),
    .A2(net260));
 sg13g2_nand2_1 _25251_ (.Y(_06458_),
    .A(\cpu.icache.r_tag[2][18] ),
    .B(net259));
 sg13g2_o21ai_1 _25252_ (.B1(_06458_),
    .Y(_02288_),
    .A1(_08577_),
    .A2(net260));
 sg13g2_nand2_1 _25253_ (.Y(_06459_),
    .A(\cpu.icache.r_tag[2][19] ),
    .B(_06455_));
 sg13g2_o21ai_1 _25254_ (.B1(_06459_),
    .Y(_02289_),
    .A1(net381),
    .A2(net260));
 sg13g2_nand2_1 _25255_ (.Y(_06460_),
    .A(\cpu.icache.r_tag[2][20] ),
    .B(net259));
 sg13g2_o21ai_1 _25256_ (.B1(_06460_),
    .Y(_02290_),
    .A1(net385),
    .A2(net260));
 sg13g2_nand2_1 _25257_ (.Y(_06461_),
    .A(\cpu.icache.r_tag[2][21] ),
    .B(net259));
 sg13g2_o21ai_1 _25258_ (.B1(_06461_),
    .Y(_02291_),
    .A1(net384),
    .A2(net260));
 sg13g2_nand2_1 _25259_ (.Y(_06462_),
    .A(\cpu.icache.r_tag[2][22] ),
    .B(net259));
 sg13g2_o21ai_1 _25260_ (.B1(_06462_),
    .Y(_02292_),
    .A1(net435),
    .A2(net260));
 sg13g2_nand2_1 _25261_ (.Y(_06463_),
    .A(\cpu.icache.r_tag[2][23] ),
    .B(net259));
 sg13g2_o21ai_1 _25262_ (.B1(_06463_),
    .Y(_02293_),
    .A1(net469),
    .A2(net260));
 sg13g2_nand2_1 _25263_ (.Y(_06464_),
    .A(\cpu.icache.r_tag[2][6] ),
    .B(net259));
 sg13g2_o21ai_1 _25264_ (.B1(_06464_),
    .Y(_02294_),
    .A1(net1047),
    .A2(net260));
 sg13g2_mux2_1 _25265_ (.A0(net956),
    .A1(\cpu.icache.r_tag[2][7] ),
    .S(net261),
    .X(_02295_));
 sg13g2_mux2_1 _25266_ (.A0(net955),
    .A1(\cpu.icache.r_tag[2][8] ),
    .S(net261),
    .X(_02296_));
 sg13g2_nand2_1 _25267_ (.Y(_06465_),
    .A(\cpu.icache.r_tag[2][9] ),
    .B(net259));
 sg13g2_o21ai_1 _25268_ (.B1(_06465_),
    .Y(_02297_),
    .A1(net958),
    .A2(net261));
 sg13g2_mux2_1 _25269_ (.A0(net954),
    .A1(\cpu.icache.r_tag[2][10] ),
    .S(net261),
    .X(_02298_));
 sg13g2_mux2_1 _25270_ (.A0(net959),
    .A1(\cpu.icache.r_tag[2][11] ),
    .S(net261),
    .X(_02299_));
 sg13g2_nand2_1 _25271_ (.Y(_06466_),
    .A(\cpu.icache.r_tag[2][12] ),
    .B(_06451_));
 sg13g2_o21ai_1 _25272_ (.B1(_06466_),
    .Y(_02300_),
    .A1(net438),
    .A2(net261));
 sg13g2_nand2_1 _25273_ (.Y(_06467_),
    .A(\cpu.icache.r_tag[2][13] ),
    .B(_06451_));
 sg13g2_o21ai_1 _25274_ (.B1(_06467_),
    .Y(_02301_),
    .A1(net386),
    .A2(net261));
 sg13g2_nand2_1 _25275_ (.Y(_06468_),
    .A(\cpu.icache.r_tag[2][14] ),
    .B(_06451_));
 sg13g2_o21ai_1 _25276_ (.B1(_06468_),
    .Y(_02302_),
    .A1(net382),
    .A2(_06452_));
 sg13g2_mux2_1 _25277_ (.A0(net957),
    .A1(\cpu.icache.r_tag[3][5] ),
    .S(net236),
    .X(_02303_));
 sg13g2_buf_1 _25278_ (.A(net262),
    .X(_06469_));
 sg13g2_buf_1 _25279_ (.A(_06363_),
    .X(_06470_));
 sg13g2_nand2_1 _25280_ (.Y(_06471_),
    .A(\cpu.icache.r_tag[3][15] ),
    .B(net258));
 sg13g2_o21ai_1 _25281_ (.B1(_06471_),
    .Y(_02304_),
    .A1(net380),
    .A2(_06469_));
 sg13g2_nand2_1 _25282_ (.Y(_06472_),
    .A(\cpu.icache.r_tag[3][16] ),
    .B(net258));
 sg13g2_o21ai_1 _25283_ (.B1(_06472_),
    .Y(_02305_),
    .A1(net383),
    .A2(net235));
 sg13g2_nand2_1 _25284_ (.Y(_06473_),
    .A(\cpu.icache.r_tag[3][17] ),
    .B(net258));
 sg13g2_o21ai_1 _25285_ (.B1(_06473_),
    .Y(_02306_),
    .A1(net437),
    .A2(net235));
 sg13g2_nand2_1 _25286_ (.Y(_06474_),
    .A(\cpu.icache.r_tag[3][18] ),
    .B(net258));
 sg13g2_o21ai_1 _25287_ (.B1(_06474_),
    .Y(_02307_),
    .A1(net436),
    .A2(net235));
 sg13g2_nand2_1 _25288_ (.Y(_06475_),
    .A(\cpu.icache.r_tag[3][19] ),
    .B(_06470_));
 sg13g2_o21ai_1 _25289_ (.B1(_06475_),
    .Y(_02308_),
    .A1(net381),
    .A2(net235));
 sg13g2_nand2_1 _25290_ (.Y(_06476_),
    .A(\cpu.icache.r_tag[3][20] ),
    .B(_06470_));
 sg13g2_o21ai_1 _25291_ (.B1(_06476_),
    .Y(_02309_),
    .A1(net385),
    .A2(_06469_));
 sg13g2_nand2_1 _25292_ (.Y(_06477_),
    .A(\cpu.icache.r_tag[3][21] ),
    .B(_06364_));
 sg13g2_o21ai_1 _25293_ (.B1(_06477_),
    .Y(_02310_),
    .A1(net384),
    .A2(net235));
 sg13g2_nand2_1 _25294_ (.Y(_06478_),
    .A(\cpu.icache.r_tag[3][22] ),
    .B(net262));
 sg13g2_o21ai_1 _25295_ (.B1(_06478_),
    .Y(_02311_),
    .A1(net435),
    .A2(net235));
 sg13g2_nand2_1 _25296_ (.Y(_06479_),
    .A(\cpu.icache.r_tag[3][23] ),
    .B(net262));
 sg13g2_o21ai_1 _25297_ (.B1(_06479_),
    .Y(_02312_),
    .A1(net469),
    .A2(net235));
 sg13g2_nand2_1 _25298_ (.Y(_06480_),
    .A(\cpu.icache.r_tag[3][6] ),
    .B(net262));
 sg13g2_o21ai_1 _25299_ (.B1(_06480_),
    .Y(_02313_),
    .A1(net1047),
    .A2(net236));
 sg13g2_mux2_1 _25300_ (.A0(net956),
    .A1(\cpu.icache.r_tag[3][7] ),
    .S(net258),
    .X(_02314_));
 sg13g2_mux2_1 _25301_ (.A0(net955),
    .A1(\cpu.icache.r_tag[3][8] ),
    .S(net258),
    .X(_02315_));
 sg13g2_nand2_1 _25302_ (.Y(_06481_),
    .A(\cpu.icache.r_tag[3][9] ),
    .B(net262));
 sg13g2_o21ai_1 _25303_ (.B1(_06481_),
    .Y(_02316_),
    .A1(net958),
    .A2(net236));
 sg13g2_mux2_1 _25304_ (.A0(net954),
    .A1(\cpu.icache.r_tag[3][10] ),
    .S(net258),
    .X(_02317_));
 sg13g2_mux2_1 _25305_ (.A0(net959),
    .A1(\cpu.icache.r_tag[3][11] ),
    .S(net258),
    .X(_02318_));
 sg13g2_nand2_1 _25306_ (.Y(_06482_),
    .A(\cpu.icache.r_tag[3][12] ),
    .B(net262));
 sg13g2_o21ai_1 _25307_ (.B1(_06482_),
    .Y(_02319_),
    .A1(net438),
    .A2(net236));
 sg13g2_nand2_1 _25308_ (.Y(_06483_),
    .A(\cpu.icache.r_tag[3][13] ),
    .B(_06364_));
 sg13g2_o21ai_1 _25309_ (.B1(_06483_),
    .Y(_02320_),
    .A1(net386),
    .A2(net236));
 sg13g2_nand2_1 _25310_ (.Y(_06484_),
    .A(\cpu.icache.r_tag[3][14] ),
    .B(net262));
 sg13g2_o21ai_1 _25311_ (.B1(_06484_),
    .Y(_02321_),
    .A1(net382),
    .A2(net236));
 sg13g2_nand2_1 _25312_ (.Y(_06485_),
    .A(net610),
    .B(_06430_));
 sg13g2_buf_1 _25313_ (.A(_06485_),
    .X(_06486_));
 sg13g2_buf_1 _25314_ (.A(_06486_),
    .X(_06487_));
 sg13g2_mux2_1 _25315_ (.A0(net957),
    .A1(\cpu.icache.r_tag[4][5] ),
    .S(net396),
    .X(_02322_));
 sg13g2_buf_1 _25316_ (.A(_06486_),
    .X(_06488_));
 sg13g2_nand2_1 _25317_ (.Y(_06489_),
    .A(\cpu.icache.r_tag[4][15] ),
    .B(net396));
 sg13g2_o21ai_1 _25318_ (.B1(_06489_),
    .Y(_02323_),
    .A1(net380),
    .A2(net395));
 sg13g2_buf_1 _25319_ (.A(_06486_),
    .X(_06490_));
 sg13g2_nand2_1 _25320_ (.Y(_06491_),
    .A(\cpu.icache.r_tag[4][16] ),
    .B(net394));
 sg13g2_o21ai_1 _25321_ (.B1(_06491_),
    .Y(_02324_),
    .A1(net383),
    .A2(net395));
 sg13g2_nand2_1 _25322_ (.Y(_06492_),
    .A(\cpu.icache.r_tag[4][17] ),
    .B(net394));
 sg13g2_o21ai_1 _25323_ (.B1(_06492_),
    .Y(_02325_),
    .A1(net437),
    .A2(net395));
 sg13g2_nand2_1 _25324_ (.Y(_06493_),
    .A(\cpu.icache.r_tag[4][18] ),
    .B(net394));
 sg13g2_o21ai_1 _25325_ (.B1(_06493_),
    .Y(_02326_),
    .A1(net436),
    .A2(net395));
 sg13g2_nand2_1 _25326_ (.Y(_06494_),
    .A(\cpu.icache.r_tag[4][19] ),
    .B(net394));
 sg13g2_o21ai_1 _25327_ (.B1(_06494_),
    .Y(_02327_),
    .A1(net381),
    .A2(_06488_));
 sg13g2_nand2_1 _25328_ (.Y(_06495_),
    .A(\cpu.icache.r_tag[4][20] ),
    .B(net394));
 sg13g2_o21ai_1 _25329_ (.B1(_06495_),
    .Y(_02328_),
    .A1(net385),
    .A2(_06488_));
 sg13g2_nand2_1 _25330_ (.Y(_06496_),
    .A(\cpu.icache.r_tag[4][21] ),
    .B(net394));
 sg13g2_o21ai_1 _25331_ (.B1(_06496_),
    .Y(_02329_),
    .A1(net384),
    .A2(net395));
 sg13g2_nand2_1 _25332_ (.Y(_06497_),
    .A(\cpu.icache.r_tag[4][22] ),
    .B(net394));
 sg13g2_o21ai_1 _25333_ (.B1(_06497_),
    .Y(_02330_),
    .A1(net435),
    .A2(net395));
 sg13g2_nand2_1 _25334_ (.Y(_06498_),
    .A(\cpu.icache.r_tag[4][23] ),
    .B(net394));
 sg13g2_o21ai_1 _25335_ (.B1(_06498_),
    .Y(_02331_),
    .A1(net469),
    .A2(net395));
 sg13g2_nand2_1 _25336_ (.Y(_06499_),
    .A(\cpu.icache.r_tag[4][6] ),
    .B(_06490_));
 sg13g2_o21ai_1 _25337_ (.B1(_06499_),
    .Y(_02332_),
    .A1(net1047),
    .A2(net395));
 sg13g2_mux2_1 _25338_ (.A0(net956),
    .A1(\cpu.icache.r_tag[4][7] ),
    .S(net396),
    .X(_02333_));
 sg13g2_mux2_1 _25339_ (.A0(net955),
    .A1(\cpu.icache.r_tag[4][8] ),
    .S(net396),
    .X(_02334_));
 sg13g2_nand2_1 _25340_ (.Y(_06500_),
    .A(\cpu.icache.r_tag[4][9] ),
    .B(_06490_));
 sg13g2_o21ai_1 _25341_ (.B1(_06500_),
    .Y(_02335_),
    .A1(net958),
    .A2(_06487_));
 sg13g2_mux2_1 _25342_ (.A0(net954),
    .A1(\cpu.icache.r_tag[4][10] ),
    .S(net396),
    .X(_02336_));
 sg13g2_mux2_1 _25343_ (.A0(net959),
    .A1(\cpu.icache.r_tag[4][11] ),
    .S(net396),
    .X(_02337_));
 sg13g2_nand2_1 _25344_ (.Y(_06501_),
    .A(\cpu.icache.r_tag[4][12] ),
    .B(_06486_));
 sg13g2_o21ai_1 _25345_ (.B1(_06501_),
    .Y(_02338_),
    .A1(net438),
    .A2(net396));
 sg13g2_nand2_1 _25346_ (.Y(_06502_),
    .A(\cpu.icache.r_tag[4][13] ),
    .B(_06486_));
 sg13g2_o21ai_1 _25347_ (.B1(_06502_),
    .Y(_02339_),
    .A1(net386),
    .A2(_06487_));
 sg13g2_nand2_1 _25348_ (.Y(_06503_),
    .A(\cpu.icache.r_tag[4][14] ),
    .B(_06486_));
 sg13g2_o21ai_1 _25349_ (.B1(_06503_),
    .Y(_02340_),
    .A1(net382),
    .A2(net396));
 sg13g2_nand2_1 _25350_ (.Y(_06504_),
    .A(net611),
    .B(_06430_));
 sg13g2_buf_1 _25351_ (.A(_06504_),
    .X(_06505_));
 sg13g2_buf_1 _25352_ (.A(_06505_),
    .X(_06506_));
 sg13g2_mux2_1 _25353_ (.A0(net957),
    .A1(\cpu.icache.r_tag[5][5] ),
    .S(net393),
    .X(_02341_));
 sg13g2_buf_1 _25354_ (.A(_06505_),
    .X(_06507_));
 sg13g2_nand2_1 _25355_ (.Y(_06508_),
    .A(\cpu.icache.r_tag[5][15] ),
    .B(_06506_));
 sg13g2_o21ai_1 _25356_ (.B1(_06508_),
    .Y(_02342_),
    .A1(net380),
    .A2(_06507_));
 sg13g2_buf_1 _25357_ (.A(_06505_),
    .X(_06509_));
 sg13g2_nand2_1 _25358_ (.Y(_06510_),
    .A(\cpu.icache.r_tag[5][16] ),
    .B(net391));
 sg13g2_o21ai_1 _25359_ (.B1(_06510_),
    .Y(_02343_),
    .A1(net383),
    .A2(net392));
 sg13g2_nand2_1 _25360_ (.Y(_06511_),
    .A(\cpu.icache.r_tag[5][17] ),
    .B(net391));
 sg13g2_o21ai_1 _25361_ (.B1(_06511_),
    .Y(_02344_),
    .A1(net437),
    .A2(net392));
 sg13g2_nand2_1 _25362_ (.Y(_06512_),
    .A(\cpu.icache.r_tag[5][18] ),
    .B(net391));
 sg13g2_o21ai_1 _25363_ (.B1(_06512_),
    .Y(_02345_),
    .A1(net436),
    .A2(net392));
 sg13g2_nand2_1 _25364_ (.Y(_06513_),
    .A(\cpu.icache.r_tag[5][19] ),
    .B(net391));
 sg13g2_o21ai_1 _25365_ (.B1(_06513_),
    .Y(_02346_),
    .A1(net381),
    .A2(_06507_));
 sg13g2_nand2_1 _25366_ (.Y(_06514_),
    .A(\cpu.icache.r_tag[5][20] ),
    .B(_06509_));
 sg13g2_o21ai_1 _25367_ (.B1(_06514_),
    .Y(_02347_),
    .A1(net385),
    .A2(net392));
 sg13g2_nand2_1 _25368_ (.Y(_06515_),
    .A(\cpu.icache.r_tag[5][21] ),
    .B(_06509_));
 sg13g2_o21ai_1 _25369_ (.B1(_06515_),
    .Y(_02348_),
    .A1(net384),
    .A2(net392));
 sg13g2_nand2_1 _25370_ (.Y(_06516_),
    .A(\cpu.icache.r_tag[5][22] ),
    .B(net391));
 sg13g2_o21ai_1 _25371_ (.B1(_06516_),
    .Y(_02349_),
    .A1(net435),
    .A2(net392));
 sg13g2_nand2_1 _25372_ (.Y(_06517_),
    .A(\cpu.icache.r_tag[5][23] ),
    .B(net391));
 sg13g2_o21ai_1 _25373_ (.B1(_06517_),
    .Y(_02350_),
    .A1(net469),
    .A2(net392));
 sg13g2_nand2_1 _25374_ (.Y(_06518_),
    .A(\cpu.icache.r_tag[5][6] ),
    .B(net391));
 sg13g2_o21ai_1 _25375_ (.B1(_06518_),
    .Y(_02351_),
    .A1(net1047),
    .A2(net392));
 sg13g2_mux2_1 _25376_ (.A0(net956),
    .A1(\cpu.icache.r_tag[5][7] ),
    .S(net393),
    .X(_02352_));
 sg13g2_mux2_1 _25377_ (.A0(net955),
    .A1(\cpu.icache.r_tag[5][8] ),
    .S(net393),
    .X(_02353_));
 sg13g2_nand2_1 _25378_ (.Y(_06519_),
    .A(\cpu.icache.r_tag[5][9] ),
    .B(net391));
 sg13g2_o21ai_1 _25379_ (.B1(_06519_),
    .Y(_02354_),
    .A1(net958),
    .A2(net393));
 sg13g2_mux2_1 _25380_ (.A0(net954),
    .A1(\cpu.icache.r_tag[5][10] ),
    .S(net393),
    .X(_02355_));
 sg13g2_mux2_1 _25381_ (.A0(net959),
    .A1(\cpu.icache.r_tag[5][11] ),
    .S(net393),
    .X(_02356_));
 sg13g2_nand2_1 _25382_ (.Y(_06520_),
    .A(\cpu.icache.r_tag[5][12] ),
    .B(_06505_));
 sg13g2_o21ai_1 _25383_ (.B1(_06520_),
    .Y(_02357_),
    .A1(net438),
    .A2(_06506_));
 sg13g2_nand2_1 _25384_ (.Y(_06521_),
    .A(\cpu.icache.r_tag[5][13] ),
    .B(_06505_));
 sg13g2_o21ai_1 _25385_ (.B1(_06521_),
    .Y(_02358_),
    .A1(net386),
    .A2(net393));
 sg13g2_nand2_1 _25386_ (.Y(_06522_),
    .A(\cpu.icache.r_tag[5][14] ),
    .B(_06505_));
 sg13g2_o21ai_1 _25387_ (.B1(_06522_),
    .Y(_02359_),
    .A1(net382),
    .A2(net393));
 sg13g2_nand2_1 _25388_ (.Y(_06523_),
    .A(net466),
    .B(_06430_));
 sg13g2_buf_1 _25389_ (.A(_06523_),
    .X(_06524_));
 sg13g2_buf_1 _25390_ (.A(_06524_),
    .X(_06525_));
 sg13g2_mux2_1 _25391_ (.A0(_04561_),
    .A1(\cpu.icache.r_tag[6][5] ),
    .S(net257),
    .X(_02360_));
 sg13g2_buf_1 _25392_ (.A(_06524_),
    .X(_06526_));
 sg13g2_nand2_1 _25393_ (.Y(_06527_),
    .A(\cpu.icache.r_tag[6][15] ),
    .B(net257));
 sg13g2_o21ai_1 _25394_ (.B1(_06527_),
    .Y(_02361_),
    .A1(net380),
    .A2(_06526_));
 sg13g2_buf_1 _25395_ (.A(_06524_),
    .X(_06528_));
 sg13g2_nand2_1 _25396_ (.Y(_06529_),
    .A(\cpu.icache.r_tag[6][16] ),
    .B(net255));
 sg13g2_o21ai_1 _25397_ (.B1(_06529_),
    .Y(_02362_),
    .A1(net383),
    .A2(net256));
 sg13g2_nand2_1 _25398_ (.Y(_06530_),
    .A(\cpu.icache.r_tag[6][17] ),
    .B(net255));
 sg13g2_o21ai_1 _25399_ (.B1(_06530_),
    .Y(_02363_),
    .A1(net437),
    .A2(net256));
 sg13g2_nand2_1 _25400_ (.Y(_06531_),
    .A(\cpu.icache.r_tag[6][18] ),
    .B(net255));
 sg13g2_o21ai_1 _25401_ (.B1(_06531_),
    .Y(_02364_),
    .A1(net436),
    .A2(net256));
 sg13g2_nand2_1 _25402_ (.Y(_06532_),
    .A(\cpu.icache.r_tag[6][19] ),
    .B(net255));
 sg13g2_o21ai_1 _25403_ (.B1(_06532_),
    .Y(_02365_),
    .A1(net381),
    .A2(net256));
 sg13g2_nand2_1 _25404_ (.Y(_06533_),
    .A(\cpu.icache.r_tag[6][20] ),
    .B(net255));
 sg13g2_o21ai_1 _25405_ (.B1(_06533_),
    .Y(_02366_),
    .A1(net385),
    .A2(net256));
 sg13g2_nand2_1 _25406_ (.Y(_06534_),
    .A(\cpu.icache.r_tag[6][21] ),
    .B(net255));
 sg13g2_o21ai_1 _25407_ (.B1(_06534_),
    .Y(_02367_),
    .A1(net384),
    .A2(net256));
 sg13g2_nand2_1 _25408_ (.Y(_06535_),
    .A(\cpu.icache.r_tag[6][22] ),
    .B(net255));
 sg13g2_o21ai_1 _25409_ (.B1(_06535_),
    .Y(_02368_),
    .A1(net435),
    .A2(net256));
 sg13g2_nand2_1 _25410_ (.Y(_06536_),
    .A(\cpu.icache.r_tag[6][23] ),
    .B(net255));
 sg13g2_o21ai_1 _25411_ (.B1(_06536_),
    .Y(_02369_),
    .A1(net469),
    .A2(net256));
 sg13g2_nand2_1 _25412_ (.Y(_06537_),
    .A(\cpu.icache.r_tag[6][6] ),
    .B(_06528_));
 sg13g2_o21ai_1 _25413_ (.B1(_06537_),
    .Y(_02370_),
    .A1(net1047),
    .A2(_06526_));
 sg13g2_mux2_1 _25414_ (.A0(_04656_),
    .A1(\cpu.icache.r_tag[6][7] ),
    .S(net257),
    .X(_02371_));
 sg13g2_mux2_1 _25415_ (.A0(_04693_),
    .A1(\cpu.icache.r_tag[6][8] ),
    .S(net257),
    .X(_02372_));
 sg13g2_nand2_1 _25416_ (.Y(_06538_),
    .A(\cpu.icache.r_tag[6][9] ),
    .B(_06528_));
 sg13g2_o21ai_1 _25417_ (.B1(_06538_),
    .Y(_02373_),
    .A1(net958),
    .A2(_06525_));
 sg13g2_mux2_1 _25418_ (.A0(_04762_),
    .A1(\cpu.icache.r_tag[6][10] ),
    .S(net257),
    .X(_02374_));
 sg13g2_mux2_1 _25419_ (.A0(_04244_),
    .A1(\cpu.icache.r_tag[6][11] ),
    .S(net257),
    .X(_02375_));
 sg13g2_nand2_1 _25420_ (.Y(_06539_),
    .A(\cpu.icache.r_tag[6][12] ),
    .B(_06524_));
 sg13g2_o21ai_1 _25421_ (.B1(_06539_),
    .Y(_02376_),
    .A1(net438),
    .A2(net257));
 sg13g2_nand2_1 _25422_ (.Y(_06540_),
    .A(\cpu.icache.r_tag[6][13] ),
    .B(_06524_));
 sg13g2_o21ai_1 _25423_ (.B1(_06540_),
    .Y(_02377_),
    .A1(net386),
    .A2(_06525_));
 sg13g2_nand2_1 _25424_ (.Y(_06541_),
    .A(\cpu.icache.r_tag[6][14] ),
    .B(_06524_));
 sg13g2_o21ai_1 _25425_ (.B1(_06541_),
    .Y(_02378_),
    .A1(_08473_),
    .A2(net257));
 sg13g2_nand2_1 _25426_ (.Y(_06542_),
    .A(net615),
    .B(_06430_));
 sg13g2_buf_1 _25427_ (.A(_06542_),
    .X(_06543_));
 sg13g2_buf_1 _25428_ (.A(_06543_),
    .X(_06544_));
 sg13g2_mux2_1 _25429_ (.A0(_04561_),
    .A1(\cpu.icache.r_tag[7][5] ),
    .S(net390),
    .X(_02379_));
 sg13g2_buf_1 _25430_ (.A(_06543_),
    .X(_06545_));
 sg13g2_nand2_1 _25431_ (.Y(_06546_),
    .A(\cpu.icache.r_tag[7][15] ),
    .B(net390));
 sg13g2_o21ai_1 _25432_ (.B1(_06546_),
    .Y(_02380_),
    .A1(net380),
    .A2(_06545_));
 sg13g2_buf_1 _25433_ (.A(_06543_),
    .X(_06547_));
 sg13g2_nand2_1 _25434_ (.Y(_06548_),
    .A(\cpu.icache.r_tag[7][16] ),
    .B(net388));
 sg13g2_o21ai_1 _25435_ (.B1(_06548_),
    .Y(_02381_),
    .A1(net383),
    .A2(net389));
 sg13g2_nand2_1 _25436_ (.Y(_06549_),
    .A(\cpu.icache.r_tag[7][17] ),
    .B(net388));
 sg13g2_o21ai_1 _25437_ (.B1(_06549_),
    .Y(_02382_),
    .A1(_08557_),
    .A2(net389));
 sg13g2_nand2_1 _25438_ (.Y(_06550_),
    .A(\cpu.icache.r_tag[7][18] ),
    .B(net388));
 sg13g2_o21ai_1 _25439_ (.B1(_06550_),
    .Y(_02383_),
    .A1(net436),
    .A2(net389));
 sg13g2_nand2_1 _25440_ (.Y(_06551_),
    .A(\cpu.icache.r_tag[7][19] ),
    .B(net388));
 sg13g2_o21ai_1 _25441_ (.B1(_06551_),
    .Y(_02384_),
    .A1(net381),
    .A2(net389));
 sg13g2_nand2_1 _25442_ (.Y(_06552_),
    .A(\cpu.icache.r_tag[7][20] ),
    .B(net388));
 sg13g2_o21ai_1 _25443_ (.B1(_06552_),
    .Y(_02385_),
    .A1(net385),
    .A2(net389));
 sg13g2_nand2_1 _25444_ (.Y(_06553_),
    .A(\cpu.icache.r_tag[7][21] ),
    .B(net388));
 sg13g2_o21ai_1 _25445_ (.B1(_06553_),
    .Y(_02386_),
    .A1(net384),
    .A2(net389));
 sg13g2_nand2_1 _25446_ (.Y(_06554_),
    .A(\cpu.icache.r_tag[7][22] ),
    .B(net388));
 sg13g2_o21ai_1 _25447_ (.B1(_06554_),
    .Y(_02387_),
    .A1(net435),
    .A2(net389));
 sg13g2_nand2_1 _25448_ (.Y(_06555_),
    .A(\cpu.icache.r_tag[7][23] ),
    .B(net388));
 sg13g2_o21ai_1 _25449_ (.B1(_06555_),
    .Y(_02388_),
    .A1(net469),
    .A2(net389));
 sg13g2_nand2_1 _25450_ (.Y(_06556_),
    .A(\cpu.icache.r_tag[7][6] ),
    .B(_06547_));
 sg13g2_o21ai_1 _25451_ (.B1(_06556_),
    .Y(_02389_),
    .A1(_08648_),
    .A2(_06545_));
 sg13g2_mux2_1 _25452_ (.A0(_04656_),
    .A1(\cpu.icache.r_tag[7][7] ),
    .S(net390),
    .X(_02390_));
 sg13g2_mux2_1 _25453_ (.A0(_04693_),
    .A1(\cpu.icache.r_tag[7][8] ),
    .S(net390),
    .X(_02391_));
 sg13g2_nand2_1 _25454_ (.Y(_06557_),
    .A(\cpu.icache.r_tag[7][9] ),
    .B(_06547_));
 sg13g2_o21ai_1 _25455_ (.B1(_06557_),
    .Y(_02392_),
    .A1(_04245_),
    .A2(_06544_));
 sg13g2_mux2_1 _25456_ (.A0(_04762_),
    .A1(\cpu.icache.r_tag[7][10] ),
    .S(net390),
    .X(_02393_));
 sg13g2_mux2_1 _25457_ (.A0(_04244_),
    .A1(\cpu.icache.r_tag[7][11] ),
    .S(net390),
    .X(_02394_));
 sg13g2_nand2_1 _25458_ (.Y(_06558_),
    .A(\cpu.icache.r_tag[7][12] ),
    .B(_06543_));
 sg13g2_o21ai_1 _25459_ (.B1(_06558_),
    .Y(_02395_),
    .A1(net438),
    .A2(net390));
 sg13g2_nand2_1 _25460_ (.Y(_06559_),
    .A(\cpu.icache.r_tag[7][13] ),
    .B(_06543_));
 sg13g2_o21ai_1 _25461_ (.B1(_06559_),
    .Y(_02396_),
    .A1(_08356_),
    .A2(net390));
 sg13g2_nand2_1 _25462_ (.Y(_06560_),
    .A(\cpu.icache.r_tag[7][14] ),
    .B(_06543_));
 sg13g2_o21ai_1 _25463_ (.B1(_06560_),
    .Y(_02397_),
    .A1(net382),
    .A2(_06544_));
 sg13g2_buf_1 _25464_ (.A(_09786_),
    .X(_06561_));
 sg13g2_nand2_1 _25465_ (.Y(_06562_),
    .A(net130),
    .B(net403));
 sg13g2_buf_2 _25466_ (.A(_06562_),
    .X(_06563_));
 sg13g2_buf_1 _25467_ (.A(_06563_),
    .X(_06564_));
 sg13g2_mux2_1 _25468_ (.A0(net880),
    .A1(\cpu.intr.r_clock_cmp[0] ),
    .S(net82),
    .X(_02407_));
 sg13g2_buf_1 _25469_ (.A(_06563_),
    .X(_06565_));
 sg13g2_mux2_1 _25470_ (.A0(_09986_),
    .A1(\cpu.intr.r_clock_cmp[10] ),
    .S(net81),
    .X(_02408_));
 sg13g2_mux2_1 _25471_ (.A0(_09991_),
    .A1(\cpu.intr.r_clock_cmp[11] ),
    .S(net81),
    .X(_02409_));
 sg13g2_nand2_1 _25472_ (.Y(_06566_),
    .A(\cpu.intr.r_clock_cmp[12] ),
    .B(_06565_));
 sg13g2_o21ai_1 _25473_ (.B1(_06566_),
    .Y(_02410_),
    .A1(_12060_),
    .A2(net82));
 sg13g2_nand2_1 _25474_ (.Y(_06567_),
    .A(\cpu.intr.r_clock_cmp[13] ),
    .B(net81));
 sg13g2_o21ai_1 _25475_ (.B1(_06567_),
    .Y(_02411_),
    .A1(_12070_),
    .A2(net82));
 sg13g2_nand2_1 _25476_ (.Y(_06568_),
    .A(\cpu.intr.r_clock_cmp[14] ),
    .B(net81));
 sg13g2_o21ai_1 _25477_ (.B1(_06568_),
    .Y(_02412_),
    .A1(_12077_),
    .A2(net82));
 sg13g2_nand2_1 _25478_ (.Y(_06569_),
    .A(\cpu.intr.r_clock_cmp[15] ),
    .B(net81));
 sg13g2_o21ai_1 _25479_ (.B1(_06569_),
    .Y(_02413_),
    .A1(_12084_),
    .A2(net82));
 sg13g2_nand2_1 _25480_ (.Y(_06570_),
    .A(_09786_),
    .B(net444));
 sg13g2_buf_1 _25481_ (.A(_06570_),
    .X(_06571_));
 sg13g2_buf_1 _25482_ (.A(_06571_),
    .X(_06572_));
 sg13g2_mux2_1 _25483_ (.A0(net880),
    .A1(\cpu.intr.r_clock_cmp[16] ),
    .S(net92),
    .X(_02414_));
 sg13g2_buf_1 _25484_ (.A(_06571_),
    .X(_06573_));
 sg13g2_mux2_1 _25485_ (.A0(net829),
    .A1(\cpu.intr.r_clock_cmp[17] ),
    .S(net91),
    .X(_02415_));
 sg13g2_nand2_1 _25486_ (.Y(_06574_),
    .A(\cpu.intr.r_clock_cmp[18] ),
    .B(net91));
 sg13g2_o21ai_1 _25487_ (.B1(_06574_),
    .Y(_02416_),
    .A1(net753),
    .A2(_06572_));
 sg13g2_nand2_1 _25488_ (.Y(_06575_),
    .A(\cpu.intr.r_clock_cmp[19] ),
    .B(_06573_));
 sg13g2_o21ai_1 _25489_ (.B1(_06575_),
    .Y(_02417_),
    .A1(net854),
    .A2(_06572_));
 sg13g2_mux2_1 _25490_ (.A0(net829),
    .A1(\cpu.intr.r_clock_cmp[1] ),
    .S(net81),
    .X(_02418_));
 sg13g2_nand2_1 _25491_ (.Y(_06576_),
    .A(\cpu.intr.r_clock_cmp[20] ),
    .B(net91));
 sg13g2_o21ai_1 _25492_ (.B1(_06576_),
    .Y(_02419_),
    .A1(net720),
    .A2(net92));
 sg13g2_mux2_1 _25493_ (.A0(net849),
    .A1(\cpu.intr.r_clock_cmp[21] ),
    .S(net91),
    .X(_02420_));
 sg13g2_mux2_1 _25494_ (.A0(net875),
    .A1(\cpu.intr.r_clock_cmp[22] ),
    .S(_06573_),
    .X(_02421_));
 sg13g2_nand2_1 _25495_ (.Y(_06577_),
    .A(\cpu.intr.r_clock_cmp[23] ),
    .B(net91));
 sg13g2_o21ai_1 _25496_ (.B1(_06577_),
    .Y(_02422_),
    .A1(net719),
    .A2(net92));
 sg13g2_mux2_1 _25497_ (.A0(_09975_),
    .A1(\cpu.intr.r_clock_cmp[24] ),
    .S(net91),
    .X(_02423_));
 sg13g2_nand2_1 _25498_ (.Y(_06578_),
    .A(\cpu.intr.r_clock_cmp[25] ),
    .B(_06571_));
 sg13g2_o21ai_1 _25499_ (.B1(_06578_),
    .Y(_02424_),
    .A1(_12157_),
    .A2(net92));
 sg13g2_mux2_1 _25500_ (.A0(_09986_),
    .A1(\cpu.intr.r_clock_cmp[26] ),
    .S(net91),
    .X(_02425_));
 sg13g2_mux2_1 _25501_ (.A0(_09991_),
    .A1(\cpu.intr.r_clock_cmp[27] ),
    .S(net91),
    .X(_02426_));
 sg13g2_nand2_1 _25502_ (.Y(_06579_),
    .A(\cpu.intr.r_clock_cmp[28] ),
    .B(_06571_));
 sg13g2_o21ai_1 _25503_ (.B1(_06579_),
    .Y(_02427_),
    .A1(_12060_),
    .A2(net92));
 sg13g2_nand2_1 _25504_ (.Y(_06580_),
    .A(\cpu.intr.r_clock_cmp[29] ),
    .B(_06571_));
 sg13g2_o21ai_1 _25505_ (.B1(_06580_),
    .Y(_02428_),
    .A1(_12070_),
    .A2(net92));
 sg13g2_nand2_1 _25506_ (.Y(_06581_),
    .A(\cpu.intr.r_clock_cmp[2] ),
    .B(_06563_));
 sg13g2_o21ai_1 _25507_ (.B1(_06581_),
    .Y(_02429_),
    .A1(net753),
    .A2(net82));
 sg13g2_nand2_1 _25508_ (.Y(_06582_),
    .A(\cpu.intr.r_clock_cmp[30] ),
    .B(_06571_));
 sg13g2_o21ai_1 _25509_ (.B1(_06582_),
    .Y(_02430_),
    .A1(_12077_),
    .A2(net92));
 sg13g2_nand2_1 _25510_ (.Y(_06583_),
    .A(\cpu.intr.r_clock_cmp[31] ),
    .B(_06571_));
 sg13g2_o21ai_1 _25511_ (.B1(_06583_),
    .Y(_02431_),
    .A1(_12084_),
    .A2(net92));
 sg13g2_nand2_1 _25512_ (.Y(_06584_),
    .A(\cpu.intr.r_clock_cmp[3] ),
    .B(_06563_));
 sg13g2_o21ai_1 _25513_ (.B1(_06584_),
    .Y(_02432_),
    .A1(net854),
    .A2(net82));
 sg13g2_nand2_1 _25514_ (.Y(_06585_),
    .A(\cpu.intr.r_clock_cmp[4] ),
    .B(_06563_));
 sg13g2_o21ai_1 _25515_ (.B1(_06585_),
    .Y(_02433_),
    .A1(net720),
    .A2(_06564_));
 sg13g2_mux2_1 _25516_ (.A0(net849),
    .A1(\cpu.intr.r_clock_cmp[5] ),
    .S(_06565_),
    .X(_02434_));
 sg13g2_mux2_1 _25517_ (.A0(net875),
    .A1(\cpu.intr.r_clock_cmp[6] ),
    .S(net81),
    .X(_02435_));
 sg13g2_nand2_1 _25518_ (.Y(_06586_),
    .A(\cpu.intr.r_clock_cmp[7] ),
    .B(_06563_));
 sg13g2_o21ai_1 _25519_ (.B1(_06586_),
    .Y(_02436_),
    .A1(net852),
    .A2(_06564_));
 sg13g2_mux2_1 _25520_ (.A0(_09975_),
    .A1(\cpu.intr.r_clock_cmp[8] ),
    .S(net81),
    .X(_02437_));
 sg13g2_nand2_1 _25521_ (.Y(_06587_),
    .A(\cpu.intr.r_clock_cmp[9] ),
    .B(_06563_));
 sg13g2_o21ai_1 _25522_ (.B1(_06587_),
    .Y(_02438_),
    .A1(_12157_),
    .A2(net82));
 sg13g2_nand2_1 _25523_ (.Y(_06588_),
    .A(_09786_),
    .B(net488));
 sg13g2_buf_1 _25524_ (.A(_06588_),
    .X(_06589_));
 sg13g2_buf_1 _25525_ (.A(_06589_),
    .X(_06590_));
 sg13g2_mux2_1 _25526_ (.A0(net880),
    .A1(\cpu.intr.r_timer_reload[0] ),
    .S(net90),
    .X(_02462_));
 sg13g2_buf_1 _25527_ (.A(_06589_),
    .X(_06591_));
 sg13g2_mux2_1 _25528_ (.A0(_09986_),
    .A1(\cpu.intr.r_timer_reload[10] ),
    .S(net89),
    .X(_02463_));
 sg13g2_mux2_1 _25529_ (.A0(_09991_),
    .A1(\cpu.intr.r_timer_reload[11] ),
    .S(net89),
    .X(_02464_));
 sg13g2_nand2_1 _25530_ (.Y(_06592_),
    .A(\cpu.intr.r_timer_reload[12] ),
    .B(net89));
 sg13g2_o21ai_1 _25531_ (.B1(_06592_),
    .Y(_02465_),
    .A1(_12060_),
    .A2(net90));
 sg13g2_nand2_1 _25532_ (.Y(_06593_),
    .A(\cpu.intr.r_timer_reload[13] ),
    .B(net89));
 sg13g2_o21ai_1 _25533_ (.B1(_06593_),
    .Y(_02466_),
    .A1(_12070_),
    .A2(net90));
 sg13g2_nand2_1 _25534_ (.Y(_06594_),
    .A(\cpu.intr.r_timer_reload[14] ),
    .B(net89));
 sg13g2_o21ai_1 _25535_ (.B1(_06594_),
    .Y(_02467_),
    .A1(_12077_),
    .A2(net90));
 sg13g2_nand2_1 _25536_ (.Y(_06595_),
    .A(\cpu.intr.r_timer_reload[15] ),
    .B(_06591_));
 sg13g2_o21ai_1 _25537_ (.B1(_06595_),
    .Y(_02468_),
    .A1(_12084_),
    .A2(net90));
 sg13g2_mux2_1 _25538_ (.A0(\cpu.intr.r_timer_reload[16] ),
    .A1(net877),
    .S(net148),
    .X(_02469_));
 sg13g2_o21ai_1 _25539_ (.B1(_09880_),
    .Y(_02470_),
    .A1(_05335_),
    .A2(net148));
 sg13g2_nand2_1 _25540_ (.Y(_06596_),
    .A(\cpu.intr.r_timer_reload[18] ),
    .B(net102));
 sg13g2_o21ai_1 _25541_ (.B1(_06596_),
    .Y(_02471_),
    .A1(net878),
    .A2(net102));
 sg13g2_inv_1 _25542_ (.Y(_06597_),
    .A(\cpu.intr.r_timer_reload[19] ));
 sg13g2_o21ai_1 _25543_ (.B1(_09891_),
    .Y(_02472_),
    .A1(_06597_),
    .A2(net148));
 sg13g2_mux2_1 _25544_ (.A0(net829),
    .A1(\cpu.intr.r_timer_reload[1] ),
    .S(net89),
    .X(_02473_));
 sg13g2_nand2_1 _25545_ (.Y(_06598_),
    .A(\cpu.intr.r_timer_reload[20] ),
    .B(_09865_));
 sg13g2_o21ai_1 _25546_ (.B1(_06598_),
    .Y(_02474_),
    .A1(net853),
    .A2(_09865_));
 sg13g2_inv_1 _25547_ (.Y(_06599_),
    .A(\cpu.intr.r_timer_reload[21] ));
 sg13g2_o21ai_1 _25548_ (.B1(_09903_),
    .Y(_02475_),
    .A1(_06599_),
    .A2(_09879_));
 sg13g2_inv_1 _25549_ (.Y(_06600_),
    .A(\cpu.intr.r_timer_reload[22] ));
 sg13g2_o21ai_1 _25550_ (.B1(_09909_),
    .Y(_02476_),
    .A1(_06600_),
    .A2(_09879_));
 sg13g2_nand2_1 _25551_ (.Y(_06601_),
    .A(\cpu.intr.r_timer_reload[23] ),
    .B(net102));
 sg13g2_o21ai_1 _25552_ (.B1(_06601_),
    .Y(_02477_),
    .A1(_12139_),
    .A2(net102));
 sg13g2_nand2_1 _25553_ (.Y(_06602_),
    .A(\cpu.intr.r_timer_reload[2] ),
    .B(_06589_));
 sg13g2_o21ai_1 _25554_ (.B1(_06602_),
    .Y(_02478_),
    .A1(net878),
    .A2(net90));
 sg13g2_nand2_1 _25555_ (.Y(_06603_),
    .A(\cpu.intr.r_timer_reload[3] ),
    .B(_06589_));
 sg13g2_o21ai_1 _25556_ (.B1(_06603_),
    .Y(_02479_),
    .A1(net854),
    .A2(_06590_));
 sg13g2_nand2_1 _25557_ (.Y(_06604_),
    .A(\cpu.intr.r_timer_reload[4] ),
    .B(_06589_));
 sg13g2_o21ai_1 _25558_ (.B1(_06604_),
    .Y(_02480_),
    .A1(net853),
    .A2(_06590_));
 sg13g2_mux2_1 _25559_ (.A0(net849),
    .A1(\cpu.intr.r_timer_reload[5] ),
    .S(net89),
    .X(_02481_));
 sg13g2_mux2_1 _25560_ (.A0(net875),
    .A1(\cpu.intr.r_timer_reload[6] ),
    .S(net89),
    .X(_02482_));
 sg13g2_nand2_1 _25561_ (.Y(_06605_),
    .A(\cpu.intr.r_timer_reload[7] ),
    .B(_06589_));
 sg13g2_o21ai_1 _25562_ (.B1(_06605_),
    .Y(_02483_),
    .A1(net852),
    .A2(net90));
 sg13g2_mux2_1 _25563_ (.A0(_09975_),
    .A1(\cpu.intr.r_timer_reload[8] ),
    .S(_06591_),
    .X(_02484_));
 sg13g2_nand2_1 _25564_ (.Y(_06606_),
    .A(\cpu.intr.r_timer_reload[9] ),
    .B(_06589_));
 sg13g2_o21ai_1 _25565_ (.B1(_06606_),
    .Y(_02485_),
    .A1(_12157_),
    .A2(net90));
 sg13g2_inv_1 _25566_ (.Y(_06607_),
    .A(_09662_));
 sg13g2_nand2b_1 _25567_ (.Y(_06608_),
    .B(_09700_),
    .A_N(_09657_));
 sg13g2_nor2_1 _25568_ (.A(_09671_),
    .B(_09659_),
    .Y(_06609_));
 sg13g2_nor4_2 _25569_ (.A(_11885_),
    .B(_11902_),
    .C(_09681_),
    .Y(_06610_),
    .D(_11883_));
 sg13g2_nor3_1 _25570_ (.A(_11903_),
    .B(_11886_),
    .C(_11901_),
    .Y(_06611_));
 sg13g2_nand3_1 _25571_ (.B(_06610_),
    .C(_06611_),
    .A(_06609_),
    .Y(_06612_));
 sg13g2_a21oi_1 _25572_ (.A1(_09163_),
    .A2(_06608_),
    .Y(_06613_),
    .B1(_06612_));
 sg13g2_buf_1 _25573_ (.A(_06613_),
    .X(_06614_));
 sg13g2_and2_1 _25574_ (.A(\cpu.qspi.r_read_delay[1][0] ),
    .B(_09693_),
    .X(_06615_));
 sg13g2_a221oi_1 _25575_ (.B2(\cpu.qspi.r_read_delay[0][0] ),
    .C1(_06615_),
    .B1(_09697_),
    .A1(\cpu.qspi.r_read_delay[2][0] ),
    .Y(_06616_),
    .A2(_09695_));
 sg13g2_nor2_1 _25576_ (.A(_09670_),
    .B(net1107),
    .Y(_06617_));
 sg13g2_nor2_1 _25577_ (.A(_09680_),
    .B(_09673_),
    .Y(_06618_));
 sg13g2_nand2_1 _25578_ (.Y(_06619_),
    .A(_06617_),
    .B(_06618_));
 sg13g2_a221oi_1 _25579_ (.B2(_06619_),
    .C1(_09678_),
    .B1(_00167_),
    .A1(_09705_),
    .Y(_06620_),
    .A2(_06607_));
 sg13g2_o21ai_1 _25580_ (.B1(_06620_),
    .Y(_06621_),
    .A1(_09724_),
    .A2(_06616_));
 sg13g2_nand2_1 _25581_ (.Y(_06622_),
    .A(net28),
    .B(_06621_));
 sg13g2_o21ai_1 _25582_ (.B1(_06622_),
    .Y(_02486_),
    .A1(_06607_),
    .A2(net28));
 sg13g2_inv_1 _25583_ (.Y(_06623_),
    .A(_09663_));
 sg13g2_and2_1 _25584_ (.A(\cpu.qspi.r_read_delay[2][1] ),
    .B(_09695_),
    .X(_06624_));
 sg13g2_a221oi_1 _25585_ (.B2(\cpu.qspi.r_read_delay[0][1] ),
    .C1(_06624_),
    .B1(_09697_),
    .A1(\cpu.qspi.r_read_delay[1][1] ),
    .Y(_06625_),
    .A2(_09693_));
 sg13g2_nor2_1 _25586_ (.A(_09705_),
    .B(_06619_),
    .Y(_06626_));
 sg13g2_xor2_1 _25587_ (.B(_09663_),
    .A(_09662_),
    .X(_06627_));
 sg13g2_nor2_1 _25588_ (.A(_06626_),
    .B(_06627_),
    .Y(_06628_));
 sg13g2_a21oi_1 _25589_ (.A1(_09724_),
    .A2(_06626_),
    .Y(_06629_),
    .B1(_06628_));
 sg13g2_o21ai_1 _25590_ (.B1(_06629_),
    .Y(_06630_),
    .A1(_09724_),
    .A2(_06625_));
 sg13g2_o21ai_1 _25591_ (.B1(_06614_),
    .Y(_06631_),
    .A1(_09678_),
    .A2(_06630_));
 sg13g2_o21ai_1 _25592_ (.B1(_06631_),
    .Y(_02487_),
    .A1(_06623_),
    .A2(net28));
 sg13g2_nor2_1 _25593_ (.A(_09662_),
    .B(_09663_),
    .Y(_06632_));
 sg13g2_xor2_1 _25594_ (.B(_06632_),
    .A(_00168_),
    .X(_06633_));
 sg13g2_and2_1 _25595_ (.A(_06617_),
    .B(_06618_),
    .X(_06634_));
 sg13g2_buf_1 _25596_ (.A(_06634_),
    .X(_06635_));
 sg13g2_o21ai_1 _25597_ (.B1(_09725_),
    .Y(_06636_),
    .A1(_09705_),
    .A2(_06635_));
 sg13g2_a22oi_1 _25598_ (.Y(_06637_),
    .B1(_06633_),
    .B2(_06636_),
    .A2(_06626_),
    .A1(_09723_));
 sg13g2_a22oi_1 _25599_ (.Y(_06638_),
    .B1(_09693_),
    .B2(\cpu.qspi.r_read_delay[1][2] ),
    .A2(_09695_),
    .A1(\cpu.qspi.r_read_delay[2][2] ));
 sg13g2_nand2_1 _25600_ (.Y(_06639_),
    .A(\cpu.qspi.r_read_delay[0][2] ),
    .B(_09697_));
 sg13g2_a21oi_1 _25601_ (.A1(_06638_),
    .A2(_06639_),
    .Y(_06640_),
    .B1(_09724_));
 sg13g2_nor3_1 _25602_ (.A(_09678_),
    .B(_06637_),
    .C(_06640_),
    .Y(_06641_));
 sg13g2_nor2_1 _25603_ (.A(_09664_),
    .B(_06614_),
    .Y(_06642_));
 sg13g2_a21oi_1 _25604_ (.A1(net28),
    .A2(_06641_),
    .Y(_02488_),
    .B1(_06642_));
 sg13g2_a21oi_1 _25605_ (.A1(_09725_),
    .A2(_06635_),
    .Y(_06643_),
    .B1(_09665_));
 sg13g2_nand2b_1 _25606_ (.Y(_06644_),
    .B(net28),
    .A_N(_06643_));
 sg13g2_nand2_1 _25607_ (.Y(_06645_),
    .A(_09725_),
    .B(_06635_));
 sg13g2_a22oi_1 _25608_ (.Y(_06646_),
    .B1(_09693_),
    .B2(\cpu.qspi.r_read_delay[1][3] ),
    .A2(_09695_),
    .A1(\cpu.qspi.r_read_delay[2][3] ));
 sg13g2_nand2_1 _25609_ (.Y(_06647_),
    .A(\cpu.qspi.r_read_delay[0][3] ),
    .B(_09697_));
 sg13g2_nand2_1 _25610_ (.Y(_06648_),
    .A(_06646_),
    .B(_06647_));
 sg13g2_a22oi_1 _25611_ (.Y(_06649_),
    .B1(_06648_),
    .B2(_09723_),
    .A2(_06645_),
    .A1(_09667_));
 sg13g2_nor2b_1 _25612_ (.A(_06649_),
    .B_N(net28),
    .Y(_06650_));
 sg13g2_a21o_1 _25613_ (.A2(_06644_),
    .A1(\cpu.qspi.r_count[3] ),
    .B1(_06650_),
    .X(_02489_));
 sg13g2_and2_1 _25614_ (.A(_09667_),
    .B(_06619_),
    .X(_06651_));
 sg13g2_nor3_1 _25615_ (.A(_09661_),
    .B(_09667_),
    .C(_06626_),
    .Y(_06652_));
 sg13g2_a21oi_1 _25616_ (.A1(_09661_),
    .A2(_06651_),
    .Y(_06653_),
    .B1(_06652_));
 sg13g2_nor2_1 _25617_ (.A(\cpu.qspi.r_count[4] ),
    .B(net28),
    .Y(_06654_));
 sg13g2_a21oi_1 _25618_ (.A1(net28),
    .A2(_06653_),
    .Y(_02490_),
    .B1(_06654_));
 sg13g2_nand2_1 _25619_ (.Y(_06655_),
    .A(_09782_),
    .B(_06227_));
 sg13g2_buf_1 _25620_ (.A(_06655_),
    .X(_06656_));
 sg13g2_nor3_1 _25621_ (.A(net410),
    .B(net575),
    .C(_06656_),
    .Y(_06657_));
 sg13g2_buf_1 _25622_ (.A(_06657_),
    .X(_06658_));
 sg13g2_nand2_1 _25623_ (.Y(_06659_),
    .A(net970),
    .B(_06658_));
 sg13g2_nand3_1 _25624_ (.B(_09782_),
    .C(_06227_),
    .A(_09039_),
    .Y(_06660_));
 sg13g2_buf_1 _25625_ (.A(_06660_),
    .X(_06661_));
 sg13g2_nand2_1 _25626_ (.Y(_06662_),
    .A(\cpu.qspi.r_read_delay[0][0] ),
    .B(_06661_));
 sg13g2_a21oi_1 _25627_ (.A1(_06659_),
    .A2(_06662_),
    .Y(_02501_),
    .B1(net606));
 sg13g2_nand2_1 _25628_ (.Y(_06663_),
    .A(net1018),
    .B(_06658_));
 sg13g2_nand2_1 _25629_ (.Y(_06664_),
    .A(\cpu.qspi.r_read_delay[0][1] ),
    .B(_06661_));
 sg13g2_a21oi_1 _25630_ (.A1(_06663_),
    .A2(_06664_),
    .Y(_02502_),
    .B1(net606));
 sg13g2_nand2_1 _25631_ (.Y(_06665_),
    .A(_09937_),
    .B(_06658_));
 sg13g2_nand2_1 _25632_ (.Y(_06666_),
    .A(\cpu.qspi.r_read_delay[0][2] ),
    .B(_06661_));
 sg13g2_nand3_1 _25633_ (.B(_06665_),
    .C(_06666_),
    .A(net687),
    .Y(_02503_));
 sg13g2_nand2_1 _25634_ (.Y(_06667_),
    .A(net1016),
    .B(_06658_));
 sg13g2_nand2_1 _25635_ (.Y(_06668_),
    .A(\cpu.qspi.r_read_delay[0][3] ),
    .B(_06661_));
 sg13g2_a21oi_1 _25636_ (.A1(_06667_),
    .A2(_06668_),
    .Y(_02504_),
    .B1(_09137_));
 sg13g2_nor2_1 _25637_ (.A(_09963_),
    .B(_06656_),
    .Y(_06669_));
 sg13g2_nand2_1 _25638_ (.Y(_06670_),
    .A(net970),
    .B(_06669_));
 sg13g2_or2_1 _25639_ (.X(_06671_),
    .B(_06656_),
    .A(_09963_));
 sg13g2_buf_1 _25640_ (.A(_06671_),
    .X(_06672_));
 sg13g2_nand2_1 _25641_ (.Y(_06673_),
    .A(\cpu.qspi.r_read_delay[1][0] ),
    .B(_06672_));
 sg13g2_buf_1 _25642_ (.A(_09136_),
    .X(_06674_));
 sg13g2_a21oi_1 _25643_ (.A1(_06670_),
    .A2(_06673_),
    .Y(_02505_),
    .B1(net556));
 sg13g2_nand2_1 _25644_ (.Y(_06675_),
    .A(net1018),
    .B(_06669_));
 sg13g2_nand2_1 _25645_ (.Y(_06676_),
    .A(\cpu.qspi.r_read_delay[1][1] ),
    .B(_06672_));
 sg13g2_a21oi_1 _25646_ (.A1(_06675_),
    .A2(_06676_),
    .Y(_02506_),
    .B1(net556));
 sg13g2_nand2_1 _25647_ (.Y(_06677_),
    .A(_09936_),
    .B(_06669_));
 sg13g2_nand2_1 _25648_ (.Y(_06678_),
    .A(\cpu.qspi.r_read_delay[1][2] ),
    .B(_06672_));
 sg13g2_nand3_1 _25649_ (.B(_06677_),
    .C(_06678_),
    .A(net687),
    .Y(_02507_));
 sg13g2_nand2_1 _25650_ (.Y(_06679_),
    .A(net1016),
    .B(_06669_));
 sg13g2_nand2_1 _25651_ (.Y(_06680_),
    .A(\cpu.qspi.r_read_delay[1][3] ),
    .B(_06672_));
 sg13g2_a21oi_1 _25652_ (.A1(_06679_),
    .A2(_06680_),
    .Y(_02508_),
    .B1(net556));
 sg13g2_nor2_1 _25653_ (.A(_04896_),
    .B(_06656_),
    .Y(_06681_));
 sg13g2_buf_1 _25654_ (.A(_06681_),
    .X(_06682_));
 sg13g2_nand2_1 _25655_ (.Y(_06683_),
    .A(net970),
    .B(_06682_));
 sg13g2_or2_1 _25656_ (.X(_06684_),
    .B(_06656_),
    .A(_04896_));
 sg13g2_buf_1 _25657_ (.A(_06684_),
    .X(_06685_));
 sg13g2_nand2_1 _25658_ (.Y(_06686_),
    .A(\cpu.qspi.r_read_delay[2][0] ),
    .B(_06685_));
 sg13g2_a21oi_1 _25659_ (.A1(_06683_),
    .A2(_06686_),
    .Y(_02509_),
    .B1(net556));
 sg13g2_nand2_1 _25660_ (.Y(_06687_),
    .A(_09929_),
    .B(_06682_));
 sg13g2_nand2_1 _25661_ (.Y(_06688_),
    .A(\cpu.qspi.r_read_delay[2][1] ),
    .B(_06685_));
 sg13g2_a21oi_1 _25662_ (.A1(_06687_),
    .A2(_06688_),
    .Y(_02510_),
    .B1(net556));
 sg13g2_nand2_1 _25663_ (.Y(_06689_),
    .A(net1017),
    .B(_06682_));
 sg13g2_nand2_1 _25664_ (.Y(_06690_),
    .A(\cpu.qspi.r_read_delay[2][2] ),
    .B(_06685_));
 sg13g2_nand3_1 _25665_ (.B(_06689_),
    .C(_06690_),
    .A(net687),
    .Y(_02511_));
 sg13g2_nand2_1 _25666_ (.Y(_06691_),
    .A(_09942_),
    .B(_06682_));
 sg13g2_nand2_1 _25667_ (.Y(_06692_),
    .A(\cpu.qspi.r_read_delay[2][3] ),
    .B(_06685_));
 sg13g2_a21oi_1 _25668_ (.A1(_06691_),
    .A2(_06692_),
    .Y(_02512_),
    .B1(net556));
 sg13g2_buf_1 _25669_ (.A(_09686_),
    .X(_06693_));
 sg13g2_buf_1 _25670_ (.A(net882),
    .X(_06694_));
 sg13g2_buf_1 _25671_ (.A(_09653_),
    .X(_06695_));
 sg13g2_mux2_1 _25672_ (.A0(net432),
    .A1(_09233_),
    .S(net129),
    .X(_06696_));
 sg13g2_nand2_1 _25673_ (.Y(_06697_),
    .A(net700),
    .B(_06696_));
 sg13g2_o21ai_1 _25674_ (.B1(_06697_),
    .Y(_06698_),
    .A1(net701),
    .A2(_08447_));
 sg13g2_mux2_1 _25675_ (.A0(_09502_),
    .A1(_09509_),
    .S(net129),
    .X(_06699_));
 sg13g2_nand2_1 _25676_ (.Y(_06700_),
    .A(net701),
    .B(_06699_));
 sg13g2_o21ai_1 _25677_ (.B1(_06700_),
    .Y(_06701_),
    .A1(net701),
    .A2(_08285_));
 sg13g2_buf_1 _25678_ (.A(_09653_),
    .X(_06702_));
 sg13g2_mux2_1 _25679_ (.A0(_00213_),
    .A1(_09531_),
    .S(net128),
    .X(_06703_));
 sg13g2_nand2_1 _25680_ (.Y(_06704_),
    .A(_09164_),
    .B(_10643_));
 sg13g2_o21ai_1 _25681_ (.B1(_06704_),
    .Y(_06705_),
    .A1(net1030),
    .A2(_06703_));
 sg13g2_nand2_1 _25682_ (.Y(_06706_),
    .A(_11902_),
    .B(_06705_));
 sg13g2_a21oi_1 _25683_ (.A1(_09681_),
    .A2(_11882_),
    .Y(_06707_),
    .B1(_11885_));
 sg13g2_buf_1 _25684_ (.A(_11991_),
    .X(_06708_));
 sg13g2_nor2b_1 _25685_ (.A(net1085),
    .B_N(_11990_),
    .Y(_06709_));
 sg13g2_a22oi_1 _25686_ (.Y(_06710_),
    .B1(_04874_),
    .B2(_12010_),
    .A2(_04843_),
    .A1(_11990_));
 sg13g2_nor2_1 _25687_ (.A(_12013_),
    .B(_06710_),
    .Y(_06711_));
 sg13g2_a21oi_1 _25688_ (.A1(_05514_),
    .A2(_06709_),
    .Y(_06712_),
    .B1(_06711_));
 sg13g2_nor2b_1 _25689_ (.A(_12123_),
    .B_N(_12010_),
    .Y(_06713_));
 sg13g2_nor2_1 _25690_ (.A(_11990_),
    .B(_06713_),
    .Y(_06714_));
 sg13g2_a22oi_1 _25691_ (.Y(_06715_),
    .B1(_05194_),
    .B2(_12010_),
    .A2(_05187_),
    .A1(_11990_));
 sg13g2_a221oi_1 _25692_ (.B2(_11990_),
    .C1(_12013_),
    .B1(_04866_),
    .A1(_12010_),
    .Y(_06716_),
    .A2(_04859_));
 sg13g2_a21oi_1 _25693_ (.A1(_12013_),
    .A2(_06715_),
    .Y(_06717_),
    .B1(_06716_));
 sg13g2_a22oi_1 _25694_ (.Y(_06718_),
    .B1(_06717_),
    .B2(net925),
    .A2(_06714_),
    .A1(_05507_));
 sg13g2_o21ai_1 _25695_ (.B1(_06718_),
    .Y(_06719_),
    .A1(_06708_),
    .A2(_06712_));
 sg13g2_nand2_1 _25696_ (.Y(_06720_),
    .A(_09673_),
    .B(_06719_));
 sg13g2_buf_1 _25697_ (.A(\cpu.qspi.r_state[0] ),
    .X(_06721_));
 sg13g2_nand2_1 _25698_ (.Y(_06722_),
    .A(net1046),
    .B(net1030));
 sg13g2_o21ai_1 _25699_ (.B1(_06722_),
    .Y(_06723_),
    .A1(net1030),
    .A2(net645));
 sg13g2_nand2_1 _25700_ (.Y(_06724_),
    .A(_06611_),
    .B(_06618_));
 sg13g2_nor2_1 _25701_ (.A(_09678_),
    .B(_06724_),
    .Y(_06725_));
 sg13g2_nor2b_1 _25702_ (.A(net1107),
    .B_N(_06610_),
    .Y(_06726_));
 sg13g2_and3_1 _25703_ (.X(_06727_),
    .A(_09720_),
    .B(_06725_),
    .C(_06726_));
 sg13g2_buf_1 _25704_ (.A(_06727_),
    .X(_06728_));
 sg13g2_a221oi_1 _25705_ (.B2(_11901_),
    .C1(_06728_),
    .B1(_06723_),
    .A1(_09707_),
    .Y(_06729_),
    .A2(_06721_));
 sg13g2_nand4_1 _25706_ (.B(_06707_),
    .C(_06720_),
    .A(_06706_),
    .Y(_06730_),
    .D(_06729_));
 sg13g2_a221oi_1 _25707_ (.B2(_11886_),
    .C1(_06730_),
    .B1(_06701_),
    .A1(_11903_),
    .Y(_06731_),
    .A2(_06698_));
 sg13g2_nand2_1 _25708_ (.Y(_06732_),
    .A(_06607_),
    .B(_09663_));
 sg13g2_mux2_1 _25709_ (.A0(_06732_),
    .A1(_09663_),
    .S(_09677_),
    .X(_06733_));
 sg13g2_nand2_1 _25710_ (.Y(_06734_),
    .A(net1107),
    .B(_09660_));
 sg13g2_a21o_1 _25711_ (.A2(_06734_),
    .A1(_00167_),
    .B1(_09663_),
    .X(_06735_));
 sg13g2_o21ai_1 _25712_ (.B1(_06735_),
    .Y(_06736_),
    .A1(net1107),
    .A2(_06733_));
 sg13g2_nand3_1 _25713_ (.B(_09662_),
    .C(_09660_),
    .A(net1107),
    .Y(_06737_));
 sg13g2_o21ai_1 _25714_ (.B1(_06737_),
    .Y(_06738_),
    .A1(_09660_),
    .A2(_06732_));
 sg13g2_nand2b_1 _25715_ (.Y(_06739_),
    .B(_09677_),
    .A_N(_09663_));
 sg13g2_a21oi_1 _25716_ (.A1(_06732_),
    .A2(_06739_),
    .Y(_06740_),
    .B1(net1107));
 sg13g2_nor3_1 _25717_ (.A(_09664_),
    .B(_06738_),
    .C(_06740_),
    .Y(_06741_));
 sg13g2_a21o_1 _25718_ (.A2(_06736_),
    .A1(_09664_),
    .B1(_06741_),
    .X(_06742_));
 sg13g2_o21ai_1 _25719_ (.B1(_06742_),
    .Y(_06743_),
    .A1(_09680_),
    .A2(net1107));
 sg13g2_xnor2_1 _25720_ (.Y(_06744_),
    .A(_09677_),
    .B(_09700_));
 sg13g2_a22oi_1 _25721_ (.Y(_06745_),
    .B1(_06744_),
    .B2(_06728_),
    .A2(_06743_),
    .A1(_06731_));
 sg13g2_and2_1 _25722_ (.A(\cpu.qspi.r_mask[1] ),
    .B(_09693_),
    .X(_06746_));
 sg13g2_a221oi_1 _25723_ (.B2(\cpu.qspi.r_mask[0] ),
    .C1(_06746_),
    .B1(_09697_),
    .A1(\cpu.qspi.r_mask[2] ),
    .Y(_06747_),
    .A2(_09695_));
 sg13g2_nor3_2 _25724_ (.A(_09670_),
    .B(_09671_),
    .C(_09659_),
    .Y(_06748_));
 sg13g2_nor2_1 _25725_ (.A(_09723_),
    .B(_09705_),
    .Y(_06749_));
 sg13g2_nand3_1 _25726_ (.B(_06748_),
    .C(_06749_),
    .A(_09658_),
    .Y(_06750_));
 sg13g2_a21oi_1 _25727_ (.A1(_11885_),
    .A2(_06747_),
    .Y(_06751_),
    .B1(_06750_));
 sg13g2_buf_2 _25728_ (.A(_06751_),
    .X(_06752_));
 sg13g2_mux2_1 _25729_ (.A0(net11),
    .A1(_06745_),
    .S(_06752_),
    .X(_02517_));
 sg13g2_mux4_1 _25730_ (.S0(_12013_),
    .A0(_05289_),
    .A1(_05582_),
    .A2(_05307_),
    .A3(_05216_),
    .S1(net925),
    .X(_06753_));
 sg13g2_mux2_1 _25731_ (.A0(_05222_),
    .A1(_05298_),
    .S(net1085),
    .X(_06754_));
 sg13g2_a22oi_1 _25732_ (.Y(_06755_),
    .B1(_06754_),
    .B2(_06708_),
    .A2(_05283_),
    .A1(_12014_));
 sg13g2_nor2b_1 _25733_ (.A(_06755_),
    .B_N(net991),
    .Y(_06756_));
 sg13g2_a221oi_1 _25734_ (.B2(net987),
    .C1(_06756_),
    .B1(_06753_),
    .A1(_05591_),
    .Y(_06757_),
    .A2(_06714_));
 sg13g2_nand2b_1 _25735_ (.Y(_06758_),
    .B(_09673_),
    .A_N(_06757_));
 sg13g2_nand2_1 _25736_ (.Y(_06759_),
    .A(_09555_),
    .B(net128));
 sg13g2_o21ai_1 _25737_ (.B1(_06759_),
    .Y(_06760_),
    .A1(_05369_),
    .A2(_06695_));
 sg13g2_nand2_1 _25738_ (.Y(_06761_),
    .A(net882),
    .B(_06760_));
 sg13g2_o21ai_1 _25739_ (.B1(_06761_),
    .Y(_06762_),
    .A1(net700),
    .A2(_10469_));
 sg13g2_buf_1 _25740_ (.A(net1030),
    .X(_06763_));
 sg13g2_mux2_1 _25741_ (.A0(_00215_),
    .A1(_09522_),
    .S(net129),
    .X(_06764_));
 sg13g2_nand2_1 _25742_ (.Y(_06765_),
    .A(net801),
    .B(_10874_));
 sg13g2_o21ai_1 _25743_ (.B1(_06765_),
    .Y(_06766_),
    .A1(net801),
    .A2(_06764_));
 sg13g2_a22oi_1 _25744_ (.Y(_06767_),
    .B1(_06766_),
    .B2(_11902_),
    .A2(_06762_),
    .A1(_11901_));
 sg13g2_mux2_1 _25745_ (.A0(net428),
    .A1(_09372_),
    .S(net128),
    .X(_06768_));
 sg13g2_nand2_1 _25746_ (.Y(_06769_),
    .A(net882),
    .B(_06768_));
 sg13g2_o21ai_1 _25747_ (.B1(_06769_),
    .Y(_06770_),
    .A1(net700),
    .A2(_08557_));
 sg13g2_mux2_1 _25748_ (.A0(_09486_),
    .A1(_09468_),
    .S(net128),
    .X(_06771_));
 sg13g2_nand2_1 _25749_ (.Y(_06772_),
    .A(_06694_),
    .B(_06771_));
 sg13g2_o21ai_1 _25750_ (.B1(_06772_),
    .Y(_06773_),
    .A1(net701),
    .A2(_08356_));
 sg13g2_a22oi_1 _25751_ (.Y(_06774_),
    .B1(_06773_),
    .B2(_11886_),
    .A2(_06770_),
    .A1(_11903_));
 sg13g2_nand4_1 _25752_ (.B(_06758_),
    .C(_06767_),
    .A(_06707_),
    .Y(_06775_),
    .D(_06774_));
 sg13g2_a21oi_1 _25753_ (.A1(_09701_),
    .A2(_06728_),
    .Y(_06776_),
    .B1(_06775_));
 sg13g2_nor2_1 _25754_ (.A(net12),
    .B(_06752_),
    .Y(_06777_));
 sg13g2_a21oi_1 _25755_ (.A1(_06752_),
    .A2(_06776_),
    .Y(_02518_),
    .B1(_06777_));
 sg13g2_inv_1 _25756_ (.Y(_06778_),
    .A(net13));
 sg13g2_nand2_1 _25757_ (.Y(_06779_),
    .A(net801),
    .B(_00272_));
 sg13g2_mux2_1 _25758_ (.A0(_00217_),
    .A1(_09540_),
    .S(net129),
    .X(_06780_));
 sg13g2_nand2_1 _25759_ (.Y(_06781_),
    .A(_06693_),
    .B(_06780_));
 sg13g2_nand3_1 _25760_ (.B(_06779_),
    .C(_06781_),
    .A(_11902_),
    .Y(_06782_));
 sg13g2_nand2_1 _25761_ (.Y(_06783_),
    .A(net691),
    .B(net1030));
 sg13g2_nand2_1 _25762_ (.Y(_06784_),
    .A(net882),
    .B(net456));
 sg13g2_a21oi_1 _25763_ (.A1(_06783_),
    .A2(_06784_),
    .Y(_06785_),
    .B1(_00169_));
 sg13g2_nand2_1 _25764_ (.Y(_06786_),
    .A(net925),
    .B(_05046_));
 sg13g2_o21ai_1 _25765_ (.B1(_06786_),
    .Y(_06787_),
    .A1(net925),
    .A2(_05421_));
 sg13g2_nand3_1 _25766_ (.B(net991),
    .C(_06787_),
    .A(_12012_),
    .Y(_06788_));
 sg13g2_mux4_1 _25767_ (.S0(net1085),
    .A0(_05651_),
    .A1(_05412_),
    .A2(_05239_),
    .A3(_05039_),
    .S1(net925),
    .X(_06789_));
 sg13g2_nand3_1 _25768_ (.B(_12010_),
    .C(_05248_),
    .A(_11991_),
    .Y(_06790_));
 sg13g2_o21ai_1 _25769_ (.B1(_06790_),
    .Y(_06791_),
    .A1(net925),
    .A2(net987));
 sg13g2_nor2_1 _25770_ (.A(net987),
    .B(net991),
    .Y(_06792_));
 sg13g2_a221oi_1 _25771_ (.B2(_12013_),
    .C1(_06792_),
    .B1(_06791_),
    .A1(net987),
    .Y(_06793_),
    .A2(_06789_));
 sg13g2_a221oi_1 _25772_ (.B2(_06793_),
    .C1(_11887_),
    .B1(_06788_),
    .A1(_05658_),
    .Y(_06794_),
    .A2(_06714_));
 sg13g2_nor4_1 _25773_ (.A(_11885_),
    .B(_06728_),
    .C(_06785_),
    .D(_06794_),
    .Y(_06795_));
 sg13g2_mux2_1 _25774_ (.A0(net431),
    .A1(_09277_),
    .S(net128),
    .X(_06796_));
 sg13g2_nand2_1 _25775_ (.Y(_06797_),
    .A(net700),
    .B(_06796_));
 sg13g2_o21ai_1 _25776_ (.B1(_06797_),
    .Y(_06798_),
    .A1(net701),
    .A2(_08577_));
 sg13g2_nand2_1 _25777_ (.Y(_06799_),
    .A(_11903_),
    .B(_06798_));
 sg13g2_mux2_1 _25778_ (.A0(net429),
    .A1(_09346_),
    .S(net128),
    .X(_06800_));
 sg13g2_nand2_1 _25779_ (.Y(_06801_),
    .A(net700),
    .B(_06800_));
 sg13g2_o21ai_1 _25780_ (.B1(_06801_),
    .Y(_06802_),
    .A1(_06693_),
    .A2(_08473_));
 sg13g2_nor2_1 _25781_ (.A(_00209_),
    .B(net129),
    .Y(_06803_));
 sg13g2_and2_1 _25782_ (.A(_09567_),
    .B(_06702_),
    .X(_06804_));
 sg13g2_o21ai_1 _25783_ (.B1(_06694_),
    .Y(_06805_),
    .A1(_06803_),
    .A2(_06804_));
 sg13g2_o21ai_1 _25784_ (.B1(_06805_),
    .Y(_06806_),
    .A1(net701),
    .A2(_10710_));
 sg13g2_a22oi_1 _25785_ (.Y(_06807_),
    .B1(_06806_),
    .B2(_11901_),
    .A2(_06802_),
    .A1(_11886_));
 sg13g2_nand4_1 _25786_ (.B(_06795_),
    .C(_06799_),
    .A(_06782_),
    .Y(_06808_),
    .D(_06807_));
 sg13g2_o21ai_1 _25787_ (.B1(_06728_),
    .Y(_06809_),
    .A1(_09677_),
    .A2(_09700_));
 sg13g2_nand3_1 _25788_ (.B(_06808_),
    .C(_06809_),
    .A(_06752_),
    .Y(_06810_));
 sg13g2_o21ai_1 _25789_ (.B1(_06810_),
    .Y(_02519_),
    .A1(_06778_),
    .A2(_06752_));
 sg13g2_inv_1 _25790_ (.Y(_06811_),
    .A(net14));
 sg13g2_mux2_1 _25791_ (.A0(_00219_),
    .A1(_09592_),
    .S(net129),
    .X(_06812_));
 sg13g2_nand2_1 _25792_ (.Y(_06813_),
    .A(net801),
    .B(_10882_));
 sg13g2_o21ai_1 _25793_ (.B1(_06813_),
    .Y(_06814_),
    .A1(net801),
    .A2(_06812_));
 sg13g2_mux2_1 _25794_ (.A0(net375),
    .A1(_09429_),
    .S(net128),
    .X(_06815_));
 sg13g2_a21oi_1 _25795_ (.A1(net700),
    .A2(_06815_),
    .Y(_06816_),
    .B1(_09688_));
 sg13g2_nand2_1 _25796_ (.Y(_06817_),
    .A(_09684_),
    .B(_11883_));
 sg13g2_nor3_1 _25797_ (.A(_09683_),
    .B(_06816_),
    .C(_06817_),
    .Y(_06818_));
 sg13g2_a21oi_1 _25798_ (.A1(_11902_),
    .A2(_06814_),
    .Y(_06819_),
    .B1(_06818_));
 sg13g2_nand2_1 _25799_ (.Y(_06820_),
    .A(_09645_),
    .B(net129));
 sg13g2_o21ai_1 _25800_ (.B1(_06820_),
    .Y(_06821_),
    .A1(_09638_),
    .A2(net129));
 sg13g2_or2_1 _25801_ (.X(_06822_),
    .B(_08494_),
    .A(net882));
 sg13g2_o21ai_1 _25802_ (.B1(_06822_),
    .Y(_06823_),
    .A1(net801),
    .A2(_06821_));
 sg13g2_a22oi_1 _25803_ (.Y(_06824_),
    .B1(_05476_),
    .B2(net987),
    .A2(_05484_),
    .A1(net991));
 sg13g2_a221oi_1 _25804_ (.B2(_12012_),
    .C1(net925),
    .B1(_06824_),
    .A1(_05084_),
    .Y(_06825_),
    .A2(_06709_));
 sg13g2_mux2_1 _25805_ (.A0(_05070_),
    .A1(_05170_),
    .S(net1085),
    .X(_06826_));
 sg13g2_mux2_1 _25806_ (.A0(_05056_),
    .A1(_05164_),
    .S(net1085),
    .X(_06827_));
 sg13g2_a22oi_1 _25807_ (.Y(_06828_),
    .B1(_06827_),
    .B2(net987),
    .A2(_06826_),
    .A1(_12011_));
 sg13g2_nor2b_1 _25808_ (.A(_06828_),
    .B_N(net925),
    .Y(_06829_));
 sg13g2_nor3_1 _25809_ (.A(_06792_),
    .B(_06825_),
    .C(_06829_),
    .Y(_06830_));
 sg13g2_a21o_1 _25810_ (.A2(_06714_),
    .A1(_05080_),
    .B1(_11887_),
    .X(_06831_));
 sg13g2_nand2_1 _25811_ (.Y(_06832_),
    .A(net692),
    .B(net1030));
 sg13g2_nand2_1 _25812_ (.Y(_06833_),
    .A(net882),
    .B(net464));
 sg13g2_a21oi_1 _25813_ (.A1(_06832_),
    .A2(_06833_),
    .Y(_06834_),
    .B1(_00169_));
 sg13g2_nor4_1 _25814_ (.A(_11885_),
    .B(_09681_),
    .C(_06728_),
    .D(_06834_),
    .Y(_06835_));
 sg13g2_o21ai_1 _25815_ (.B1(_06835_),
    .Y(_06836_),
    .A1(_06830_),
    .A2(_06831_));
 sg13g2_a21oi_1 _25816_ (.A1(_11903_),
    .A2(_06823_),
    .Y(_06837_),
    .B1(_06836_));
 sg13g2_nand2_1 _25817_ (.Y(_06838_),
    .A(_09580_),
    .B(net128));
 sg13g2_o21ai_1 _25818_ (.B1(_06838_),
    .Y(_06839_),
    .A1(_00211_),
    .A2(_06695_));
 sg13g2_nand2_1 _25819_ (.Y(_06840_),
    .A(net700),
    .B(_06839_));
 sg13g2_o21ai_1 _25820_ (.B1(_06840_),
    .Y(_06841_),
    .A1(net701),
    .A2(_10740_));
 sg13g2_mux2_1 _25821_ (.A0(net427),
    .A1(_09384_),
    .S(_06702_),
    .X(_06842_));
 sg13g2_nand2_1 _25822_ (.Y(_06843_),
    .A(net700),
    .B(_06842_));
 sg13g2_o21ai_1 _25823_ (.B1(_06843_),
    .Y(_06844_),
    .A1(net701),
    .A2(_08515_));
 sg13g2_a22oi_1 _25824_ (.Y(_06845_),
    .B1(_06844_),
    .B2(_11886_),
    .A2(_06841_),
    .A1(_11901_));
 sg13g2_nand3_1 _25825_ (.B(_06837_),
    .C(_06845_),
    .A(_06819_),
    .Y(_06846_));
 sg13g2_nand3_1 _25826_ (.B(_06809_),
    .C(_06846_),
    .A(_06752_),
    .Y(_06847_));
 sg13g2_o21ai_1 _25827_ (.B1(_06847_),
    .Y(_02520_),
    .A1(_06811_),
    .A2(_06752_));
 sg13g2_nand2_1 _25828_ (.Y(_06848_),
    .A(net637),
    .B(net645));
 sg13g2_nor2_1 _25829_ (.A(_09031_),
    .B(_09048_),
    .Y(_06849_));
 sg13g2_nand3_1 _25830_ (.B(net644),
    .C(_06849_),
    .A(net848),
    .Y(_06850_));
 sg13g2_buf_1 _25831_ (.A(_06850_),
    .X(_06851_));
 sg13g2_nor2_1 _25832_ (.A(_06848_),
    .B(_06851_),
    .Y(_06852_));
 sg13g2_buf_4 _25833_ (.X(_06853_),
    .A(_06852_));
 sg13g2_mux2_1 _25834_ (.A0(\cpu.spi.r_clk_count[0][0] ),
    .A1(net877),
    .S(_06853_),
    .X(_02525_));
 sg13g2_mux2_1 _25835_ (.A0(\cpu.spi.r_clk_count[0][1] ),
    .A1(net855),
    .S(_06853_),
    .X(_02526_));
 sg13g2_mux2_1 _25836_ (.A0(\cpu.spi.r_clk_count[0][2] ),
    .A1(net876),
    .S(_06853_),
    .X(_02527_));
 sg13g2_mux2_1 _25837_ (.A0(\cpu.spi.r_clk_count[0][3] ),
    .A1(net1016),
    .S(_06853_),
    .X(_02528_));
 sg13g2_mux2_1 _25838_ (.A0(\cpu.spi.r_clk_count[0][4] ),
    .A1(net1022),
    .S(_06853_),
    .X(_02529_));
 sg13g2_mux2_1 _25839_ (.A0(\cpu.spi.r_clk_count[0][5] ),
    .A1(net986),
    .S(_06853_),
    .X(_02530_));
 sg13g2_mux2_1 _25840_ (.A0(\cpu.spi.r_clk_count[0][6] ),
    .A1(net974),
    .S(_06853_),
    .X(_02531_));
 sg13g2_mux2_1 _25841_ (.A0(\cpu.spi.r_clk_count[0][7] ),
    .A1(net1019),
    .S(_06853_),
    .X(_02532_));
 sg13g2_nor2_1 _25842_ (.A(_04913_),
    .B(_06851_),
    .Y(_06854_));
 sg13g2_buf_4 _25843_ (.X(_06855_),
    .A(_06854_));
 sg13g2_mux2_1 _25844_ (.A0(\cpu.spi.r_clk_count[1][0] ),
    .A1(net877),
    .S(_06855_),
    .X(_02533_));
 sg13g2_mux2_1 _25845_ (.A0(\cpu.spi.r_clk_count[1][1] ),
    .A1(net855),
    .S(_06855_),
    .X(_02534_));
 sg13g2_mux2_1 _25846_ (.A0(\cpu.spi.r_clk_count[1][2] ),
    .A1(net876),
    .S(_06855_),
    .X(_02535_));
 sg13g2_mux2_1 _25847_ (.A0(\cpu.spi.r_clk_count[1][3] ),
    .A1(net1016),
    .S(_06855_),
    .X(_02536_));
 sg13g2_mux2_1 _25848_ (.A0(\cpu.spi.r_clk_count[1][4] ),
    .A1(net1022),
    .S(_06855_),
    .X(_02537_));
 sg13g2_mux2_1 _25849_ (.A0(\cpu.spi.r_clk_count[1][5] ),
    .A1(net986),
    .S(_06855_),
    .X(_02538_));
 sg13g2_mux2_1 _25850_ (.A0(\cpu.spi.r_clk_count[1][6] ),
    .A1(_12136_),
    .S(_06855_),
    .X(_02539_));
 sg13g2_mux2_1 _25851_ (.A0(\cpu.spi.r_clk_count[1][7] ),
    .A1(net1019),
    .S(_06855_),
    .X(_02540_));
 sg13g2_nor3_1 _25852_ (.A(_09031_),
    .B(_09048_),
    .C(_06848_),
    .Y(_06856_));
 sg13g2_nor2_1 _25853_ (.A(net848),
    .B(net410),
    .Y(_06857_));
 sg13g2_nand2_1 _25854_ (.Y(_06858_),
    .A(_06856_),
    .B(_06857_));
 sg13g2_buf_1 _25855_ (.A(_06858_),
    .X(_06859_));
 sg13g2_mux2_1 _25856_ (.A0(net880),
    .A1(_04957_),
    .S(net88),
    .X(_02541_));
 sg13g2_mux2_1 _25857_ (.A0(net829),
    .A1(_05328_),
    .S(net88),
    .X(_02542_));
 sg13g2_nand2_1 _25858_ (.Y(_06860_),
    .A(_05379_),
    .B(net88));
 sg13g2_o21ai_1 _25859_ (.B1(_06860_),
    .Y(_02543_),
    .A1(net878),
    .A2(net88));
 sg13g2_nand2_1 _25860_ (.Y(_06861_),
    .A(_05458_),
    .B(net88));
 sg13g2_o21ai_1 _25861_ (.B1(_06861_),
    .Y(_02544_),
    .A1(net854),
    .A2(net88));
 sg13g2_nand2_1 _25862_ (.Y(_06862_),
    .A(_05522_),
    .B(_06858_));
 sg13g2_o21ai_1 _25863_ (.B1(_06862_),
    .Y(_02545_),
    .A1(net853),
    .A2(net88));
 sg13g2_mux2_1 _25864_ (.A0(net849),
    .A1(_05620_),
    .S(_06859_),
    .X(_02546_));
 sg13g2_mux2_1 _25865_ (.A0(net875),
    .A1(_05678_),
    .S(net88),
    .X(_02547_));
 sg13g2_nand2_1 _25866_ (.Y(_06863_),
    .A(_05123_),
    .B(_06858_));
 sg13g2_o21ai_1 _25867_ (.B1(_06863_),
    .Y(_02548_),
    .A1(net852),
    .A2(_06859_));
 sg13g2_buf_1 _25868_ (.A(_00204_),
    .X(_06864_));
 sg13g2_nor4_1 _25869_ (.A(\cpu.spi.r_state[5] ),
    .B(net1110),
    .C(_09127_),
    .D(_11906_),
    .Y(_06865_));
 sg13g2_buf_1 _25870_ (.A(_06865_),
    .X(_06866_));
 sg13g2_nand2_1 _25871_ (.Y(_06867_),
    .A(_06864_),
    .B(net623));
 sg13g2_buf_2 _25872_ (.A(_06867_),
    .X(_06868_));
 sg13g2_buf_1 _25873_ (.A(_06868_),
    .X(_06869_));
 sg13g2_nor2_1 _25874_ (.A(net728),
    .B(_04957_),
    .Y(_06870_));
 sg13g2_a21oi_1 _25875_ (.A1(net728),
    .A2(_00281_),
    .Y(_06871_),
    .B1(_06870_));
 sg13g2_buf_1 _25876_ (.A(net995),
    .X(_06872_));
 sg13g2_mux2_1 _25877_ (.A0(_00281_),
    .A1(_00280_),
    .S(net800),
    .X(_06873_));
 sg13g2_nor2_1 _25878_ (.A(net859),
    .B(_06873_),
    .Y(_06874_));
 sg13g2_a21oi_1 _25879_ (.A1(net859),
    .A2(_06871_),
    .Y(_06875_),
    .B1(_06874_));
 sg13g2_nand2_1 _25880_ (.Y(_06876_),
    .A(net304),
    .B(_06875_));
 sg13g2_nor2_1 _25881_ (.A(_09085_),
    .B(_06866_),
    .Y(_06877_));
 sg13g2_nand2b_1 _25882_ (.Y(_06878_),
    .B(_09054_),
    .A_N(_09085_));
 sg13g2_o21ai_1 _25883_ (.B1(_06878_),
    .Y(_06879_),
    .A1(_09054_),
    .A2(_06875_));
 sg13g2_a22oi_1 _25884_ (.Y(_06880_),
    .B1(_06879_),
    .B2(net856),
    .A2(_06877_),
    .A1(_06876_));
 sg13g2_nand2b_1 _25885_ (.Y(_06881_),
    .B(_11948_),
    .A_N(\cpu.spi.r_clk_count[0][0] ));
 sg13g2_o21ai_1 _25886_ (.B1(_06881_),
    .Y(_06882_),
    .A1(net501),
    .A2(_04957_));
 sg13g2_mux2_1 _25887_ (.A0(\cpu.spi.r_clk_count[0][0] ),
    .A1(\cpu.spi.r_clk_count[1][0] ),
    .S(net585),
    .X(_06883_));
 sg13g2_nor2_1 _25888_ (.A(_11946_),
    .B(_06883_),
    .Y(_06884_));
 sg13g2_a21oi_1 _25889_ (.A1(_11946_),
    .A2(_06882_),
    .Y(_06885_),
    .B1(_06884_));
 sg13g2_nor2_1 _25890_ (.A(_06885_),
    .B(_06869_),
    .Y(_06886_));
 sg13g2_a21oi_1 _25891_ (.A1(net439),
    .A2(_06880_),
    .Y(_06887_),
    .B1(_06886_));
 sg13g2_inv_1 _25892_ (.Y(_06888_),
    .A(_09132_));
 sg13g2_and2_1 _25893_ (.A(_06888_),
    .B(net623),
    .X(_06889_));
 sg13g2_nor2_1 _25894_ (.A(_06864_),
    .B(net379),
    .Y(_06890_));
 sg13g2_nor2_1 _25895_ (.A(_09043_),
    .B(_09094_),
    .Y(_06891_));
 sg13g2_o21ai_1 _25896_ (.B1(_09162_),
    .Y(_06892_),
    .A1(_09056_),
    .A2(_06891_));
 sg13g2_a221oi_1 _25897_ (.B2(_09108_),
    .C1(_06892_),
    .B1(_06890_),
    .A1(_06864_),
    .Y(_06893_),
    .A2(_06889_));
 sg13g2_buf_1 _25898_ (.A(_06893_),
    .X(_06894_));
 sg13g2_mux2_1 _25899_ (.A0(_09085_),
    .A1(_06887_),
    .S(_06894_),
    .X(_02549_));
 sg13g2_nand2b_1 _25900_ (.Y(_06895_),
    .B(_11947_),
    .A_N(\cpu.spi.r_clk_count[0][1] ));
 sg13g2_o21ai_1 _25901_ (.B1(_06895_),
    .Y(_06896_),
    .A1(_11947_),
    .A2(_05328_));
 sg13g2_mux2_1 _25902_ (.A0(\cpu.spi.r_clk_count[0][1] ),
    .A1(\cpu.spi.r_clk_count[1][1] ),
    .S(net585),
    .X(_06897_));
 sg13g2_nor2_1 _25903_ (.A(net857),
    .B(_06897_),
    .Y(_06898_));
 sg13g2_a21oi_1 _25904_ (.A1(net857),
    .A2(_06896_),
    .Y(_06899_),
    .B1(_06898_));
 sg13g2_o21ai_1 _25905_ (.B1(_09085_),
    .Y(_06900_),
    .A1(_06868_),
    .A2(_06899_));
 sg13g2_o21ai_1 _25906_ (.B1(net31),
    .Y(_06901_),
    .A1(_09056_),
    .A2(_06900_));
 sg13g2_nor2_1 _25907_ (.A(_06868_),
    .B(_06899_),
    .Y(_06902_));
 sg13g2_mux2_1 _25908_ (.A0(_00286_),
    .A1(_00285_),
    .S(_06872_),
    .X(_06903_));
 sg13g2_nor2_1 _25909_ (.A(_11918_),
    .B(_05328_),
    .Y(_06904_));
 sg13g2_a21oi_1 _25910_ (.A1(net800),
    .A2(_00286_),
    .Y(_06905_),
    .B1(_06904_));
 sg13g2_nand2_1 _25911_ (.Y(_06906_),
    .A(net996),
    .B(_06905_));
 sg13g2_o21ai_1 _25912_ (.B1(_06906_),
    .Y(_06907_),
    .A1(net859),
    .A2(_06903_));
 sg13g2_nand2_1 _25913_ (.Y(_06908_),
    .A(_09108_),
    .B(_06907_));
 sg13g2_o21ai_1 _25914_ (.B1(_06908_),
    .Y(_06909_),
    .A1(net103),
    .A2(_09087_));
 sg13g2_nand2_1 _25915_ (.Y(_06910_),
    .A(_09085_),
    .B(\cpu.spi.r_count[1] ));
 sg13g2_a21oi_1 _25916_ (.A1(_09087_),
    .A2(_06910_),
    .Y(_06911_),
    .B1(_06866_));
 sg13g2_o21ai_1 _25917_ (.B1(_06911_),
    .Y(_06912_),
    .A1(net378),
    .A2(_06907_));
 sg13g2_nand2_1 _25918_ (.Y(_06913_),
    .A(_06868_),
    .B(_06912_));
 sg13g2_a21oi_1 _25919_ (.A1(_09098_),
    .A2(_06909_),
    .Y(_06914_),
    .B1(_06913_));
 sg13g2_nor2_1 _25920_ (.A(_06902_),
    .B(_06914_),
    .Y(_06915_));
 sg13g2_a22oi_1 _25921_ (.Y(_06916_),
    .B1(_06915_),
    .B2(net31),
    .A2(_06901_),
    .A1(\cpu.spi.r_count[1] ));
 sg13g2_inv_1 _25922_ (.Y(_02550_),
    .A(_06916_));
 sg13g2_nor2_1 _25923_ (.A(net800),
    .B(_05379_),
    .Y(_06917_));
 sg13g2_a21oi_1 _25924_ (.A1(net728),
    .A2(_00095_),
    .Y(_06918_),
    .B1(_06917_));
 sg13g2_mux2_1 _25925_ (.A0(_00095_),
    .A1(_00094_),
    .S(_11929_),
    .X(_06919_));
 sg13g2_nor2_1 _25926_ (.A(net996),
    .B(_06919_),
    .Y(_06920_));
 sg13g2_a21oi_1 _25927_ (.A1(net859),
    .A2(_06918_),
    .Y(_06921_),
    .B1(_06920_));
 sg13g2_nand2_1 _25928_ (.Y(_06922_),
    .A(net304),
    .B(_06921_));
 sg13g2_xor2_1 _25929_ (.B(_09087_),
    .A(_09084_),
    .X(_06923_));
 sg13g2_nor2_1 _25930_ (.A(net623),
    .B(_06923_),
    .Y(_06924_));
 sg13g2_nand2b_1 _25931_ (.Y(_06925_),
    .B(net103),
    .A_N(_06921_));
 sg13g2_o21ai_1 _25932_ (.B1(_06925_),
    .Y(_06926_),
    .A1(net103),
    .A2(_06923_));
 sg13g2_a22oi_1 _25933_ (.Y(_06927_),
    .B1(_06926_),
    .B2(net856),
    .A2(_06924_),
    .A1(_06922_));
 sg13g2_nand2b_1 _25934_ (.Y(_06928_),
    .B(net501),
    .A_N(\cpu.spi.r_clk_count[0][2] ));
 sg13g2_o21ai_1 _25935_ (.B1(_06928_),
    .Y(_06929_),
    .A1(net501),
    .A2(_05379_));
 sg13g2_mux2_1 _25936_ (.A0(\cpu.spi.r_clk_count[0][2] ),
    .A1(\cpu.spi.r_clk_count[1][2] ),
    .S(net520),
    .X(_06930_));
 sg13g2_nor2_1 _25937_ (.A(net727),
    .B(_06930_),
    .Y(_06931_));
 sg13g2_a21oi_1 _25938_ (.A1(net640),
    .A2(_06929_),
    .Y(_06932_),
    .B1(_06931_));
 sg13g2_nor2_1 _25939_ (.A(net439),
    .B(_06932_),
    .Y(_06933_));
 sg13g2_a21oi_1 _25940_ (.A1(net439),
    .A2(_06927_),
    .Y(_06934_),
    .B1(_06933_));
 sg13g2_mux2_1 _25941_ (.A0(_09084_),
    .A1(_06934_),
    .S(net31),
    .X(_02551_));
 sg13g2_nor2_1 _25942_ (.A(_09084_),
    .B(_09087_),
    .Y(_06935_));
 sg13g2_xnor2_1 _25943_ (.Y(_06936_),
    .A(\cpu.spi.r_count[3] ),
    .B(_06935_));
 sg13g2_nor2_1 _25944_ (.A(net623),
    .B(_06936_),
    .Y(_06937_));
 sg13g2_nor2_1 _25945_ (.A(net800),
    .B(_05458_),
    .Y(_06938_));
 sg13g2_a21oi_1 _25946_ (.A1(net728),
    .A2(_00105_),
    .Y(_06939_),
    .B1(_06938_));
 sg13g2_nand2_1 _25947_ (.Y(_06940_),
    .A(net858),
    .B(_00104_));
 sg13g2_o21ai_1 _25948_ (.B1(_06940_),
    .Y(_06941_),
    .A1(net858),
    .A2(_05460_));
 sg13g2_nor2_1 _25949_ (.A(net996),
    .B(_06941_),
    .Y(_06942_));
 sg13g2_a21oi_1 _25950_ (.A1(net859),
    .A2(_06939_),
    .Y(_06943_),
    .B1(_06942_));
 sg13g2_nand2_1 _25951_ (.Y(_06944_),
    .A(net379),
    .B(_06943_));
 sg13g2_nand2b_1 _25952_ (.Y(_06945_),
    .B(net103),
    .A_N(_06943_));
 sg13g2_o21ai_1 _25953_ (.B1(_06945_),
    .Y(_06946_),
    .A1(net103),
    .A2(_06936_));
 sg13g2_a22oi_1 _25954_ (.Y(_06947_),
    .B1(_06946_),
    .B2(net856),
    .A2(_06944_),
    .A1(_06937_));
 sg13g2_nand2b_1 _25955_ (.Y(_06948_),
    .B(net501),
    .A_N(\cpu.spi.r_clk_count[0][3] ));
 sg13g2_o21ai_1 _25956_ (.B1(_06948_),
    .Y(_06949_),
    .A1(net501),
    .A2(_05458_));
 sg13g2_mux2_1 _25957_ (.A0(\cpu.spi.r_clk_count[0][3] ),
    .A1(\cpu.spi.r_clk_count[1][3] ),
    .S(net520),
    .X(_06950_));
 sg13g2_nor2_1 _25958_ (.A(net727),
    .B(_06950_),
    .Y(_06951_));
 sg13g2_a21oi_1 _25959_ (.A1(net640),
    .A2(_06949_),
    .Y(_06952_),
    .B1(_06951_));
 sg13g2_nor2_1 _25960_ (.A(net439),
    .B(_06952_),
    .Y(_06953_));
 sg13g2_a21oi_1 _25961_ (.A1(net439),
    .A2(_06947_),
    .Y(_06954_),
    .B1(_06953_));
 sg13g2_mux2_1 _25962_ (.A0(\cpu.spi.r_count[3] ),
    .A1(_06954_),
    .S(net31),
    .X(_02552_));
 sg13g2_xnor2_1 _25963_ (.Y(_06955_),
    .A(\cpu.spi.r_count[4] ),
    .B(_09088_));
 sg13g2_nor2_1 _25964_ (.A(net623),
    .B(_06955_),
    .Y(_06956_));
 sg13g2_nor2_1 _25965_ (.A(net800),
    .B(_05522_),
    .Y(_06957_));
 sg13g2_a21oi_1 _25966_ (.A1(net728),
    .A2(_00115_),
    .Y(_06958_),
    .B1(_06957_));
 sg13g2_nand2_1 _25967_ (.Y(_06959_),
    .A(net858),
    .B(_00114_));
 sg13g2_o21ai_1 _25968_ (.B1(_06959_),
    .Y(_06960_),
    .A1(net858),
    .A2(_05523_));
 sg13g2_nor2_1 _25969_ (.A(net996),
    .B(_06960_),
    .Y(_06961_));
 sg13g2_a21oi_1 _25970_ (.A1(net859),
    .A2(_06958_),
    .Y(_06962_),
    .B1(_06961_));
 sg13g2_nand2_1 _25971_ (.Y(_06963_),
    .A(net379),
    .B(_06962_));
 sg13g2_nand2b_1 _25972_ (.Y(_06964_),
    .B(_09108_),
    .A_N(_06962_));
 sg13g2_o21ai_1 _25973_ (.B1(_06964_),
    .Y(_06965_),
    .A1(net103),
    .A2(_06955_));
 sg13g2_a22oi_1 _25974_ (.Y(_06966_),
    .B1(_06965_),
    .B2(net856),
    .A2(_06963_),
    .A1(_06956_));
 sg13g2_nand2b_1 _25975_ (.Y(_06967_),
    .B(net520),
    .A_N(\cpu.spi.r_clk_count[0][4] ));
 sg13g2_o21ai_1 _25976_ (.B1(_06967_),
    .Y(_06968_),
    .A1(net501),
    .A2(_05522_));
 sg13g2_mux2_1 _25977_ (.A0(\cpu.spi.r_clk_count[0][4] ),
    .A1(\cpu.spi.r_clk_count[1][4] ),
    .S(net520),
    .X(_06969_));
 sg13g2_nor2_1 _25978_ (.A(net727),
    .B(_06969_),
    .Y(_06970_));
 sg13g2_a21oi_1 _25979_ (.A1(net640),
    .A2(_06968_),
    .Y(_06971_),
    .B1(_06970_));
 sg13g2_nor2_1 _25980_ (.A(net439),
    .B(_06971_),
    .Y(_06972_));
 sg13g2_a21oi_1 _25981_ (.A1(net439),
    .A2(_06966_),
    .Y(_06973_),
    .B1(_06972_));
 sg13g2_mux2_1 _25982_ (.A0(\cpu.spi.r_count[4] ),
    .A1(_06973_),
    .S(net31),
    .X(_02553_));
 sg13g2_nor2_1 _25983_ (.A(net800),
    .B(_05620_),
    .Y(_06974_));
 sg13g2_a21oi_1 _25984_ (.A1(net800),
    .A2(_00121_),
    .Y(_06975_),
    .B1(_06974_));
 sg13g2_nand2_1 _25985_ (.Y(_06976_),
    .A(net995),
    .B(_00120_));
 sg13g2_o21ai_1 _25986_ (.B1(_06976_),
    .Y(_06977_),
    .A1(_11929_),
    .A2(_05621_));
 sg13g2_nor2_1 _25987_ (.A(net996),
    .B(_06977_),
    .Y(_06978_));
 sg13g2_a21oi_1 _25988_ (.A1(net859),
    .A2(_06975_),
    .Y(_06979_),
    .B1(_06978_));
 sg13g2_nand2_1 _25989_ (.Y(_06980_),
    .A(net304),
    .B(_06979_));
 sg13g2_xnor2_1 _25990_ (.Y(_06981_),
    .A(\cpu.spi.r_count[5] ),
    .B(_09089_));
 sg13g2_nor2_1 _25991_ (.A(net623),
    .B(_06981_),
    .Y(_06982_));
 sg13g2_nand2b_1 _25992_ (.Y(_06983_),
    .B(_09108_),
    .A_N(_06979_));
 sg13g2_o21ai_1 _25993_ (.B1(_06983_),
    .Y(_06984_),
    .A1(net103),
    .A2(_06981_));
 sg13g2_a22oi_1 _25994_ (.Y(_06985_),
    .B1(_06984_),
    .B2(net856),
    .A2(_06982_),
    .A1(_06980_));
 sg13g2_nand2b_1 _25995_ (.Y(_06986_),
    .B(net520),
    .A_N(\cpu.spi.r_clk_count[0][5] ));
 sg13g2_o21ai_1 _25996_ (.B1(_06986_),
    .Y(_06987_),
    .A1(net501),
    .A2(_05620_));
 sg13g2_mux2_1 _25997_ (.A0(\cpu.spi.r_clk_count[0][5] ),
    .A1(\cpu.spi.r_clk_count[1][5] ),
    .S(net520),
    .X(_06988_));
 sg13g2_nor2_1 _25998_ (.A(net727),
    .B(_06988_),
    .Y(_06989_));
 sg13g2_a21oi_1 _25999_ (.A1(net640),
    .A2(_06987_),
    .Y(_06990_),
    .B1(_06989_));
 sg13g2_nor2_1 _26000_ (.A(_06868_),
    .B(_06990_),
    .Y(_06991_));
 sg13g2_a21oi_1 _26001_ (.A1(_06869_),
    .A2(_06985_),
    .Y(_06992_),
    .B1(_06991_));
 sg13g2_mux2_1 _26002_ (.A0(\cpu.spi.r_count[5] ),
    .A1(_06992_),
    .S(net31),
    .X(_02554_));
 sg13g2_nor2_1 _26003_ (.A(net858),
    .B(_05678_),
    .Y(_06993_));
 sg13g2_a21oi_1 _26004_ (.A1(net800),
    .A2(_00132_),
    .Y(_06994_),
    .B1(_06993_));
 sg13g2_nand2_1 _26005_ (.Y(_06995_),
    .A(net995),
    .B(_00131_));
 sg13g2_o21ai_1 _26006_ (.B1(_06995_),
    .Y(_06996_),
    .A1(net858),
    .A2(_05679_));
 sg13g2_nor2_1 _26007_ (.A(net996),
    .B(_06996_),
    .Y(_06997_));
 sg13g2_a21oi_1 _26008_ (.A1(net859),
    .A2(_06994_),
    .Y(_06998_),
    .B1(_06997_));
 sg13g2_nand2_1 _26009_ (.Y(_06999_),
    .A(net304),
    .B(_06998_));
 sg13g2_xnor2_1 _26010_ (.Y(_07000_),
    .A(\cpu.spi.r_count[6] ),
    .B(_09090_));
 sg13g2_nor2_1 _26011_ (.A(net623),
    .B(_07000_),
    .Y(_07001_));
 sg13g2_nand2b_1 _26012_ (.Y(_07002_),
    .B(_09108_),
    .A_N(_06998_));
 sg13g2_o21ai_1 _26013_ (.B1(_07002_),
    .Y(_07003_),
    .A1(net103),
    .A2(_07000_));
 sg13g2_a22oi_1 _26014_ (.Y(_07004_),
    .B1(_07003_),
    .B2(_11965_),
    .A2(_07001_),
    .A1(_06999_));
 sg13g2_nand2b_1 _26015_ (.Y(_07005_),
    .B(net520),
    .A_N(\cpu.spi.r_clk_count[0][6] ));
 sg13g2_o21ai_1 _26016_ (.B1(_07005_),
    .Y(_07006_),
    .A1(net501),
    .A2(_05678_));
 sg13g2_mux2_1 _26017_ (.A0(\cpu.spi.r_clk_count[0][6] ),
    .A1(\cpu.spi.r_clk_count[1][6] ),
    .S(net520),
    .X(_07007_));
 sg13g2_nor2_1 _26018_ (.A(net727),
    .B(_07007_),
    .Y(_07008_));
 sg13g2_a21oi_1 _26019_ (.A1(net640),
    .A2(_07006_),
    .Y(_07009_),
    .B1(_07008_));
 sg13g2_nor2_1 _26020_ (.A(_06868_),
    .B(_07009_),
    .Y(_07010_));
 sg13g2_a21oi_1 _26021_ (.A1(net439),
    .A2(_07004_),
    .Y(_07011_),
    .B1(_07010_));
 sg13g2_mux2_1 _26022_ (.A0(\cpu.spi.r_count[6] ),
    .A1(_07011_),
    .S(net31),
    .X(_02555_));
 sg13g2_nand2b_1 _26023_ (.Y(_07012_),
    .B(net585),
    .A_N(\cpu.spi.r_clk_count[0][7] ));
 sg13g2_o21ai_1 _26024_ (.B1(_07012_),
    .Y(_07013_),
    .A1(net585),
    .A2(_05123_));
 sg13g2_mux2_1 _26025_ (.A0(\cpu.spi.r_clk_count[0][7] ),
    .A1(\cpu.spi.r_clk_count[1][7] ),
    .S(net646),
    .X(_07014_));
 sg13g2_nor2_1 _26026_ (.A(net857),
    .B(_07014_),
    .Y(_07015_));
 sg13g2_a21oi_1 _26027_ (.A1(net857),
    .A2(_07013_),
    .Y(_07016_),
    .B1(_07015_));
 sg13g2_nor2_1 _26028_ (.A(_06868_),
    .B(_07016_),
    .Y(_07017_));
 sg13g2_nor3_1 _26029_ (.A(_09056_),
    .B(_09092_),
    .C(_07017_),
    .Y(_07018_));
 sg13g2_nand2b_1 _26030_ (.Y(_07019_),
    .B(net31),
    .A_N(_07018_));
 sg13g2_nor2_1 _26031_ (.A(net995),
    .B(_05123_),
    .Y(_07020_));
 sg13g2_a21oi_1 _26032_ (.A1(net858),
    .A2(_00143_),
    .Y(_07021_),
    .B1(_07020_));
 sg13g2_nand2_1 _26033_ (.Y(_07022_),
    .A(_11917_),
    .B(_00142_));
 sg13g2_o21ai_1 _26034_ (.B1(_07022_),
    .Y(_07023_),
    .A1(net995),
    .A2(_05124_));
 sg13g2_nor2_1 _26035_ (.A(_11912_),
    .B(_07023_),
    .Y(_07024_));
 sg13g2_a21oi_1 _26036_ (.A1(net996),
    .A2(_07021_),
    .Y(_07025_),
    .B1(_07024_));
 sg13g2_nand2_1 _26037_ (.Y(_07026_),
    .A(_09054_),
    .B(net379));
 sg13g2_o21ai_1 _26038_ (.B1(_07026_),
    .Y(_07027_),
    .A1(_09054_),
    .A2(_07025_));
 sg13g2_nor2_1 _26039_ (.A(_09083_),
    .B(_07025_),
    .Y(_07028_));
 sg13g2_nor2b_1 _26040_ (.A(_09092_),
    .B_N(_09083_),
    .Y(_07029_));
 sg13g2_a21oi_1 _26041_ (.A1(_09092_),
    .A2(_07028_),
    .Y(_07030_),
    .B1(_07029_));
 sg13g2_o21ai_1 _26042_ (.B1(_06868_),
    .Y(_07031_),
    .A1(net623),
    .A2(_07030_));
 sg13g2_a21oi_1 _26043_ (.A1(_09098_),
    .A2(_07027_),
    .Y(_07032_),
    .B1(_07031_));
 sg13g2_nor2_1 _26044_ (.A(_07017_),
    .B(_07032_),
    .Y(_07033_));
 sg13g2_a22oi_1 _26045_ (.Y(_07034_),
    .B1(_07033_),
    .B2(_06894_),
    .A2(_07019_),
    .A1(_09083_));
 sg13g2_inv_1 _26046_ (.Y(_02556_),
    .A(_07034_));
 sg13g2_mux4_1 _26047_ (.S0(_05541_),
    .A0(_08991_),
    .A1(_09004_),
    .A2(_08996_),
    .A3(_09002_),
    .S1(\cpu.gpio.r_spi_miso_src[1][2] ),
    .X(_07035_));
 sg13g2_nand2_1 _26048_ (.Y(_07036_),
    .A(_08985_),
    .B(_05541_));
 sg13g2_nand2b_1 _26049_ (.Y(_07037_),
    .B(_08982_),
    .A_N(_05541_));
 sg13g2_nand3_1 _26050_ (.B(_07036_),
    .C(_07037_),
    .A(_06245_),
    .Y(_07038_));
 sg13g2_o21ai_1 _26051_ (.B1(_07038_),
    .Y(_07039_),
    .A1(_06245_),
    .A2(_07035_));
 sg13g2_nand2b_1 _26052_ (.Y(_07040_),
    .B(_05541_),
    .A_N(_08993_));
 sg13g2_o21ai_1 _26053_ (.B1(_07040_),
    .Y(_07041_),
    .A1(_09005_),
    .A2(_05541_));
 sg13g2_a21o_1 _26054_ (.A2(_07041_),
    .A1(\cpu.gpio.r_spi_miso_src[1][1] ),
    .B1(_00137_),
    .X(_07042_));
 sg13g2_mux4_1 _26055_ (.S0(_05541_),
    .A0(_09000_),
    .A1(_08980_),
    .A2(_08998_),
    .A3(_08987_),
    .S1(\cpu.gpio.r_spi_miso_src[1][2] ),
    .X(_07043_));
 sg13g2_nor3_1 _26056_ (.A(_06243_),
    .B(_06245_),
    .C(_07043_),
    .Y(_07044_));
 sg13g2_a221oi_1 _26057_ (.B2(_06245_),
    .C1(_07044_),
    .B1(_07042_),
    .A1(_06243_),
    .Y(_07045_),
    .A2(_07039_));
 sg13g2_mux4_1 _26058_ (.S0(_04965_),
    .A0(_09000_),
    .A1(_08980_),
    .A2(_08998_),
    .A3(_08987_),
    .S1(\cpu.gpio.r_spi_miso_src[0][2] ),
    .X(_07046_));
 sg13g2_nand2_1 _26059_ (.Y(_07047_),
    .A(_08993_),
    .B(_04965_));
 sg13g2_nand2b_1 _26060_ (.Y(_07048_),
    .B(_09005_),
    .A_N(_04965_));
 sg13g2_nand3_1 _26061_ (.B(_07047_),
    .C(_07048_),
    .A(_06242_),
    .Y(_07049_));
 sg13g2_o21ai_1 _26062_ (.B1(_07049_),
    .Y(_07050_),
    .A1(_06242_),
    .A2(_07046_));
 sg13g2_mux2_1 _26063_ (.A0(_08982_),
    .A1(_08985_),
    .S(_04965_),
    .X(_07051_));
 sg13g2_o21ai_1 _26064_ (.B1(_05364_),
    .Y(_07052_),
    .A1(_06241_),
    .A2(_07051_));
 sg13g2_mux4_1 _26065_ (.S0(_04965_),
    .A0(_08991_),
    .A1(_09004_),
    .A2(_08996_),
    .A3(_09002_),
    .S1(\cpu.gpio.r_spi_miso_src[0][2] ),
    .X(_07053_));
 sg13g2_nor3_1 _26066_ (.A(_06241_),
    .B(_06242_),
    .C(_07053_),
    .Y(_07054_));
 sg13g2_a221oi_1 _26067_ (.B2(_06242_),
    .C1(_07054_),
    .B1(_07052_),
    .A1(_06241_),
    .Y(_07055_),
    .A2(_07050_));
 sg13g2_mux2_1 _26068_ (.A0(_07045_),
    .A1(_07055_),
    .S(_11923_),
    .X(_07056_));
 sg13g2_nor3_1 _26069_ (.A(_09114_),
    .B(_09117_),
    .C(_11970_),
    .Y(_07057_));
 sg13g2_nand3_1 _26070_ (.B(_09117_),
    .C(_11970_),
    .A(_09114_),
    .Y(_07058_));
 sg13g2_nand2b_1 _26071_ (.Y(_07059_),
    .B(_07058_),
    .A_N(_07057_));
 sg13g2_nand3_1 _26072_ (.B(_09094_),
    .C(_07059_),
    .A(net901),
    .Y(_07060_));
 sg13g2_buf_4 _26073_ (.X(_07061_),
    .A(_07060_));
 sg13g2_mux2_1 _26074_ (.A0(_07056_),
    .A1(_09073_),
    .S(_07061_),
    .X(_02560_));
 sg13g2_mux2_1 _26075_ (.A0(_09073_),
    .A1(_09072_),
    .S(_07061_),
    .X(_02561_));
 sg13g2_mux2_1 _26076_ (.A0(_09072_),
    .A1(_09076_),
    .S(_07061_),
    .X(_02562_));
 sg13g2_mux2_1 _26077_ (.A0(_09076_),
    .A1(_09070_),
    .S(_07061_),
    .X(_02563_));
 sg13g2_mux2_1 _26078_ (.A0(_09070_),
    .A1(_09078_),
    .S(_07061_),
    .X(_02564_));
 sg13g2_mux2_1 _26079_ (.A0(_09078_),
    .A1(_09077_),
    .S(_07061_),
    .X(_02565_));
 sg13g2_mux2_1 _26080_ (.A0(_09077_),
    .A1(_09071_),
    .S(_07061_),
    .X(_02566_));
 sg13g2_mux2_1 _26081_ (.A0(_09071_),
    .A1(\cpu.spi.r_in[7] ),
    .S(_07061_),
    .X(_02567_));
 sg13g2_nor3_2 _26082_ (.A(net575),
    .B(net448),
    .C(_06851_),
    .Y(_07062_));
 sg13g2_mux2_1 _26083_ (.A0(\cpu.spi.r_mode[0][0] ),
    .A1(net877),
    .S(_07062_),
    .X(_02569_));
 sg13g2_mux2_1 _26084_ (.A0(_11927_),
    .A1(net855),
    .S(_07062_),
    .X(_02570_));
 sg13g2_nor3_2 _26085_ (.A(net575),
    .B(net566),
    .C(_06851_),
    .Y(_07063_));
 sg13g2_mux2_1 _26086_ (.A0(\cpu.spi.r_mode[1][0] ),
    .A1(net877),
    .S(_07063_),
    .X(_02571_));
 sg13g2_mux2_1 _26087_ (.A0(_11928_),
    .A1(net855),
    .S(_07063_),
    .X(_02572_));
 sg13g2_nand4_1 _26088_ (.B(net566),
    .C(_06849_),
    .A(net673),
    .Y(_07064_),
    .D(_06857_));
 sg13g2_buf_1 _26089_ (.A(_07064_),
    .X(_07065_));
 sg13g2_mux2_1 _26090_ (.A0(net880),
    .A1(\cpu.spi.r_mode[2][0] ),
    .S(_07065_),
    .X(_02573_));
 sg13g2_mux2_1 _26091_ (.A0(net829),
    .A1(_11933_),
    .S(_07065_),
    .X(_02574_));
 sg13g2_nor2_1 _26092_ (.A(_09044_),
    .B(_11936_),
    .Y(_07066_));
 sg13g2_buf_2 _26093_ (.A(_07066_),
    .X(_07067_));
 sg13g2_a22oi_1 _26094_ (.Y(_07068_),
    .B1(_07067_),
    .B2(_06888_),
    .A2(_11973_),
    .A1(net1110));
 sg13g2_nand4_1 _26095_ (.B(_09162_),
    .C(_11977_),
    .A(_09056_),
    .Y(_07069_),
    .D(_07068_));
 sg13g2_buf_1 _26096_ (.A(_07069_),
    .X(_07070_));
 sg13g2_buf_1 _26097_ (.A(_09125_),
    .X(_07071_));
 sg13g2_buf_1 _26098_ (.A(_11970_),
    .X(_07072_));
 sg13g2_nand2b_1 _26099_ (.Y(_07073_),
    .B(_00202_),
    .A_N(net555));
 sg13g2_nor2_1 _26100_ (.A(_09125_),
    .B(_06864_),
    .Y(_07074_));
 sg13g2_a221oi_1 _26101_ (.B2(_07074_),
    .C1(_11959_),
    .B1(_07073_),
    .A1(net799),
    .Y(_07075_),
    .A2(net1024));
 sg13g2_nand2_1 _26102_ (.Y(_07076_),
    .A(\cpu.spi.r_out[0] ),
    .B(net67));
 sg13g2_o21ai_1 _26103_ (.B1(_07076_),
    .Y(_02575_),
    .A1(net67),
    .A2(_07075_));
 sg13g2_mux2_1 _26104_ (.A0(_00162_),
    .A1(_00202_),
    .S(net555),
    .X(_07077_));
 sg13g2_a22oi_1 _26105_ (.Y(_07078_),
    .B1(_07067_),
    .B2(net1023),
    .A2(net726),
    .A1(\cpu.spi.r_out[0] ));
 sg13g2_o21ai_1 _26106_ (.B1(_07078_),
    .Y(_07079_),
    .A1(net799),
    .A2(_07077_));
 sg13g2_mux2_1 _26107_ (.A0(_07079_),
    .A1(\cpu.spi.r_out[1] ),
    .S(_07070_),
    .X(_02576_));
 sg13g2_mux2_1 _26108_ (.A0(_00163_),
    .A1(_00162_),
    .S(net555),
    .X(_07080_));
 sg13g2_a22oi_1 _26109_ (.Y(_07081_),
    .B1(_07067_),
    .B2(net1017),
    .A2(net726),
    .A1(\cpu.spi.r_out[1] ));
 sg13g2_o21ai_1 _26110_ (.B1(_07081_),
    .Y(_07082_),
    .A1(net799),
    .A2(_07080_));
 sg13g2_mux2_1 _26111_ (.A0(_07082_),
    .A1(\cpu.spi.r_out[2] ),
    .S(net67),
    .X(_02577_));
 sg13g2_mux2_1 _26112_ (.A0(_00266_),
    .A1(_00163_),
    .S(net555),
    .X(_07083_));
 sg13g2_a22oi_1 _26113_ (.Y(_07084_),
    .B1(_07067_),
    .B2(_09890_),
    .A2(net726),
    .A1(\cpu.spi.r_out[2] ));
 sg13g2_o21ai_1 _26114_ (.B1(_07084_),
    .Y(_07085_),
    .A1(net799),
    .A2(_07083_));
 sg13g2_mux2_1 _26115_ (.A0(_07085_),
    .A1(\cpu.spi.r_out[3] ),
    .S(net67),
    .X(_02578_));
 sg13g2_mux2_1 _26116_ (.A0(_00164_),
    .A1(_00266_),
    .S(net555),
    .X(_07086_));
 sg13g2_a22oi_1 _26117_ (.Y(_07087_),
    .B1(_07067_),
    .B2(net1105),
    .A2(net726),
    .A1(\cpu.spi.r_out[3] ));
 sg13g2_o21ai_1 _26118_ (.B1(_07087_),
    .Y(_07088_),
    .A1(net799),
    .A2(_07086_));
 sg13g2_mux2_1 _26119_ (.A0(_07088_),
    .A1(\cpu.spi.r_out[4] ),
    .S(net67),
    .X(_02579_));
 sg13g2_mux2_1 _26120_ (.A0(_00165_),
    .A1(_00164_),
    .S(net555),
    .X(_07089_));
 sg13g2_a22oi_1 _26121_ (.Y(_07090_),
    .B1(_07067_),
    .B2(_09901_),
    .A2(net726),
    .A1(\cpu.spi.r_out[4] ));
 sg13g2_o21ai_1 _26122_ (.B1(_07090_),
    .Y(_07091_),
    .A1(net799),
    .A2(_07089_));
 sg13g2_mux2_1 _26123_ (.A0(_07091_),
    .A1(\cpu.spi.r_out[5] ),
    .S(net67),
    .X(_02580_));
 sg13g2_inv_1 _26124_ (.Y(_07092_),
    .A(_00166_));
 sg13g2_nand2_1 _26125_ (.Y(_07093_),
    .A(_00165_),
    .B(net555));
 sg13g2_o21ai_1 _26126_ (.B1(_07093_),
    .Y(_07094_),
    .A1(_07092_),
    .A2(net555));
 sg13g2_a22oi_1 _26127_ (.Y(_07095_),
    .B1(_07067_),
    .B2(_09907_),
    .A2(_11959_),
    .A1(\cpu.spi.r_out[5] ));
 sg13g2_o21ai_1 _26128_ (.B1(_07095_),
    .Y(_07096_),
    .A1(_07071_),
    .A2(_07094_));
 sg13g2_mux2_1 _26129_ (.A0(_07096_),
    .A1(\cpu.spi.r_out[6] ),
    .S(net67),
    .X(_02581_));
 sg13g2_buf_1 _26130_ (.A(_00260_),
    .X(_07097_));
 sg13g2_nor2_1 _26131_ (.A(_07097_),
    .B(_07072_),
    .Y(_07098_));
 sg13g2_a21oi_1 _26132_ (.A1(_07092_),
    .A2(_07072_),
    .Y(_07099_),
    .B1(_07098_));
 sg13g2_a22oi_1 _26133_ (.Y(_07100_),
    .B1(_07067_),
    .B2(net1104),
    .A2(net726),
    .A1(\cpu.spi.r_out[6] ));
 sg13g2_o21ai_1 _26134_ (.B1(_07100_),
    .Y(_07101_),
    .A1(_07071_),
    .A2(_07099_));
 sg13g2_mux2_1 _26135_ (.A0(_07101_),
    .A1(\cpu.spi.r_out[7] ),
    .S(net67),
    .X(_02582_));
 sg13g2_nor4_2 _26136_ (.A(_06888_),
    .B(net778),
    .C(_09040_),
    .Y(_07102_),
    .D(_09048_));
 sg13g2_mux2_1 _26137_ (.A0(net728),
    .A1(net448),
    .S(_07102_),
    .X(_02585_));
 sg13g2_nand2_1 _26138_ (.Y(_07103_),
    .A(net579),
    .B(_07102_));
 sg13g2_o21ai_1 _26139_ (.B1(_07103_),
    .Y(_02586_),
    .A1(_11926_),
    .A2(_07102_));
 sg13g2_mux2_1 _26140_ (.A0(\cpu.spi.r_src[0] ),
    .A1(net876),
    .S(_07062_),
    .X(_02587_));
 sg13g2_mux2_1 _26141_ (.A0(\cpu.spi.r_src[1] ),
    .A1(net876),
    .S(_07063_),
    .X(_02588_));
 sg13g2_nand2_1 _26142_ (.Y(_07104_),
    .A(_11915_),
    .B(_07065_));
 sg13g2_o21ai_1 _26143_ (.B1(_07104_),
    .Y(_02589_),
    .A1(net878),
    .A2(_07065_));
 sg13g2_nand2b_1 _26144_ (.Y(_07105_),
    .B(_05127_),
    .A_N(_09048_));
 sg13g2_buf_1 _26145_ (.A(_07105_),
    .X(_07106_));
 sg13g2_buf_1 _26146_ (.A(_07106_),
    .X(_07107_));
 sg13g2_mux2_1 _26147_ (.A0(net880),
    .A1(\cpu.spi.r_timeout[0] ),
    .S(_07107_),
    .X(_02590_));
 sg13g2_mux2_1 _26148_ (.A0(net829),
    .A1(\cpu.spi.r_timeout[1] ),
    .S(_07107_),
    .X(_02591_));
 sg13g2_nand2_1 _26149_ (.Y(_07108_),
    .A(\cpu.spi.r_timeout[2] ),
    .B(net87));
 sg13g2_o21ai_1 _26150_ (.B1(_07108_),
    .Y(_02592_),
    .A1(net878),
    .A2(net87));
 sg13g2_nand2_1 _26151_ (.Y(_07109_),
    .A(\cpu.spi.r_timeout[3] ),
    .B(net87));
 sg13g2_o21ai_1 _26152_ (.B1(_07109_),
    .Y(_02593_),
    .A1(net854),
    .A2(net87));
 sg13g2_nand2_1 _26153_ (.Y(_07110_),
    .A(\cpu.spi.r_timeout[4] ),
    .B(_07106_));
 sg13g2_o21ai_1 _26154_ (.B1(_07110_),
    .Y(_02594_),
    .A1(net853),
    .A2(net87));
 sg13g2_mux2_1 _26155_ (.A0(net849),
    .A1(\cpu.spi.r_timeout[5] ),
    .S(net87),
    .X(_02595_));
 sg13g2_mux2_1 _26156_ (.A0(net875),
    .A1(\cpu.spi.r_timeout[6] ),
    .S(net87),
    .X(_02596_));
 sg13g2_nand2_1 _26157_ (.Y(_07111_),
    .A(\cpu.spi.r_timeout[7] ),
    .B(_07106_));
 sg13g2_o21ai_1 _26158_ (.B1(_07111_),
    .Y(_02597_),
    .A1(net852),
    .A2(net87));
 sg13g2_inv_1 _26159_ (.Y(_07112_),
    .A(\cpu.spi.r_timeout_count[0] ));
 sg13g2_mux2_1 _26160_ (.A0(_09114_),
    .A1(_09054_),
    .S(_09044_),
    .X(_07113_));
 sg13g2_nor2_1 _26161_ (.A(_09082_),
    .B(_09112_),
    .Y(_07114_));
 sg13g2_nor2_1 _26162_ (.A(_09114_),
    .B(_07114_),
    .Y(_07115_));
 sg13g2_nor4_1 _26163_ (.A(_11910_),
    .B(_09061_),
    .C(_09082_),
    .D(_09113_),
    .Y(_07116_));
 sg13g2_nor4_1 _26164_ (.A(net897),
    .B(_07113_),
    .C(_07115_),
    .D(_07116_),
    .Y(_07117_));
 sg13g2_buf_2 _26165_ (.A(_07117_),
    .X(_07118_));
 sg13g2_buf_1 _26166_ (.A(_07118_),
    .X(_07119_));
 sg13g2_mux2_1 _26167_ (.A0(_00263_),
    .A1(\cpu.spi.r_timeout[0] ),
    .S(net1033),
    .X(_07120_));
 sg13g2_nand2_1 _26168_ (.Y(_07121_),
    .A(net66),
    .B(_07120_));
 sg13g2_o21ai_1 _26169_ (.B1(_07121_),
    .Y(_02598_),
    .A1(_07112_),
    .A2(net66));
 sg13g2_o21ai_1 _26170_ (.B1(net66),
    .Y(_07122_),
    .A1(_07112_),
    .A2(net899));
 sg13g2_nor2_1 _26171_ (.A(\cpu.spi.r_timeout_count[0] ),
    .B(\cpu.spi.r_timeout_count[1] ),
    .Y(_07123_));
 sg13g2_mux2_1 _26172_ (.A0(\cpu.spi.r_timeout[1] ),
    .A1(_07123_),
    .S(net799),
    .X(_07124_));
 sg13g2_a22oi_1 _26173_ (.Y(_07125_),
    .B1(_07124_),
    .B2(net66),
    .A2(_07122_),
    .A1(\cpu.spi.r_timeout_count[1] ));
 sg13g2_inv_1 _26174_ (.Y(_02599_),
    .A(_07125_));
 sg13g2_o21ai_1 _26175_ (.B1(_07118_),
    .Y(_07126_),
    .A1(net899),
    .A2(_07123_));
 sg13g2_mux2_1 _26176_ (.A0(\cpu.spi.r_timeout[2] ),
    .A1(_09062_),
    .S(net799),
    .X(_07127_));
 sg13g2_a22oi_1 _26177_ (.Y(_07128_),
    .B1(_07127_),
    .B2(net66),
    .A2(_07126_),
    .A1(\cpu.spi.r_timeout_count[2] ));
 sg13g2_inv_1 _26178_ (.Y(_02600_),
    .A(_07128_));
 sg13g2_o21ai_1 _26179_ (.B1(_07118_),
    .Y(_07129_),
    .A1(net899),
    .A2(_09062_));
 sg13g2_nand2b_1 _26180_ (.Y(_07130_),
    .B(_09062_),
    .A_N(\cpu.spi.r_timeout_count[3] ));
 sg13g2_nand2_1 _26181_ (.Y(_07131_),
    .A(net856),
    .B(\cpu.spi.r_timeout[3] ));
 sg13g2_o21ai_1 _26182_ (.B1(_07131_),
    .Y(_07132_),
    .A1(net899),
    .A2(_07130_));
 sg13g2_a22oi_1 _26183_ (.Y(_07133_),
    .B1(_07132_),
    .B2(net66),
    .A2(_07129_),
    .A1(\cpu.spi.r_timeout_count[3] ));
 sg13g2_inv_1 _26184_ (.Y(_02601_),
    .A(_07133_));
 sg13g2_o21ai_1 _26185_ (.B1(_07118_),
    .Y(_07134_),
    .A1(net899),
    .A2(_09063_));
 sg13g2_nand2_1 _26186_ (.Y(_07135_),
    .A(net1033),
    .B(\cpu.spi.r_timeout[4] ));
 sg13g2_o21ai_1 _26187_ (.B1(_07135_),
    .Y(_07136_),
    .A1(net899),
    .A2(_09064_));
 sg13g2_a22oi_1 _26188_ (.Y(_07137_),
    .B1(_07136_),
    .B2(net66),
    .A2(_07134_),
    .A1(\cpu.spi.r_timeout_count[4] ));
 sg13g2_inv_1 _26189_ (.Y(_02602_),
    .A(_07137_));
 sg13g2_nor2_1 _26190_ (.A(\cpu.spi.r_timeout_count[4] ),
    .B(_07130_),
    .Y(_07138_));
 sg13g2_o21ai_1 _26191_ (.B1(_07118_),
    .Y(_07139_),
    .A1(net899),
    .A2(_07138_));
 sg13g2_mux2_1 _26192_ (.A0(\cpu.spi.r_timeout[5] ),
    .A1(_09065_),
    .S(_09125_),
    .X(_07140_));
 sg13g2_a22oi_1 _26193_ (.Y(_07141_),
    .B1(_07140_),
    .B2(_07119_),
    .A2(_07139_),
    .A1(\cpu.spi.r_timeout_count[5] ));
 sg13g2_inv_1 _26194_ (.Y(_02603_),
    .A(_07141_));
 sg13g2_o21ai_1 _26195_ (.B1(_07118_),
    .Y(_07142_),
    .A1(net856),
    .A2(_09065_));
 sg13g2_nand2_1 _26196_ (.Y(_07143_),
    .A(net1033),
    .B(\cpu.spi.r_timeout[6] ));
 sg13g2_o21ai_1 _26197_ (.B1(_07143_),
    .Y(_07144_),
    .A1(_09099_),
    .A2(_09067_));
 sg13g2_a22oi_1 _26198_ (.Y(_07145_),
    .B1(_07144_),
    .B2(net66),
    .A2(_07142_),
    .A1(\cpu.spi.r_timeout_count[6] ));
 sg13g2_inv_1 _26199_ (.Y(_02604_),
    .A(_07145_));
 sg13g2_inv_1 _26200_ (.Y(_07146_),
    .A(_09067_));
 sg13g2_o21ai_1 _26201_ (.B1(_07118_),
    .Y(_07147_),
    .A1(net856),
    .A2(_07146_));
 sg13g2_nor3_1 _26202_ (.A(\cpu.spi.r_timeout_count[7] ),
    .B(net1033),
    .C(_09067_),
    .Y(_07148_));
 sg13g2_a21o_1 _26203_ (.A2(\cpu.spi.r_timeout[7] ),
    .A1(net899),
    .B1(_07148_),
    .X(_07149_));
 sg13g2_a22oi_1 _26204_ (.Y(_07150_),
    .B1(_07149_),
    .B2(_07119_),
    .A2(_07147_),
    .A1(\cpu.spi.r_timeout_count[7] ));
 sg13g2_inv_1 _26205_ (.Y(_02605_),
    .A(_07150_));
 sg13g2_buf_1 _26206_ (.A(\cpu.uart.r_rcnt[0] ),
    .X(_07151_));
 sg13g2_nor2_1 _26207_ (.A(_07151_),
    .B(\cpu.uart.r_rcnt[1] ),
    .Y(_07152_));
 sg13g2_nand2_1 _26208_ (.Y(_07153_),
    .A(net252),
    .B(_07152_));
 sg13g2_nor2_1 _26209_ (.A(net897),
    .B(_07153_),
    .Y(_07154_));
 sg13g2_buf_2 _26210_ (.A(\cpu.uart.r_rstate[3] ),
    .X(_07155_));
 sg13g2_buf_1 _26211_ (.A(_07155_),
    .X(_07156_));
 sg13g2_buf_1 _26212_ (.A(\cpu.uart.r_rstate[1] ),
    .X(_07157_));
 sg13g2_buf_1 _26213_ (.A(\cpu.uart.r_rstate[2] ),
    .X(_07158_));
 sg13g2_nor2_2 _26214_ (.A(net1071),
    .B(_07158_),
    .Y(_07159_));
 sg13g2_buf_2 _26215_ (.A(\cpu.uart.r_rstate[0] ),
    .X(_07160_));
 sg13g2_inv_1 _26216_ (.Y(_07161_),
    .A(_07160_));
 sg13g2_nand3_1 _26217_ (.B(net924),
    .C(_07159_),
    .A(_07161_),
    .Y(_07162_));
 sg13g2_o21ai_1 _26218_ (.B1(_07162_),
    .Y(_07163_),
    .A1(net924),
    .A2(_07159_));
 sg13g2_and2_1 _26219_ (.A(_07154_),
    .B(_07163_),
    .X(_07164_));
 sg13g2_buf_2 _26220_ (.A(_07164_),
    .X(_07165_));
 sg13g2_mux2_1 _26221_ (.A0(\cpu.uart.r_ib[0] ),
    .A1(\cpu.uart.r_ib[1] ),
    .S(_07165_),
    .X(_02618_));
 sg13g2_mux2_1 _26222_ (.A0(\cpu.uart.r_ib[1] ),
    .A1(\cpu.uart.r_ib[2] ),
    .S(_07165_),
    .X(_02619_));
 sg13g2_mux2_1 _26223_ (.A0(\cpu.uart.r_ib[2] ),
    .A1(\cpu.uart.r_ib[3] ),
    .S(_07165_),
    .X(_02620_));
 sg13g2_mux2_1 _26224_ (.A0(\cpu.uart.r_ib[3] ),
    .A1(\cpu.uart.r_ib[4] ),
    .S(_07165_),
    .X(_02621_));
 sg13g2_mux2_1 _26225_ (.A0(\cpu.uart.r_ib[4] ),
    .A1(\cpu.uart.r_ib[5] ),
    .S(_07165_),
    .X(_02622_));
 sg13g2_mux2_1 _26226_ (.A0(\cpu.uart.r_ib[5] ),
    .A1(\cpu.uart.r_ib[6] ),
    .S(_07165_),
    .X(_02623_));
 sg13g2_xor2_1 _26227_ (.B(\cpu.uart.r_r ),
    .A(\cpu.uart.r_r_invert ),
    .X(_07166_));
 sg13g2_mux2_1 _26228_ (.A0(\cpu.uart.r_ib[6] ),
    .A1(_07166_),
    .S(_07165_),
    .X(_02624_));
 sg13g2_and4_1 _26229_ (.A(_07160_),
    .B(net924),
    .C(_07154_),
    .D(_07159_),
    .X(_07167_));
 sg13g2_buf_1 _26230_ (.A(_07167_),
    .X(_07168_));
 sg13g2_mux2_1 _26231_ (.A0(\cpu.uart.r_in[0] ),
    .A1(\cpu.uart.r_ib[0] ),
    .S(net127),
    .X(_02625_));
 sg13g2_mux2_1 _26232_ (.A0(\cpu.uart.r_in[1] ),
    .A1(\cpu.uart.r_ib[1] ),
    .S(net127),
    .X(_02626_));
 sg13g2_mux2_1 _26233_ (.A0(\cpu.uart.r_in[2] ),
    .A1(\cpu.uart.r_ib[2] ),
    .S(net127),
    .X(_02627_));
 sg13g2_mux2_1 _26234_ (.A0(\cpu.uart.r_in[3] ),
    .A1(\cpu.uart.r_ib[3] ),
    .S(net127),
    .X(_02628_));
 sg13g2_mux2_1 _26235_ (.A0(\cpu.uart.r_in[4] ),
    .A1(\cpu.uart.r_ib[4] ),
    .S(net127),
    .X(_02629_));
 sg13g2_mux2_1 _26236_ (.A0(\cpu.uart.r_in[5] ),
    .A1(\cpu.uart.r_ib[5] ),
    .S(net127),
    .X(_02630_));
 sg13g2_mux2_1 _26237_ (.A0(\cpu.uart.r_in[6] ),
    .A1(\cpu.uart.r_ib[6] ),
    .S(net127),
    .X(_02631_));
 sg13g2_mux2_1 _26238_ (.A0(\cpu.uart.r_in[7] ),
    .A1(_07166_),
    .S(_07168_),
    .X(_02632_));
 sg13g2_buf_1 _26239_ (.A(\cpu.uart.r_xstate[1] ),
    .X(_07169_));
 sg13g2_buf_1 _26240_ (.A(\cpu.uart.r_xstate[3] ),
    .X(_07170_));
 sg13g2_buf_1 _26241_ (.A(_07170_),
    .X(_07171_));
 sg13g2_buf_1 _26242_ (.A(\cpu.uart.r_xstate[2] ),
    .X(_07172_));
 sg13g2_buf_1 _26243_ (.A(_07172_),
    .X(_07173_));
 sg13g2_nor3_1 _26244_ (.A(_07169_),
    .B(net923),
    .C(_07173_),
    .Y(_07174_));
 sg13g2_buf_1 _26245_ (.A(\cpu.uart.r_xstate[0] ),
    .X(_07175_));
 sg13g2_inv_1 _26246_ (.Y(_07176_),
    .A(_07175_));
 sg13g2_nor2_1 _26247_ (.A(net1037),
    .B(net965),
    .Y(_07177_));
 sg13g2_and3_1 _26248_ (.X(_07178_),
    .A(net994),
    .B(_07177_),
    .C(_06227_));
 sg13g2_buf_1 _26249_ (.A(_07178_),
    .X(_07179_));
 sg13g2_nand2_1 _26250_ (.Y(_07180_),
    .A(_07176_),
    .B(_07179_));
 sg13g2_nand2_1 _26251_ (.Y(_07181_),
    .A(net402),
    .B(_07179_));
 sg13g2_nand3_1 _26252_ (.B(_07177_),
    .C(_06227_),
    .A(_11938_),
    .Y(_07182_));
 sg13g2_nor2_1 _26253_ (.A(net1070),
    .B(net1069),
    .Y(_07183_));
 sg13g2_nor2_1 _26254_ (.A(_07170_),
    .B(net922),
    .Y(_07184_));
 sg13g2_and2_1 _26255_ (.A(_07183_),
    .B(_07184_),
    .X(_07185_));
 sg13g2_buf_1 _26256_ (.A(_07185_),
    .X(_07186_));
 sg13g2_inv_1 _26257_ (.Y(_07187_),
    .A(_07186_));
 sg13g2_nor2b_1 _26258_ (.A(_07172_),
    .B_N(_07170_),
    .Y(_07188_));
 sg13g2_and2_1 _26259_ (.A(net1070),
    .B(_07188_),
    .X(_07189_));
 sg13g2_buf_1 _26260_ (.A(_07189_),
    .X(_07190_));
 sg13g2_nand2_1 _26261_ (.Y(_07191_),
    .A(net1069),
    .B(_07190_));
 sg13g2_o21ai_1 _26262_ (.B1(_07191_),
    .Y(_07192_),
    .A1(_07182_),
    .A2(_07187_));
 sg13g2_and2_1 _26263_ (.A(net1070),
    .B(\cpu.uart.r_xstate[0] ),
    .X(_07193_));
 sg13g2_buf_1 _26264_ (.A(_07193_),
    .X(_07194_));
 sg13g2_nand2_1 _26265_ (.Y(_07195_),
    .A(_07171_),
    .B(_07194_));
 sg13g2_buf_1 _26266_ (.A(\cpu.uart.r_xcnt[0] ),
    .X(_07196_));
 sg13g2_nor2_1 _26267_ (.A(_07196_),
    .B(\cpu.uart.r_xcnt[1] ),
    .Y(_07197_));
 sg13g2_nand2_1 _26268_ (.Y(_07198_),
    .A(_09743_),
    .B(_07197_));
 sg13g2_buf_1 _26269_ (.A(_07198_),
    .X(_07199_));
 sg13g2_a21o_1 _26270_ (.A2(_07199_),
    .A1(net923),
    .B1(net1070),
    .X(_07200_));
 sg13g2_a21oi_1 _26271_ (.A1(_07195_),
    .A2(_07200_),
    .Y(_07201_),
    .B1(_07173_));
 sg13g2_nor2_1 _26272_ (.A(net923),
    .B(_07199_),
    .Y(_07202_));
 sg13g2_o21ai_1 _26273_ (.B1(net1039),
    .Y(_07203_),
    .A1(_07201_),
    .A2(_07202_));
 sg13g2_a221oi_1 _26274_ (.B2(_07192_),
    .C1(_07203_),
    .B1(_07181_),
    .A1(_07174_),
    .Y(_07204_),
    .A2(_07180_));
 sg13g2_buf_1 _26275_ (.A(_07204_),
    .X(_07205_));
 sg13g2_buf_1 _26276_ (.A(_07205_),
    .X(_07206_));
 sg13g2_nor2_1 _26277_ (.A(_07169_),
    .B(net922),
    .Y(_07207_));
 sg13g2_xnor2_1 _26278_ (.Y(_07208_),
    .A(net923),
    .B(_07207_));
 sg13g2_buf_1 _26279_ (.A(_07208_),
    .X(_07209_));
 sg13g2_buf_1 _26280_ (.A(_07209_),
    .X(_07210_));
 sg13g2_nor2b_1 _26281_ (.A(_07209_),
    .B_N(_09859_),
    .Y(_07211_));
 sg13g2_a21oi_1 _26282_ (.A1(\cpu.uart.r_out[1] ),
    .A2(_07210_),
    .Y(_07212_),
    .B1(_07211_));
 sg13g2_nor2_1 _26283_ (.A(\cpu.uart.r_out[0] ),
    .B(net74),
    .Y(_07213_));
 sg13g2_a21oi_1 _26284_ (.A1(net74),
    .A2(_07212_),
    .Y(_02633_),
    .B1(_07213_));
 sg13g2_nor2b_1 _26285_ (.A(_07209_),
    .B_N(_09870_),
    .Y(_07214_));
 sg13g2_a21oi_1 _26286_ (.A1(\cpu.uart.r_out[2] ),
    .A2(net554),
    .Y(_07215_),
    .B1(_07214_));
 sg13g2_nor2_1 _26287_ (.A(\cpu.uart.r_out[1] ),
    .B(_07206_),
    .Y(_07216_));
 sg13g2_a21oi_1 _26288_ (.A1(net74),
    .A2(_07215_),
    .Y(_02634_),
    .B1(_07216_));
 sg13g2_nor2_1 _26289_ (.A(net878),
    .B(net554),
    .Y(_07217_));
 sg13g2_a21oi_1 _26290_ (.A1(\cpu.uart.r_out[3] ),
    .A2(net554),
    .Y(_07218_),
    .B1(_07217_));
 sg13g2_nor2_1 _26291_ (.A(\cpu.uart.r_out[2] ),
    .B(_07205_),
    .Y(_07219_));
 sg13g2_a21oi_1 _26292_ (.A1(net74),
    .A2(_07218_),
    .Y(_02635_),
    .B1(_07219_));
 sg13g2_nor2_1 _26293_ (.A(_12111_),
    .B(net554),
    .Y(_07220_));
 sg13g2_a21oi_1 _26294_ (.A1(\cpu.uart.r_out[4] ),
    .A2(net554),
    .Y(_07221_),
    .B1(_07220_));
 sg13g2_nor2_1 _26295_ (.A(\cpu.uart.r_out[3] ),
    .B(_07205_),
    .Y(_07222_));
 sg13g2_a21oi_1 _26296_ (.A1(net74),
    .A2(_07221_),
    .Y(_02636_),
    .B1(_07222_));
 sg13g2_nor2_1 _26297_ (.A(_12120_),
    .B(_07209_),
    .Y(_07223_));
 sg13g2_a21oi_1 _26298_ (.A1(\cpu.uart.r_out[5] ),
    .A2(net554),
    .Y(_07224_),
    .B1(_07223_));
 sg13g2_nor2_1 _26299_ (.A(\cpu.uart.r_out[4] ),
    .B(_07205_),
    .Y(_07225_));
 sg13g2_a21oi_1 _26300_ (.A1(net74),
    .A2(_07224_),
    .Y(_02637_),
    .B1(_07225_));
 sg13g2_nor2b_1 _26301_ (.A(_07209_),
    .B_N(_09901_),
    .Y(_07226_));
 sg13g2_a21oi_1 _26302_ (.A1(\cpu.uart.r_out[6] ),
    .A2(net554),
    .Y(_07227_),
    .B1(_07226_));
 sg13g2_nor2_1 _26303_ (.A(\cpu.uart.r_out[5] ),
    .B(_07205_),
    .Y(_07228_));
 sg13g2_a21oi_1 _26304_ (.A1(net74),
    .A2(_07227_),
    .Y(_02638_),
    .B1(_07228_));
 sg13g2_nor2b_1 _26305_ (.A(_07209_),
    .B_N(_09907_),
    .Y(_07229_));
 sg13g2_a21oi_1 _26306_ (.A1(\cpu.uart.r_out[7] ),
    .A2(net554),
    .Y(_07230_),
    .B1(_07229_));
 sg13g2_nor2_1 _26307_ (.A(\cpu.uart.r_out[6] ),
    .B(_07205_),
    .Y(_07231_));
 sg13g2_a21oi_1 _26308_ (.A1(net74),
    .A2(_07230_),
    .Y(_02639_),
    .B1(_07231_));
 sg13g2_nor2_1 _26309_ (.A(_07097_),
    .B(_07210_),
    .Y(_07232_));
 sg13g2_mux2_1 _26310_ (.A0(\cpu.uart.r_out[7] ),
    .A1(_07232_),
    .S(_07206_),
    .X(_02640_));
 sg13g2_nand2_1 _26311_ (.Y(_07233_),
    .A(_07157_),
    .B(_07155_));
 sg13g2_inv_1 _26312_ (.Y(_07234_),
    .A(_07233_));
 sg13g2_nor4_1 _26313_ (.A(net1071),
    .B(_07158_),
    .C(_07155_),
    .D(_09743_),
    .Y(_07235_));
 sg13g2_o21ai_1 _26314_ (.B1(_07160_),
    .Y(_07236_),
    .A1(_07234_),
    .A2(_07235_));
 sg13g2_nor4_1 _26315_ (.A(_07160_),
    .B(net1071),
    .C(_07158_),
    .D(_07155_),
    .Y(_07237_));
 sg13g2_nand2_1 _26316_ (.Y(_07238_),
    .A(_07166_),
    .B(_07237_));
 sg13g2_buf_1 _26317_ (.A(_07158_),
    .X(_07239_));
 sg13g2_nor2b_1 _26318_ (.A(_09743_),
    .B_N(net1071),
    .Y(_07240_));
 sg13g2_o21ai_1 _26319_ (.B1(_07155_),
    .Y(_07241_),
    .A1(net921),
    .A2(_07240_));
 sg13g2_nand3_1 _26320_ (.B(_07238_),
    .C(_07241_),
    .A(_07236_),
    .Y(_07242_));
 sg13g2_nor2b_1 _26321_ (.A(_07155_),
    .B_N(_07166_),
    .Y(_07243_));
 sg13g2_nor2_1 _26322_ (.A(_07161_),
    .B(net1071),
    .Y(_07244_));
 sg13g2_a22oi_1 _26323_ (.Y(_07245_),
    .B1(_07243_),
    .B2(_07244_),
    .A2(_07234_),
    .A1(_07161_));
 sg13g2_nor3_1 _26324_ (.A(net921),
    .B(_07153_),
    .C(_07245_),
    .Y(_07246_));
 sg13g2_xor2_1 _26325_ (.B(_07159_),
    .A(net924),
    .X(_07247_));
 sg13g2_o21ai_1 _26326_ (.B1(net901),
    .Y(_07248_),
    .A1(_09744_),
    .A2(_07247_));
 sg13g2_nor3_2 _26327_ (.A(_07242_),
    .B(_07246_),
    .C(_07248_),
    .Y(_07249_));
 sg13g2_and2_1 _26328_ (.A(_07160_),
    .B(net1071),
    .X(_07250_));
 sg13g2_buf_1 _26329_ (.A(_07250_),
    .X(_07251_));
 sg13g2_o21ai_1 _26330_ (.B1(net924),
    .Y(_07252_),
    .A1(_07239_),
    .A2(_07251_));
 sg13g2_nor2b_1 _26331_ (.A(_07237_),
    .B_N(_07252_),
    .Y(_07253_));
 sg13g2_nand3_1 _26332_ (.B(_07249_),
    .C(_07253_),
    .A(_07151_),
    .Y(_07254_));
 sg13g2_o21ai_1 _26333_ (.B1(_07254_),
    .Y(_07255_),
    .A1(_07151_),
    .A2(_07249_));
 sg13g2_inv_1 _26334_ (.Y(_02643_),
    .A(_07255_));
 sg13g2_nand2_1 _26335_ (.Y(_07256_),
    .A(_07151_),
    .B(_07253_));
 sg13g2_nand2_1 _26336_ (.Y(_07257_),
    .A(_07249_),
    .B(_07256_));
 sg13g2_nand2_1 _26337_ (.Y(_07258_),
    .A(\cpu.uart.r_rcnt[1] ),
    .B(_07257_));
 sg13g2_nand3_1 _26338_ (.B(_07249_),
    .C(_07253_),
    .A(_07152_),
    .Y(_07259_));
 sg13g2_nand2_1 _26339_ (.Y(_02644_),
    .A(_07258_),
    .B(_07259_));
 sg13g2_buf_1 _26340_ (.A(\cpu.gpio.genblk1[3].srcs_o[1] ),
    .X(_07260_));
 sg13g2_and2_1 _26341_ (.A(_07170_),
    .B(_07172_),
    .X(_07261_));
 sg13g2_buf_1 _26342_ (.A(_07261_),
    .X(_07262_));
 sg13g2_and2_1 _26343_ (.A(_07183_),
    .B(_07262_),
    .X(_07263_));
 sg13g2_buf_1 _26344_ (.A(_07263_),
    .X(_07264_));
 sg13g2_nor4_1 _26345_ (.A(net778),
    .B(_07190_),
    .C(_07186_),
    .D(_07264_),
    .Y(_07265_));
 sg13g2_nand2_1 _26346_ (.Y(_07266_),
    .A(\cpu.uart.r_out[0] ),
    .B(_07209_));
 sg13g2_xor2_1 _26347_ (.B(_07266_),
    .A(\cpu.uart.r_x_invert ),
    .X(_07267_));
 sg13g2_nor2_1 _26348_ (.A(_00259_),
    .B(_07265_),
    .Y(_07268_));
 sg13g2_a21oi_1 _26349_ (.A1(_07265_),
    .A2(_07267_),
    .Y(_07269_),
    .B1(_07268_));
 sg13g2_nor2_2 _26350_ (.A(_07181_),
    .B(_07191_),
    .Y(_07270_));
 sg13g2_nor2b_1 _26351_ (.A(_07170_),
    .B_N(_07172_),
    .Y(_07271_));
 sg13g2_nor2_1 _26352_ (.A(_07188_),
    .B(_07271_),
    .Y(_07272_));
 sg13g2_a22oi_1 _26353_ (.Y(_07273_),
    .B1(_07272_),
    .B2(_07176_),
    .A2(_07184_),
    .A1(_09743_));
 sg13g2_nor2_1 _26354_ (.A(net1070),
    .B(_07273_),
    .Y(_07274_));
 sg13g2_a21oi_1 _26355_ (.A1(_07195_),
    .A2(_07199_),
    .Y(_07275_),
    .B1(net922));
 sg13g2_nor3_1 _26356_ (.A(_07202_),
    .B(_07274_),
    .C(_07275_),
    .Y(_07276_));
 sg13g2_o21ai_1 _26357_ (.B1(net783),
    .Y(_07277_),
    .A1(_07270_),
    .A2(_07276_));
 sg13g2_mux2_1 _26358_ (.A0(net1068),
    .A1(_07269_),
    .S(_07277_),
    .X(_02649_));
 sg13g2_nand2_1 _26359_ (.Y(_07278_),
    .A(_07171_),
    .B(net922));
 sg13g2_o21ai_1 _26360_ (.B1(_07278_),
    .Y(_07279_),
    .A1(net1069),
    .A2(net252));
 sg13g2_nand2_1 _26361_ (.Y(_07280_),
    .A(net1070),
    .B(_07279_));
 sg13g2_o21ai_1 _26362_ (.B1(net252),
    .Y(_07281_),
    .A1(net1069),
    .A2(net923));
 sg13g2_a21o_1 _26363_ (.A2(_07190_),
    .A1(_07175_),
    .B1(_07264_),
    .X(_07282_));
 sg13g2_nand2b_1 _26364_ (.Y(_07283_),
    .B(net252),
    .A_N(_07197_));
 sg13g2_a21oi_1 _26365_ (.A1(net1069),
    .A2(_07262_),
    .Y(_07284_),
    .B1(net897));
 sg13g2_o21ai_1 _26366_ (.B1(_07284_),
    .Y(_07285_),
    .A1(net923),
    .A2(net252));
 sg13g2_a221oi_1 _26367_ (.B2(_07283_),
    .C1(_07285_),
    .B1(_07282_),
    .A1(_07207_),
    .Y(_07286_),
    .A2(_07281_));
 sg13g2_nand3b_1 _26368_ (.B(_07280_),
    .C(_07286_),
    .Y(_07287_),
    .A_N(_07270_));
 sg13g2_buf_1 _26369_ (.A(_07287_),
    .X(_07288_));
 sg13g2_nor2_1 _26370_ (.A(_07183_),
    .B(_07278_),
    .Y(_07289_));
 sg13g2_or2_1 _26371_ (.X(_07290_),
    .B(_07289_),
    .A(_07174_));
 sg13g2_inv_1 _26372_ (.Y(_07291_),
    .A(_07290_));
 sg13g2_nand2b_1 _26373_ (.Y(_07292_),
    .B(_07291_),
    .A_N(_07288_));
 sg13g2_nand2_1 _26374_ (.Y(_07293_),
    .A(_07196_),
    .B(_07292_));
 sg13g2_o21ai_1 _26375_ (.B1(_07293_),
    .Y(_02652_),
    .A1(_07196_),
    .A2(_07288_));
 sg13g2_a21o_1 _26376_ (.A2(_07291_),
    .A1(_07196_),
    .B1(_07288_),
    .X(_07294_));
 sg13g2_o21ai_1 _26377_ (.B1(\cpu.uart.r_xcnt[1] ),
    .Y(_07295_),
    .A1(_07196_),
    .A2(_07292_));
 sg13g2_o21ai_1 _26378_ (.B1(_07295_),
    .Y(_02653_),
    .A1(\cpu.uart.r_xcnt[1] ),
    .A2(_07294_));
 sg13g2_nor3_1 _26379_ (.A(_09046_),
    .B(net583),
    .C(net674),
    .Y(_07296_));
 sg13g2_buf_1 _26380_ (.A(_07296_),
    .X(_07297_));
 sg13g2_nand3_1 _26381_ (.B(_10008_),
    .C(_10013_),
    .A(_10002_),
    .Y(_07298_));
 sg13g2_nor3_1 _26382_ (.A(_09977_),
    .B(_10004_),
    .C(_07298_),
    .Y(_07299_));
 sg13g2_nand2_1 _26383_ (.Y(_07300_),
    .A(net130),
    .B(_09923_));
 sg13g2_buf_2 _26384_ (.A(_07300_),
    .X(_07301_));
 sg13g2_o21ai_1 _26385_ (.B1(_07301_),
    .Y(_07302_),
    .A1(net159),
    .A2(_07299_));
 sg13g2_nand2_1 _26386_ (.Y(_07303_),
    .A(_04916_),
    .B(_07302_));
 sg13g2_buf_1 _26387_ (.A(_09968_),
    .X(_07304_));
 sg13g2_nor2b_1 _26388_ (.A(_04916_),
    .B_N(_07299_),
    .Y(_07305_));
 sg13g2_a22oi_1 _26389_ (.Y(_07306_),
    .B1(_07305_),
    .B2(net101),
    .A2(_07304_),
    .A1(_09860_));
 sg13g2_nand2_1 _26390_ (.Y(_02439_),
    .A(_07303_),
    .B(_07306_));
 sg13g2_a21o_1 _26391_ (.A2(_07299_),
    .A1(_04916_),
    .B1(net159),
    .X(_07307_));
 sg13g2_a21oi_1 _26392_ (.A1(_07301_),
    .A2(_07307_),
    .Y(_07308_),
    .B1(_05339_));
 sg13g2_nand2_1 _26393_ (.Y(_07309_),
    .A(_04916_),
    .B(_05339_));
 sg13g2_nor2_1 _26394_ (.A(_07298_),
    .B(_07309_),
    .Y(_07310_));
 sg13g2_nand2_1 _26395_ (.Y(_07311_),
    .A(_10009_),
    .B(_07310_));
 sg13g2_nor2_1 _26396_ (.A(net159),
    .B(_07311_),
    .Y(_07312_));
 sg13g2_nand2_1 _26397_ (.Y(_07313_),
    .A(net130),
    .B(net423));
 sg13g2_nor2_1 _26398_ (.A(net1018),
    .B(_07313_),
    .Y(_07314_));
 sg13g2_nor3_1 _26399_ (.A(_07308_),
    .B(_07312_),
    .C(_07314_),
    .Y(_02440_));
 sg13g2_a21oi_1 _26400_ (.A1(_09933_),
    .A2(_07311_),
    .Y(_07315_),
    .B1(_09925_));
 sg13g2_nor2_1 _26401_ (.A(_05388_),
    .B(_07315_),
    .Y(_07316_));
 sg13g2_a221oi_1 _26402_ (.B2(_05388_),
    .C1(_07316_),
    .B1(_07312_),
    .A1(_09883_),
    .Y(_02441_),
    .A2(_07304_));
 sg13g2_nand3_1 _26403_ (.B(_10005_),
    .C(_07310_),
    .A(_05388_),
    .Y(_07317_));
 sg13g2_buf_1 _26404_ (.A(_07317_),
    .X(_07318_));
 sg13g2_a21oi_1 _26405_ (.A1(_09933_),
    .A2(_07318_),
    .Y(_07319_),
    .B1(_09958_));
 sg13g2_nand2b_1 _26406_ (.Y(_07320_),
    .B(_07319_),
    .A_N(_05434_));
 sg13g2_o21ai_1 _26407_ (.B1(_05434_),
    .Y(_07321_),
    .A1(net159),
    .A2(_07318_));
 sg13g2_a22oi_1 _26408_ (.Y(_02442_),
    .B1(_07320_),
    .B2(_07321_),
    .A2(net86),
    .A1(net721));
 sg13g2_and4_1 _26409_ (.A(_05388_),
    .B(_05434_),
    .C(_10009_),
    .D(_07310_),
    .X(_07322_));
 sg13g2_and2_1 _26410_ (.A(_05555_),
    .B(_07322_),
    .X(_07323_));
 sg13g2_buf_1 _26411_ (.A(_07323_),
    .X(_07324_));
 sg13g2_or2_1 _26412_ (.X(_07325_),
    .B(_07322_),
    .A(_07297_));
 sg13g2_a21oi_1 _26413_ (.A1(_07301_),
    .A2(_07325_),
    .Y(_07326_),
    .B1(_05555_));
 sg13g2_a221oi_1 _26414_ (.B2(_09934_),
    .C1(_07326_),
    .B1(_07324_),
    .A1(net853),
    .Y(_02443_),
    .A2(net86));
 sg13g2_nand2_1 _26415_ (.Y(_07327_),
    .A(_05434_),
    .B(_05555_));
 sg13g2_nor2_1 _26416_ (.A(_07318_),
    .B(_07327_),
    .Y(_07328_));
 sg13g2_o21ai_1 _26417_ (.B1(_07301_),
    .Y(_07329_),
    .A1(_07297_),
    .A2(_07328_));
 sg13g2_nand2_1 _26418_ (.Y(_07330_),
    .A(net1073),
    .B(_07329_));
 sg13g2_nor3_1 _26419_ (.A(net1073),
    .B(_07318_),
    .C(_07327_),
    .Y(_07331_));
 sg13g2_a22oi_1 _26420_ (.Y(_07332_),
    .B1(_07331_),
    .B2(_09919_),
    .A2(_09968_),
    .A1(net1021));
 sg13g2_nand2_1 _26421_ (.Y(_02444_),
    .A(_07330_),
    .B(_07332_));
 sg13g2_inv_1 _26422_ (.Y(_07333_),
    .A(_05668_));
 sg13g2_nand2_1 _26423_ (.Y(_07334_),
    .A(net1073),
    .B(_07324_));
 sg13g2_a21oi_1 _26424_ (.A1(net101),
    .A2(_07334_),
    .Y(_07335_),
    .B1(net98));
 sg13g2_nor2_1 _26425_ (.A(_05668_),
    .B(_07334_),
    .Y(_07336_));
 sg13g2_a22oi_1 _26426_ (.Y(_07337_),
    .B1(_07336_),
    .B2(net101),
    .A2(_09968_),
    .A1(net1020));
 sg13g2_o21ai_1 _26427_ (.B1(_07337_),
    .Y(_02445_),
    .A1(_07333_),
    .A2(_07335_));
 sg13g2_and4_1 _26428_ (.A(net1073),
    .B(_05668_),
    .C(net99),
    .D(_07328_),
    .X(_07338_));
 sg13g2_nand3_1 _26429_ (.B(_05668_),
    .C(_07328_),
    .A(net1073),
    .Y(_07339_));
 sg13g2_a21oi_1 _26430_ (.A1(net99),
    .A2(_07339_),
    .Y(_07340_),
    .B1(_09925_));
 sg13g2_nor2_1 _26431_ (.A(_05115_),
    .B(_07340_),
    .Y(_07341_));
 sg13g2_a221oi_1 _26432_ (.B2(_05115_),
    .C1(_07341_),
    .B1(_07338_),
    .A1(net852),
    .Y(_02446_),
    .A2(net86));
 sg13g2_nand4_1 _26433_ (.B(_05668_),
    .C(_05115_),
    .A(net1073),
    .Y(_07342_),
    .D(_07324_));
 sg13g2_a21oi_1 _26434_ (.A1(_09918_),
    .A2(_07342_),
    .Y(_07343_),
    .B1(_09925_));
 sg13g2_nor2_1 _26435_ (.A(_05720_),
    .B(_07343_),
    .Y(_07344_));
 sg13g2_nand4_1 _26436_ (.B(_05668_),
    .C(_05115_),
    .A(net1073),
    .Y(_07345_),
    .D(_05720_));
 sg13g2_inv_1 _26437_ (.Y(_07346_),
    .A(_07345_));
 sg13g2_and2_1 _26438_ (.A(_07324_),
    .B(_07346_),
    .X(_07347_));
 sg13g2_buf_1 _26439_ (.A(_07347_),
    .X(_07348_));
 sg13g2_nor2b_1 _26440_ (.A(_07296_),
    .B_N(_07348_),
    .Y(_07349_));
 sg13g2_nor2_1 _26441_ (.A(_09975_),
    .B(_07313_),
    .Y(_07350_));
 sg13g2_nor3_1 _26442_ (.A(_07344_),
    .B(_07349_),
    .C(_07350_),
    .Y(_02447_));
 sg13g2_or2_1 _26443_ (.X(_07351_),
    .B(_07348_),
    .A(_07296_));
 sg13g2_a21oi_1 _26444_ (.A1(_07301_),
    .A2(_07351_),
    .Y(_07352_),
    .B1(_05733_));
 sg13g2_a221oi_1 _26445_ (.B2(_05733_),
    .C1(_07352_),
    .B1(_07349_),
    .A1(_12157_),
    .Y(_02448_),
    .A2(net86));
 sg13g2_a21o_1 _26446_ (.A2(_07348_),
    .A1(_05733_),
    .B1(net159),
    .X(_07353_));
 sg13g2_a21oi_1 _26447_ (.A1(_07301_),
    .A2(_07353_),
    .Y(_07354_),
    .B1(_05029_));
 sg13g2_nand3_1 _26448_ (.B(_05029_),
    .C(_07349_),
    .A(_05733_),
    .Y(_07355_));
 sg13g2_o21ai_1 _26449_ (.B1(_07355_),
    .Y(_07356_),
    .A1(_09986_),
    .A2(_07313_));
 sg13g2_nor2_1 _26450_ (.A(_07354_),
    .B(_07356_),
    .Y(_02449_));
 sg13g2_inv_1 _26451_ (.Y(_07357_),
    .A(_05154_));
 sg13g2_and4_1 _26452_ (.A(_05733_),
    .B(_05029_),
    .C(_07328_),
    .D(_07346_),
    .X(_07358_));
 sg13g2_buf_1 _26453_ (.A(_07358_),
    .X(_07359_));
 sg13g2_o21ai_1 _26454_ (.B1(_07301_),
    .Y(_07360_),
    .A1(net159),
    .A2(_07359_));
 sg13g2_nand3_1 _26455_ (.B(net99),
    .C(_07359_),
    .A(_05154_),
    .Y(_07361_));
 sg13g2_o21ai_1 _26456_ (.B1(_07361_),
    .Y(_07362_),
    .A1(_09991_),
    .A2(_07313_));
 sg13g2_a21oi_1 _26457_ (.A1(_07357_),
    .A2(_07360_),
    .Y(_02450_),
    .B1(_07362_));
 sg13g2_nand4_1 _26458_ (.B(_05029_),
    .C(_05154_),
    .A(_05733_),
    .Y(_07363_),
    .D(_07348_));
 sg13g2_a21oi_1 _26459_ (.A1(_09918_),
    .A2(_07363_),
    .Y(_07364_),
    .B1(_09925_));
 sg13g2_inv_1 _26460_ (.Y(_07365_),
    .A(_07363_));
 sg13g2_nand3_1 _26461_ (.B(net99),
    .C(_07365_),
    .A(_05178_),
    .Y(_07366_));
 sg13g2_o21ai_1 _26462_ (.B1(_07366_),
    .Y(_07367_),
    .A1(_05178_),
    .A2(_07364_));
 sg13g2_a21oi_1 _26463_ (.A1(_12060_),
    .A2(net86),
    .Y(_02451_),
    .B1(_07367_));
 sg13g2_nand3_1 _26464_ (.B(_05178_),
    .C(_07359_),
    .A(_05154_),
    .Y(_07368_));
 sg13g2_a21oi_1 _26465_ (.A1(_09918_),
    .A2(_07368_),
    .Y(_07369_),
    .B1(_09925_));
 sg13g2_inv_1 _26466_ (.Y(_07370_),
    .A(_07368_));
 sg13g2_nand3_1 _26467_ (.B(net99),
    .C(_07370_),
    .A(_05208_),
    .Y(_07371_));
 sg13g2_o21ai_1 _26468_ (.B1(_07371_),
    .Y(_07372_),
    .A1(_05208_),
    .A2(_07369_));
 sg13g2_a21oi_1 _26469_ (.A1(_12070_),
    .A2(net86),
    .Y(_02452_),
    .B1(_07372_));
 sg13g2_nand3_1 _26470_ (.B(_05208_),
    .C(_07365_),
    .A(_05178_),
    .Y(_07373_));
 sg13g2_a21oi_1 _26471_ (.A1(net99),
    .A2(_07373_),
    .Y(_07374_),
    .B1(net98));
 sg13g2_nand2b_1 _26472_ (.Y(_07375_),
    .B(_07374_),
    .A_N(_05231_));
 sg13g2_o21ai_1 _26473_ (.B1(_05231_),
    .Y(_07376_),
    .A1(net159),
    .A2(_07373_));
 sg13g2_a22oi_1 _26474_ (.Y(_02453_),
    .B1(_07375_),
    .B2(_07376_),
    .A2(net86),
    .A1(_12077_));
 sg13g2_nand3_1 _26475_ (.B(_05231_),
    .C(_07370_),
    .A(_05208_),
    .Y(_07377_));
 sg13g2_a21oi_1 _26476_ (.A1(net99),
    .A2(_07377_),
    .Y(_07378_),
    .B1(_09925_));
 sg13g2_nand2b_1 _26477_ (.Y(_07379_),
    .B(_07378_),
    .A_N(_05262_));
 sg13g2_o21ai_1 _26478_ (.B1(_05262_),
    .Y(_07380_),
    .A1(net159),
    .A2(_07377_));
 sg13g2_a22oi_1 _26479_ (.Y(_02454_),
    .B1(_07379_),
    .B2(_07380_),
    .A2(net86),
    .A1(_12084_));
 sg13g2_nor2_1 _26480_ (.A(\cpu.r_clk_invert ),
    .B(net684),
    .Y(_07381_));
 sg13g2_a21oi_1 _26481_ (.A1(_08987_),
    .A2(net684),
    .Y(_02521_),
    .B1(_07381_));
 sg13g2_nand2b_1 _26482_ (.Y(_07382_),
    .B(net901),
    .A_N(\cpu.d_flush_all ));
 sg13g2_buf_2 _26483_ (.A(_07382_),
    .X(_07383_));
 sg13g2_nor2b_1 _26484_ (.A(\cpu.dcache.r_valid[0] ),
    .B_N(_12145_),
    .Y(_07384_));
 sg13g2_nand4_1 _26485_ (.B(_03058_),
    .C(_12094_),
    .A(_09182_),
    .Y(_07385_),
    .D(_11993_));
 sg13g2_buf_2 _26486_ (.A(_07385_),
    .X(_07386_));
 sg13g2_nor2_1 _26487_ (.A(_12008_),
    .B(_07386_),
    .Y(_07387_));
 sg13g2_nor3_1 _26488_ (.A(_07383_),
    .B(_07384_),
    .C(_07387_),
    .Y(_00718_));
 sg13g2_nor2_1 _26489_ (.A(\cpu.dcache.r_valid[1] ),
    .B(net294),
    .Y(_07388_));
 sg13g2_nor2_1 _26490_ (.A(_12212_),
    .B(_07386_),
    .Y(_07389_));
 sg13g2_nor3_1 _26491_ (.A(_07383_),
    .B(_07388_),
    .C(_07389_),
    .Y(_00719_));
 sg13g2_nor2_1 _26492_ (.A(\cpu.dcache.r_valid[2] ),
    .B(net362),
    .Y(_07390_));
 sg13g2_nor2_1 _26493_ (.A(_12337_),
    .B(_07386_),
    .Y(_07391_));
 sg13g2_nor3_1 _26494_ (.A(_07383_),
    .B(_07390_),
    .C(_07391_),
    .Y(_00720_));
 sg13g2_nor2_1 _26495_ (.A(\cpu.dcache.r_valid[3] ),
    .B(net221),
    .Y(_07392_));
 sg13g2_nor2_1 _26496_ (.A(_12463_),
    .B(_07386_),
    .Y(_07393_));
 sg13g2_nor3_1 _26497_ (.A(_07383_),
    .B(_07392_),
    .C(_07393_),
    .Y(_00721_));
 sg13g2_inv_1 _26498_ (.Y(_07394_),
    .A(\cpu.dcache.r_valid[4] ));
 sg13g2_inv_1 _26499_ (.Y(_07395_),
    .A(_07386_));
 sg13g2_a221oi_1 _26500_ (.B2(_09916_),
    .C1(_07383_),
    .B1(_07395_),
    .A1(_07394_),
    .Y(_00722_),
    .A2(net412));
 sg13g2_nor2_1 _26501_ (.A(\cpu.dcache.r_valid[5] ),
    .B(net360),
    .Y(_07396_));
 sg13g2_nor2_1 _26502_ (.A(_02698_),
    .B(_07386_),
    .Y(_07397_));
 sg13g2_nor3_1 _26503_ (.A(_07383_),
    .B(_07396_),
    .C(_07397_),
    .Y(_00723_));
 sg13g2_nor2_1 _26504_ (.A(\cpu.dcache.r_valid[6] ),
    .B(_02895_),
    .Y(_07398_));
 sg13g2_nor2_1 _26505_ (.A(_02822_),
    .B(_07386_),
    .Y(_07399_));
 sg13g2_nor3_1 _26506_ (.A(_07383_),
    .B(_07398_),
    .C(_07399_),
    .Y(_00724_));
 sg13g2_nor2_1 _26507_ (.A(\cpu.dcache.r_valid[7] ),
    .B(_03011_),
    .Y(_07400_));
 sg13g2_nor2_1 _26508_ (.A(net672),
    .B(_07386_),
    .Y(_07401_));
 sg13g2_nor3_1 _26509_ (.A(_07383_),
    .B(_07400_),
    .C(_07401_),
    .Y(_00725_));
 sg13g2_nor3_1 _26510_ (.A(net1102),
    .B(net1015),
    .C(_10022_),
    .Y(_07402_));
 sg13g2_nand2_1 _26511_ (.Y(_07403_),
    .A(_04775_),
    .B(_07402_));
 sg13g2_buf_1 _26512_ (.A(_07403_),
    .X(_07404_));
 sg13g2_nand2_1 _26513_ (.Y(_07405_),
    .A(_08134_),
    .B(net474));
 sg13g2_o21ai_1 _26514_ (.B1(_07405_),
    .Y(_07406_),
    .A1(_03717_),
    .A2(net474));
 sg13g2_and3_1 _26515_ (.X(_00773_),
    .A(net290),
    .B(_09118_),
    .C(_07406_));
 sg13g2_and4_1 _26516_ (.A(_03598_),
    .B(_10205_),
    .C(\cpu.dec.do_flush_all ),
    .D(_11900_),
    .X(_00905_));
 sg13g2_and4_1 _26517_ (.A(net961),
    .B(_10327_),
    .C(\cpu.dec.do_flush_all ),
    .D(_11900_),
    .X(_00923_));
 sg13g2_nand2_1 _26518_ (.Y(_07407_),
    .A(net729),
    .B(_04003_));
 sg13g2_nor2_1 _26519_ (.A(net801),
    .B(net729),
    .Y(_07408_));
 sg13g2_a21oi_1 _26520_ (.A1(net290),
    .A2(_07407_),
    .Y(_07409_),
    .B1(_07408_));
 sg13g2_nor3_1 _26521_ (.A(_11503_),
    .B(_10722_),
    .C(_10371_),
    .Y(_07410_));
 sg13g2_nand3_1 _26522_ (.B(net729),
    .C(_07410_),
    .A(net961),
    .Y(_07411_));
 sg13g2_mux2_1 _26523_ (.A0(_10238_),
    .A1(_08966_),
    .S(_07411_),
    .X(_07412_));
 sg13g2_nor2_1 _26524_ (.A(_08190_),
    .B(net474),
    .Y(_07413_));
 sg13g2_a21oi_1 _26525_ (.A1(net474),
    .A2(_07412_),
    .Y(_07414_),
    .B1(_07413_));
 sg13g2_nor3_1 _26526_ (.A(_09124_),
    .B(_07409_),
    .C(_07414_),
    .Y(_00924_));
 sg13g2_nand3b_1 _26527_ (.B(_08180_),
    .C(net729),
    .Y(_07415_),
    .A_N(_00277_));
 sg13g2_nor2_1 _26528_ (.A(_11505_),
    .B(_08127_),
    .Y(_07416_));
 sg13g2_a21oi_1 _26529_ (.A1(_11494_),
    .A2(net291),
    .Y(_07417_),
    .B1(_04832_));
 sg13g2_o21ai_1 _26530_ (.B1(_09655_),
    .Y(_07418_),
    .A1(_09122_),
    .A2(net643));
 sg13g2_nand2_1 _26531_ (.Y(_07419_),
    .A(_08129_),
    .B(_07418_));
 sg13g2_nand2_1 _26532_ (.Y(_07420_),
    .A(net783),
    .B(_07419_));
 sg13g2_a221oi_1 _26533_ (.B2(_07417_),
    .C1(_07420_),
    .B1(_07416_),
    .A1(_08128_),
    .Y(_01042_),
    .A2(_07415_));
 sg13g2_a21o_1 _26534_ (.A2(net291),
    .A1(_11494_),
    .B1(_04832_),
    .X(_07421_));
 sg13g2_nor2_1 _26535_ (.A(_11505_),
    .B(_08125_),
    .Y(_07422_));
 sg13g2_a221oi_1 _26536_ (.B2(_07422_),
    .C1(_07420_),
    .B1(_07421_),
    .A1(_08126_),
    .Y(_01043_),
    .A2(_07415_));
 sg13g2_inv_1 _26537_ (.Y(_07423_),
    .A(\cpu.icache.r_valid[0] ));
 sg13g2_nand2b_1 _26538_ (.Y(_07424_),
    .B(_08963_),
    .A_N(\cpu.ex.i_flush_all ));
 sg13g2_buf_2 _26539_ (.A(_07424_),
    .X(_07425_));
 sg13g2_a21oi_1 _26540_ (.A1(_07423_),
    .A2(net309),
    .Y(_02398_),
    .B1(_07425_));
 sg13g2_nor2_1 _26541_ (.A(\cpu.icache.r_valid[1] ),
    .B(_06333_),
    .Y(_07426_));
 sg13g2_nor2_1 _26542_ (.A(_07425_),
    .B(_07426_),
    .Y(_02399_));
 sg13g2_nor2_1 _26543_ (.A(\cpu.icache.r_valid[2] ),
    .B(_06350_),
    .Y(_07427_));
 sg13g2_nor2_1 _26544_ (.A(_07425_),
    .B(_07427_),
    .Y(_02400_));
 sg13g2_inv_1 _26545_ (.Y(_07428_),
    .A(\cpu.icache.r_valid[3] ));
 sg13g2_a21oi_1 _26546_ (.A1(_07428_),
    .A2(net235),
    .Y(_02401_),
    .B1(_07425_));
 sg13g2_nor2_1 _26547_ (.A(\cpu.icache.r_valid[4] ),
    .B(_06375_),
    .Y(_07429_));
 sg13g2_nor2_1 _26548_ (.A(_07425_),
    .B(_07429_),
    .Y(_02402_));
 sg13g2_nor2_1 _26549_ (.A(\cpu.icache.r_valid[5] ),
    .B(_06390_),
    .Y(_07430_));
 sg13g2_nor2_1 _26550_ (.A(_07425_),
    .B(_07430_),
    .Y(_02403_));
 sg13g2_inv_1 _26551_ (.Y(_07431_),
    .A(\cpu.icache.r_valid[6] ));
 sg13g2_a21oi_1 _26552_ (.A1(_07431_),
    .A2(_06399_),
    .Y(_02404_),
    .B1(_07425_));
 sg13g2_nor2_1 _26553_ (.A(\cpu.icache.r_valid[7] ),
    .B(_06410_),
    .Y(_07432_));
 sg13g2_nor2_1 _26554_ (.A(_07425_),
    .B(_07432_),
    .Y(_02405_));
 sg13g2_nand3_1 _26555_ (.B(net130),
    .C(net355),
    .A(net1106),
    .Y(_07433_));
 sg13g2_nand2_1 _26556_ (.Y(_07434_),
    .A(_08975_),
    .B(_07433_));
 sg13g2_nand3_1 _26557_ (.B(net130),
    .C(net357),
    .A(net1106),
    .Y(_07435_));
 sg13g2_a21oi_1 _26558_ (.A1(_07434_),
    .A2(_07435_),
    .Y(_00294_),
    .B1(net556));
 sg13g2_nor2_1 _26559_ (.A(_03058_),
    .B(net1086),
    .Y(_07436_));
 sg13g2_nor2b_1 _26560_ (.A(_07436_),
    .B_N(_00292_),
    .Y(_00563_));
 sg13g2_nor2_1 _26561_ (.A(_12014_),
    .B(_12053_),
    .Y(_07437_));
 sg13g2_nor2_1 _26562_ (.A(_07436_),
    .B(_07437_),
    .Y(_00564_));
 sg13g2_xor2_1 _26563_ (.B(_11993_),
    .A(net991),
    .X(_07438_));
 sg13g2_nor2_1 _26564_ (.A(_07436_),
    .B(_07438_),
    .Y(_00565_));
 sg13g2_nor2_1 _26565_ (.A(_09052_),
    .B(net474),
    .Y(_07439_));
 sg13g2_a21oi_1 _26566_ (.A1(net920),
    .A2(_07404_),
    .Y(_07440_),
    .B1(_07439_));
 sg13g2_nor2_1 _26567_ (.A(net607),
    .B(_07440_),
    .Y(_00774_));
 sg13g2_a21oi_2 _26568_ (.B1(net214),
    .Y(_07441_),
    .A2(_04128_),
    .A1(_11497_));
 sg13g2_and2_1 _26569_ (.A(net789),
    .B(_07441_),
    .X(_07442_));
 sg13g2_nor2_1 _26570_ (.A(_10181_),
    .B(_09144_),
    .Y(_07443_));
 sg13g2_a21oi_1 _26571_ (.A1(_07410_),
    .A2(_07443_),
    .Y(_07444_),
    .B1(net789));
 sg13g2_nor2_1 _26572_ (.A(_09122_),
    .B(_07444_),
    .Y(_07445_));
 sg13g2_nor2_1 _26573_ (.A(_03700_),
    .B(_07445_),
    .Y(_07446_));
 sg13g2_nor2_1 _26574_ (.A(_10181_),
    .B(_07446_),
    .Y(_07447_));
 sg13g2_a21oi_1 _26575_ (.A1(_08190_),
    .A2(_07446_),
    .Y(_07448_),
    .B1(_07447_));
 sg13g2_nor2_1 _26576_ (.A(_07441_),
    .B(_07448_),
    .Y(_07449_));
 sg13g2_buf_1 _26577_ (.A(net783),
    .X(_07450_));
 sg13g2_o21ai_1 _26578_ (.B1(_07450_),
    .Y(_00775_),
    .A1(_07442_),
    .A2(_07449_));
 sg13g2_mux2_1 _26579_ (.A0(net965),
    .A1(_10753_),
    .S(net474),
    .X(_07451_));
 sg13g2_and2_1 _26580_ (.A(_08965_),
    .B(_07451_),
    .X(_00776_));
 sg13g2_o21ai_1 _26581_ (.B1(_06763_),
    .Y(_07452_),
    .A1(_08260_),
    .A2(_08923_));
 sg13g2_nor3_1 _26582_ (.A(\cpu.ex.r_branch_stall ),
    .B(_11495_),
    .C(_03590_),
    .Y(_07453_));
 sg13g2_nand3_1 _26583_ (.B(net729),
    .C(_07453_),
    .A(_08180_),
    .Y(_07454_));
 sg13g2_nand3_1 _26584_ (.B(_07419_),
    .C(_07454_),
    .A(_11621_),
    .Y(_07455_));
 sg13g2_nand3_1 _26585_ (.B(_11502_),
    .C(_07455_),
    .A(net1119),
    .Y(_07456_));
 sg13g2_a21o_1 _26586_ (.A2(_07456_),
    .A1(net68),
    .B1(_06763_),
    .X(_07457_));
 sg13g2_nand3_1 _26587_ (.B(_07452_),
    .C(_07457_),
    .A(_08965_),
    .Y(_00921_));
 sg13g2_nand2_1 _26588_ (.Y(_07458_),
    .A(_09182_),
    .B(net1031));
 sg13g2_nand3_1 _26589_ (.B(\cpu.dec.do_flush_write ),
    .C(_04132_),
    .A(net961),
    .Y(_07459_));
 sg13g2_a21oi_1 _26590_ (.A1(_07458_),
    .A2(_07459_),
    .Y(_00922_),
    .B1(net556));
 sg13g2_nand2_1 _26591_ (.Y(_07460_),
    .A(\cpu.dec.io ),
    .B(_04132_));
 sg13g2_nand2_1 _26592_ (.Y(_07461_),
    .A(_03057_),
    .B(net1031));
 sg13g2_a21oi_1 _26593_ (.A1(_07460_),
    .A2(_07461_),
    .Y(_00925_),
    .B1(_06674_));
 sg13g2_nor2_1 _26594_ (.A(net673),
    .B(net474),
    .Y(_07462_));
 sg13g2_a21oi_1 _26595_ (.A1(_10238_),
    .A2(net474),
    .Y(_07463_),
    .B1(_07462_));
 sg13g2_mux2_1 _26596_ (.A0(_07463_),
    .A1(_08967_),
    .S(_07441_),
    .X(_07464_));
 sg13g2_nor2_1 _26597_ (.A(net607),
    .B(_07464_),
    .Y(_00972_));
 sg13g2_inv_1 _26598_ (.Y(_07465_),
    .A(_11528_));
 sg13g2_a22oi_1 _26599_ (.Y(_07466_),
    .B1(_07465_),
    .B2(net1122),
    .A2(_04132_),
    .A1(_11495_));
 sg13g2_nor2_1 _26600_ (.A(net607),
    .B(_07466_),
    .Y(_00973_));
 sg13g2_nor2_2 _26601_ (.A(_08189_),
    .B(_05813_),
    .Y(_07467_));
 sg13g2_mux2_1 _26602_ (.A0(_10382_),
    .A1(_09106_),
    .S(_07467_),
    .X(_07468_));
 sg13g2_nand2_1 _26603_ (.Y(_07469_),
    .A(net290),
    .B(_07468_));
 sg13g2_a21oi_1 _26604_ (.A1(_11497_),
    .A2(_07469_),
    .Y(_01048_),
    .B1(_06674_));
 sg13g2_mux2_1 _26605_ (.A0(_10080_),
    .A1(_11988_),
    .S(_07467_),
    .X(_07470_));
 sg13g2_nand2_1 _26606_ (.Y(_07471_),
    .A(_04439_),
    .B(_07470_));
 sg13g2_o21ai_1 _26607_ (.B1(_07471_),
    .Y(_07472_),
    .A1(_09183_),
    .A2(_04439_));
 sg13g2_nor2_1 _26608_ (.A(net607),
    .B(_07472_),
    .Y(_01049_));
 sg13g2_nand2_1 _26609_ (.Y(_07473_),
    .A(net575),
    .B(_07467_));
 sg13g2_o21ai_1 _26610_ (.B1(_07473_),
    .Y(_07474_),
    .A1(_10232_),
    .A2(_07467_));
 sg13g2_nor2_1 _26611_ (.A(_08131_),
    .B(_10119_),
    .Y(_07475_));
 sg13g2_a21oi_1 _26612_ (.A1(_08220_),
    .A2(_07474_),
    .Y(_07476_),
    .B1(_07475_));
 sg13g2_nor2_1 _26613_ (.A(net607),
    .B(_07476_),
    .Y(_01050_));
 sg13g2_nand2_1 _26614_ (.Y(_07477_),
    .A(_00267_),
    .B(_05902_));
 sg13g2_nor4_2 _26615_ (.A(net944),
    .B(net950),
    .C(net948),
    .Y(_07478_),
    .D(_07477_));
 sg13g2_nor2b_1 _26616_ (.A(_00235_),
    .B_N(_05798_),
    .Y(_07479_));
 sg13g2_o21ai_1 _26617_ (.B1(_07479_),
    .Y(_07480_),
    .A1(_08190_),
    .A2(_00233_));
 sg13g2_a21o_1 _26618_ (.A2(_07480_),
    .A1(_05797_),
    .B1(_11496_),
    .X(_07481_));
 sg13g2_buf_1 _26619_ (.A(_07481_),
    .X(_07482_));
 sg13g2_nand2b_1 _26620_ (.Y(_07483_),
    .B(_05797_),
    .A_N(_07482_));
 sg13g2_buf_1 _26621_ (.A(_07483_),
    .X(_07484_));
 sg13g2_a21oi_1 _26622_ (.A1(_03465_),
    .A2(_10205_),
    .Y(_07485_),
    .B1(_05797_));
 sg13g2_nor2_1 _26623_ (.A(_07482_),
    .B(_07485_),
    .Y(_07486_));
 sg13g2_buf_2 _26624_ (.A(_07486_),
    .X(_07487_));
 sg13g2_o21ai_1 _26625_ (.B1(_07487_),
    .Y(_07488_),
    .A1(_07478_),
    .A2(net158));
 sg13g2_nor2_1 _26626_ (.A(_09875_),
    .B(net158),
    .Y(_07489_));
 sg13g2_buf_2 _26627_ (.A(_07489_),
    .X(_07490_));
 sg13g2_buf_1 _26628_ (.A(_07490_),
    .X(_07491_));
 sg13g2_a22oi_1 _26629_ (.Y(_07492_),
    .B1(net85),
    .B2(_07478_),
    .A2(_07488_),
    .A1(\cpu.genblk1.mmu.r_valid_d[0] ));
 sg13g2_nor2_1 _26630_ (.A(_09130_),
    .B(_07492_),
    .Y(_01051_));
 sg13g2_nor3_2 _26631_ (.A(net827),
    .B(_11985_),
    .C(net708),
    .Y(_07493_));
 sg13g2_nor2_1 _26632_ (.A(_11188_),
    .B(_07477_),
    .Y(_07494_));
 sg13g2_a21oi_1 _26633_ (.A1(net1072),
    .A2(_05902_),
    .Y(_07495_),
    .B1(_05837_));
 sg13g2_a21o_1 _26634_ (.A2(_07494_),
    .A1(net950),
    .B1(_07495_),
    .X(_07496_));
 sg13g2_a22oi_1 _26635_ (.Y(_07497_),
    .B1(_07496_),
    .B2(_10080_),
    .A2(_07494_),
    .A1(_05914_));
 sg13g2_buf_2 _26636_ (.A(_07497_),
    .X(_07498_));
 sg13g2_nor2_2 _26637_ (.A(net158),
    .B(_07498_),
    .Y(_07499_));
 sg13g2_buf_1 _26638_ (.A(net158),
    .X(_07500_));
 sg13g2_buf_1 _26639_ (.A(_07487_),
    .X(_07501_));
 sg13g2_o21ai_1 _26640_ (.B1(net125),
    .Y(_07502_),
    .A1(_05868_),
    .A2(_07500_));
 sg13g2_a22oi_1 _26641_ (.Y(_07503_),
    .B1(_07502_),
    .B2(\cpu.genblk1.mmu.r_valid_d[10] ),
    .A2(_07499_),
    .A1(_07493_));
 sg13g2_nor2_1 _26642_ (.A(_09130_),
    .B(_07503_),
    .Y(_01052_));
 sg13g2_buf_1 _26643_ (.A(_09129_),
    .X(_07504_));
 sg13g2_o21ai_1 _26644_ (.B1(net125),
    .Y(_07505_),
    .A1(_05873_),
    .A2(net126));
 sg13g2_a22oi_1 _26645_ (.Y(_07506_),
    .B1(_07505_),
    .B2(\cpu.genblk1.mmu.r_valid_d[11] ),
    .A2(_07490_),
    .A1(_05873_));
 sg13g2_nor2_1 _26646_ (.A(net553),
    .B(_07506_),
    .Y(_01053_));
 sg13g2_nand2_1 _26647_ (.Y(_07507_),
    .A(_05824_),
    .B(_04844_));
 sg13g2_nor3_1 _26648_ (.A(_05816_),
    .B(net951),
    .C(_07507_),
    .Y(_07508_));
 sg13g2_buf_2 _26649_ (.A(_07508_),
    .X(_07509_));
 sg13g2_nor3_1 _26650_ (.A(_05816_),
    .B(_05811_),
    .C(_05823_),
    .Y(_07510_));
 sg13g2_o21ai_1 _26651_ (.B1(net1072),
    .Y(_07511_),
    .A1(_05827_),
    .A2(_07510_));
 sg13g2_buf_1 _26652_ (.A(_07511_),
    .X(_07512_));
 sg13g2_nor2_1 _26653_ (.A(_07498_),
    .B(_07512_),
    .Y(_07513_));
 sg13g2_o21ai_1 _26654_ (.B1(net125),
    .Y(_07514_),
    .A1(net126),
    .A2(_07513_));
 sg13g2_a22oi_1 _26655_ (.Y(_07515_),
    .B1(_07514_),
    .B2(\cpu.genblk1.mmu.r_valid_d[12] ),
    .A2(_07509_),
    .A1(_07499_));
 sg13g2_nor2_1 _26656_ (.A(net553),
    .B(_07515_),
    .Y(_01054_));
 sg13g2_or2_1 _26657_ (.X(_07516_),
    .B(_05885_),
    .A(_05823_));
 sg13g2_buf_1 _26658_ (.A(_07516_),
    .X(_07517_));
 sg13g2_nor2_2 _26659_ (.A(_07498_),
    .B(_07517_),
    .Y(_07518_));
 sg13g2_o21ai_1 _26660_ (.B1(net125),
    .Y(_07519_),
    .A1(net126),
    .A2(_07518_));
 sg13g2_a22oi_1 _26661_ (.Y(_07520_),
    .B1(_07519_),
    .B2(\cpu.genblk1.mmu.r_valid_d[13] ),
    .A2(_07518_),
    .A1(_07491_));
 sg13g2_nor2_1 _26662_ (.A(_07504_),
    .B(_07520_),
    .Y(_01055_));
 sg13g2_nor2_1 _26663_ (.A(net708),
    .B(_07507_),
    .Y(_07521_));
 sg13g2_buf_2 _26664_ (.A(_07521_),
    .X(_07522_));
 sg13g2_nor2_1 _26665_ (.A(_06010_),
    .B(_07498_),
    .Y(_07523_));
 sg13g2_o21ai_1 _26666_ (.B1(net125),
    .Y(_07524_),
    .A1(net126),
    .A2(_07523_));
 sg13g2_a22oi_1 _26667_ (.Y(_07525_),
    .B1(_07524_),
    .B2(\cpu.genblk1.mmu.r_valid_d[14] ),
    .A2(_07522_),
    .A1(_07499_));
 sg13g2_nor2_1 _26668_ (.A(net553),
    .B(_07525_),
    .Y(_01056_));
 sg13g2_nor2_2 _26669_ (.A(_05839_),
    .B(_07498_),
    .Y(_07526_));
 sg13g2_o21ai_1 _26670_ (.B1(net125),
    .Y(_07527_),
    .A1(_07500_),
    .A2(_07526_));
 sg13g2_a22oi_1 _26671_ (.Y(_07528_),
    .B1(_07527_),
    .B2(\cpu.genblk1.mmu.r_valid_d[15] ),
    .A2(_07526_),
    .A1(_07491_));
 sg13g2_nor2_1 _26672_ (.A(net553),
    .B(_07528_),
    .Y(_01057_));
 sg13g2_a21oi_1 _26673_ (.A1(_05803_),
    .A2(_05851_),
    .Y(_07529_),
    .B1(_11985_));
 sg13g2_and2_1 _26674_ (.A(_06072_),
    .B(_07529_),
    .X(_07530_));
 sg13g2_buf_1 _26675_ (.A(_07530_),
    .X(_07531_));
 sg13g2_nor2_1 _26676_ (.A(_10327_),
    .B(_05795_),
    .Y(_07532_));
 sg13g2_nor2b_1 _26677_ (.A(_07532_),
    .B_N(_03465_),
    .Y(_07533_));
 sg13g2_buf_1 _26678_ (.A(_07533_),
    .X(_07534_));
 sg13g2_buf_1 _26679_ (.A(net552),
    .X(_07535_));
 sg13g2_o21ai_1 _26680_ (.B1(_05839_),
    .Y(_07536_),
    .A1(_05851_),
    .A2(_05903_));
 sg13g2_nand2_1 _26681_ (.Y(_07537_),
    .A(net1072),
    .B(_07536_));
 sg13g2_nor2_1 _26682_ (.A(_07498_),
    .B(_07537_),
    .Y(_07538_));
 sg13g2_a21oi_1 _26683_ (.A1(_03465_),
    .A2(_10458_),
    .Y(_07539_),
    .B1(_05797_));
 sg13g2_nor2_1 _26684_ (.A(_07482_),
    .B(_07539_),
    .Y(_07540_));
 sg13g2_buf_2 _26685_ (.A(_07540_),
    .X(_07541_));
 sg13g2_buf_1 _26686_ (.A(_07541_),
    .X(_07542_));
 sg13g2_o21ai_1 _26687_ (.B1(net124),
    .Y(_07543_),
    .A1(net473),
    .A2(_07538_));
 sg13g2_a22oi_1 _26688_ (.Y(_07544_),
    .B1(_07543_),
    .B2(\cpu.genblk1.mmu.r_valid_d[16] ),
    .A2(_07531_),
    .A1(_07499_));
 sg13g2_nor2_1 _26689_ (.A(net553),
    .B(_07544_),
    .Y(_01058_));
 sg13g2_nor4_1 _26690_ (.A(_10079_),
    .B(net950),
    .C(net948),
    .D(net1072),
    .Y(_07545_));
 sg13g2_nand3_1 _26691_ (.B(net948),
    .C(net1072),
    .A(net944),
    .Y(_07546_));
 sg13g2_nand2b_1 _26692_ (.Y(_07547_),
    .B(_07546_),
    .A_N(_07545_));
 sg13g2_nand2b_1 _26693_ (.Y(_07548_),
    .B(net950),
    .A_N(net1072));
 sg13g2_a21oi_1 _26694_ (.A1(_05902_),
    .A2(_07548_),
    .Y(_07549_),
    .B1(_05913_));
 sg13g2_a22oi_1 _26695_ (.Y(_07550_),
    .B1(_07549_),
    .B2(_05951_),
    .A2(_07547_),
    .A1(_05902_));
 sg13g2_buf_1 _26696_ (.A(_07550_),
    .X(_07551_));
 sg13g2_nor3_2 _26697_ (.A(net827),
    .B(_05885_),
    .C(net551),
    .Y(_07552_));
 sg13g2_o21ai_1 _26698_ (.B1(net124),
    .Y(_07553_),
    .A1(net473),
    .A2(_07552_));
 sg13g2_a22oi_1 _26699_ (.Y(_07554_),
    .B1(_07553_),
    .B2(\cpu.genblk1.mmu.r_valid_d[17] ),
    .A2(_07552_),
    .A1(net85));
 sg13g2_nor2_1 _26700_ (.A(net553),
    .B(_07554_),
    .Y(_01059_));
 sg13g2_nor2_1 _26701_ (.A(net552),
    .B(_07482_),
    .Y(_07555_));
 sg13g2_buf_2 _26702_ (.A(_07555_),
    .X(_07556_));
 sg13g2_nor2b_1 _26703_ (.A(net551),
    .B_N(_07493_),
    .Y(_07557_));
 sg13g2_o21ai_1 _26704_ (.B1(net124),
    .Y(_07558_),
    .A1(net473),
    .A2(_05916_));
 sg13g2_a22oi_1 _26705_ (.Y(_07559_),
    .B1(_07558_),
    .B2(\cpu.genblk1.mmu.r_valid_d[18] ),
    .A2(_07557_),
    .A1(_07556_));
 sg13g2_nor2_1 _26706_ (.A(net553),
    .B(_07559_),
    .Y(_01060_));
 sg13g2_o21ai_1 _26707_ (.B1(net124),
    .Y(_07560_),
    .A1(net473),
    .A2(_05925_));
 sg13g2_a22oi_1 _26708_ (.Y(_07561_),
    .B1(_07560_),
    .B2(\cpu.genblk1.mmu.r_valid_d[19] ),
    .A2(_07490_),
    .A1(_05925_));
 sg13g2_nor2_1 _26709_ (.A(net553),
    .B(_07561_),
    .Y(_01061_));
 sg13g2_nor2_1 _26710_ (.A(_05913_),
    .B(net1072),
    .Y(_07562_));
 sg13g2_a22oi_1 _26711_ (.Y(_07563_),
    .B1(_05914_),
    .B2(_07562_),
    .A2(_05878_),
    .A1(net1072));
 sg13g2_inv_1 _26712_ (.Y(_07564_),
    .A(_07563_));
 sg13g2_a22oi_1 _26713_ (.Y(_07565_),
    .B1(_07564_),
    .B2(_05902_),
    .A2(_07549_),
    .A1(_10080_));
 sg13g2_buf_1 _26714_ (.A(_07565_),
    .X(_07566_));
 sg13g2_nor3_2 _26715_ (.A(_05828_),
    .B(_05885_),
    .C(net472),
    .Y(_07567_));
 sg13g2_o21ai_1 _26716_ (.B1(_07501_),
    .Y(_07568_),
    .A1(net126),
    .A2(_07567_));
 sg13g2_a22oi_1 _26717_ (.Y(_07569_),
    .B1(_07568_),
    .B2(\cpu.genblk1.mmu.r_valid_d[1] ),
    .A2(_07567_),
    .A1(net85));
 sg13g2_nor2_1 _26718_ (.A(_07504_),
    .B(_07569_),
    .Y(_01062_));
 sg13g2_buf_1 _26719_ (.A(_09129_),
    .X(_07570_));
 sg13g2_inv_1 _26720_ (.Y(_07571_),
    .A(_07551_));
 sg13g2_and2_1 _26721_ (.A(_07556_),
    .B(_07509_),
    .X(_07572_));
 sg13g2_buf_1 _26722_ (.A(_07572_),
    .X(_07573_));
 sg13g2_nor2_1 _26723_ (.A(_07512_),
    .B(net551),
    .Y(_07574_));
 sg13g2_o21ai_1 _26724_ (.B1(net124),
    .Y(_07575_),
    .A1(net473),
    .A2(_07574_));
 sg13g2_a22oi_1 _26725_ (.Y(_07576_),
    .B1(_07575_),
    .B2(\cpu.genblk1.mmu.r_valid_d[20] ),
    .A2(_07573_),
    .A1(_07571_));
 sg13g2_nor2_1 _26726_ (.A(net550),
    .B(_07576_),
    .Y(_01063_));
 sg13g2_nor2_2 _26727_ (.A(_07517_),
    .B(net551),
    .Y(_07577_));
 sg13g2_o21ai_1 _26728_ (.B1(net124),
    .Y(_07578_),
    .A1(net473),
    .A2(_07577_));
 sg13g2_a22oi_1 _26729_ (.Y(_07579_),
    .B1(_07578_),
    .B2(\cpu.genblk1.mmu.r_valid_d[21] ),
    .A2(_07577_),
    .A1(net85));
 sg13g2_nor2_1 _26730_ (.A(net550),
    .B(_07579_),
    .Y(_01064_));
 sg13g2_nor4_1 _26731_ (.A(net552),
    .B(net708),
    .C(_07482_),
    .D(_07507_),
    .Y(_07580_));
 sg13g2_nor2_1 _26732_ (.A(_06010_),
    .B(net551),
    .Y(_07581_));
 sg13g2_o21ai_1 _26733_ (.B1(net124),
    .Y(_07582_),
    .A1(net473),
    .A2(_07581_));
 sg13g2_a22oi_1 _26734_ (.Y(_07583_),
    .B1(_07582_),
    .B2(\cpu.genblk1.mmu.r_valid_d[22] ),
    .A2(_07580_),
    .A1(_07571_));
 sg13g2_nor2_1 _26735_ (.A(net550),
    .B(_07583_),
    .Y(_01065_));
 sg13g2_nor2_2 _26736_ (.A(_05839_),
    .B(_05900_),
    .Y(_07584_));
 sg13g2_o21ai_1 _26737_ (.B1(net124),
    .Y(_07585_),
    .A1(net473),
    .A2(_07584_));
 sg13g2_a22oi_1 _26738_ (.Y(_07586_),
    .B1(_07585_),
    .B2(\cpu.genblk1.mmu.r_valid_d[23] ),
    .A2(_07584_),
    .A1(net85));
 sg13g2_nor2_1 _26739_ (.A(net550),
    .B(_07586_),
    .Y(_01066_));
 sg13g2_nor2_1 _26740_ (.A(_07537_),
    .B(net551),
    .Y(_07587_));
 sg13g2_o21ai_1 _26741_ (.B1(_07541_),
    .Y(_07588_),
    .A1(net552),
    .A2(_07587_));
 sg13g2_nand2_1 _26742_ (.Y(_07589_),
    .A(_07556_),
    .B(_07531_));
 sg13g2_nor2_1 _26743_ (.A(net551),
    .B(_07589_),
    .Y(_07590_));
 sg13g2_a21oi_1 _26744_ (.A1(\cpu.genblk1.mmu.r_valid_d[24] ),
    .A2(_07588_),
    .Y(_07591_),
    .B1(_07590_));
 sg13g2_nor2_1 _26745_ (.A(net550),
    .B(_07591_),
    .Y(_01067_));
 sg13g2_a21oi_1 _26746_ (.A1(_05951_),
    .A2(_07496_),
    .Y(_07592_),
    .B1(_07478_));
 sg13g2_buf_2 _26747_ (.A(_07592_),
    .X(_07593_));
 sg13g2_nor3_2 _26748_ (.A(_05828_),
    .B(_05885_),
    .C(_07593_),
    .Y(_07594_));
 sg13g2_o21ai_1 _26749_ (.B1(_07542_),
    .Y(_07595_),
    .A1(_07535_),
    .A2(_07594_));
 sg13g2_a22oi_1 _26750_ (.Y(_07596_),
    .B1(_07595_),
    .B2(\cpu.genblk1.mmu.r_valid_d[25] ),
    .A2(_07594_),
    .A1(net85));
 sg13g2_nor2_1 _26751_ (.A(net550),
    .B(_07596_),
    .Y(_01068_));
 sg13g2_o21ai_1 _26752_ (.B1(_07541_),
    .Y(_07597_),
    .A1(net552),
    .A2(_05961_));
 sg13g2_nor2b_1 _26753_ (.A(_07593_),
    .B_N(_07493_),
    .Y(_07598_));
 sg13g2_a22oi_1 _26754_ (.Y(_07599_),
    .B1(_07598_),
    .B2(_07556_),
    .A2(_07597_),
    .A1(\cpu.genblk1.mmu.r_valid_d[26] ));
 sg13g2_nor2_1 _26755_ (.A(_07570_),
    .B(_07599_),
    .Y(_01069_));
 sg13g2_o21ai_1 _26756_ (.B1(_07542_),
    .Y(_07600_),
    .A1(_07535_),
    .A2(_05967_));
 sg13g2_a22oi_1 _26757_ (.Y(_07601_),
    .B1(_07600_),
    .B2(\cpu.genblk1.mmu.r_valid_d[27] ),
    .A2(_07490_),
    .A1(_05967_));
 sg13g2_nor2_1 _26758_ (.A(net550),
    .B(_07601_),
    .Y(_01070_));
 sg13g2_inv_1 _26759_ (.Y(_07602_),
    .A(_07593_));
 sg13g2_nor2_1 _26760_ (.A(_07512_),
    .B(_07593_),
    .Y(_07603_));
 sg13g2_o21ai_1 _26761_ (.B1(_07541_),
    .Y(_07604_),
    .A1(_07534_),
    .A2(_07603_));
 sg13g2_a22oi_1 _26762_ (.Y(_07605_),
    .B1(_07604_),
    .B2(\cpu.genblk1.mmu.r_valid_d[28] ),
    .A2(_07602_),
    .A1(_07573_));
 sg13g2_nor2_1 _26763_ (.A(_07570_),
    .B(_07605_),
    .Y(_01071_));
 sg13g2_nor2_2 _26764_ (.A(_07517_),
    .B(_07593_),
    .Y(_07606_));
 sg13g2_o21ai_1 _26765_ (.B1(_07541_),
    .Y(_07607_),
    .A1(net552),
    .A2(_07606_));
 sg13g2_a22oi_1 _26766_ (.Y(_07608_),
    .B1(_07607_),
    .B2(\cpu.genblk1.mmu.r_valid_d[29] ),
    .A2(_07606_),
    .A1(net85));
 sg13g2_nor2_1 _26767_ (.A(net550),
    .B(_07608_),
    .Y(_01072_));
 sg13g2_buf_1 _26768_ (.A(_09129_),
    .X(_07609_));
 sg13g2_nor3_1 _26769_ (.A(net827),
    .B(_05865_),
    .C(net472),
    .Y(_07610_));
 sg13g2_o21ai_1 _26770_ (.B1(_07487_),
    .Y(_07611_),
    .A1(net158),
    .A2(_07610_));
 sg13g2_and2_1 _26771_ (.A(_04844_),
    .B(_07610_),
    .X(_07612_));
 sg13g2_a22oi_1 _26772_ (.Y(_07613_),
    .B1(_07612_),
    .B2(_07556_),
    .A2(_07611_),
    .A1(\cpu.genblk1.mmu.r_valid_d[2] ));
 sg13g2_nor2_1 _26773_ (.A(net549),
    .B(_07613_),
    .Y(_01073_));
 sg13g2_nor2_1 _26774_ (.A(_06010_),
    .B(_07593_),
    .Y(_07614_));
 sg13g2_o21ai_1 _26775_ (.B1(_07541_),
    .Y(_07615_),
    .A1(_07534_),
    .A2(_07614_));
 sg13g2_a22oi_1 _26776_ (.Y(_07616_),
    .B1(_07615_),
    .B2(\cpu.genblk1.mmu.r_valid_d[30] ),
    .A2(_07602_),
    .A1(_07580_));
 sg13g2_nor2_1 _26777_ (.A(_07609_),
    .B(_07616_),
    .Y(_01074_));
 sg13g2_nor2_2 _26778_ (.A(_05839_),
    .B(_07593_),
    .Y(_07617_));
 sg13g2_o21ai_1 _26779_ (.B1(_07541_),
    .Y(_07618_),
    .A1(net552),
    .A2(_07617_));
 sg13g2_a22oi_1 _26780_ (.Y(_07619_),
    .B1(_07618_),
    .B2(\cpu.genblk1.mmu.r_valid_d[31] ),
    .A2(_07617_),
    .A1(net85));
 sg13g2_nor2_1 _26781_ (.A(_07609_),
    .B(_07619_),
    .Y(_01075_));
 sg13g2_nor2b_2 _26782_ (.A(net472),
    .B_N(_05827_),
    .Y(_07620_));
 sg13g2_o21ai_1 _26783_ (.B1(_07501_),
    .Y(_07621_),
    .A1(net126),
    .A2(_07620_));
 sg13g2_a22oi_1 _26784_ (.Y(_07622_),
    .B1(_07621_),
    .B2(\cpu.genblk1.mmu.r_valid_d[3] ),
    .A2(_07620_),
    .A1(_07490_));
 sg13g2_nor2_1 _26785_ (.A(net549),
    .B(_07622_),
    .Y(_01076_));
 sg13g2_inv_1 _26786_ (.Y(_07623_),
    .A(net472));
 sg13g2_nor2_1 _26787_ (.A(_07512_),
    .B(net472),
    .Y(_07624_));
 sg13g2_o21ai_1 _26788_ (.B1(net125),
    .Y(_07625_),
    .A1(net158),
    .A2(_07624_));
 sg13g2_a22oi_1 _26789_ (.Y(_07626_),
    .B1(_07625_),
    .B2(\cpu.genblk1.mmu.r_valid_d[4] ),
    .A2(_07573_),
    .A1(_07623_));
 sg13g2_nor2_1 _26790_ (.A(net549),
    .B(_07626_),
    .Y(_01077_));
 sg13g2_o21ai_1 _26791_ (.B1(net125),
    .Y(_07627_),
    .A1(_06004_),
    .A2(net126));
 sg13g2_a22oi_1 _26792_ (.Y(_07628_),
    .B1(_07627_),
    .B2(\cpu.genblk1.mmu.r_valid_d[5] ),
    .A2(_07490_),
    .A1(_06004_));
 sg13g2_nor2_1 _26793_ (.A(net549),
    .B(_07628_),
    .Y(_01078_));
 sg13g2_o21ai_1 _26794_ (.B1(_07487_),
    .Y(_07629_),
    .A1(_06011_),
    .A2(net158));
 sg13g2_nor2b_1 _26795_ (.A(net472),
    .B_N(_07522_),
    .Y(_07630_));
 sg13g2_a22oi_1 _26796_ (.Y(_07631_),
    .B1(_07630_),
    .B2(_07556_),
    .A2(_07629_),
    .A1(\cpu.genblk1.mmu.r_valid_d[6] ));
 sg13g2_nor2_1 _26797_ (.A(net549),
    .B(_07631_),
    .Y(_01079_));
 sg13g2_o21ai_1 _26798_ (.B1(_07487_),
    .Y(_07632_),
    .A1(_06016_),
    .A2(net126));
 sg13g2_a22oi_1 _26799_ (.Y(_07633_),
    .B1(_07632_),
    .B2(\cpu.genblk1.mmu.r_valid_d[7] ),
    .A2(_07490_),
    .A1(_06016_));
 sg13g2_nor2_1 _26800_ (.A(net549),
    .B(_07633_),
    .Y(_01080_));
 sg13g2_nor2_1 _26801_ (.A(_07537_),
    .B(_07566_),
    .Y(_07634_));
 sg13g2_o21ai_1 _26802_ (.B1(_07487_),
    .Y(_07635_),
    .A1(_07484_),
    .A2(_07634_));
 sg13g2_nor2_1 _26803_ (.A(net472),
    .B(_07589_),
    .Y(_07636_));
 sg13g2_a21oi_1 _26804_ (.A1(\cpu.genblk1.mmu.r_valid_d[8] ),
    .A2(_07635_),
    .Y(_07637_),
    .B1(_07636_));
 sg13g2_nor2_1 _26805_ (.A(net549),
    .B(_07637_),
    .Y(_01081_));
 sg13g2_nor3_2 _26806_ (.A(net827),
    .B(_05885_),
    .C(_07498_),
    .Y(_07638_));
 sg13g2_o21ai_1 _26807_ (.B1(_07487_),
    .Y(_07639_),
    .A1(net158),
    .A2(_07638_));
 sg13g2_a22oi_1 _26808_ (.Y(_07640_),
    .B1(_07639_),
    .B2(\cpu.genblk1.mmu.r_valid_d[9] ),
    .A2(_07638_),
    .A1(_07490_));
 sg13g2_nor2_1 _26809_ (.A(net549),
    .B(_07640_),
    .Y(_01082_));
 sg13g2_buf_1 _26810_ (.A(_09129_),
    .X(_07641_));
 sg13g2_nand2_1 _26811_ (.Y(_07642_),
    .A(_08189_),
    .B(_00233_));
 sg13g2_a21oi_1 _26812_ (.A1(_07479_),
    .A2(_07642_),
    .Y(_07643_),
    .B1(_07533_));
 sg13g2_nand2b_1 _26813_ (.Y(_07644_),
    .B(_08259_),
    .A_N(_07643_));
 sg13g2_buf_1 _26814_ (.A(_07644_),
    .X(_07645_));
 sg13g2_nand2b_1 _26815_ (.Y(_07646_),
    .B(_05797_),
    .A_N(_07645_));
 sg13g2_buf_1 _26816_ (.A(_07646_),
    .X(_07647_));
 sg13g2_nor2b_1 _26817_ (.A(_10327_),
    .B_N(_03465_),
    .Y(_07648_));
 sg13g2_a21oi_1 _26818_ (.A1(_05795_),
    .A2(_07648_),
    .Y(_07649_),
    .B1(_07645_));
 sg13g2_buf_2 _26819_ (.A(_07649_),
    .X(_07650_));
 sg13g2_o21ai_1 _26820_ (.B1(_07650_),
    .Y(_07651_),
    .A1(_07478_),
    .A2(net188));
 sg13g2_nor2_1 _26821_ (.A(_09875_),
    .B(_07647_),
    .Y(_07652_));
 sg13g2_buf_2 _26822_ (.A(_07652_),
    .X(_07653_));
 sg13g2_buf_1 _26823_ (.A(_07653_),
    .X(_07654_));
 sg13g2_a22oi_1 _26824_ (.Y(_07655_),
    .B1(net108),
    .B2(_07478_),
    .A2(_07651_),
    .A1(\cpu.genblk1.mmu.r_valid_i[0] ));
 sg13g2_nor2_1 _26825_ (.A(net548),
    .B(_07655_),
    .Y(_01083_));
 sg13g2_nor2_1 _26826_ (.A(_07498_),
    .B(net188),
    .Y(_07656_));
 sg13g2_buf_1 _26827_ (.A(net188),
    .X(_07657_));
 sg13g2_buf_1 _26828_ (.A(_07650_),
    .X(_07658_));
 sg13g2_o21ai_1 _26829_ (.B1(net156),
    .Y(_07659_),
    .A1(_05868_),
    .A2(net157));
 sg13g2_a22oi_1 _26830_ (.Y(_07660_),
    .B1(_07659_),
    .B2(\cpu.genblk1.mmu.r_valid_i[10] ),
    .A2(_07656_),
    .A1(_07493_));
 sg13g2_nor2_1 _26831_ (.A(net548),
    .B(_07660_),
    .Y(_01084_));
 sg13g2_o21ai_1 _26832_ (.B1(net156),
    .Y(_07661_),
    .A1(_05873_),
    .A2(net157));
 sg13g2_a22oi_1 _26833_ (.Y(_07662_),
    .B1(_07661_),
    .B2(\cpu.genblk1.mmu.r_valid_i[11] ),
    .A2(_07654_),
    .A1(_05873_));
 sg13g2_nor2_1 _26834_ (.A(net548),
    .B(_07662_),
    .Y(_01085_));
 sg13g2_o21ai_1 _26835_ (.B1(net156),
    .Y(_07663_),
    .A1(_07513_),
    .A2(_07657_));
 sg13g2_a22oi_1 _26836_ (.Y(_07664_),
    .B1(_07663_),
    .B2(\cpu.genblk1.mmu.r_valid_i[12] ),
    .A2(_07656_),
    .A1(_07509_));
 sg13g2_nor2_1 _26837_ (.A(_07641_),
    .B(_07664_),
    .Y(_01086_));
 sg13g2_o21ai_1 _26838_ (.B1(net156),
    .Y(_07665_),
    .A1(_07518_),
    .A2(net157));
 sg13g2_a22oi_1 _26839_ (.Y(_07666_),
    .B1(_07665_),
    .B2(\cpu.genblk1.mmu.r_valid_i[13] ),
    .A2(_07654_),
    .A1(_07518_));
 sg13g2_nor2_1 _26840_ (.A(_07641_),
    .B(_07666_),
    .Y(_01087_));
 sg13g2_o21ai_1 _26841_ (.B1(_07658_),
    .Y(_07667_),
    .A1(_07523_),
    .A2(net157));
 sg13g2_a22oi_1 _26842_ (.Y(_07668_),
    .B1(_07667_),
    .B2(\cpu.genblk1.mmu.r_valid_i[14] ),
    .A2(_07656_),
    .A1(_07522_));
 sg13g2_nor2_1 _26843_ (.A(net548),
    .B(_07668_),
    .Y(_01088_));
 sg13g2_o21ai_1 _26844_ (.B1(_07658_),
    .Y(_07669_),
    .A1(_07526_),
    .A2(net157));
 sg13g2_a22oi_1 _26845_ (.Y(_07670_),
    .B1(_07669_),
    .B2(\cpu.genblk1.mmu.r_valid_i[15] ),
    .A2(net108),
    .A1(_07526_));
 sg13g2_nor2_1 _26846_ (.A(net548),
    .B(_07670_),
    .Y(_01089_));
 sg13g2_a21oi_1 _26847_ (.A1(_03465_),
    .A2(_10427_),
    .Y(_07671_),
    .B1(_05797_));
 sg13g2_nor2_1 _26848_ (.A(_07645_),
    .B(_07671_),
    .Y(_07672_));
 sg13g2_buf_2 _26849_ (.A(_07672_),
    .X(_07673_));
 sg13g2_buf_1 _26850_ (.A(_07673_),
    .X(_07674_));
 sg13g2_o21ai_1 _26851_ (.B1(_07674_),
    .Y(_07675_),
    .A1(_07538_),
    .A2(_07657_));
 sg13g2_a22oi_1 _26852_ (.Y(_07676_),
    .B1(_07675_),
    .B2(\cpu.genblk1.mmu.r_valid_i[16] ),
    .A2(_07656_),
    .A1(_07531_));
 sg13g2_nor2_1 _26853_ (.A(net548),
    .B(_07676_),
    .Y(_01090_));
 sg13g2_o21ai_1 _26854_ (.B1(net155),
    .Y(_07677_),
    .A1(_07552_),
    .A2(net157));
 sg13g2_a22oi_1 _26855_ (.Y(_07678_),
    .B1(_07677_),
    .B2(\cpu.genblk1.mmu.r_valid_i[17] ),
    .A2(net108),
    .A1(_07552_));
 sg13g2_nor2_1 _26856_ (.A(net548),
    .B(_07678_),
    .Y(_01091_));
 sg13g2_nor2_1 _26857_ (.A(net552),
    .B(_07645_),
    .Y(_07679_));
 sg13g2_o21ai_1 _26858_ (.B1(net155),
    .Y(_07680_),
    .A1(_05916_),
    .A2(net157));
 sg13g2_a22oi_1 _26859_ (.Y(_07681_),
    .B1(_07680_),
    .B2(\cpu.genblk1.mmu.r_valid_i[18] ),
    .A2(_07679_),
    .A1(_07557_));
 sg13g2_nor2_1 _26860_ (.A(net548),
    .B(_07681_),
    .Y(_01092_));
 sg13g2_buf_1 _26861_ (.A(_09129_),
    .X(_07682_));
 sg13g2_o21ai_1 _26862_ (.B1(net155),
    .Y(_07683_),
    .A1(_05925_),
    .A2(net157));
 sg13g2_a22oi_1 _26863_ (.Y(_07684_),
    .B1(_07683_),
    .B2(\cpu.genblk1.mmu.r_valid_i[19] ),
    .A2(net108),
    .A1(_05925_));
 sg13g2_nor2_1 _26864_ (.A(net547),
    .B(_07684_),
    .Y(_01093_));
 sg13g2_buf_1 _26865_ (.A(net188),
    .X(_07685_));
 sg13g2_o21ai_1 _26866_ (.B1(net156),
    .Y(_07686_),
    .A1(_07567_),
    .A2(net154));
 sg13g2_a22oi_1 _26867_ (.Y(_07687_),
    .B1(_07686_),
    .B2(\cpu.genblk1.mmu.r_valid_i[1] ),
    .A2(net108),
    .A1(_07567_));
 sg13g2_nor2_1 _26868_ (.A(net547),
    .B(_07687_),
    .Y(_01094_));
 sg13g2_nor2_1 _26869_ (.A(net551),
    .B(net188),
    .Y(_07688_));
 sg13g2_o21ai_1 _26870_ (.B1(net155),
    .Y(_07689_),
    .A1(_07574_),
    .A2(net154));
 sg13g2_a22oi_1 _26871_ (.Y(_07690_),
    .B1(_07689_),
    .B2(\cpu.genblk1.mmu.r_valid_i[20] ),
    .A2(_07688_),
    .A1(_07509_));
 sg13g2_nor2_1 _26872_ (.A(net547),
    .B(_07690_),
    .Y(_01095_));
 sg13g2_o21ai_1 _26873_ (.B1(net155),
    .Y(_07691_),
    .A1(_07577_),
    .A2(net154));
 sg13g2_a22oi_1 _26874_ (.Y(_07692_),
    .B1(_07691_),
    .B2(\cpu.genblk1.mmu.r_valid_i[21] ),
    .A2(net108),
    .A1(_07577_));
 sg13g2_nor2_1 _26875_ (.A(net547),
    .B(_07692_),
    .Y(_01096_));
 sg13g2_o21ai_1 _26876_ (.B1(net155),
    .Y(_07693_),
    .A1(_07581_),
    .A2(net154));
 sg13g2_a22oi_1 _26877_ (.Y(_07694_),
    .B1(_07693_),
    .B2(\cpu.genblk1.mmu.r_valid_i[22] ),
    .A2(_07688_),
    .A1(_07522_));
 sg13g2_nor2_1 _26878_ (.A(net547),
    .B(_07694_),
    .Y(_01097_));
 sg13g2_o21ai_1 _26879_ (.B1(net155),
    .Y(_07695_),
    .A1(_07584_),
    .A2(net154));
 sg13g2_a22oi_1 _26880_ (.Y(_07696_),
    .B1(_07695_),
    .B2(\cpu.genblk1.mmu.r_valid_i[23] ),
    .A2(net108),
    .A1(_07584_));
 sg13g2_nor2_1 _26881_ (.A(net547),
    .B(_07696_),
    .Y(_01098_));
 sg13g2_o21ai_1 _26882_ (.B1(net155),
    .Y(_07697_),
    .A1(_07587_),
    .A2(net154));
 sg13g2_a22oi_1 _26883_ (.Y(_07698_),
    .B1(_07697_),
    .B2(\cpu.genblk1.mmu.r_valid_i[24] ),
    .A2(_07688_),
    .A1(_07531_));
 sg13g2_nor2_1 _26884_ (.A(_07682_),
    .B(_07698_),
    .Y(_01099_));
 sg13g2_o21ai_1 _26885_ (.B1(_07674_),
    .Y(_07699_),
    .A1(_07594_),
    .A2(net154));
 sg13g2_a22oi_1 _26886_ (.Y(_07700_),
    .B1(_07699_),
    .B2(\cpu.genblk1.mmu.r_valid_i[25] ),
    .A2(net108),
    .A1(_07594_));
 sg13g2_nor2_1 _26887_ (.A(net547),
    .B(_07700_),
    .Y(_01100_));
 sg13g2_nor2_1 _26888_ (.A(_07593_),
    .B(net188),
    .Y(_07701_));
 sg13g2_o21ai_1 _26889_ (.B1(_07673_),
    .Y(_07702_),
    .A1(_05961_),
    .A2(_07685_));
 sg13g2_a22oi_1 _26890_ (.Y(_07703_),
    .B1(_07702_),
    .B2(\cpu.genblk1.mmu.r_valid_i[26] ),
    .A2(_07701_),
    .A1(_07493_));
 sg13g2_nor2_1 _26891_ (.A(_07682_),
    .B(_07703_),
    .Y(_01101_));
 sg13g2_o21ai_1 _26892_ (.B1(_07673_),
    .Y(_07704_),
    .A1(_05967_),
    .A2(net154));
 sg13g2_a22oi_1 _26893_ (.Y(_07705_),
    .B1(_07704_),
    .B2(\cpu.genblk1.mmu.r_valid_i[27] ),
    .A2(_07653_),
    .A1(_05967_));
 sg13g2_nor2_1 _26894_ (.A(net547),
    .B(_07705_),
    .Y(_01102_));
 sg13g2_buf_1 _26895_ (.A(_09129_),
    .X(_07706_));
 sg13g2_o21ai_1 _26896_ (.B1(_07673_),
    .Y(_07707_),
    .A1(_07603_),
    .A2(_07685_));
 sg13g2_a22oi_1 _26897_ (.Y(_07708_),
    .B1(_07707_),
    .B2(\cpu.genblk1.mmu.r_valid_i[28] ),
    .A2(_07701_),
    .A1(_07509_));
 sg13g2_nor2_1 _26898_ (.A(net546),
    .B(_07708_),
    .Y(_01103_));
 sg13g2_buf_1 _26899_ (.A(_07647_),
    .X(_07709_));
 sg13g2_o21ai_1 _26900_ (.B1(_07673_),
    .Y(_07710_),
    .A1(_07606_),
    .A2(_07709_));
 sg13g2_a22oi_1 _26901_ (.Y(_07711_),
    .B1(_07710_),
    .B2(\cpu.genblk1.mmu.r_valid_i[29] ),
    .A2(_07653_),
    .A1(_07606_));
 sg13g2_nor2_1 _26902_ (.A(_07706_),
    .B(_07711_),
    .Y(_01104_));
 sg13g2_o21ai_1 _26903_ (.B1(net156),
    .Y(_07712_),
    .A1(_07610_),
    .A2(net153));
 sg13g2_a22oi_1 _26904_ (.Y(_07713_),
    .B1(_07712_),
    .B2(\cpu.genblk1.mmu.r_valid_i[2] ),
    .A2(_07679_),
    .A1(_07612_));
 sg13g2_nor2_1 _26905_ (.A(net546),
    .B(_07713_),
    .Y(_01105_));
 sg13g2_o21ai_1 _26906_ (.B1(_07673_),
    .Y(_07714_),
    .A1(_07614_),
    .A2(_07709_));
 sg13g2_a22oi_1 _26907_ (.Y(_07715_),
    .B1(_07714_),
    .B2(\cpu.genblk1.mmu.r_valid_i[30] ),
    .A2(_07701_),
    .A1(_07522_));
 sg13g2_nor2_1 _26908_ (.A(net546),
    .B(_07715_),
    .Y(_01106_));
 sg13g2_o21ai_1 _26909_ (.B1(_07673_),
    .Y(_07716_),
    .A1(_07617_),
    .A2(net153));
 sg13g2_a22oi_1 _26910_ (.Y(_07717_),
    .B1(_07716_),
    .B2(\cpu.genblk1.mmu.r_valid_i[31] ),
    .A2(_07653_),
    .A1(_07617_));
 sg13g2_nor2_1 _26911_ (.A(_07706_),
    .B(_07717_),
    .Y(_01107_));
 sg13g2_o21ai_1 _26912_ (.B1(net156),
    .Y(_07718_),
    .A1(_07620_),
    .A2(net153));
 sg13g2_a22oi_1 _26913_ (.Y(_07719_),
    .B1(_07718_),
    .B2(\cpu.genblk1.mmu.r_valid_i[3] ),
    .A2(_07653_),
    .A1(_07620_));
 sg13g2_nor2_1 _26914_ (.A(net546),
    .B(_07719_),
    .Y(_01108_));
 sg13g2_nor2_1 _26915_ (.A(net472),
    .B(net188),
    .Y(_07720_));
 sg13g2_o21ai_1 _26916_ (.B1(net156),
    .Y(_07721_),
    .A1(_07624_),
    .A2(net153));
 sg13g2_a22oi_1 _26917_ (.Y(_07722_),
    .B1(_07721_),
    .B2(\cpu.genblk1.mmu.r_valid_i[4] ),
    .A2(_07720_),
    .A1(_07509_));
 sg13g2_nor2_1 _26918_ (.A(net546),
    .B(_07722_),
    .Y(_01109_));
 sg13g2_o21ai_1 _26919_ (.B1(_07650_),
    .Y(_07723_),
    .A1(_06004_),
    .A2(net153));
 sg13g2_a22oi_1 _26920_ (.Y(_07724_),
    .B1(_07723_),
    .B2(\cpu.genblk1.mmu.r_valid_i[5] ),
    .A2(_07653_),
    .A1(_06004_));
 sg13g2_nor2_1 _26921_ (.A(net546),
    .B(_07724_),
    .Y(_01110_));
 sg13g2_o21ai_1 _26922_ (.B1(_07650_),
    .Y(_07725_),
    .A1(_06011_),
    .A2(net153));
 sg13g2_a22oi_1 _26923_ (.Y(_07726_),
    .B1(_07725_),
    .B2(\cpu.genblk1.mmu.r_valid_i[6] ),
    .A2(_07720_),
    .A1(_07522_));
 sg13g2_nor2_1 _26924_ (.A(net546),
    .B(_07726_),
    .Y(_01111_));
 sg13g2_o21ai_1 _26925_ (.B1(_07650_),
    .Y(_07727_),
    .A1(_06016_),
    .A2(net153));
 sg13g2_a22oi_1 _26926_ (.Y(_07728_),
    .B1(_07727_),
    .B2(\cpu.genblk1.mmu.r_valid_i[7] ),
    .A2(_07653_),
    .A1(_06016_));
 sg13g2_nor2_1 _26927_ (.A(net546),
    .B(_07728_),
    .Y(_01112_));
 sg13g2_buf_2 _26928_ (.A(_09136_),
    .X(_07729_));
 sg13g2_o21ai_1 _26929_ (.B1(_07650_),
    .Y(_07730_),
    .A1(_07634_),
    .A2(net153));
 sg13g2_a22oi_1 _26930_ (.Y(_07731_),
    .B1(_07730_),
    .B2(\cpu.genblk1.mmu.r_valid_i[8] ),
    .A2(_07720_),
    .A1(_07531_));
 sg13g2_nor2_1 _26931_ (.A(_07729_),
    .B(_07731_),
    .Y(_01113_));
 sg13g2_o21ai_1 _26932_ (.B1(_07650_),
    .Y(_07732_),
    .A1(_07638_),
    .A2(net188));
 sg13g2_a22oi_1 _26933_ (.Y(_07733_),
    .B1(_07732_),
    .B2(\cpu.genblk1.mmu.r_valid_i[9] ),
    .A2(_07653_),
    .A1(_07638_));
 sg13g2_nor2_1 _26934_ (.A(_07729_),
    .B(_07733_),
    .Y(_01114_));
 sg13g2_and2_1 _26935_ (.A(_05089_),
    .B(_06229_),
    .X(_07734_));
 sg13g2_buf_2 _26936_ (.A(_07734_),
    .X(_07735_));
 sg13g2_nand2_1 _26937_ (.Y(_07736_),
    .A(net970),
    .B(_07735_));
 sg13g2_nand2_1 _26938_ (.Y(_07737_),
    .A(_05089_),
    .B(_06229_));
 sg13g2_buf_2 _26939_ (.A(_07737_),
    .X(_07738_));
 sg13g2_nand2_1 _26940_ (.Y(_07739_),
    .A(_08990_),
    .B(_07738_));
 sg13g2_buf_1 _26941_ (.A(_09136_),
    .X(_07740_));
 sg13g2_a21oi_1 _26942_ (.A1(_07736_),
    .A2(_07739_),
    .Y(_01915_),
    .B1(net544));
 sg13g2_nand2_1 _26943_ (.Y(_07741_),
    .A(_09929_),
    .B(_07735_));
 sg13g2_nand2_1 _26944_ (.Y(_07742_),
    .A(\cpu.gpio.r_enable_in[1] ),
    .B(_07738_));
 sg13g2_a21oi_1 _26945_ (.A1(_07741_),
    .A2(_07742_),
    .Y(_01916_),
    .B1(net544));
 sg13g2_nand2_1 _26946_ (.Y(_07743_),
    .A(_09936_),
    .B(_07735_));
 sg13g2_nand2_1 _26947_ (.Y(_07744_),
    .A(\cpu.gpio.r_enable_in[2] ),
    .B(_07738_));
 sg13g2_a21oi_1 _26948_ (.A1(_07743_),
    .A2(_07744_),
    .Y(_01917_),
    .B1(net544));
 sg13g2_nand2_1 _26949_ (.Y(_07745_),
    .A(_09942_),
    .B(_07735_));
 sg13g2_nand2_1 _26950_ (.Y(_07746_),
    .A(\cpu.gpio.r_enable_in[3] ),
    .B(_07738_));
 sg13g2_a21oi_1 _26951_ (.A1(_07745_),
    .A2(_07746_),
    .Y(_01918_),
    .B1(net544));
 sg13g2_nand2_1 _26952_ (.Y(_07747_),
    .A(net1105),
    .B(_07735_));
 sg13g2_nand2_1 _26953_ (.Y(_07748_),
    .A(_08995_),
    .B(_07738_));
 sg13g2_a21oi_1 _26954_ (.A1(_07747_),
    .A2(_07748_),
    .Y(_01919_),
    .B1(net544));
 sg13g2_nand2_1 _26955_ (.Y(_07749_),
    .A(net1021),
    .B(_07735_));
 sg13g2_nand2_1 _26956_ (.Y(_07750_),
    .A(_09001_),
    .B(_07738_));
 sg13g2_a21oi_1 _26957_ (.A1(_07749_),
    .A2(_07750_),
    .Y(_01920_),
    .B1(_07740_));
 sg13g2_nand2_1 _26958_ (.Y(_07751_),
    .A(net1020),
    .B(_07735_));
 sg13g2_nand2_1 _26959_ (.Y(_07752_),
    .A(_08997_),
    .B(_07738_));
 sg13g2_a21oi_1 _26960_ (.A1(_07751_),
    .A2(_07752_),
    .Y(_01921_),
    .B1(_07740_));
 sg13g2_nand2_1 _26961_ (.Y(_07753_),
    .A(net1104),
    .B(_07735_));
 sg13g2_nand2_1 _26962_ (.Y(_07754_),
    .A(\cpu.gpio.r_enable_in[7] ),
    .B(_07738_));
 sg13g2_a21oi_1 _26963_ (.A1(_07753_),
    .A2(_07754_),
    .Y(_01922_),
    .B1(net544));
 sg13g2_buf_1 _26964_ (.A(_06229_),
    .X(_07755_));
 sg13g2_nand3_1 _26965_ (.B(net287),
    .C(net107),
    .A(_09895_),
    .Y(_07756_));
 sg13g2_nand2_1 _26966_ (.Y(_07757_),
    .A(net287),
    .B(net107));
 sg13g2_nand2_1 _26967_ (.Y(_07758_),
    .A(\cpu.gpio.r_enable_io[4] ),
    .B(_07757_));
 sg13g2_a21oi_1 _26968_ (.A1(_07756_),
    .A2(_07758_),
    .Y(_01923_),
    .B1(net544));
 sg13g2_nand3_1 _26969_ (.B(net287),
    .C(net107),
    .A(_09902_),
    .Y(_07759_));
 sg13g2_nand2_1 _26970_ (.Y(_07760_),
    .A(_08984_),
    .B(_07757_));
 sg13g2_a21oi_1 _26971_ (.A1(_07759_),
    .A2(_07760_),
    .Y(_01924_),
    .B1(net544));
 sg13g2_nand3_1 _26972_ (.B(_05459_),
    .C(net107),
    .A(net1020),
    .Y(_07761_));
 sg13g2_nand2_1 _26973_ (.Y(_07762_),
    .A(\cpu.gpio.r_enable_io[6] ),
    .B(_07757_));
 sg13g2_buf_1 _26974_ (.A(_09136_),
    .X(_07763_));
 sg13g2_a21oi_1 _26975_ (.A1(_07761_),
    .A2(_07762_),
    .Y(_01925_),
    .B1(net543));
 sg13g2_nand3_1 _26976_ (.B(_05459_),
    .C(net107),
    .A(_09910_),
    .Y(_07764_));
 sg13g2_nand2_1 _26977_ (.Y(_07765_),
    .A(_08992_),
    .B(_07757_));
 sg13g2_a21oi_1 _26978_ (.A1(_07764_),
    .A2(_07765_),
    .Y(_01926_),
    .B1(net543));
 sg13g2_nand3_1 _26979_ (.B(_05024_),
    .C(_06229_),
    .A(net830),
    .Y(_07766_));
 sg13g2_buf_2 _26980_ (.A(_07766_),
    .X(_07767_));
 sg13g2_nand2_1 _26981_ (.Y(_07768_),
    .A(net7),
    .B(_07767_));
 sg13g2_o21ai_1 _26982_ (.B1(_07768_),
    .Y(_07769_),
    .A1(net853),
    .A2(_07767_));
 sg13g2_and2_1 _26983_ (.A(net687),
    .B(_07769_),
    .X(_01927_));
 sg13g2_mux2_1 _26984_ (.A0(_09901_),
    .A1(net8),
    .S(_07767_),
    .X(_07770_));
 sg13g2_and2_1 _26985_ (.A(net648),
    .B(_07770_),
    .X(_01928_));
 sg13g2_mux2_1 _26986_ (.A0(_09907_),
    .A1(net9),
    .S(_07767_),
    .X(_07771_));
 sg13g2_and2_1 _26987_ (.A(net648),
    .B(_07771_),
    .X(_01929_));
 sg13g2_nand2_1 _26988_ (.Y(_07772_),
    .A(net10),
    .B(_07767_));
 sg13g2_o21ai_1 _26989_ (.B1(_07772_),
    .Y(_07773_),
    .A1(net852),
    .A2(_07767_));
 sg13g2_and2_1 _26990_ (.A(net648),
    .B(_07773_),
    .X(_01930_));
 sg13g2_nand2_1 _26991_ (.Y(_07774_),
    .A(_04980_),
    .B(_06229_));
 sg13g2_buf_2 _26992_ (.A(_07774_),
    .X(_07775_));
 sg13g2_nor2_1 _26993_ (.A(net1024),
    .B(_07775_),
    .Y(_07776_));
 sg13g2_a21oi_1 _26994_ (.A1(_04980_),
    .A2(_07755_),
    .Y(_07777_),
    .B1(_04977_));
 sg13g2_o21ai_1 _26995_ (.B1(net622),
    .Y(_01976_),
    .A1(_07776_),
    .A2(_07777_));
 sg13g2_buf_1 _26996_ (.A(\cpu.gpio.r_src_o[6][1] ),
    .X(_07778_));
 sg13g2_mux2_1 _26997_ (.A0(net1023),
    .A1(_07778_),
    .S(_07775_),
    .X(_07779_));
 sg13g2_and2_1 _26998_ (.A(net648),
    .B(_07779_),
    .X(_01977_));
 sg13g2_nand2_1 _26999_ (.Y(_07780_),
    .A(\cpu.gpio.r_src_o[6][2] ),
    .B(_07775_));
 sg13g2_o21ai_1 _27000_ (.B1(_07780_),
    .Y(_07781_),
    .A1(net878),
    .A2(_07775_));
 sg13g2_and2_1 _27001_ (.A(net648),
    .B(_07781_),
    .X(_01978_));
 sg13g2_nand2_1 _27002_ (.Y(_07782_),
    .A(\cpu.gpio.r_src_o[6][3] ),
    .B(_07775_));
 sg13g2_o21ai_1 _27003_ (.B1(_07782_),
    .Y(_07783_),
    .A1(net854),
    .A2(_07775_));
 sg13g2_and2_1 _27004_ (.A(net648),
    .B(_07783_),
    .X(_01979_));
 sg13g2_nand3_1 _27005_ (.B(_05365_),
    .C(net107),
    .A(net1024),
    .Y(_07784_));
 sg13g2_nand2_1 _27006_ (.Y(_07785_),
    .A(_05365_),
    .B(net107));
 sg13g2_nand2_1 _27007_ (.Y(_07786_),
    .A(_04967_),
    .B(_07785_));
 sg13g2_a21oi_1 _27008_ (.A1(_07784_),
    .A2(_07786_),
    .Y(_01984_),
    .B1(net543));
 sg13g2_nand3_1 _27009_ (.B(_05365_),
    .C(_07755_),
    .A(net1018),
    .Y(_07787_));
 sg13g2_nand2_1 _27010_ (.Y(_07788_),
    .A(\cpu.gpio.r_uart_rx_src[1] ),
    .B(_07785_));
 sg13g2_a21oi_1 _27011_ (.A1(_07787_),
    .A2(_07788_),
    .Y(_01985_),
    .B1(_07763_));
 sg13g2_nand3_1 _27012_ (.B(_05365_),
    .C(net107),
    .A(net1017),
    .Y(_07789_));
 sg13g2_nand2_1 _27013_ (.Y(_07790_),
    .A(\cpu.gpio.r_uart_rx_src[2] ),
    .B(_07785_));
 sg13g2_a21oi_1 _27014_ (.A1(_07789_),
    .A2(_07790_),
    .Y(_01986_),
    .B1(_07763_));
 sg13g2_and2_1 _27015_ (.A(\cpu.i_wstrobe_d ),
    .B(_00293_),
    .X(_02243_));
 sg13g2_nor2_1 _27016_ (.A(_06272_),
    .B(_06285_),
    .Y(_07791_));
 sg13g2_nor2_1 _27017_ (.A(_06299_),
    .B(_07791_),
    .Y(_02244_));
 sg13g2_xor2_1 _27018_ (.B(_06300_),
    .A(\cpu.icache.r_offset[2] ),
    .X(_07792_));
 sg13g2_nor2_1 _27019_ (.A(_06299_),
    .B(_07792_),
    .Y(_02245_));
 sg13g2_nand4_1 _27020_ (.B(_09870_),
    .C(_06561_),
    .A(net644),
    .Y(_07793_),
    .D(_04887_));
 sg13g2_xnor2_1 _27021_ (.Y(_07794_),
    .A(\cpu.intr.r_clock_cmp[17] ),
    .B(_05339_));
 sg13g2_xnor2_1 _27022_ (.Y(_07795_),
    .A(\cpu.intr.r_clock_cmp[1] ),
    .B(_09931_));
 sg13g2_xnor2_1 _27023_ (.Y(_07796_),
    .A(\cpu.intr.r_clock_cmp[13] ),
    .B(_10002_));
 sg13g2_xnor2_1 _27024_ (.Y(_07797_),
    .A(\cpu.intr.r_clock_cmp[5] ),
    .B(_09953_));
 sg13g2_nand4_1 _27025_ (.B(_07795_),
    .C(_07796_),
    .A(_07794_),
    .Y(_07798_),
    .D(_07797_));
 sg13g2_xnor2_1 _27026_ (.Y(_07799_),
    .A(\cpu.intr.r_clock_cmp[26] ),
    .B(_05029_));
 sg13g2_xnor2_1 _27027_ (.Y(_07800_),
    .A(\cpu.intr.r_clock_cmp[0] ),
    .B(_09930_));
 sg13g2_xnor2_1 _27028_ (.Y(_07801_),
    .A(\cpu.intr.r_clock_cmp[28] ),
    .B(_05178_));
 sg13g2_xnor2_1 _27029_ (.Y(_07802_),
    .A(\cpu.intr.r_clock_cmp[7] ),
    .B(_09970_));
 sg13g2_nand4_1 _27030_ (.B(_07800_),
    .C(_07801_),
    .A(_07799_),
    .Y(_07803_),
    .D(_07802_));
 sg13g2_xnor2_1 _27031_ (.Y(_07804_),
    .A(\cpu.intr.r_clock_cmp[3] ),
    .B(_09943_));
 sg13g2_xnor2_1 _27032_ (.Y(_07805_),
    .A(\cpu.intr.r_clock_cmp[24] ),
    .B(_05720_));
 sg13g2_xnor2_1 _27033_ (.Y(_07806_),
    .A(\cpu.intr.r_clock_cmp[11] ),
    .B(_09992_));
 sg13g2_xnor2_1 _27034_ (.Y(_07807_),
    .A(\cpu.intr.r_clock_cmp[29] ),
    .B(_05208_));
 sg13g2_nand4_1 _27035_ (.B(_07805_),
    .C(_07806_),
    .A(_07804_),
    .Y(_07808_),
    .D(_07807_));
 sg13g2_xnor2_1 _27036_ (.Y(_07809_),
    .A(\cpu.intr.r_clock_cmp[30] ),
    .B(_05231_));
 sg13g2_xnor2_1 _27037_ (.Y(_07810_),
    .A(\cpu.intr.r_clock_cmp[21] ),
    .B(net1073));
 sg13g2_xnor2_1 _27038_ (.Y(_07811_),
    .A(\cpu.intr.r_clock_cmp[23] ),
    .B(_05115_));
 sg13g2_xnor2_1 _27039_ (.Y(_07812_),
    .A(\cpu.intr.r_clock_cmp[8] ),
    .B(_09976_));
 sg13g2_nand4_1 _27040_ (.B(_07810_),
    .C(_07811_),
    .A(_07809_),
    .Y(_07813_),
    .D(_07812_));
 sg13g2_nor4_1 _27041_ (.A(_07798_),
    .B(_07803_),
    .C(_07808_),
    .D(_07813_),
    .Y(_07814_));
 sg13g2_xnor2_1 _27042_ (.Y(_07815_),
    .A(\cpu.intr.r_clock_cmp[9] ),
    .B(_09982_));
 sg13g2_xnor2_1 _27043_ (.Y(_07816_),
    .A(\cpu.intr.r_clock_cmp[27] ),
    .B(_05154_));
 sg13g2_xnor2_1 _27044_ (.Y(_07817_),
    .A(\cpu.intr.r_clock_cmp[31] ),
    .B(_05262_));
 sg13g2_xnor2_1 _27045_ (.Y(_07818_),
    .A(\cpu.intr.r_clock_cmp[14] ),
    .B(_10008_));
 sg13g2_nand4_1 _27046_ (.B(_07816_),
    .C(_07817_),
    .A(_07815_),
    .Y(_07819_),
    .D(_07818_));
 sg13g2_xnor2_1 _27047_ (.Y(_07820_),
    .A(\cpu.intr.r_clock_cmp[4] ),
    .B(_09948_));
 sg13g2_xnor2_1 _27048_ (.Y(_07821_),
    .A(\cpu.intr.r_clock_cmp[25] ),
    .B(_05733_));
 sg13g2_xnor2_1 _27049_ (.Y(_07822_),
    .A(\cpu.intr.r_clock_cmp[19] ),
    .B(_05434_));
 sg13g2_xnor2_1 _27050_ (.Y(_07823_),
    .A(\cpu.intr.r_clock_cmp[12] ),
    .B(_09998_));
 sg13g2_nand4_1 _27051_ (.B(_07821_),
    .C(_07822_),
    .A(_07820_),
    .Y(_07824_),
    .D(_07823_));
 sg13g2_xnor2_1 _27052_ (.Y(_07825_),
    .A(\cpu.intr.r_clock_cmp[6] ),
    .B(_09959_));
 sg13g2_xnor2_1 _27053_ (.Y(_07826_),
    .A(\cpu.intr.r_clock_cmp[18] ),
    .B(_05388_));
 sg13g2_xnor2_1 _27054_ (.Y(_07827_),
    .A(\cpu.intr.r_clock_cmp[20] ),
    .B(_05555_));
 sg13g2_xnor2_1 _27055_ (.Y(_07828_),
    .A(\cpu.intr.r_clock_cmp[16] ),
    .B(_04916_));
 sg13g2_nand4_1 _27056_ (.B(_07826_),
    .C(_07827_),
    .A(_07825_),
    .Y(_07829_),
    .D(_07828_));
 sg13g2_xnor2_1 _27057_ (.Y(_07830_),
    .A(\cpu.intr.r_clock_cmp[2] ),
    .B(_09938_));
 sg13g2_xnor2_1 _27058_ (.Y(_07831_),
    .A(\cpu.intr.r_clock_cmp[22] ),
    .B(_05668_));
 sg13g2_xnor2_1 _27059_ (.Y(_07832_),
    .A(\cpu.intr.r_clock_cmp[15] ),
    .B(_10013_));
 sg13g2_xnor2_1 _27060_ (.Y(_07833_),
    .A(\cpu.intr.r_clock_cmp[10] ),
    .B(_09987_));
 sg13g2_nand4_1 _27061_ (.B(_07831_),
    .C(_07832_),
    .A(_07830_),
    .Y(_07834_),
    .D(_07833_));
 sg13g2_nor4_1 _27062_ (.A(_07819_),
    .B(_07824_),
    .C(_07829_),
    .D(_07834_),
    .Y(_07835_));
 sg13g2_nor2_1 _27063_ (.A(net575),
    .B(_07793_),
    .Y(_07836_));
 sg13g2_a221oi_1 _27064_ (.B2(_07835_),
    .C1(_07836_),
    .B1(_07814_),
    .A1(_08968_),
    .Y(_07837_),
    .A2(_07793_));
 sg13g2_nor2_1 _27065_ (.A(net545),
    .B(_07837_),
    .Y(_02406_));
 sg13g2_and2_1 _27066_ (.A(net130),
    .B(net289),
    .X(_07838_));
 sg13g2_buf_1 _27067_ (.A(_07838_),
    .X(_07839_));
 sg13g2_nand2_1 _27068_ (.Y(_07840_),
    .A(net970),
    .B(_07839_));
 sg13g2_nand2_1 _27069_ (.Y(_07841_),
    .A(net130),
    .B(net289));
 sg13g2_buf_1 _27070_ (.A(_07841_),
    .X(_07842_));
 sg13g2_nand2_1 _27071_ (.Y(_07843_),
    .A(\cpu.intr.r_enable[0] ),
    .B(_07842_));
 sg13g2_a21oi_1 _27072_ (.A1(_07840_),
    .A2(_07843_),
    .Y(_02455_),
    .B1(net543));
 sg13g2_nand2_1 _27073_ (.Y(_07844_),
    .A(net1018),
    .B(_07839_));
 sg13g2_nand2_1 _27074_ (.Y(_07845_),
    .A(\cpu.intr.r_enable[1] ),
    .B(_07842_));
 sg13g2_a21oi_1 _27075_ (.A1(_07844_),
    .A2(_07845_),
    .Y(_02456_),
    .B1(net543));
 sg13g2_nand2_1 _27076_ (.Y(_07846_),
    .A(net1017),
    .B(_07839_));
 sg13g2_nand2_1 _27077_ (.Y(_07847_),
    .A(_08970_),
    .B(_07842_));
 sg13g2_a21oi_1 _27078_ (.A1(_07846_),
    .A2(_07847_),
    .Y(_02457_),
    .B1(net543));
 sg13g2_nand2_1 _27079_ (.Y(_07848_),
    .A(net1106),
    .B(_07839_));
 sg13g2_nand2_1 _27080_ (.Y(_07849_),
    .A(\cpu.intr.r_enable[3] ),
    .B(_07842_));
 sg13g2_a21oi_1 _27081_ (.A1(_07848_),
    .A2(_07849_),
    .Y(_02458_),
    .B1(net543));
 sg13g2_nand2_1 _27082_ (.Y(_07850_),
    .A(net1105),
    .B(_07839_));
 sg13g2_nand2_1 _27083_ (.Y(_07851_),
    .A(_09008_),
    .B(_07842_));
 sg13g2_a21oi_1 _27084_ (.A1(_07850_),
    .A2(_07851_),
    .Y(_02459_),
    .B1(net543));
 sg13g2_nand2_1 _27085_ (.Y(_07852_),
    .A(net1021),
    .B(_07839_));
 sg13g2_nand2_1 _27086_ (.Y(_07853_),
    .A(\cpu.intr.r_enable[5] ),
    .B(_07842_));
 sg13g2_buf_1 _27087_ (.A(_09136_),
    .X(_07854_));
 sg13g2_a21oi_1 _27088_ (.A1(_07852_),
    .A2(_07853_),
    .Y(_02460_),
    .B1(net542));
 sg13g2_nand3_1 _27089_ (.B(net130),
    .C(net355),
    .A(net1017),
    .Y(_07855_));
 sg13g2_nand3_1 _27090_ (.B(_06561_),
    .C(net357),
    .A(_09881_),
    .Y(_07856_));
 sg13g2_nand2_1 _27091_ (.Y(_07857_),
    .A(_09819_),
    .B(_07856_));
 sg13g2_a21oi_1 _27092_ (.A1(_08969_),
    .A2(_07855_),
    .Y(_07858_),
    .B1(_07857_));
 sg13g2_nor2_1 _27093_ (.A(net545),
    .B(_07858_),
    .Y(_02461_));
 sg13g2_and2_1 _27094_ (.A(_09658_),
    .B(_06725_),
    .X(_07859_));
 sg13g2_nand4_1 _27095_ (.B(_06749_),
    .C(_06726_),
    .A(_09704_),
    .Y(_07860_),
    .D(_07859_));
 sg13g2_buf_1 _27096_ (.A(_07860_),
    .X(_07861_));
 sg13g2_o21ai_1 _27097_ (.B1(net783),
    .Y(_07862_),
    .A1(_06748_),
    .A2(_07861_));
 sg13g2_nor2b_1 _27098_ (.A(_09697_),
    .B_N(_09720_),
    .Y(_07863_));
 sg13g2_o21ai_1 _27099_ (.B1(net19),
    .Y(_07864_),
    .A1(_07861_),
    .A2(_07863_));
 sg13g2_nand2b_1 _27100_ (.Y(_02491_),
    .B(_07864_),
    .A_N(_07862_));
 sg13g2_nand3b_1 _27101_ (.B(_06721_),
    .C(_09660_),
    .Y(_07865_),
    .A_N(_09720_));
 sg13g2_a21o_1 _27102_ (.A2(_07865_),
    .A1(_06748_),
    .B1(_07861_),
    .X(_07866_));
 sg13g2_nand2_1 _27103_ (.Y(_07867_),
    .A(_09720_),
    .B(_06748_));
 sg13g2_nor2_1 _27104_ (.A(_09693_),
    .B(_07867_),
    .Y(_07868_));
 sg13g2_o21ai_1 _27105_ (.B1(net20),
    .Y(_07869_),
    .A1(_07861_),
    .A2(_07868_));
 sg13g2_nand3_1 _27106_ (.B(_07866_),
    .C(_07869_),
    .A(net687),
    .Y(_02492_));
 sg13g2_nor2b_1 _27107_ (.A(_09695_),
    .B_N(_09720_),
    .Y(_07870_));
 sg13g2_buf_1 _27108_ (.A(\cpu.gpio.genblk1[3].srcs_o[11] ),
    .X(_07871_));
 sg13g2_o21ai_1 _27109_ (.B1(_07871_),
    .Y(_07872_),
    .A1(_07861_),
    .A2(_07870_));
 sg13g2_nand2b_1 _27110_ (.Y(_02493_),
    .B(_07872_),
    .A_N(_07862_));
 sg13g2_nor3_1 _27111_ (.A(_09163_),
    .B(_09671_),
    .C(_06721_),
    .Y(_07873_));
 sg13g2_nand3_1 _27112_ (.B(_06617_),
    .C(_07873_),
    .A(_06610_),
    .Y(_07874_));
 sg13g2_nor3_1 _27113_ (.A(_09678_),
    .B(_06724_),
    .C(_07874_),
    .Y(_07875_));
 sg13g2_a21oi_1 _27114_ (.A1(_06749_),
    .A2(_07875_),
    .Y(_07876_),
    .B1(_09660_));
 sg13g2_nor2_1 _27115_ (.A(net545),
    .B(_07876_),
    .Y(_02494_));
 sg13g2_nand2_1 _27116_ (.Y(_07877_),
    .A(net1104),
    .B(_06658_));
 sg13g2_nand2_1 _27117_ (.Y(_07878_),
    .A(\cpu.qspi.r_mask[0] ),
    .B(_06661_));
 sg13g2_a21oi_1 _27118_ (.A1(_07877_),
    .A2(_07878_),
    .Y(_02495_),
    .B1(_07854_));
 sg13g2_nor3_1 _27119_ (.A(net993),
    .B(_04925_),
    .C(_06656_),
    .Y(_07879_));
 sg13g2_inv_1 _27120_ (.Y(_07880_),
    .A(_07097_));
 sg13g2_a22oi_1 _27121_ (.Y(_07881_),
    .B1(_07879_),
    .B2(_07880_),
    .A2(_06672_),
    .A1(\cpu.qspi.r_mask[1] ));
 sg13g2_nand2_1 _27122_ (.Y(_02496_),
    .A(net622),
    .B(_07881_));
 sg13g2_nor2_1 _27123_ (.A(_07097_),
    .B(_06685_),
    .Y(_07882_));
 sg13g2_a21oi_1 _27124_ (.A1(\cpu.qspi.r_mask[2] ),
    .A2(_06685_),
    .Y(_07883_),
    .B1(_07882_));
 sg13g2_nor2_1 _27125_ (.A(net545),
    .B(_07883_),
    .Y(_02497_));
 sg13g2_nand2_1 _27126_ (.Y(_07884_),
    .A(\cpu.qspi.r_quad[0] ),
    .B(_06661_));
 sg13g2_nand2_1 _27127_ (.Y(_07885_),
    .A(_09908_),
    .B(_06658_));
 sg13g2_nand3_1 _27128_ (.B(_07884_),
    .C(_07885_),
    .A(net687),
    .Y(_02498_));
 sg13g2_a22oi_1 _27129_ (.Y(_07886_),
    .B1(_07879_),
    .B2(_07092_),
    .A2(_06672_),
    .A1(\cpu.qspi.r_quad[1] ));
 sg13g2_nor2_1 _27130_ (.A(net545),
    .B(_07886_),
    .Y(_02499_));
 sg13g2_nand2_1 _27131_ (.Y(_07887_),
    .A(_00166_),
    .B(_06682_));
 sg13g2_o21ai_1 _27132_ (.B1(_07887_),
    .Y(_07888_),
    .A1(\cpu.qspi.r_quad[2] ),
    .A2(_06682_));
 sg13g2_nand2_1 _27133_ (.Y(_02500_),
    .A(net622),
    .B(_07888_));
 sg13g2_or2_1 _27134_ (.X(_07889_),
    .B(_06656_),
    .A(_04891_));
 sg13g2_buf_1 _27135_ (.A(_07889_),
    .X(_07890_));
 sg13g2_mux2_1 _27136_ (.A0(net1024),
    .A1(_09684_),
    .S(_07890_),
    .X(_07891_));
 sg13g2_nand2b_1 _27137_ (.Y(_02513_),
    .B(net622),
    .A_N(_07891_));
 sg13g2_mux2_1 _27138_ (.A0(net1023),
    .A1(_09683_),
    .S(_07890_),
    .X(_07892_));
 sg13g2_nand2b_1 _27139_ (.Y(_02514_),
    .B(_07450_),
    .A_N(_07892_));
 sg13g2_or2_1 _27140_ (.X(_07893_),
    .B(_09705_),
    .A(_11885_));
 sg13g2_nor2_1 _27141_ (.A(_11883_),
    .B(_06721_),
    .Y(_07894_));
 sg13g2_nand2_1 _27142_ (.Y(_07895_),
    .A(_06609_),
    .B(_07894_));
 sg13g2_o21ai_1 _27143_ (.B1(_07894_),
    .Y(_07896_),
    .A1(_07893_),
    .A2(_07895_));
 sg13g2_nand2b_1 _27144_ (.Y(_07897_),
    .B(_11885_),
    .A_N(_06747_));
 sg13g2_nor3_1 _27145_ (.A(_11902_),
    .B(_09723_),
    .C(_09681_),
    .Y(_07898_));
 sg13g2_and4_1 _27146_ (.A(_06617_),
    .B(_07859_),
    .C(_07897_),
    .D(_07898_),
    .X(_07899_));
 sg13g2_buf_1 _27147_ (.A(_07899_),
    .X(_07900_));
 sg13g2_mux2_1 _27148_ (.A0(net3),
    .A1(_07896_),
    .S(_07900_),
    .X(_07901_));
 sg13g2_and2_1 _27149_ (.A(_11884_),
    .B(_07901_),
    .X(_02515_));
 sg13g2_nand2b_1 _27150_ (.Y(_07902_),
    .B(net6),
    .A_N(_07900_));
 sg13g2_nor3_1 _27151_ (.A(_09700_),
    .B(_07893_),
    .C(_07895_),
    .Y(_07903_));
 sg13g2_o21ai_1 _27152_ (.B1(_07900_),
    .Y(_07904_),
    .A1(_11883_),
    .A2(_07903_));
 sg13g2_a21oi_1 _27153_ (.A1(_07902_),
    .A2(_07904_),
    .Y(_02516_),
    .B1(_07854_));
 sg13g2_nor3_1 _27154_ (.A(net1034),
    .B(_09044_),
    .C(_09132_),
    .Y(_07905_));
 sg13g2_a221oi_1 _27155_ (.B2(net1034),
    .C1(_07905_),
    .B1(_09113_),
    .A1(net1033),
    .Y(_07906_),
    .A2(_09054_));
 sg13g2_buf_1 _27156_ (.A(_07906_),
    .X(_07907_));
 sg13g2_nand3_1 _27157_ (.B(net1034),
    .C(_07907_),
    .A(_09059_),
    .Y(_07908_));
 sg13g2_o21ai_1 _27158_ (.B1(_07908_),
    .Y(_07909_),
    .A1(_09059_),
    .A2(_07907_));
 sg13g2_nand2_1 _27159_ (.Y(_02522_),
    .A(net622),
    .B(_07909_));
 sg13g2_inv_1 _27160_ (.Y(_07910_),
    .A(_11910_));
 sg13g2_nand2_1 _27161_ (.Y(_07911_),
    .A(_09059_),
    .B(_07910_));
 sg13g2_a21oi_1 _27162_ (.A1(_07907_),
    .A2(_07911_),
    .Y(_07912_),
    .B1(_09060_));
 sg13g2_inv_1 _27163_ (.Y(_07913_),
    .A(_09059_));
 sg13g2_and4_1 _27164_ (.A(_07913_),
    .B(_09060_),
    .C(_07910_),
    .D(_07907_),
    .X(_07914_));
 sg13g2_o21ai_1 _27165_ (.B1(net622),
    .Y(_02523_),
    .A1(_07912_),
    .A2(_07914_));
 sg13g2_nor2_1 _27166_ (.A(_09059_),
    .B(_09060_),
    .Y(_07915_));
 sg13g2_or2_1 _27167_ (.X(_07916_),
    .B(_07915_),
    .A(_11910_));
 sg13g2_a21oi_1 _27168_ (.A1(_07907_),
    .A2(_07916_),
    .Y(_07917_),
    .B1(\cpu.spi.r_bits[2] ));
 sg13g2_and4_1 _27169_ (.A(\cpu.spi.r_bits[2] ),
    .B(_07910_),
    .C(_07915_),
    .D(_07907_),
    .X(_07918_));
 sg13g2_o21ai_1 _27170_ (.B1(net622),
    .Y(_02524_),
    .A1(_07917_),
    .A2(_07918_));
 sg13g2_buf_1 _27171_ (.A(\cpu.gpio.genblk1[3].srcs_o[6] ),
    .X(_07919_));
 sg13g2_inv_1 _27172_ (.Y(_07920_),
    .A(net1066));
 sg13g2_a21oi_1 _27173_ (.A1(_09043_),
    .A2(_09054_),
    .Y(_07921_),
    .B1(_06864_));
 sg13g2_or2_1 _27174_ (.X(_07922_),
    .B(_09127_),
    .A(_09044_));
 sg13g2_buf_1 _27175_ (.A(_07922_),
    .X(_07923_));
 sg13g2_nand2_1 _27176_ (.Y(_07924_),
    .A(net379),
    .B(_07923_));
 sg13g2_nor3_1 _27177_ (.A(net1110),
    .B(_09093_),
    .C(_07923_),
    .Y(_07925_));
 sg13g2_a21oi_1 _27178_ (.A1(net996),
    .A2(_06872_),
    .Y(_07926_),
    .B1(net378));
 sg13g2_nor3_1 _27179_ (.A(_00256_),
    .B(_07925_),
    .C(_07926_),
    .Y(_07927_));
 sg13g2_a21oi_1 _27180_ (.A1(_00256_),
    .A2(_07924_),
    .Y(_07928_),
    .B1(_07927_));
 sg13g2_nand2b_1 _27181_ (.Y(_07929_),
    .B(_07928_),
    .A_N(_07921_));
 sg13g2_buf_1 _27182_ (.A(_07929_),
    .X(_07930_));
 sg13g2_nor3_1 _27183_ (.A(_11914_),
    .B(net728),
    .C(_07930_),
    .Y(_07931_));
 sg13g2_inv_1 _27184_ (.Y(_07932_),
    .A(_07930_));
 sg13g2_a21oi_1 _27185_ (.A1(_07923_),
    .A2(_07932_),
    .Y(_07933_),
    .B1(_09136_));
 sg13g2_o21ai_1 _27186_ (.B1(_07933_),
    .Y(_02557_),
    .A1(_07920_),
    .A2(_07931_));
 sg13g2_nand2_1 _27187_ (.Y(_07934_),
    .A(_11926_),
    .B(_11930_));
 sg13g2_buf_1 _27188_ (.A(\cpu.gpio.genblk1[3].srcs_o[7] ),
    .X(_07935_));
 sg13g2_o21ai_1 _27189_ (.B1(net1065),
    .Y(_07936_),
    .A1(_07930_),
    .A2(_07934_));
 sg13g2_nand2_1 _27190_ (.Y(_02558_),
    .A(_07933_),
    .B(_07936_));
 sg13g2_buf_1 _27191_ (.A(\cpu.gpio.genblk1[3].srcs_o[8] ),
    .X(_07937_));
 sg13g2_inv_1 _27192_ (.Y(_07938_),
    .A(net1064));
 sg13g2_nor3_1 _27193_ (.A(_11926_),
    .B(_11930_),
    .C(_07930_),
    .Y(_07939_));
 sg13g2_o21ai_1 _27194_ (.B1(_07933_),
    .Y(_02559_),
    .A1(_07938_),
    .A2(_07939_));
 sg13g2_or2_1 _27195_ (.X(_07940_),
    .B(_09043_),
    .A(_06864_));
 sg13g2_o21ai_1 _27196_ (.B1(_09160_),
    .Y(_07941_),
    .A1(_09108_),
    .A2(_07940_));
 sg13g2_nand2_1 _27197_ (.Y(_07942_),
    .A(_09082_),
    .B(net379));
 sg13g2_a21oi_1 _27198_ (.A1(net1034),
    .A2(_07942_),
    .Y(_07943_),
    .B1(_07905_));
 sg13g2_nor2b_1 _27199_ (.A(_07941_),
    .B_N(_07943_),
    .Y(_07944_));
 sg13g2_mux2_1 _27200_ (.A0(_08976_),
    .A1(_09058_),
    .S(_07944_),
    .X(_07945_));
 sg13g2_and2_1 _27201_ (.A(net648),
    .B(_07945_),
    .X(_02568_));
 sg13g2_nor3_1 _27202_ (.A(net1034),
    .B(_09132_),
    .C(_07923_),
    .Y(_07946_));
 sg13g2_a21oi_1 _27203_ (.A1(net1034),
    .A2(_07942_),
    .Y(_07947_),
    .B1(_07946_));
 sg13g2_nor2b_1 _27204_ (.A(_07941_),
    .B_N(_07947_),
    .Y(_07948_));
 sg13g2_nand3b_1 _27205_ (.B(_09056_),
    .C(_07948_),
    .Y(_07949_),
    .A_N(_09127_));
 sg13g2_o21ai_1 _27206_ (.B1(_07949_),
    .Y(_07950_),
    .A1(\cpu.spi.r_ready ),
    .A2(_09095_));
 sg13g2_nor2_1 _27207_ (.A(\cpu.spi.r_ready ),
    .B(_07948_),
    .Y(_07951_));
 sg13g2_a21oi_1 _27208_ (.A1(_09114_),
    .A2(_07950_),
    .Y(_07952_),
    .B1(_07951_));
 sg13g2_nand2b_1 _27209_ (.Y(_02583_),
    .B(net622),
    .A_N(_07952_));
 sg13g2_and2_1 _27210_ (.A(_09056_),
    .B(_07943_),
    .X(_07953_));
 sg13g2_nand2b_1 _27211_ (.Y(_07954_),
    .B(\cpu.spi.r_searching ),
    .A_N(_07953_));
 sg13g2_nand3b_1 _27212_ (.B(_09040_),
    .C(_07953_),
    .Y(_07955_),
    .A_N(_06864_));
 sg13g2_a21oi_1 _27213_ (.A1(_07954_),
    .A2(_07955_),
    .Y(_02584_),
    .B1(net542));
 sg13g2_buf_1 _27214_ (.A(_07179_),
    .X(_07956_));
 sg13g2_and2_1 _27215_ (.A(_04890_),
    .B(net106),
    .X(_07957_));
 sg13g2_buf_2 _27216_ (.A(_07957_),
    .X(_07958_));
 sg13g2_nand2_1 _27217_ (.Y(_07959_),
    .A(_02832_),
    .B(_07958_));
 sg13g2_nand2_1 _27218_ (.Y(_07960_),
    .A(_04890_),
    .B(_07179_));
 sg13g2_buf_2 _27219_ (.A(_07960_),
    .X(_07961_));
 sg13g2_nand2_1 _27220_ (.Y(_07962_),
    .A(\cpu.uart.r_div_value[0] ),
    .B(_07961_));
 sg13g2_nand3_1 _27221_ (.B(_07959_),
    .C(_07962_),
    .A(net687),
    .Y(_02606_));
 sg13g2_nand3_1 _27222_ (.B(net355),
    .C(net106),
    .A(net1017),
    .Y(_07963_));
 sg13g2_nand2_1 _27223_ (.Y(_07964_),
    .A(net355),
    .B(_07956_));
 sg13g2_nand2_1 _27224_ (.Y(_07965_),
    .A(_09766_),
    .B(_07964_));
 sg13g2_a21oi_1 _27225_ (.A1(_07963_),
    .A2(_07965_),
    .Y(_02607_),
    .B1(net542));
 sg13g2_nand3_1 _27226_ (.B(net355),
    .C(_07956_),
    .A(net1106),
    .Y(_07966_));
 sg13g2_nand2_1 _27227_ (.Y(_07967_),
    .A(\cpu.uart.r_div_value[11] ),
    .B(_07964_));
 sg13g2_a21oi_1 _27228_ (.A1(_07966_),
    .A2(_07967_),
    .Y(_02608_),
    .B1(net542));
 sg13g2_nand2_1 _27229_ (.Y(_07968_),
    .A(net1018),
    .B(_07958_));
 sg13g2_nand2_1 _27230_ (.Y(_07969_),
    .A(\cpu.uart.r_div_value[1] ),
    .B(_07961_));
 sg13g2_a21oi_1 _27231_ (.A1(_07968_),
    .A2(_07969_),
    .Y(_02609_),
    .B1(net542));
 sg13g2_nand2_1 _27232_ (.Y(_07970_),
    .A(net1017),
    .B(_07958_));
 sg13g2_nand2_1 _27233_ (.Y(_07971_),
    .A(\cpu.uart.r_div_value[2] ),
    .B(_07961_));
 sg13g2_a21oi_1 _27234_ (.A1(_07970_),
    .A2(_07971_),
    .Y(_02610_),
    .B1(net542));
 sg13g2_nand2_1 _27235_ (.Y(_07972_),
    .A(net1106),
    .B(_07958_));
 sg13g2_nand2_1 _27236_ (.Y(_07973_),
    .A(\cpu.uart.r_div_value[3] ),
    .B(_07961_));
 sg13g2_a21oi_1 _27237_ (.A1(_07972_),
    .A2(_07973_),
    .Y(_02611_),
    .B1(net542));
 sg13g2_nand2_1 _27238_ (.Y(_07974_),
    .A(net1105),
    .B(_07958_));
 sg13g2_nand2_1 _27239_ (.Y(_07975_),
    .A(\cpu.uart.r_div_value[4] ),
    .B(_07961_));
 sg13g2_a21oi_1 _27240_ (.A1(_07974_),
    .A2(_07975_),
    .Y(_02612_),
    .B1(net542));
 sg13g2_nand2_1 _27241_ (.Y(_07976_),
    .A(_09902_),
    .B(_07958_));
 sg13g2_nand2_1 _27242_ (.Y(_07977_),
    .A(\cpu.uart.r_div_value[5] ),
    .B(_07961_));
 sg13g2_a21oi_1 _27243_ (.A1(_07976_),
    .A2(_07977_),
    .Y(_02613_),
    .B1(net647));
 sg13g2_nand2_1 _27244_ (.Y(_07978_),
    .A(_09908_),
    .B(_07958_));
 sg13g2_nand2_1 _27245_ (.Y(_07979_),
    .A(\cpu.uart.r_div_value[6] ),
    .B(_07961_));
 sg13g2_a21oi_1 _27246_ (.A1(_07978_),
    .A2(_07979_),
    .Y(_02614_),
    .B1(net647));
 sg13g2_nand2_1 _27247_ (.Y(_07980_),
    .A(net1104),
    .B(_07958_));
 sg13g2_nand2_1 _27248_ (.Y(_07981_),
    .A(\cpu.uart.r_div_value[7] ),
    .B(_07961_));
 sg13g2_a21oi_1 _27249_ (.A1(_07980_),
    .A2(_07981_),
    .Y(_02615_),
    .B1(net647));
 sg13g2_nand3_1 _27250_ (.B(net355),
    .C(net106),
    .A(net1024),
    .Y(_07982_));
 sg13g2_nand2_1 _27251_ (.Y(_07983_),
    .A(\cpu.uart.r_div_value[8] ),
    .B(_07964_));
 sg13g2_a21oi_1 _27252_ (.A1(_07982_),
    .A2(_07983_),
    .Y(_02616_),
    .B1(net647));
 sg13g2_nand3_1 _27253_ (.B(net355),
    .C(net106),
    .A(net1023),
    .Y(_07984_));
 sg13g2_nand2_1 _27254_ (.Y(_07985_),
    .A(\cpu.uart.r_div_value[9] ),
    .B(_07964_));
 sg13g2_a21oi_1 _27255_ (.A1(_07984_),
    .A2(_07985_),
    .Y(_02617_),
    .B1(_11904_));
 sg13g2_nand3_1 _27256_ (.B(_07177_),
    .C(_06857_),
    .A(_08187_),
    .Y(_07986_));
 sg13g2_nor4_1 _27257_ (.A(net966),
    .B(net575),
    .C(net676),
    .D(_07986_),
    .Y(_07987_));
 sg13g2_nand2_1 _27258_ (.Y(_07988_),
    .A(_08973_),
    .B(net901));
 sg13g2_a21oi_1 _27259_ (.A1(_09017_),
    .A2(_07987_),
    .Y(_07989_),
    .B1(_07988_));
 sg13g2_nand3_1 _27260_ (.B(_04924_),
    .C(net106),
    .A(net1023),
    .Y(_07990_));
 sg13g2_a21o_1 _27261_ (.A2(_07990_),
    .A1(_07989_),
    .B1(net127),
    .X(_02641_));
 sg13g2_nand3_1 _27262_ (.B(net404),
    .C(net106),
    .A(net1023),
    .Y(_07991_));
 sg13g2_nand2_1 _27263_ (.Y(_07992_),
    .A(net404),
    .B(net106));
 sg13g2_nand2_1 _27264_ (.Y(_07993_),
    .A(\cpu.uart.r_r_invert ),
    .B(_07992_));
 sg13g2_a21oi_1 _27265_ (.A1(_07991_),
    .A2(_07993_),
    .Y(_02642_),
    .B1(net647));
 sg13g2_a21oi_1 _27266_ (.A1(_07160_),
    .A2(_09743_),
    .Y(_07994_),
    .B1(_07155_));
 sg13g2_a21oi_1 _27267_ (.A1(_07161_),
    .A2(net252),
    .Y(_07995_),
    .B1(_07233_));
 sg13g2_a221oi_1 _27268_ (.B2(_07994_),
    .C1(_07995_),
    .B1(_07159_),
    .A1(net921),
    .Y(_07996_),
    .A2(_07155_));
 sg13g2_a21oi_1 _27269_ (.A1(_07153_),
    .A2(_07996_),
    .Y(_07997_),
    .B1(_07242_));
 sg13g2_buf_2 _27270_ (.A(_07997_),
    .X(_07998_));
 sg13g2_o21ai_1 _27271_ (.B1(_07998_),
    .Y(_07999_),
    .A1(net921),
    .A2(_07233_));
 sg13g2_xnor2_1 _27272_ (.Y(_08000_),
    .A(_07161_),
    .B(_07999_));
 sg13g2_nor2_1 _27273_ (.A(net545),
    .B(_08000_),
    .Y(_02645_));
 sg13g2_o21ai_1 _27274_ (.B1(_07998_),
    .Y(_08001_),
    .A1(_07160_),
    .A2(net924));
 sg13g2_nand2_1 _27275_ (.Y(_08002_),
    .A(net1071),
    .B(_08001_));
 sg13g2_nand2b_1 _27276_ (.Y(_08003_),
    .B(net921),
    .A_N(net924));
 sg13g2_o21ai_1 _27277_ (.B1(_08003_),
    .Y(_08004_),
    .A1(net921),
    .A2(_07243_));
 sg13g2_nand3_1 _27278_ (.B(_07998_),
    .C(_08004_),
    .A(_07244_),
    .Y(_08005_));
 sg13g2_a21oi_1 _27279_ (.A1(_08002_),
    .A2(_08005_),
    .Y(_02646_),
    .B1(net647));
 sg13g2_nand2_1 _27280_ (.Y(_08006_),
    .A(_07160_),
    .B(net1071));
 sg13g2_nor3_1 _27281_ (.A(_07239_),
    .B(_07156_),
    .C(_08006_),
    .Y(_08007_));
 sg13g2_o21ai_1 _27282_ (.B1(_07998_),
    .Y(_08008_),
    .A1(net924),
    .A2(_07251_));
 sg13g2_a22oi_1 _27283_ (.Y(_08009_),
    .B1(_08008_),
    .B2(net921),
    .A2(_08007_),
    .A1(_07998_));
 sg13g2_nor2_1 _27284_ (.A(net545),
    .B(_08009_),
    .Y(_02647_));
 sg13g2_a21oi_1 _27285_ (.A1(_07251_),
    .A2(_07998_),
    .Y(_08010_),
    .B1(_07156_));
 sg13g2_nor2b_1 _27286_ (.A(net921),
    .B_N(_07157_),
    .Y(_08011_));
 sg13g2_a21oi_1 _27287_ (.A1(_07998_),
    .A2(_08011_),
    .Y(_08012_),
    .B1(_09136_));
 sg13g2_nor2b_1 _27288_ (.A(_08010_),
    .B_N(_08012_),
    .Y(_02648_));
 sg13g2_and2_1 _27289_ (.A(net252),
    .B(_07197_),
    .X(_08013_));
 sg13g2_and2_1 _27290_ (.A(_07176_),
    .B(_07190_),
    .X(_08014_));
 sg13g2_o21ai_1 _27291_ (.B1(_08014_),
    .Y(_08015_),
    .A1(_08972_),
    .A2(_08013_));
 sg13g2_o21ai_1 _27292_ (.B1(net598),
    .Y(_08016_),
    .A1(_00202_),
    .A2(_04896_));
 sg13g2_nor2_1 _27293_ (.A(net676),
    .B(_07187_),
    .Y(_08017_));
 sg13g2_a21o_1 _27294_ (.A2(net289),
    .A1(_09859_),
    .B1(_05340_),
    .X(_08018_));
 sg13g2_a22oi_1 _27295_ (.Y(_08019_),
    .B1(_08018_),
    .B2(_07190_),
    .A2(_08017_),
    .A1(_08016_));
 sg13g2_o21ai_1 _27296_ (.B1(_08972_),
    .Y(_08020_),
    .A1(_07182_),
    .A2(_08019_));
 sg13g2_a21oi_1 _27297_ (.A1(_08015_),
    .A2(_08020_),
    .Y(_02650_),
    .B1(net647));
 sg13g2_nand3_1 _27298_ (.B(net404),
    .C(net106),
    .A(net1024),
    .Y(_08021_));
 sg13g2_nand2_1 _27299_ (.Y(_08022_),
    .A(\cpu.uart.r_x_invert ),
    .B(_07992_));
 sg13g2_a21oi_1 _27300_ (.A1(_08021_),
    .A2(_08022_),
    .Y(_02651_),
    .B1(net647));
 sg13g2_a21oi_1 _27301_ (.A1(_05340_),
    .A2(_07179_),
    .Y(_08023_),
    .B1(_07191_));
 sg13g2_or2_1 _27302_ (.X(_08024_),
    .B(_08023_),
    .A(_07264_));
 sg13g2_a221oi_1 _27303_ (.B2(_07199_),
    .C1(_07276_),
    .B1(_08024_),
    .A1(_07181_),
    .Y(_08025_),
    .A2(_07186_));
 sg13g2_buf_2 _27304_ (.A(_08025_),
    .X(_08026_));
 sg13g2_nand2_1 _27305_ (.Y(_08027_),
    .A(_07278_),
    .B(_08026_));
 sg13g2_a21oi_1 _27306_ (.A1(_08013_),
    .A2(_07270_),
    .Y(_08028_),
    .B1(_08027_));
 sg13g2_o21ai_1 _27307_ (.B1(net779),
    .Y(_08029_),
    .A1(net1069),
    .A2(_08026_));
 sg13g2_a21oi_1 _27308_ (.A1(net1069),
    .A2(_08028_),
    .Y(_02654_),
    .B1(_08029_));
 sg13g2_o21ai_1 _27309_ (.B1(_08026_),
    .Y(_08030_),
    .A1(net1069),
    .A2(_07262_));
 sg13g2_nor3_1 _27310_ (.A(net1070),
    .B(_07176_),
    .C(_08027_),
    .Y(_08031_));
 sg13g2_a21oi_1 _27311_ (.A1(net1070),
    .A2(_08030_),
    .Y(_08032_),
    .B1(_08031_));
 sg13g2_nor2_1 _27312_ (.A(net545),
    .B(_08032_),
    .Y(_02655_));
 sg13g2_inv_1 _27313_ (.Y(_08033_),
    .A(_08026_));
 sg13g2_nand3b_1 _27314_ (.B(_07194_),
    .C(_08026_),
    .Y(_08034_),
    .A_N(net922));
 sg13g2_nand2b_1 _27315_ (.Y(_08035_),
    .B(net922),
    .A_N(_07194_));
 sg13g2_a21oi_1 _27316_ (.A1(_08034_),
    .A2(_08035_),
    .Y(_08036_),
    .B1(net923));
 sg13g2_a221oi_1 _27317_ (.B2(net922),
    .C1(_08036_),
    .B1(_08033_),
    .A1(_07199_),
    .Y(_08037_),
    .A2(_07270_));
 sg13g2_nor2_1 _27318_ (.A(net606),
    .B(_08037_),
    .Y(_02656_));
 sg13g2_a22oi_1 _27319_ (.Y(_08038_),
    .B1(_07271_),
    .B2(_07194_),
    .A2(_07270_),
    .A1(_07199_));
 sg13g2_inv_1 _27320_ (.Y(_08039_),
    .A(_08038_));
 sg13g2_o21ai_1 _27321_ (.B1(_08026_),
    .Y(_08040_),
    .A1(net922),
    .A2(_07194_));
 sg13g2_a22oi_1 _27322_ (.Y(_08041_),
    .B1(_08040_),
    .B2(net923),
    .A2(_08039_),
    .A1(_08026_));
 sg13g2_nor2_1 _27323_ (.A(net606),
    .B(_08041_),
    .Y(_02657_));
 sg13g2_nand2b_1 _27324_ (.Y(\cpu.ex.genblk3.c_supmode ),
    .B(_07445_),
    .A_N(_07441_));
 sg13g2_nor4_1 _27325_ (.A(_09723_),
    .B(_09659_),
    .C(_06724_),
    .D(_07874_),
    .Y(_08042_));
 sg13g2_nor2b_1 _27326_ (.A(_09705_),
    .B_N(_08042_),
    .Y(_08043_));
 sg13g2_a22oi_1 _27327_ (.Y(_08044_),
    .B1(_09677_),
    .B2(_08043_),
    .A2(net600),
    .A1(_09673_));
 sg13g2_inv_1 _27328_ (.Y(\cpu.qspi.c_rstrobe_d ),
    .A(_08044_));
 sg13g2_nor2_1 _27329_ (.A(_09678_),
    .B(net600),
    .Y(_08045_));
 sg13g2_a22oi_1 _27330_ (.Y(_08046_),
    .B1(_08042_),
    .B2(_08045_),
    .A2(net600),
    .A1(_09670_));
 sg13g2_nor2_1 _27331_ (.A(net801),
    .B(_08046_),
    .Y(\cpu.qspi.c_wstrobe_d ));
 sg13g2_nor2_1 _27332_ (.A(_00173_),
    .B(_08046_),
    .Y(\cpu.qspi.c_wstrobe_i ));
 sg13g2_mux4_1 _27333_ (.S0(_04967_),
    .A0(_08991_),
    .A1(_09004_),
    .A2(_09000_),
    .A3(_08980_),
    .S1(\cpu.gpio.r_uart_rx_src[1] ),
    .X(_08047_));
 sg13g2_mux4_1 _27334_ (.S0(_04967_),
    .A0(_08996_),
    .A1(_09002_),
    .A2(_08998_),
    .A3(_08987_),
    .S1(\cpu.gpio.r_uart_rx_src[1] ),
    .X(_08048_));
 sg13g2_mux2_1 _27335_ (.A0(_08047_),
    .A1(_08048_),
    .S(\cpu.gpio.r_uart_rx_src[2] ),
    .X(\cpu.gpio.uart_rx ));
 sg13g2_mux4_1 _27336_ (.S0(_04971_),
    .A0(net1090),
    .A1(net1091),
    .A2(net1066),
    .A3(net1065),
    .S1(_05315_),
    .X(_08049_));
 sg13g2_mux4_1 _27337_ (.S0(_04971_),
    .A0(\cpu.gpio.genblk2[4].srcs_io[0] ),
    .A1(net1068),
    .A2(_11981_),
    .A3(_11964_),
    .S1(_05315_),
    .X(_08050_));
 sg13g2_nor2b_1 _27338_ (.A(_05368_),
    .B_N(_08050_),
    .Y(_08051_));
 sg13g2_a21oi_1 _27339_ (.A1(_05368_),
    .A2(_08049_),
    .Y(_08052_),
    .B1(_08051_));
 sg13g2_nand2b_1 _27340_ (.Y(_08053_),
    .B(net1064),
    .A_N(_04971_));
 sg13g2_nand3_1 _27341_ (.B(_05315_),
    .C(net1067),
    .A(_04971_),
    .Y(_08054_));
 sg13g2_o21ai_1 _27342_ (.B1(_08054_),
    .Y(_08055_),
    .A1(_05315_),
    .A2(_08053_));
 sg13g2_nand3_1 _27343_ (.B(_00171_),
    .C(_08055_),
    .A(_05453_),
    .Y(_08056_));
 sg13g2_o21ai_1 _27344_ (.B1(_08056_),
    .Y(net15),
    .A1(_05453_),
    .A2(_08052_));
 sg13g2_mux4_1 _27345_ (.S0(_05535_),
    .A0(net1090),
    .A1(net1091),
    .A2(net1066),
    .A3(net1065),
    .S1(_05607_),
    .X(_08057_));
 sg13g2_mux4_1 _27346_ (.S0(_05535_),
    .A0(\cpu.gpio.genblk2[5].srcs_io[0] ),
    .A1(net1068),
    .A2(net1088),
    .A3(net1089),
    .S1(_05607_),
    .X(_08058_));
 sg13g2_nor2b_1 _27347_ (.A(_05693_),
    .B_N(_08058_),
    .Y(_08059_));
 sg13g2_a21oi_1 _27348_ (.A1(_05693_),
    .A2(_08057_),
    .Y(_08060_),
    .B1(_08059_));
 sg13g2_nand2b_1 _27349_ (.Y(_08061_),
    .B(net1064),
    .A_N(_05535_));
 sg13g2_nand3_1 _27350_ (.B(_05607_),
    .C(net1067),
    .A(_05535_),
    .Y(_08062_));
 sg13g2_o21ai_1 _27351_ (.B1(_08062_),
    .Y(_08063_),
    .A1(_05607_),
    .A2(_08061_));
 sg13g2_nand3_1 _27352_ (.B(_00170_),
    .C(_08063_),
    .A(_05105_),
    .Y(_08064_));
 sg13g2_o21ai_1 _27353_ (.B1(_08064_),
    .Y(net16),
    .A1(_05105_),
    .A2(_08060_));
 sg13g2_mux4_1 _27354_ (.S0(_04975_),
    .A0(net1090),
    .A1(net1091),
    .A2(net1066),
    .A3(net1065),
    .S1(_06250_),
    .X(_08065_));
 sg13g2_mux4_1 _27355_ (.S0(_04975_),
    .A0(\cpu.gpio.genblk2[6].srcs_io[0] ),
    .A1(net1068),
    .A2(net1088),
    .A3(net1089),
    .S1(_06250_),
    .X(_08066_));
 sg13g2_nor2b_1 _27356_ (.A(\cpu.gpio.r_src_io[6][2] ),
    .B_N(_08066_),
    .Y(_08067_));
 sg13g2_a21oi_1 _27357_ (.A1(\cpu.gpio.r_src_io[6][2] ),
    .A2(_08065_),
    .Y(_08068_),
    .B1(_08067_));
 sg13g2_nand2b_1 _27358_ (.Y(_08069_),
    .B(net1064),
    .A_N(_04975_));
 sg13g2_nand3_1 _27359_ (.B(net1067),
    .C(_06250_),
    .A(_04975_),
    .Y(_08070_));
 sg13g2_o21ai_1 _27360_ (.B1(_08070_),
    .Y(_08071_),
    .A1(_06250_),
    .A2(_08069_));
 sg13g2_nand3_1 _27361_ (.B(\cpu.gpio.r_src_io[6][3] ),
    .C(_08071_),
    .A(_00096_),
    .Y(_08072_));
 sg13g2_o21ai_1 _27362_ (.B1(_08072_),
    .Y(net17),
    .A1(\cpu.gpio.r_src_io[6][3] ),
    .A2(_08068_));
 sg13g2_mux4_1 _27363_ (.S0(_05537_),
    .A0(net1090),
    .A1(_11956_),
    .A2(_07919_),
    .A3(net1065),
    .S1(_06251_),
    .X(_08073_));
 sg13g2_mux4_1 _27364_ (.S0(_05537_),
    .A0(\cpu.gpio.genblk2[7].srcs_io[0] ),
    .A1(net1068),
    .A2(_11981_),
    .A3(_11964_),
    .S1(_06251_),
    .X(_08074_));
 sg13g2_nor2b_1 _27365_ (.A(\cpu.gpio.r_src_io[7][2] ),
    .B_N(_08074_),
    .Y(_08075_));
 sg13g2_a21oi_1 _27366_ (.A1(\cpu.gpio.r_src_io[7][2] ),
    .A2(_08073_),
    .Y(_08076_),
    .B1(_08075_));
 sg13g2_nand2b_1 _27367_ (.Y(_08077_),
    .B(_07937_),
    .A_N(_05537_));
 sg13g2_nand3_1 _27368_ (.B(net1067),
    .C(_06251_),
    .A(_05537_),
    .Y(_08078_));
 sg13g2_o21ai_1 _27369_ (.B1(_08078_),
    .Y(_08079_),
    .A1(_06251_),
    .A2(_08077_));
 sg13g2_nand3_1 _27370_ (.B(\cpu.gpio.r_src_io[7][3] ),
    .C(_08079_),
    .A(_00133_),
    .Y(_08080_));
 sg13g2_o21ai_1 _27371_ (.B1(_08080_),
    .Y(net18),
    .A1(\cpu.gpio.r_src_io[7][3] ),
    .A2(_08076_));
 sg13g2_xor2_1 _27372_ (.B(clknet_leaf_76_clk),
    .A(\cpu.r_clk_invert ),
    .X(net21));
 sg13g2_mux4_1 _27373_ (.S0(_05531_),
    .A0(net1090),
    .A1(net1091),
    .A2(net1066),
    .A3(_07935_),
    .S1(_06253_),
    .X(_08081_));
 sg13g2_mux4_1 _27374_ (.S0(_05531_),
    .A0(\cpu.gpio.genblk1[3].srcs_o[0] ),
    .A1(_07260_),
    .A2(net1088),
    .A3(net1089),
    .S1(_06253_),
    .X(_08082_));
 sg13g2_nor2b_1 _27375_ (.A(\cpu.gpio.r_src_o[3][2] ),
    .B_N(_08082_),
    .Y(_08083_));
 sg13g2_a21oi_1 _27376_ (.A1(\cpu.gpio.r_src_o[3][2] ),
    .A2(_08081_),
    .Y(_08084_),
    .B1(_08083_));
 sg13g2_nand2b_1 _27377_ (.Y(_08085_),
    .B(net1064),
    .A_N(_05531_));
 sg13g2_nand3_1 _27378_ (.B(net1067),
    .C(_06253_),
    .A(_05531_),
    .Y(_08086_));
 sg13g2_o21ai_1 _27379_ (.B1(_08086_),
    .Y(_08087_),
    .A1(_06253_),
    .A2(_08085_));
 sg13g2_nand3_1 _27380_ (.B(\cpu.gpio.r_src_o[3][3] ),
    .C(_08087_),
    .A(_00136_),
    .Y(_08088_));
 sg13g2_o21ai_1 _27381_ (.B1(_08088_),
    .Y(net22),
    .A1(\cpu.gpio.r_src_o[3][3] ),
    .A2(_08084_));
 sg13g2_mux4_1 _27382_ (.S0(_04982_),
    .A0(_11962_),
    .A1(_11956_),
    .A2(net1066),
    .A3(_07935_),
    .S1(_06256_),
    .X(_08089_));
 sg13g2_mux4_1 _27383_ (.S0(_04982_),
    .A0(\cpu.gpio.genblk1[4].srcs_o[0] ),
    .A1(net1068),
    .A2(net1088),
    .A3(net1089),
    .S1(_06256_),
    .X(_08090_));
 sg13g2_nor2b_1 _27384_ (.A(\cpu.gpio.r_src_o[4][2] ),
    .B_N(_08090_),
    .Y(_08091_));
 sg13g2_a21oi_1 _27385_ (.A1(\cpu.gpio.r_src_o[4][2] ),
    .A2(_08089_),
    .Y(_08092_),
    .B1(_08091_));
 sg13g2_nand2b_1 _27386_ (.Y(_08093_),
    .B(net1064),
    .A_N(_04982_));
 sg13g2_nand3_1 _27387_ (.B(net1067),
    .C(_06256_),
    .A(_04982_),
    .Y(_08094_));
 sg13g2_o21ai_1 _27388_ (.B1(_08094_),
    .Y(_08095_),
    .A1(_06256_),
    .A2(_08093_));
 sg13g2_nand3_1 _27389_ (.B(\cpu.gpio.r_src_o[4][3] ),
    .C(_08095_),
    .A(_00098_),
    .Y(_08096_));
 sg13g2_o21ai_1 _27390_ (.B1(_08096_),
    .Y(net23),
    .A1(\cpu.gpio.r_src_o[4][3] ),
    .A2(_08092_));
 sg13g2_mux4_1 _27391_ (.S0(_05538_),
    .A0(net1090),
    .A1(net1091),
    .A2(net1066),
    .A3(net1065),
    .S1(_06260_),
    .X(_08097_));
 sg13g2_mux4_1 _27392_ (.S0(_05538_),
    .A0(\cpu.gpio.genblk1[5].srcs_o[0] ),
    .A1(net1068),
    .A2(net1088),
    .A3(net1089),
    .S1(_06260_),
    .X(_08098_));
 sg13g2_nor2b_1 _27393_ (.A(\cpu.gpio.r_src_o[5][2] ),
    .B_N(_08098_),
    .Y(_08099_));
 sg13g2_a21oi_1 _27394_ (.A1(\cpu.gpio.r_src_o[5][2] ),
    .A2(_08097_),
    .Y(_08100_),
    .B1(_08099_));
 sg13g2_nand2b_1 _27395_ (.Y(_08101_),
    .B(net1064),
    .A_N(_05538_));
 sg13g2_nand3_1 _27396_ (.B(net1067),
    .C(_06260_),
    .A(_05538_),
    .Y(_08102_));
 sg13g2_o21ai_1 _27397_ (.B1(_08102_),
    .Y(_08103_),
    .A1(_06260_),
    .A2(_08101_));
 sg13g2_nand3_1 _27398_ (.B(\cpu.gpio.r_src_o[5][3] ),
    .C(_08103_),
    .A(_00135_),
    .Y(_08104_));
 sg13g2_o21ai_1 _27399_ (.B1(_08104_),
    .Y(net24),
    .A1(\cpu.gpio.r_src_o[5][3] ),
    .A2(_08100_));
 sg13g2_mux4_1 _27400_ (.S0(_04977_),
    .A0(net1090),
    .A1(net1091),
    .A2(net1066),
    .A3(net1065),
    .S1(_07778_),
    .X(_08105_));
 sg13g2_mux4_1 _27401_ (.S0(_04977_),
    .A0(\cpu.gpio.genblk1[6].srcs_o[0] ),
    .A1(net1068),
    .A2(net1088),
    .A3(net1089),
    .S1(_07778_),
    .X(_08106_));
 sg13g2_nor2b_1 _27402_ (.A(\cpu.gpio.r_src_o[6][2] ),
    .B_N(_08106_),
    .Y(_08107_));
 sg13g2_a21oi_1 _27403_ (.A1(\cpu.gpio.r_src_o[6][2] ),
    .A2(_08105_),
    .Y(_08108_),
    .B1(_08107_));
 sg13g2_nand2b_1 _27404_ (.Y(_08109_),
    .B(net1064),
    .A_N(_04977_));
 sg13g2_nand3_1 _27405_ (.B(net1067),
    .C(_07778_),
    .A(_04977_),
    .Y(_08110_));
 sg13g2_o21ai_1 _27406_ (.B1(_08110_),
    .Y(_08111_),
    .A1(_07778_),
    .A2(_08109_));
 sg13g2_nand3_1 _27407_ (.B(\cpu.gpio.r_src_o[6][3] ),
    .C(_08111_),
    .A(_00097_),
    .Y(_08112_));
 sg13g2_o21ai_1 _27408_ (.B1(_08112_),
    .Y(net25),
    .A1(\cpu.gpio.r_src_o[6][3] ),
    .A2(_08108_));
 sg13g2_mux4_1 _27409_ (.S0(_05530_),
    .A0(_11962_),
    .A1(net1091),
    .A2(_07919_),
    .A3(net1065),
    .S1(_06263_),
    .X(_08113_));
 sg13g2_mux4_1 _27410_ (.S0(_05530_),
    .A0(\cpu.gpio.genblk1[7].srcs_o[0] ),
    .A1(_07260_),
    .A2(net1088),
    .A3(net1089),
    .S1(_06263_),
    .X(_08114_));
 sg13g2_nor2b_1 _27411_ (.A(\cpu.gpio.r_src_o[7][2] ),
    .B_N(_08114_),
    .Y(_08115_));
 sg13g2_a21oi_1 _27412_ (.A1(\cpu.gpio.r_src_o[7][2] ),
    .A2(_08113_),
    .Y(_08116_),
    .B1(_08115_));
 sg13g2_nand2b_1 _27413_ (.Y(_08117_),
    .B(_07937_),
    .A_N(_05530_));
 sg13g2_nand3_1 _27414_ (.B(_07871_),
    .C(_06263_),
    .A(_05530_),
    .Y(_08118_));
 sg13g2_o21ai_1 _27415_ (.B1(_08118_),
    .Y(_08119_),
    .A1(_06263_),
    .A2(_08117_));
 sg13g2_nand3_1 _27416_ (.B(\cpu.gpio.r_src_o[7][3] ),
    .C(_08119_),
    .A(_00134_),
    .Y(_08120_));
 sg13g2_o21ai_1 _27417_ (.B1(_08120_),
    .Y(net26),
    .A1(\cpu.gpio.r_src_o[7][3] ),
    .A2(_08116_));
 sg13g2_dfrbp_1 _27418_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1124),
    .D(_00294_),
    .Q_N(_14820_),
    .Q(\cpu.intr.r_swi ));
 sg13g2_dfrbp_1 _27419_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1125),
    .D(_00295_),
    .Q_N(_14819_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[5] ));
 sg13g2_dfrbp_1 _27420_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1126),
    .D(_00296_),
    .Q_N(_14818_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[4] ));
 sg13g2_dfrbp_1 _27421_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1127),
    .D(_00297_),
    .Q_N(_14817_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[3] ));
 sg13g2_dfrbp_1 _27422_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1128),
    .D(_00298_),
    .Q_N(_14816_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[2] ));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_1 _27424_ (.A(net6),
    .X(net4));
 sg13g2_buf_1 _27425_ (.A(net6),
    .X(net5));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1129),
    .D(_00299_),
    .Q_N(_14815_),
    .Q(\cpu.dcache.r_data[0][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1130),
    .D(_00300_),
    .Q_N(_00093_),
    .Q(\cpu.dcache.r_data[0][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1131),
    .D(_00301_),
    .Q_N(_00103_),
    .Q(\cpu.dcache.r_data[0][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1132),
    .D(_00302_),
    .Q_N(_00113_),
    .Q(\cpu.dcache.r_data[0][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1133),
    .D(_00303_),
    .Q_N(_00119_),
    .Q(\cpu.dcache.r_data[0][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1134),
    .D(_00304_),
    .Q_N(_00130_),
    .Q(\cpu.dcache.r_data[0][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1135),
    .D(_00305_),
    .Q_N(_00141_),
    .Q(\cpu.dcache.r_data[0][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1136),
    .D(_00306_),
    .Q_N(_14814_),
    .Q(\cpu.dcache.r_data[0][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1137),
    .D(_00307_),
    .Q_N(_00282_),
    .Q(\cpu.dcache.r_data[0][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1138),
    .D(_00308_),
    .Q_N(_00091_),
    .Q(\cpu.dcache.r_data[0][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][19]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1139),
    .D(_00309_),
    .Q_N(_00101_),
    .Q(\cpu.dcache.r_data[0][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1140),
    .D(_00310_),
    .Q_N(_14813_),
    .Q(\cpu.dcache.r_data[0][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][20]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1141),
    .D(_00311_),
    .Q_N(_00111_),
    .Q(\cpu.dcache.r_data[0][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][21]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1142),
    .D(_00312_),
    .Q_N(_00117_),
    .Q(\cpu.dcache.r_data[0][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][22]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1143),
    .D(_00313_),
    .Q_N(_00128_),
    .Q(\cpu.dcache.r_data[0][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][23]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1144),
    .D(_00314_),
    .Q_N(_00139_),
    .Q(\cpu.dcache.r_data[0][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][24]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1145),
    .D(_00315_),
    .Q_N(_00278_),
    .Q(\cpu.dcache.r_data[0][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][25]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1146),
    .D(_00316_),
    .Q_N(_00283_),
    .Q(\cpu.dcache.r_data[0][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][26]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1147),
    .D(_00317_),
    .Q_N(_00092_),
    .Q(\cpu.dcache.r_data[0][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][27]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1148),
    .D(_00318_),
    .Q_N(_00102_),
    .Q(\cpu.dcache.r_data[0][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][28]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1149),
    .D(_00319_),
    .Q_N(_00112_),
    .Q(\cpu.dcache.r_data[0][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][29]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1150),
    .D(_00320_),
    .Q_N(_00118_),
    .Q(\cpu.dcache.r_data[0][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1151),
    .D(_00321_),
    .Q_N(_14812_),
    .Q(\cpu.dcache.r_data[0][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][30]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1152),
    .D(_00322_),
    .Q_N(_00129_),
    .Q(\cpu.dcache.r_data[0][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][31]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1153),
    .D(_00323_),
    .Q_N(_00140_),
    .Q(\cpu.dcache.r_data[0][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1154),
    .D(_00324_),
    .Q_N(_14811_),
    .Q(\cpu.dcache.r_data[0][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1155),
    .D(_00325_),
    .Q_N(_00110_),
    .Q(\cpu.dcache.r_data[0][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1156),
    .D(_00326_),
    .Q_N(_00116_),
    .Q(\cpu.dcache.r_data[0][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1157),
    .D(_00327_),
    .Q_N(_00127_),
    .Q(\cpu.dcache.r_data[0][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1158),
    .D(_00328_),
    .Q_N(_00138_),
    .Q(\cpu.dcache.r_data[0][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1159),
    .D(_00329_),
    .Q_N(_00279_),
    .Q(\cpu.dcache.r_data[0][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1160),
    .D(_00330_),
    .Q_N(_00284_),
    .Q(\cpu.dcache.r_data[0][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1161),
    .D(_00331_),
    .Q_N(_14810_),
    .Q(\cpu.dcache.r_data[1][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1162),
    .D(_00332_),
    .Q_N(_14809_),
    .Q(\cpu.dcache.r_data[1][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1163),
    .D(_00333_),
    .Q_N(_14808_),
    .Q(\cpu.dcache.r_data[1][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1164),
    .D(_00334_),
    .Q_N(_14807_),
    .Q(\cpu.dcache.r_data[1][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1165),
    .D(_00335_),
    .Q_N(_14806_),
    .Q(\cpu.dcache.r_data[1][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1166),
    .D(_00336_),
    .Q_N(_14805_),
    .Q(\cpu.dcache.r_data[1][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1167),
    .D(_00337_),
    .Q_N(_14804_),
    .Q(\cpu.dcache.r_data[1][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1168),
    .D(_00338_),
    .Q_N(_14803_),
    .Q(\cpu.dcache.r_data[1][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1169),
    .D(_00339_),
    .Q_N(_14802_),
    .Q(\cpu.dcache.r_data[1][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1170),
    .D(_00340_),
    .Q_N(_14801_),
    .Q(\cpu.dcache.r_data[1][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][19]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1171),
    .D(_00341_),
    .Q_N(_14800_),
    .Q(\cpu.dcache.r_data[1][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1172),
    .D(_00342_),
    .Q_N(_14799_),
    .Q(\cpu.dcache.r_data[1][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][20]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1173),
    .D(_00343_),
    .Q_N(_14798_),
    .Q(\cpu.dcache.r_data[1][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][21]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1174),
    .D(_00344_),
    .Q_N(_14797_),
    .Q(\cpu.dcache.r_data[1][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][22]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1175),
    .D(_00345_),
    .Q_N(_14796_),
    .Q(\cpu.dcache.r_data[1][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][23]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1176),
    .D(_00346_),
    .Q_N(_14795_),
    .Q(\cpu.dcache.r_data[1][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][24]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1177),
    .D(_00347_),
    .Q_N(_14794_),
    .Q(\cpu.dcache.r_data[1][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][25]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1178),
    .D(_00348_),
    .Q_N(_14793_),
    .Q(\cpu.dcache.r_data[1][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][26]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1179),
    .D(_00349_),
    .Q_N(_14792_),
    .Q(\cpu.dcache.r_data[1][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][27]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1180),
    .D(_00350_),
    .Q_N(_14791_),
    .Q(\cpu.dcache.r_data[1][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][28]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1181),
    .D(_00351_),
    .Q_N(_14790_),
    .Q(\cpu.dcache.r_data[1][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][29]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1182),
    .D(_00352_),
    .Q_N(_14789_),
    .Q(\cpu.dcache.r_data[1][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1183),
    .D(_00353_),
    .Q_N(_14788_),
    .Q(\cpu.dcache.r_data[1][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][30]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1184),
    .D(_00354_),
    .Q_N(_14787_),
    .Q(\cpu.dcache.r_data[1][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][31]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1185),
    .D(_00355_),
    .Q_N(_14786_),
    .Q(\cpu.dcache.r_data[1][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1186),
    .D(_00356_),
    .Q_N(_14785_),
    .Q(\cpu.dcache.r_data[1][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1187),
    .D(_00357_),
    .Q_N(_14784_),
    .Q(\cpu.dcache.r_data[1][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1188),
    .D(_00358_),
    .Q_N(_14783_),
    .Q(\cpu.dcache.r_data[1][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1189),
    .D(_00359_),
    .Q_N(_14782_),
    .Q(\cpu.dcache.r_data[1][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1190),
    .D(_00360_),
    .Q_N(_14781_),
    .Q(\cpu.dcache.r_data[1][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1191),
    .D(_00361_),
    .Q_N(_14780_),
    .Q(\cpu.dcache.r_data[1][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1192),
    .D(_00362_),
    .Q_N(_14779_),
    .Q(\cpu.dcache.r_data[1][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1193),
    .D(_00363_),
    .Q_N(_14778_),
    .Q(\cpu.dcache.r_data[2][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1194),
    .D(_00364_),
    .Q_N(_14777_),
    .Q(\cpu.dcache.r_data[2][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1195),
    .D(_00365_),
    .Q_N(_14776_),
    .Q(\cpu.dcache.r_data[2][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1196),
    .D(_00366_),
    .Q_N(_14775_),
    .Q(\cpu.dcache.r_data[2][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1197),
    .D(_00367_),
    .Q_N(_14774_),
    .Q(\cpu.dcache.r_data[2][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1198),
    .D(_00368_),
    .Q_N(_14773_),
    .Q(\cpu.dcache.r_data[2][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1199),
    .D(_00369_),
    .Q_N(_14772_),
    .Q(\cpu.dcache.r_data[2][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1200),
    .D(_00370_),
    .Q_N(_14771_),
    .Q(\cpu.dcache.r_data[2][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1201),
    .D(_00371_),
    .Q_N(_14770_),
    .Q(\cpu.dcache.r_data[2][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1202),
    .D(_00372_),
    .Q_N(_14769_),
    .Q(\cpu.dcache.r_data[2][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][19]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1203),
    .D(_00373_),
    .Q_N(_14768_),
    .Q(\cpu.dcache.r_data[2][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1204),
    .D(_00374_),
    .Q_N(_14767_),
    .Q(\cpu.dcache.r_data[2][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][20]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1205),
    .D(_00375_),
    .Q_N(_14766_),
    .Q(\cpu.dcache.r_data[2][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][21]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1206),
    .D(_00376_),
    .Q_N(_14765_),
    .Q(\cpu.dcache.r_data[2][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][22]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1207),
    .D(_00377_),
    .Q_N(_14764_),
    .Q(\cpu.dcache.r_data[2][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][23]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1208),
    .D(_00378_),
    .Q_N(_14763_),
    .Q(\cpu.dcache.r_data[2][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][24]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1209),
    .D(_00379_),
    .Q_N(_14762_),
    .Q(\cpu.dcache.r_data[2][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][25]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1210),
    .D(_00380_),
    .Q_N(_14761_),
    .Q(\cpu.dcache.r_data[2][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][26]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1211),
    .D(_00381_),
    .Q_N(_14760_),
    .Q(\cpu.dcache.r_data[2][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][27]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1212),
    .D(_00382_),
    .Q_N(_14759_),
    .Q(\cpu.dcache.r_data[2][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][28]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1213),
    .D(_00383_),
    .Q_N(_14758_),
    .Q(\cpu.dcache.r_data[2][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][29]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1214),
    .D(_00384_),
    .Q_N(_14757_),
    .Q(\cpu.dcache.r_data[2][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1215),
    .D(_00385_),
    .Q_N(_14756_),
    .Q(\cpu.dcache.r_data[2][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][30]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1216),
    .D(_00386_),
    .Q_N(_14755_),
    .Q(\cpu.dcache.r_data[2][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][31]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1217),
    .D(_00387_),
    .Q_N(_14754_),
    .Q(\cpu.dcache.r_data[2][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1218),
    .D(_00388_),
    .Q_N(_14753_),
    .Q(\cpu.dcache.r_data[2][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1219),
    .D(_00389_),
    .Q_N(_14752_),
    .Q(\cpu.dcache.r_data[2][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1220),
    .D(_00390_),
    .Q_N(_14751_),
    .Q(\cpu.dcache.r_data[2][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1221),
    .D(_00391_),
    .Q_N(_14750_),
    .Q(\cpu.dcache.r_data[2][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1222),
    .D(_00392_),
    .Q_N(_14749_),
    .Q(\cpu.dcache.r_data[2][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1223),
    .D(_00393_),
    .Q_N(_14748_),
    .Q(\cpu.dcache.r_data[2][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1224),
    .D(_00394_),
    .Q_N(_14747_),
    .Q(\cpu.dcache.r_data[2][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1225),
    .D(_00395_),
    .Q_N(_14746_),
    .Q(\cpu.dcache.r_data[3][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1226),
    .D(_00396_),
    .Q_N(_14745_),
    .Q(\cpu.dcache.r_data[3][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1227),
    .D(_00397_),
    .Q_N(_14744_),
    .Q(\cpu.dcache.r_data[3][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1228),
    .D(_00398_),
    .Q_N(_14743_),
    .Q(\cpu.dcache.r_data[3][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1229),
    .D(_00399_),
    .Q_N(_14742_),
    .Q(\cpu.dcache.r_data[3][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1230),
    .D(_00400_),
    .Q_N(_14741_),
    .Q(\cpu.dcache.r_data[3][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1231),
    .D(_00401_),
    .Q_N(_14740_),
    .Q(\cpu.dcache.r_data[3][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1232),
    .D(_00402_),
    .Q_N(_14739_),
    .Q(\cpu.dcache.r_data[3][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1233),
    .D(_00403_),
    .Q_N(_14738_),
    .Q(\cpu.dcache.r_data[3][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1234),
    .D(_00404_),
    .Q_N(_14737_),
    .Q(\cpu.dcache.r_data[3][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][19]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1235),
    .D(_00405_),
    .Q_N(_14736_),
    .Q(\cpu.dcache.r_data[3][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1236),
    .D(_00406_),
    .Q_N(_14735_),
    .Q(\cpu.dcache.r_data[3][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][20]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1237),
    .D(_00407_),
    .Q_N(_14734_),
    .Q(\cpu.dcache.r_data[3][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][21]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1238),
    .D(_00408_),
    .Q_N(_14733_),
    .Q(\cpu.dcache.r_data[3][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][22]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1239),
    .D(_00409_),
    .Q_N(_14732_),
    .Q(\cpu.dcache.r_data[3][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][23]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1240),
    .D(_00410_),
    .Q_N(_14731_),
    .Q(\cpu.dcache.r_data[3][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][24]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1241),
    .D(_00411_),
    .Q_N(_14730_),
    .Q(\cpu.dcache.r_data[3][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][25]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1242),
    .D(_00412_),
    .Q_N(_14729_),
    .Q(\cpu.dcache.r_data[3][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][26]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1243),
    .D(_00413_),
    .Q_N(_14728_),
    .Q(\cpu.dcache.r_data[3][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][27]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1244),
    .D(_00414_),
    .Q_N(_14727_),
    .Q(\cpu.dcache.r_data[3][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][28]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1245),
    .D(_00415_),
    .Q_N(_14726_),
    .Q(\cpu.dcache.r_data[3][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][29]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1246),
    .D(_00416_),
    .Q_N(_14725_),
    .Q(\cpu.dcache.r_data[3][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1247),
    .D(_00417_),
    .Q_N(_14724_),
    .Q(\cpu.dcache.r_data[3][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][30]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1248),
    .D(_00418_),
    .Q_N(_14723_),
    .Q(\cpu.dcache.r_data[3][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][31]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1249),
    .D(_00419_),
    .Q_N(_14722_),
    .Q(\cpu.dcache.r_data[3][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1250),
    .D(_00420_),
    .Q_N(_14721_),
    .Q(\cpu.dcache.r_data[3][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1251),
    .D(_00421_),
    .Q_N(_14720_),
    .Q(\cpu.dcache.r_data[3][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1252),
    .D(_00422_),
    .Q_N(_14719_),
    .Q(\cpu.dcache.r_data[3][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1253),
    .D(_00423_),
    .Q_N(_14718_),
    .Q(\cpu.dcache.r_data[3][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1254),
    .D(_00424_),
    .Q_N(_14717_),
    .Q(\cpu.dcache.r_data[3][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1255),
    .D(_00425_),
    .Q_N(_14716_),
    .Q(\cpu.dcache.r_data[3][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1256),
    .D(_00426_),
    .Q_N(_14715_),
    .Q(\cpu.dcache.r_data[3][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1257),
    .D(_00427_),
    .Q_N(_14714_),
    .Q(\cpu.dcache.r_data[4][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1258),
    .D(_00428_),
    .Q_N(_14713_),
    .Q(\cpu.dcache.r_data[4][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1259),
    .D(_00429_),
    .Q_N(_14712_),
    .Q(\cpu.dcache.r_data[4][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1260),
    .D(_00430_),
    .Q_N(_14711_),
    .Q(\cpu.dcache.r_data[4][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1261),
    .D(_00431_),
    .Q_N(_14710_),
    .Q(\cpu.dcache.r_data[4][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1262),
    .D(_00432_),
    .Q_N(_14709_),
    .Q(\cpu.dcache.r_data[4][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1263),
    .D(_00433_),
    .Q_N(_14708_),
    .Q(\cpu.dcache.r_data[4][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1264),
    .D(_00434_),
    .Q_N(_14707_),
    .Q(\cpu.dcache.r_data[4][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1265),
    .D(_00435_),
    .Q_N(_14706_),
    .Q(\cpu.dcache.r_data[4][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1266),
    .D(_00436_),
    .Q_N(_14705_),
    .Q(\cpu.dcache.r_data[4][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][19]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1267),
    .D(_00437_),
    .Q_N(_14704_),
    .Q(\cpu.dcache.r_data[4][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1268),
    .D(_00438_),
    .Q_N(_14703_),
    .Q(\cpu.dcache.r_data[4][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][20]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1269),
    .D(_00439_),
    .Q_N(_14702_),
    .Q(\cpu.dcache.r_data[4][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][21]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1270),
    .D(_00440_),
    .Q_N(_14701_),
    .Q(\cpu.dcache.r_data[4][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][22]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1271),
    .D(_00441_),
    .Q_N(_14700_),
    .Q(\cpu.dcache.r_data[4][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][23]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1272),
    .D(_00442_),
    .Q_N(_14699_),
    .Q(\cpu.dcache.r_data[4][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][24]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1273),
    .D(_00443_),
    .Q_N(_14698_),
    .Q(\cpu.dcache.r_data[4][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][25]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1274),
    .D(_00444_),
    .Q_N(_14697_),
    .Q(\cpu.dcache.r_data[4][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][26]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1275),
    .D(_00445_),
    .Q_N(_14696_),
    .Q(\cpu.dcache.r_data[4][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][27]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1276),
    .D(_00446_),
    .Q_N(_14695_),
    .Q(\cpu.dcache.r_data[4][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][28]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1277),
    .D(_00447_),
    .Q_N(_14694_),
    .Q(\cpu.dcache.r_data[4][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][29]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1278),
    .D(_00448_),
    .Q_N(_14693_),
    .Q(\cpu.dcache.r_data[4][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1279),
    .D(_00449_),
    .Q_N(_14692_),
    .Q(\cpu.dcache.r_data[4][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][30]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1280),
    .D(_00450_),
    .Q_N(_14691_),
    .Q(\cpu.dcache.r_data[4][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][31]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1281),
    .D(_00451_),
    .Q_N(_14690_),
    .Q(\cpu.dcache.r_data[4][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1282),
    .D(_00452_),
    .Q_N(_14689_),
    .Q(\cpu.dcache.r_data[4][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1283),
    .D(_00453_),
    .Q_N(_14688_),
    .Q(\cpu.dcache.r_data[4][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1284),
    .D(_00454_),
    .Q_N(_14687_),
    .Q(\cpu.dcache.r_data[4][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1285),
    .D(_00455_),
    .Q_N(_14686_),
    .Q(\cpu.dcache.r_data[4][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1286),
    .D(_00456_),
    .Q_N(_14685_),
    .Q(\cpu.dcache.r_data[4][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1287),
    .D(_00457_),
    .Q_N(_14684_),
    .Q(\cpu.dcache.r_data[4][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1288),
    .D(_00458_),
    .Q_N(_14683_),
    .Q(\cpu.dcache.r_data[4][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1289),
    .D(_00459_),
    .Q_N(_14682_),
    .Q(\cpu.dcache.r_data[5][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1290),
    .D(_00460_),
    .Q_N(_14681_),
    .Q(\cpu.dcache.r_data[5][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1291),
    .D(_00461_),
    .Q_N(_14680_),
    .Q(\cpu.dcache.r_data[5][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1292),
    .D(_00462_),
    .Q_N(_14679_),
    .Q(\cpu.dcache.r_data[5][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1293),
    .D(_00463_),
    .Q_N(_14678_),
    .Q(\cpu.dcache.r_data[5][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1294),
    .D(_00464_),
    .Q_N(_14677_),
    .Q(\cpu.dcache.r_data[5][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1295),
    .D(_00465_),
    .Q_N(_14676_),
    .Q(\cpu.dcache.r_data[5][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1296),
    .D(_00466_),
    .Q_N(_14675_),
    .Q(\cpu.dcache.r_data[5][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1297),
    .D(_00467_),
    .Q_N(_14674_),
    .Q(\cpu.dcache.r_data[5][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1298),
    .D(_00468_),
    .Q_N(_14673_),
    .Q(\cpu.dcache.r_data[5][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][19]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1299),
    .D(_00469_),
    .Q_N(_14672_),
    .Q(\cpu.dcache.r_data[5][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1300),
    .D(_00470_),
    .Q_N(_14671_),
    .Q(\cpu.dcache.r_data[5][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][20]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1301),
    .D(_00471_),
    .Q_N(_14670_),
    .Q(\cpu.dcache.r_data[5][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][21]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1302),
    .D(_00472_),
    .Q_N(_14669_),
    .Q(\cpu.dcache.r_data[5][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][22]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1303),
    .D(_00473_),
    .Q_N(_14668_),
    .Q(\cpu.dcache.r_data[5][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][23]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1304),
    .D(_00474_),
    .Q_N(_14667_),
    .Q(\cpu.dcache.r_data[5][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][24]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1305),
    .D(_00475_),
    .Q_N(_14666_),
    .Q(\cpu.dcache.r_data[5][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][25]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1306),
    .D(_00476_),
    .Q_N(_14665_),
    .Q(\cpu.dcache.r_data[5][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][26]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1307),
    .D(_00477_),
    .Q_N(_14664_),
    .Q(\cpu.dcache.r_data[5][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][27]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1308),
    .D(_00478_),
    .Q_N(_14663_),
    .Q(\cpu.dcache.r_data[5][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][28]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1309),
    .D(_00479_),
    .Q_N(_14662_),
    .Q(\cpu.dcache.r_data[5][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][29]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1310),
    .D(_00480_),
    .Q_N(_14661_),
    .Q(\cpu.dcache.r_data[5][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1311),
    .D(_00481_),
    .Q_N(_14660_),
    .Q(\cpu.dcache.r_data[5][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][30]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1312),
    .D(_00482_),
    .Q_N(_14659_),
    .Q(\cpu.dcache.r_data[5][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][31]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1313),
    .D(_00483_),
    .Q_N(_14658_),
    .Q(\cpu.dcache.r_data[5][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1314),
    .D(_00484_),
    .Q_N(_14657_),
    .Q(\cpu.dcache.r_data[5][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1315),
    .D(_00485_),
    .Q_N(_14656_),
    .Q(\cpu.dcache.r_data[5][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1316),
    .D(_00486_),
    .Q_N(_14655_),
    .Q(\cpu.dcache.r_data[5][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1317),
    .D(_00487_),
    .Q_N(_14654_),
    .Q(\cpu.dcache.r_data[5][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1318),
    .D(_00488_),
    .Q_N(_14653_),
    .Q(\cpu.dcache.r_data[5][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1319),
    .D(_00489_),
    .Q_N(_14652_),
    .Q(\cpu.dcache.r_data[5][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1320),
    .D(_00490_),
    .Q_N(_14651_),
    .Q(\cpu.dcache.r_data[5][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1321),
    .D(_00491_),
    .Q_N(_14650_),
    .Q(\cpu.dcache.r_data[6][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1322),
    .D(_00492_),
    .Q_N(_14649_),
    .Q(\cpu.dcache.r_data[6][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1323),
    .D(_00493_),
    .Q_N(_14648_),
    .Q(\cpu.dcache.r_data[6][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1324),
    .D(_00494_),
    .Q_N(_14647_),
    .Q(\cpu.dcache.r_data[6][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1325),
    .D(_00495_),
    .Q_N(_14646_),
    .Q(\cpu.dcache.r_data[6][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1326),
    .D(_00496_),
    .Q_N(_14645_),
    .Q(\cpu.dcache.r_data[6][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1327),
    .D(_00497_),
    .Q_N(_14644_),
    .Q(\cpu.dcache.r_data[6][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1328),
    .D(_00498_),
    .Q_N(_14643_),
    .Q(\cpu.dcache.r_data[6][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1329),
    .D(_00499_),
    .Q_N(_14642_),
    .Q(\cpu.dcache.r_data[6][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1330),
    .D(_00500_),
    .Q_N(_14641_),
    .Q(\cpu.dcache.r_data[6][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][19]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1331),
    .D(_00501_),
    .Q_N(_14640_),
    .Q(\cpu.dcache.r_data[6][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1332),
    .D(_00502_),
    .Q_N(_14639_),
    .Q(\cpu.dcache.r_data[6][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][20]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1333),
    .D(_00503_),
    .Q_N(_14638_),
    .Q(\cpu.dcache.r_data[6][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][21]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1334),
    .D(_00504_),
    .Q_N(_14637_),
    .Q(\cpu.dcache.r_data[6][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][22]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1335),
    .D(_00505_),
    .Q_N(_14636_),
    .Q(\cpu.dcache.r_data[6][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][23]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1336),
    .D(_00506_),
    .Q_N(_14635_),
    .Q(\cpu.dcache.r_data[6][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][24]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1337),
    .D(_00507_),
    .Q_N(_14634_),
    .Q(\cpu.dcache.r_data[6][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][25]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1338),
    .D(_00508_),
    .Q_N(_14633_),
    .Q(\cpu.dcache.r_data[6][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][26]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1339),
    .D(_00509_),
    .Q_N(_14632_),
    .Q(\cpu.dcache.r_data[6][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][27]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1340),
    .D(_00510_),
    .Q_N(_14631_),
    .Q(\cpu.dcache.r_data[6][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][28]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1341),
    .D(_00511_),
    .Q_N(_14630_),
    .Q(\cpu.dcache.r_data[6][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][29]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1342),
    .D(_00512_),
    .Q_N(_14629_),
    .Q(\cpu.dcache.r_data[6][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1343),
    .D(_00513_),
    .Q_N(_14628_),
    .Q(\cpu.dcache.r_data[6][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][30]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1344),
    .D(_00514_),
    .Q_N(_14627_),
    .Q(\cpu.dcache.r_data[6][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][31]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1345),
    .D(_00515_),
    .Q_N(_14626_),
    .Q(\cpu.dcache.r_data[6][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1346),
    .D(_00516_),
    .Q_N(_14625_),
    .Q(\cpu.dcache.r_data[6][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1347),
    .D(_00517_),
    .Q_N(_14624_),
    .Q(\cpu.dcache.r_data[6][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1348),
    .D(_00518_),
    .Q_N(_14623_),
    .Q(\cpu.dcache.r_data[6][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1349),
    .D(_00519_),
    .Q_N(_14622_),
    .Q(\cpu.dcache.r_data[6][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1350),
    .D(_00520_),
    .Q_N(_14621_),
    .Q(\cpu.dcache.r_data[6][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1351),
    .D(_00521_),
    .Q_N(_14620_),
    .Q(\cpu.dcache.r_data[6][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1352),
    .D(_00522_),
    .Q_N(_14619_),
    .Q(\cpu.dcache.r_data[6][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1353),
    .D(_00523_),
    .Q_N(_14618_),
    .Q(\cpu.dcache.r_data[7][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1354),
    .D(_00524_),
    .Q_N(_14617_),
    .Q(\cpu.dcache.r_data[7][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1355),
    .D(_00525_),
    .Q_N(_14616_),
    .Q(\cpu.dcache.r_data[7][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1356),
    .D(_00526_),
    .Q_N(_14615_),
    .Q(\cpu.dcache.r_data[7][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1357),
    .D(_00527_),
    .Q_N(_14614_),
    .Q(\cpu.dcache.r_data[7][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1358),
    .D(_00528_),
    .Q_N(_14613_),
    .Q(\cpu.dcache.r_data[7][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1359),
    .D(_00529_),
    .Q_N(_14612_),
    .Q(\cpu.dcache.r_data[7][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1360),
    .D(_00530_),
    .Q_N(_14611_),
    .Q(\cpu.dcache.r_data[7][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1361),
    .D(_00531_),
    .Q_N(_14610_),
    .Q(\cpu.dcache.r_data[7][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1362),
    .D(_00532_),
    .Q_N(_14609_),
    .Q(\cpu.dcache.r_data[7][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][19]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1363),
    .D(_00533_),
    .Q_N(_14608_),
    .Q(\cpu.dcache.r_data[7][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1364),
    .D(_00534_),
    .Q_N(_14607_),
    .Q(\cpu.dcache.r_data[7][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][20]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1365),
    .D(_00535_),
    .Q_N(_14606_),
    .Q(\cpu.dcache.r_data[7][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][21]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1366),
    .D(_00536_),
    .Q_N(_14605_),
    .Q(\cpu.dcache.r_data[7][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][22]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1367),
    .D(_00537_),
    .Q_N(_14604_),
    .Q(\cpu.dcache.r_data[7][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][23]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1368),
    .D(_00538_),
    .Q_N(_14603_),
    .Q(\cpu.dcache.r_data[7][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][24]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1369),
    .D(_00539_),
    .Q_N(_14602_),
    .Q(\cpu.dcache.r_data[7][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][25]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1370),
    .D(_00540_),
    .Q_N(_14601_),
    .Q(\cpu.dcache.r_data[7][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][26]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1371),
    .D(_00541_),
    .Q_N(_14600_),
    .Q(\cpu.dcache.r_data[7][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][27]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1372),
    .D(_00542_),
    .Q_N(_14599_),
    .Q(\cpu.dcache.r_data[7][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][28]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1373),
    .D(_00543_),
    .Q_N(_14598_),
    .Q(\cpu.dcache.r_data[7][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][29]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1374),
    .D(_00544_),
    .Q_N(_14597_),
    .Q(\cpu.dcache.r_data[7][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1375),
    .D(_00545_),
    .Q_N(_14596_),
    .Q(\cpu.dcache.r_data[7][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][30]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1376),
    .D(_00546_),
    .Q_N(_14595_),
    .Q(\cpu.dcache.r_data[7][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][31]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1377),
    .D(_00547_),
    .Q_N(_14594_),
    .Q(\cpu.dcache.r_data[7][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1378),
    .D(_00548_),
    .Q_N(_14593_),
    .Q(\cpu.dcache.r_data[7][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1379),
    .D(_00549_),
    .Q_N(_14592_),
    .Q(\cpu.dcache.r_data[7][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1380),
    .D(_00550_),
    .Q_N(_14591_),
    .Q(\cpu.dcache.r_data[7][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1381),
    .D(_00551_),
    .Q_N(_14590_),
    .Q(\cpu.dcache.r_data[7][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1382),
    .D(_00552_),
    .Q_N(_14589_),
    .Q(\cpu.dcache.r_data[7][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1383),
    .D(_00553_),
    .Q_N(_14588_),
    .Q(\cpu.dcache.r_data[7][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1384),
    .D(_00554_),
    .Q_N(_14587_),
    .Q(\cpu.dcache.r_data[7][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[0]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1385),
    .D(_00555_),
    .Q_N(_14586_),
    .Q(\cpu.dcache.r_dirty[0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[1]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1386),
    .D(_00556_),
    .Q_N(_14585_),
    .Q(\cpu.dcache.r_dirty[1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[2]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1387),
    .D(_00557_),
    .Q_N(_14584_),
    .Q(\cpu.dcache.r_dirty[2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[3]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1388),
    .D(_00558_),
    .Q_N(_14583_),
    .Q(\cpu.dcache.r_dirty[3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[4]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1389),
    .D(_00559_),
    .Q_N(_14582_),
    .Q(\cpu.dcache.r_dirty[4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[5]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1390),
    .D(_00560_),
    .Q_N(_14581_),
    .Q(\cpu.dcache.r_dirty[5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[6]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1391),
    .D(_00561_),
    .Q_N(_14580_),
    .Q(\cpu.dcache.r_dirty[6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[7]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1392),
    .D(_00562_),
    .Q_N(_14579_),
    .Q(\cpu.dcache.r_dirty[7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_offset[0]$_SDFF_PN0_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1393),
    .D(_00563_),
    .Q_N(_00292_),
    .Q(\cpu.dcache.r_offset[0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_offset[1]$_SDFF_PN0_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1394),
    .D(_00564_),
    .Q_N(_14578_),
    .Q(\cpu.dcache.r_offset[1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_offset[2]$_SDFF_PN0_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1395),
    .D(_00565_),
    .Q_N(_00255_),
    .Q(\cpu.dcache.r_offset[2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1396),
    .D(_00566_),
    .Q_N(_00208_),
    .Q(\cpu.dcache.r_tag[0][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1397),
    .D(_00567_),
    .Q_N(_00224_),
    .Q(\cpu.dcache.r_tag[0][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1398),
    .D(_00568_),
    .Q_N(_00225_),
    .Q(\cpu.dcache.r_tag[0][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1399),
    .D(_00569_),
    .Q_N(_00226_),
    .Q(\cpu.dcache.r_tag[0][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1400),
    .D(_00570_),
    .Q_N(_00227_),
    .Q(\cpu.dcache.r_tag[0][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1401),
    .D(_00571_),
    .Q_N(_00228_),
    .Q(\cpu.dcache.r_tag[0][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1402),
    .D(_00572_),
    .Q_N(_14577_),
    .Q(\cpu.dcache.r_tag[0][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1403),
    .D(_00573_),
    .Q_N(_14576_),
    .Q(\cpu.dcache.r_tag[0][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1404),
    .D(_00574_),
    .Q_N(_14575_),
    .Q(\cpu.dcache.r_tag[0][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1405),
    .D(_00575_),
    .Q_N(_00229_),
    .Q(\cpu.dcache.r_tag[0][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1406),
    .D(_00576_),
    .Q_N(_00210_),
    .Q(\cpu.dcache.r_tag[0][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1407),
    .D(_00577_),
    .Q_N(_00212_),
    .Q(\cpu.dcache.r_tag[0][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1408),
    .D(_00578_),
    .Q_N(_00214_),
    .Q(\cpu.dcache.r_tag[0][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1409),
    .D(_00579_),
    .Q_N(_00216_),
    .Q(\cpu.dcache.r_tag[0][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1410),
    .D(_00580_),
    .Q_N(_00218_),
    .Q(\cpu.dcache.r_tag[0][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1411),
    .D(_00581_),
    .Q_N(_00220_),
    .Q(\cpu.dcache.r_tag[0][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1412),
    .D(_00582_),
    .Q_N(_00221_),
    .Q(\cpu.dcache.r_tag[0][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1413),
    .D(_00583_),
    .Q_N(_00222_),
    .Q(\cpu.dcache.r_tag[0][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1414),
    .D(_00584_),
    .Q_N(_00223_),
    .Q(\cpu.dcache.r_tag[0][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1415),
    .D(_00585_),
    .Q_N(_14574_),
    .Q(\cpu.dcache.r_tag[1][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1416),
    .D(_00586_),
    .Q_N(_14573_),
    .Q(\cpu.dcache.r_tag[1][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1417),
    .D(_00587_),
    .Q_N(_14572_),
    .Q(\cpu.dcache.r_tag[1][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1418),
    .D(_00588_),
    .Q_N(_14571_),
    .Q(\cpu.dcache.r_tag[1][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1419),
    .D(_00589_),
    .Q_N(_14570_),
    .Q(\cpu.dcache.r_tag[1][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1420),
    .D(_00590_),
    .Q_N(_14569_),
    .Q(\cpu.dcache.r_tag[1][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1421),
    .D(_00591_),
    .Q_N(_14568_),
    .Q(\cpu.dcache.r_tag[1][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1422),
    .D(_00592_),
    .Q_N(_14567_),
    .Q(\cpu.dcache.r_tag[1][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1423),
    .D(_00593_),
    .Q_N(_14566_),
    .Q(\cpu.dcache.r_tag[1][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1424),
    .D(_00594_),
    .Q_N(_14565_),
    .Q(\cpu.dcache.r_tag[1][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1425),
    .D(_00595_),
    .Q_N(_14564_),
    .Q(\cpu.dcache.r_tag[1][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1426),
    .D(_00596_),
    .Q_N(_14563_),
    .Q(\cpu.dcache.r_tag[1][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1427),
    .D(_00597_),
    .Q_N(_14562_),
    .Q(\cpu.dcache.r_tag[1][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1428),
    .D(_00598_),
    .Q_N(_14561_),
    .Q(\cpu.dcache.r_tag[1][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1429),
    .D(_00599_),
    .Q_N(_14560_),
    .Q(\cpu.dcache.r_tag[1][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1430),
    .D(_00600_),
    .Q_N(_14559_),
    .Q(\cpu.dcache.r_tag[1][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1431),
    .D(_00601_),
    .Q_N(_14558_),
    .Q(\cpu.dcache.r_tag[1][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1432),
    .D(_00602_),
    .Q_N(_14557_),
    .Q(\cpu.dcache.r_tag[1][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1433),
    .D(_00603_),
    .Q_N(_14556_),
    .Q(\cpu.dcache.r_tag[1][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1434),
    .D(_00604_),
    .Q_N(_14555_),
    .Q(\cpu.dcache.r_tag[2][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1435),
    .D(_00605_),
    .Q_N(_14554_),
    .Q(\cpu.dcache.r_tag[2][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1436),
    .D(_00606_),
    .Q_N(_14553_),
    .Q(\cpu.dcache.r_tag[2][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1437),
    .D(_00607_),
    .Q_N(_14552_),
    .Q(\cpu.dcache.r_tag[2][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1438),
    .D(_00608_),
    .Q_N(_14551_),
    .Q(\cpu.dcache.r_tag[2][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1439),
    .D(_00609_),
    .Q_N(_14550_),
    .Q(\cpu.dcache.r_tag[2][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1440),
    .D(_00610_),
    .Q_N(_14549_),
    .Q(\cpu.dcache.r_tag[2][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1441),
    .D(_00611_),
    .Q_N(_14548_),
    .Q(\cpu.dcache.r_tag[2][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1442),
    .D(_00612_),
    .Q_N(_14547_),
    .Q(\cpu.dcache.r_tag[2][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1443),
    .D(_00613_),
    .Q_N(_14546_),
    .Q(\cpu.dcache.r_tag[2][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1444),
    .D(_00614_),
    .Q_N(_14545_),
    .Q(\cpu.dcache.r_tag[2][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1445),
    .D(_00615_),
    .Q_N(_14544_),
    .Q(\cpu.dcache.r_tag[2][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1446),
    .D(_00616_),
    .Q_N(_14543_),
    .Q(\cpu.dcache.r_tag[2][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1447),
    .D(_00617_),
    .Q_N(_14542_),
    .Q(\cpu.dcache.r_tag[2][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1448),
    .D(_00618_),
    .Q_N(_14541_),
    .Q(\cpu.dcache.r_tag[2][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1449),
    .D(_00619_),
    .Q_N(_14540_),
    .Q(\cpu.dcache.r_tag[2][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1450),
    .D(_00620_),
    .Q_N(_14539_),
    .Q(\cpu.dcache.r_tag[2][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1451),
    .D(_00621_),
    .Q_N(_14538_),
    .Q(\cpu.dcache.r_tag[2][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1452),
    .D(_00622_),
    .Q_N(_14537_),
    .Q(\cpu.dcache.r_tag[2][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1453),
    .D(_00623_),
    .Q_N(_14536_),
    .Q(\cpu.dcache.r_tag[3][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1454),
    .D(_00624_),
    .Q_N(_14535_),
    .Q(\cpu.dcache.r_tag[3][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1455),
    .D(_00625_),
    .Q_N(_14534_),
    .Q(\cpu.dcache.r_tag[3][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1456),
    .D(_00626_),
    .Q_N(_14533_),
    .Q(\cpu.dcache.r_tag[3][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1457),
    .D(_00627_),
    .Q_N(_14532_),
    .Q(\cpu.dcache.r_tag[3][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1458),
    .D(_00628_),
    .Q_N(_14531_),
    .Q(\cpu.dcache.r_tag[3][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1459),
    .D(_00629_),
    .Q_N(_14530_),
    .Q(\cpu.dcache.r_tag[3][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1460),
    .D(_00630_),
    .Q_N(_14529_),
    .Q(\cpu.dcache.r_tag[3][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1461),
    .D(_00631_),
    .Q_N(_14528_),
    .Q(\cpu.dcache.r_tag[3][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1462),
    .D(_00632_),
    .Q_N(_14527_),
    .Q(\cpu.dcache.r_tag[3][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1463),
    .D(_00633_),
    .Q_N(_14526_),
    .Q(\cpu.dcache.r_tag[3][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1464),
    .D(_00634_),
    .Q_N(_14525_),
    .Q(\cpu.dcache.r_tag[3][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1465),
    .D(_00635_),
    .Q_N(_14524_),
    .Q(\cpu.dcache.r_tag[3][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1466),
    .D(_00636_),
    .Q_N(_14523_),
    .Q(\cpu.dcache.r_tag[3][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1467),
    .D(_00637_),
    .Q_N(_14522_),
    .Q(\cpu.dcache.r_tag[3][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1468),
    .D(_00638_),
    .Q_N(_14521_),
    .Q(\cpu.dcache.r_tag[3][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1469),
    .D(_00639_),
    .Q_N(_14520_),
    .Q(\cpu.dcache.r_tag[3][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1470),
    .D(_00640_),
    .Q_N(_14519_),
    .Q(\cpu.dcache.r_tag[3][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1471),
    .D(_00641_),
    .Q_N(_14518_),
    .Q(\cpu.dcache.r_tag[3][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1472),
    .D(_00642_),
    .Q_N(_14517_),
    .Q(\cpu.dcache.r_tag[4][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1473),
    .D(_00643_),
    .Q_N(_14516_),
    .Q(\cpu.dcache.r_tag[4][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1474),
    .D(_00644_),
    .Q_N(_14515_),
    .Q(\cpu.dcache.r_tag[4][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1475),
    .D(_00645_),
    .Q_N(_14514_),
    .Q(\cpu.dcache.r_tag[4][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1476),
    .D(_00646_),
    .Q_N(_14513_),
    .Q(\cpu.dcache.r_tag[4][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1477),
    .D(_00647_),
    .Q_N(_14512_),
    .Q(\cpu.dcache.r_tag[4][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1478),
    .D(_00648_),
    .Q_N(_14511_),
    .Q(\cpu.dcache.r_tag[4][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1479),
    .D(_00649_),
    .Q_N(_14510_),
    .Q(\cpu.dcache.r_tag[4][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1480),
    .D(_00650_),
    .Q_N(_14509_),
    .Q(\cpu.dcache.r_tag[4][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1481),
    .D(_00651_),
    .Q_N(_14508_),
    .Q(\cpu.dcache.r_tag[4][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1482),
    .D(_00652_),
    .Q_N(_14507_),
    .Q(\cpu.dcache.r_tag[4][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1483),
    .D(_00653_),
    .Q_N(_14506_),
    .Q(\cpu.dcache.r_tag[4][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1484),
    .D(_00654_),
    .Q_N(_14505_),
    .Q(\cpu.dcache.r_tag[4][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1485),
    .D(_00655_),
    .Q_N(_14504_),
    .Q(\cpu.dcache.r_tag[4][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1486),
    .D(_00656_),
    .Q_N(_14503_),
    .Q(\cpu.dcache.r_tag[4][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1487),
    .D(_00657_),
    .Q_N(_14502_),
    .Q(\cpu.dcache.r_tag[4][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1488),
    .D(_00658_),
    .Q_N(_14501_),
    .Q(\cpu.dcache.r_tag[4][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1489),
    .D(_00659_),
    .Q_N(_14500_),
    .Q(\cpu.dcache.r_tag[4][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1490),
    .D(_00660_),
    .Q_N(_14499_),
    .Q(\cpu.dcache.r_tag[4][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1491),
    .D(_00661_),
    .Q_N(_14498_),
    .Q(\cpu.dcache.r_tag[5][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1492),
    .D(_00662_),
    .Q_N(_14497_),
    .Q(\cpu.dcache.r_tag[5][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1493),
    .D(_00663_),
    .Q_N(_14496_),
    .Q(\cpu.dcache.r_tag[5][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1494),
    .D(_00664_),
    .Q_N(_14495_),
    .Q(\cpu.dcache.r_tag[5][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1495),
    .D(_00665_),
    .Q_N(_14494_),
    .Q(\cpu.dcache.r_tag[5][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1496),
    .D(_00666_),
    .Q_N(_14493_),
    .Q(\cpu.dcache.r_tag[5][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1497),
    .D(_00667_),
    .Q_N(_14492_),
    .Q(\cpu.dcache.r_tag[5][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1498),
    .D(_00668_),
    .Q_N(_14491_),
    .Q(\cpu.dcache.r_tag[5][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1499),
    .D(_00669_),
    .Q_N(_14490_),
    .Q(\cpu.dcache.r_tag[5][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1500),
    .D(_00670_),
    .Q_N(_14489_),
    .Q(\cpu.dcache.r_tag[5][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1501),
    .D(_00671_),
    .Q_N(_14488_),
    .Q(\cpu.dcache.r_tag[5][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1502),
    .D(_00672_),
    .Q_N(_14487_),
    .Q(\cpu.dcache.r_tag[5][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1503),
    .D(_00673_),
    .Q_N(_14486_),
    .Q(\cpu.dcache.r_tag[5][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1504),
    .D(_00674_),
    .Q_N(_14485_),
    .Q(\cpu.dcache.r_tag[5][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1505),
    .D(_00675_),
    .Q_N(_14484_),
    .Q(\cpu.dcache.r_tag[5][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1506),
    .D(_00676_),
    .Q_N(_14483_),
    .Q(\cpu.dcache.r_tag[5][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1507),
    .D(_00677_),
    .Q_N(_14482_),
    .Q(\cpu.dcache.r_tag[5][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1508),
    .D(_00678_),
    .Q_N(_14481_),
    .Q(\cpu.dcache.r_tag[5][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1509),
    .D(_00679_),
    .Q_N(_14480_),
    .Q(\cpu.dcache.r_tag[5][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1510),
    .D(_00680_),
    .Q_N(_14479_),
    .Q(\cpu.dcache.r_tag[6][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1511),
    .D(_00681_),
    .Q_N(_14478_),
    .Q(\cpu.dcache.r_tag[6][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1512),
    .D(_00682_),
    .Q_N(_14477_),
    .Q(\cpu.dcache.r_tag[6][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1513),
    .D(_00683_),
    .Q_N(_14476_),
    .Q(\cpu.dcache.r_tag[6][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1514),
    .D(_00684_),
    .Q_N(_14475_),
    .Q(\cpu.dcache.r_tag[6][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1515),
    .D(_00685_),
    .Q_N(_14474_),
    .Q(\cpu.dcache.r_tag[6][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1516),
    .D(_00686_),
    .Q_N(_14473_),
    .Q(\cpu.dcache.r_tag[6][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1517),
    .D(_00687_),
    .Q_N(_14472_),
    .Q(\cpu.dcache.r_tag[6][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1518),
    .D(_00688_),
    .Q_N(_14471_),
    .Q(\cpu.dcache.r_tag[6][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1519),
    .D(_00689_),
    .Q_N(_14470_),
    .Q(\cpu.dcache.r_tag[6][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1520),
    .D(_00690_),
    .Q_N(_14469_),
    .Q(\cpu.dcache.r_tag[6][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1521),
    .D(_00691_),
    .Q_N(_14468_),
    .Q(\cpu.dcache.r_tag[6][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1522),
    .D(_00692_),
    .Q_N(_14467_),
    .Q(\cpu.dcache.r_tag[6][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1523),
    .D(_00693_),
    .Q_N(_14466_),
    .Q(\cpu.dcache.r_tag[6][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1524),
    .D(_00694_),
    .Q_N(_14465_),
    .Q(\cpu.dcache.r_tag[6][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1525),
    .D(_00695_),
    .Q_N(_14464_),
    .Q(\cpu.dcache.r_tag[6][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1526),
    .D(_00696_),
    .Q_N(_14463_),
    .Q(\cpu.dcache.r_tag[6][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1527),
    .D(_00697_),
    .Q_N(_14462_),
    .Q(\cpu.dcache.r_tag[6][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1528),
    .D(_00698_),
    .Q_N(_14461_),
    .Q(\cpu.dcache.r_tag[6][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1529),
    .D(_00699_),
    .Q_N(_14460_),
    .Q(\cpu.dcache.r_tag[7][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1530),
    .D(_00700_),
    .Q_N(_14459_),
    .Q(\cpu.dcache.r_tag[7][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1531),
    .D(_00701_),
    .Q_N(_14458_),
    .Q(\cpu.dcache.r_tag[7][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1532),
    .D(_00702_),
    .Q_N(_14457_),
    .Q(\cpu.dcache.r_tag[7][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1533),
    .D(_00703_),
    .Q_N(_14456_),
    .Q(\cpu.dcache.r_tag[7][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1534),
    .D(_00704_),
    .Q_N(_14455_),
    .Q(\cpu.dcache.r_tag[7][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1535),
    .D(_00705_),
    .Q_N(_14454_),
    .Q(\cpu.dcache.r_tag[7][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1536),
    .D(_00706_),
    .Q_N(_14453_),
    .Q(\cpu.dcache.r_tag[7][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1537),
    .D(_00707_),
    .Q_N(_14452_),
    .Q(\cpu.dcache.r_tag[7][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1538),
    .D(_00708_),
    .Q_N(_14451_),
    .Q(\cpu.dcache.r_tag[7][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1539),
    .D(_00709_),
    .Q_N(_14450_),
    .Q(\cpu.dcache.r_tag[7][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1540),
    .D(_00710_),
    .Q_N(_14449_),
    .Q(\cpu.dcache.r_tag[7][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1541),
    .D(_00711_),
    .Q_N(_14448_),
    .Q(\cpu.dcache.r_tag[7][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1542),
    .D(_00712_),
    .Q_N(_14447_),
    .Q(\cpu.dcache.r_tag[7][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1543),
    .D(_00713_),
    .Q_N(_14446_),
    .Q(\cpu.dcache.r_tag[7][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1544),
    .D(_00714_),
    .Q_N(_14445_),
    .Q(\cpu.dcache.r_tag[7][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1545),
    .D(_00715_),
    .Q_N(_14444_),
    .Q(\cpu.dcache.r_tag[7][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1546),
    .D(_00716_),
    .Q_N(_14443_),
    .Q(\cpu.dcache.r_tag[7][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1547),
    .D(_00717_),
    .Q_N(_14442_),
    .Q(\cpu.dcache.r_tag[7][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1548),
    .D(_00718_),
    .Q_N(_14441_),
    .Q(\cpu.dcache.r_valid[0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1549),
    .D(_00719_),
    .Q_N(_14440_),
    .Q(\cpu.dcache.r_valid[1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1550),
    .D(_00720_),
    .Q_N(_14439_),
    .Q(\cpu.dcache.r_valid[2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1551),
    .D(_00721_),
    .Q_N(_14438_),
    .Q(\cpu.dcache.r_valid[3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1552),
    .D(_00722_),
    .Q_N(_14437_),
    .Q(\cpu.dcache.r_valid[4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1553),
    .D(_00723_),
    .Q_N(_14436_),
    .Q(\cpu.dcache.r_valid[5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1554),
    .D(_00724_),
    .Q_N(_14435_),
    .Q(\cpu.dcache.r_valid[6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1555),
    .D(_00725_),
    .Q_N(_14434_),
    .Q(\cpu.dcache.r_valid[7] ));
 sg13g2_dfrbp_1 \cpu.dec.r_br$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1556),
    .D(_00726_),
    .Q_N(_14433_),
    .Q(\cpu.br ));
 sg13g2_dfrbp_1 \cpu.dec.r_cond[0]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1557),
    .D(_00727_),
    .Q_N(_14432_),
    .Q(\cpu.cond[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_cond[1]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1558),
    .D(_00728_),
    .Q_N(_14431_),
    .Q(\cpu.cond[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_cond[2]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1559),
    .D(_00729_),
    .Q_N(_00252_),
    .Q(\cpu.cond[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_div$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1560),
    .D(_00730_),
    .Q_N(_14430_),
    .Q(\cpu.dec.div ));
 sg13g2_dfrbp_1 \cpu.dec.r_flush_all$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1561),
    .D(_00731_),
    .Q_N(_14429_),
    .Q(\cpu.dec.do_flush_all ));
 sg13g2_dfrbp_1 \cpu.dec.r_flush_write$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1562),
    .D(_00732_),
    .Q_N(_14428_),
    .Q(\cpu.dec.do_flush_write ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[0]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1563),
    .D(_00733_),
    .Q_N(_14427_),
    .Q(\cpu.dec.imm[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[10]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1564),
    .D(_00734_),
    .Q_N(_14426_),
    .Q(\cpu.dec.imm[10] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[11]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1565),
    .D(_00735_),
    .Q_N(_14425_),
    .Q(\cpu.dec.imm[11] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[12]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1566),
    .D(_00736_),
    .Q_N(_14424_),
    .Q(\cpu.dec.imm[12] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[13]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1567),
    .D(_00737_),
    .Q_N(_14423_),
    .Q(\cpu.dec.imm[13] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[14]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1568),
    .D(_00738_),
    .Q_N(_14422_),
    .Q(\cpu.dec.imm[14] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[15]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1569),
    .D(_00739_),
    .Q_N(_14421_),
    .Q(\cpu.dec.imm[15] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[1]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1570),
    .D(_00740_),
    .Q_N(_14420_),
    .Q(\cpu.dec.imm[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[2]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1571),
    .D(_00741_),
    .Q_N(_14419_),
    .Q(\cpu.dec.imm[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[3]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1572),
    .D(_00742_),
    .Q_N(_14418_),
    .Q(\cpu.dec.imm[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[4]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1573),
    .D(_00743_),
    .Q_N(_14417_),
    .Q(\cpu.dec.imm[4] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[5]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1574),
    .D(_00744_),
    .Q_N(_14416_),
    .Q(\cpu.dec.imm[5] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[6]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1575),
    .D(_00745_),
    .Q_N(_14415_),
    .Q(\cpu.dec.imm[6] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[7]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1576),
    .D(_00746_),
    .Q_N(_14414_),
    .Q(\cpu.dec.imm[7] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[8]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1577),
    .D(_00747_),
    .Q_N(_14413_),
    .Q(\cpu.dec.imm[8] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[9]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1578),
    .D(_00748_),
    .Q_N(_14412_),
    .Q(\cpu.dec.imm[9] ));
 sg13g2_dfrbp_1 \cpu.dec.r_inv_mmu$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1579),
    .D(_00749_),
    .Q_N(_14411_),
    .Q(\cpu.dec.do_inv_mmu ));
 sg13g2_dfrbp_1 \cpu.dec.r_io$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1580),
    .D(_00750_),
    .Q_N(_14410_),
    .Q(\cpu.dec.io ));
 sg13g2_dfrbp_1 \cpu.dec.r_jmp$_SDFFCE_PP0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1581),
    .D(_00751_),
    .Q_N(_00236_),
    .Q(\cpu.dec.jmp ));
 sg13g2_dfrbp_1 \cpu.dec.r_load$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1582),
    .D(_00752_),
    .Q_N(_14409_),
    .Q(\cpu.dec.load ));
 sg13g2_dfrbp_1 \cpu.dec.r_mult$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1583),
    .D(_00753_),
    .Q_N(_14408_),
    .Q(\cpu.dec.mult ));
 sg13g2_dfrbp_1 \cpu.dec.r_needs_rs2$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1584),
    .D(_00754_),
    .Q_N(_14821_),
    .Q(\cpu.dec.needs_rs2 ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[10]$_DFF_P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1585),
    .D(_00011_),
    .Q_N(_14822_),
    .Q(\cpu.dec.r_op[10] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[1]$_DFF_P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1586),
    .D(_00012_),
    .Q_N(_14823_),
    .Q(\cpu.dec.r_op[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[2]$_DFF_P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1587),
    .D(_00013_),
    .Q_N(_14824_),
    .Q(\cpu.dec.r_op[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[3]$_DFF_P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1588),
    .D(_00014_),
    .Q_N(_14825_),
    .Q(\cpu.dec.r_op[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[4]$_DFF_P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1589),
    .D(_00015_),
    .Q_N(_14826_),
    .Q(\cpu.dec.r_op[4] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[5]$_DFF_P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1590),
    .D(_00016_),
    .Q_N(_14827_),
    .Q(\cpu.dec.r_op[5] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[6]$_DFF_P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1591),
    .D(_00017_),
    .Q_N(_14828_),
    .Q(\cpu.dec.r_op[6] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[7]$_DFF_P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1592),
    .D(_00018_),
    .Q_N(_14829_),
    .Q(\cpu.dec.r_op[7] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[8]$_DFF_P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1593),
    .D(_00019_),
    .Q_N(_14830_),
    .Q(\cpu.dec.r_op[8] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[9]$_DFF_P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1594),
    .D(_00020_),
    .Q_N(_14407_),
    .Q(\cpu.dec.r_op[9] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[0]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1595),
    .D(_00755_),
    .Q_N(_14406_),
    .Q(\cpu.dec.r_rd[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[1]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1596),
    .D(_00756_),
    .Q_N(_14405_),
    .Q(\cpu.dec.r_rd[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[2]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1597),
    .D(_00757_),
    .Q_N(_14404_),
    .Q(\cpu.dec.r_rd[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[3]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1598),
    .D(_00758_),
    .Q_N(_14831_),
    .Q(\cpu.dec.r_rd[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_ready$_DFF_P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1599),
    .D(_00052_),
    .Q_N(_14403_),
    .Q(\cpu.dec.iready ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[0]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1600),
    .D(_00759_),
    .Q_N(_14402_),
    .Q(\cpu.dec.r_rs1[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[1]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1601),
    .D(_00760_),
    .Q_N(_14401_),
    .Q(\cpu.dec.r_rs1[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[2]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1602),
    .D(_00761_),
    .Q_N(_14400_),
    .Q(\cpu.dec.r_rs1[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[3]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1603),
    .D(_00762_),
    .Q_N(_14399_),
    .Q(\cpu.dec.r_rs1[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[0]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1604),
    .D(_00763_),
    .Q_N(_14398_),
    .Q(\cpu.dec.r_rs2[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[1]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1605),
    .D(_00764_),
    .Q_N(_14397_),
    .Q(\cpu.dec.r_rs2[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[2]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1606),
    .D(_00765_),
    .Q_N(_14396_),
    .Q(\cpu.dec.r_rs2[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[3]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1607),
    .D(_00766_),
    .Q_N(_14395_),
    .Q(\cpu.dec.r_rs2[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2_pc$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1608),
    .D(_00767_),
    .Q_N(_14394_),
    .Q(\cpu.dec.r_rs2_pc ));
 sg13g2_dfrbp_1 \cpu.dec.r_set_cc$_SDFFCE_PP0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1609),
    .D(_00768_),
    .Q_N(_14393_),
    .Q(\cpu.dec.r_set_cc ));
 sg13g2_dfrbp_1 \cpu.dec.r_store$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1610),
    .D(_00769_),
    .Q_N(_00277_),
    .Q(\cpu.dec.r_store ));
 sg13g2_dfrbp_1 \cpu.dec.r_swapsp$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1611),
    .D(_00770_),
    .Q_N(_14392_),
    .Q(\cpu.dec.r_swapsp ));
 sg13g2_dfrbp_1 \cpu.dec.r_sys_call$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1612),
    .D(_00771_),
    .Q_N(_00253_),
    .Q(\cpu.dec.r_sys_call ));
 sg13g2_dfrbp_1 \cpu.dec.r_trap$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1613),
    .D(_00772_),
    .Q_N(_14391_),
    .Q(\cpu.dec.r_trap ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_mmu_d_proxy$_SDFFE_PP0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1614),
    .D(_00773_),
    .Q_N(_14390_),
    .Q(\cpu.ex.genblk3.r_mmu_d_proxy ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_mmu_enable$_SDFFE_PN0P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1615),
    .D(_00774_),
    .Q_N(_00176_),
    .Q(\cpu.ex.genblk3.r_mmu_enable ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_prev_supmode$_SDFFE_PN1P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1616),
    .D(_00775_),
    .Q_N(_14832_),
    .Q(\cpu.ex.genblk3.r_prev_supmode ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_supmode$_DFF_P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1617),
    .D(\cpu.ex.genblk3.c_supmode ),
    .Q_N(_00177_),
    .Q(\cpu.dec.supmode ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_user_io$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1618),
    .D(_00776_),
    .Q_N(_14389_),
    .Q(\cpu.dec.user_io ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[0]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1619),
    .D(_00777_),
    .Q_N(_14388_),
    .Q(\cpu.ex.r_10[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[10]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1620),
    .D(_00778_),
    .Q_N(_14387_),
    .Q(\cpu.ex.r_10[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[11]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1621),
    .D(_00779_),
    .Q_N(_14386_),
    .Q(\cpu.ex.r_10[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[12]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1622),
    .D(_00780_),
    .Q_N(_14385_),
    .Q(\cpu.ex.r_10[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[13]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1623),
    .D(_00781_),
    .Q_N(_14384_),
    .Q(\cpu.ex.r_10[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[14]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1624),
    .D(_00782_),
    .Q_N(_14383_),
    .Q(\cpu.ex.r_10[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[15]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1625),
    .D(_00783_),
    .Q_N(_14382_),
    .Q(\cpu.ex.r_10[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[1]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1626),
    .D(_00784_),
    .Q_N(_14381_),
    .Q(\cpu.ex.r_10[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[2]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1627),
    .D(_00785_),
    .Q_N(_14380_),
    .Q(\cpu.ex.r_10[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[3]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1628),
    .D(_00786_),
    .Q_N(_14379_),
    .Q(\cpu.ex.r_10[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[4]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1629),
    .D(_00787_),
    .Q_N(_14378_),
    .Q(\cpu.ex.r_10[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[5]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1630),
    .D(_00788_),
    .Q_N(_14377_),
    .Q(\cpu.ex.r_10[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[6]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1631),
    .D(_00789_),
    .Q_N(_14376_),
    .Q(\cpu.ex.r_10[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[7]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1632),
    .D(_00790_),
    .Q_N(_14375_),
    .Q(\cpu.ex.r_10[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[8]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1633),
    .D(_00791_),
    .Q_N(_14374_),
    .Q(\cpu.ex.r_10[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[9]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1634),
    .D(_00792_),
    .Q_N(_14373_),
    .Q(\cpu.ex.r_10[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[0]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1635),
    .D(_00793_),
    .Q_N(_14372_),
    .Q(\cpu.ex.r_11[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[10]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1636),
    .D(_00794_),
    .Q_N(_14371_),
    .Q(\cpu.ex.r_11[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[11]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1637),
    .D(_00795_),
    .Q_N(_14370_),
    .Q(\cpu.ex.r_11[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[12]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1638),
    .D(_00796_),
    .Q_N(_14369_),
    .Q(\cpu.ex.r_11[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[13]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1639),
    .D(_00797_),
    .Q_N(_14368_),
    .Q(\cpu.ex.r_11[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[14]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1640),
    .D(_00798_),
    .Q_N(_14367_),
    .Q(\cpu.ex.r_11[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[15]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1641),
    .D(_00799_),
    .Q_N(_14366_),
    .Q(\cpu.ex.r_11[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[1]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1642),
    .D(_00800_),
    .Q_N(_14365_),
    .Q(\cpu.ex.r_11[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[2]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1643),
    .D(_00801_),
    .Q_N(_14364_),
    .Q(\cpu.ex.r_11[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[3]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1644),
    .D(_00802_),
    .Q_N(_14363_),
    .Q(\cpu.ex.r_11[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[4]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1645),
    .D(_00803_),
    .Q_N(_14362_),
    .Q(\cpu.ex.r_11[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[5]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1646),
    .D(_00804_),
    .Q_N(_14361_),
    .Q(\cpu.ex.r_11[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[6]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1647),
    .D(_00805_),
    .Q_N(_14360_),
    .Q(\cpu.ex.r_11[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[7]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1648),
    .D(_00806_),
    .Q_N(_14359_),
    .Q(\cpu.ex.r_11[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[8]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1649),
    .D(_00807_),
    .Q_N(_14358_),
    .Q(\cpu.ex.r_11[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[9]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1650),
    .D(_00808_),
    .Q_N(_14357_),
    .Q(\cpu.ex.r_11[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[0]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1651),
    .D(_00809_),
    .Q_N(_14356_),
    .Q(\cpu.ex.r_12[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[10]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1652),
    .D(_00810_),
    .Q_N(_14355_),
    .Q(\cpu.ex.r_12[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[11]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1653),
    .D(_00811_),
    .Q_N(_14354_),
    .Q(\cpu.ex.r_12[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[12]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1654),
    .D(_00812_),
    .Q_N(_14353_),
    .Q(\cpu.ex.r_12[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[13]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1655),
    .D(_00813_),
    .Q_N(_14352_),
    .Q(\cpu.ex.r_12[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[14]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1656),
    .D(_00814_),
    .Q_N(_14351_),
    .Q(\cpu.ex.r_12[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[15]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1657),
    .D(_00815_),
    .Q_N(_14350_),
    .Q(\cpu.ex.r_12[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[1]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1658),
    .D(_00816_),
    .Q_N(_14349_),
    .Q(\cpu.ex.r_12[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[2]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1659),
    .D(_00817_),
    .Q_N(_14348_),
    .Q(\cpu.ex.r_12[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[3]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1660),
    .D(_00818_),
    .Q_N(_14347_),
    .Q(\cpu.ex.r_12[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[4]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1661),
    .D(_00819_),
    .Q_N(_14346_),
    .Q(\cpu.ex.r_12[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[5]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1662),
    .D(_00820_),
    .Q_N(_14345_),
    .Q(\cpu.ex.r_12[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[6]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1663),
    .D(_00821_),
    .Q_N(_14344_),
    .Q(\cpu.ex.r_12[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[7]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1664),
    .D(_00822_),
    .Q_N(_14343_),
    .Q(\cpu.ex.r_12[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[8]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1665),
    .D(_00823_),
    .Q_N(_14342_),
    .Q(\cpu.ex.r_12[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[9]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1666),
    .D(_00824_),
    .Q_N(_14341_),
    .Q(\cpu.ex.r_12[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[0]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1667),
    .D(_00825_),
    .Q_N(_14340_),
    .Q(\cpu.ex.r_13[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[10]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1668),
    .D(_00826_),
    .Q_N(_14339_),
    .Q(\cpu.ex.r_13[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[11]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1669),
    .D(_00827_),
    .Q_N(_14338_),
    .Q(\cpu.ex.r_13[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[12]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1670),
    .D(_00828_),
    .Q_N(_14337_),
    .Q(\cpu.ex.r_13[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[13]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1671),
    .D(_00829_),
    .Q_N(_14336_),
    .Q(\cpu.ex.r_13[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[14]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1672),
    .D(_00830_),
    .Q_N(_14335_),
    .Q(\cpu.ex.r_13[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[15]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1673),
    .D(_00831_),
    .Q_N(_14334_),
    .Q(\cpu.ex.r_13[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[1]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1674),
    .D(_00832_),
    .Q_N(_14333_),
    .Q(\cpu.ex.r_13[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[2]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1675),
    .D(_00833_),
    .Q_N(_14332_),
    .Q(\cpu.ex.r_13[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[3]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1676),
    .D(_00834_),
    .Q_N(_14331_),
    .Q(\cpu.ex.r_13[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[4]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1677),
    .D(_00835_),
    .Q_N(_14330_),
    .Q(\cpu.ex.r_13[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[5]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1678),
    .D(_00836_),
    .Q_N(_14329_),
    .Q(\cpu.ex.r_13[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[6]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1679),
    .D(_00837_),
    .Q_N(_14328_),
    .Q(\cpu.ex.r_13[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[7]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1680),
    .D(_00838_),
    .Q_N(_14327_),
    .Q(\cpu.ex.r_13[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[8]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1681),
    .D(_00839_),
    .Q_N(_14326_),
    .Q(\cpu.ex.r_13[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[9]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1682),
    .D(_00840_),
    .Q_N(_14325_),
    .Q(\cpu.ex.r_13[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[0]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1683),
    .D(_00841_),
    .Q_N(_14324_),
    .Q(\cpu.ex.r_14[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[10]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1684),
    .D(_00842_),
    .Q_N(_14323_),
    .Q(\cpu.ex.r_14[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[11]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1685),
    .D(_00843_),
    .Q_N(_14322_),
    .Q(\cpu.ex.r_14[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[12]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1686),
    .D(_00844_),
    .Q_N(_14321_),
    .Q(\cpu.ex.r_14[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[13]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1687),
    .D(_00845_),
    .Q_N(_14320_),
    .Q(\cpu.ex.r_14[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[14]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1688),
    .D(_00846_),
    .Q_N(_14319_),
    .Q(\cpu.ex.r_14[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[15]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1689),
    .D(_00847_),
    .Q_N(_14318_),
    .Q(\cpu.ex.r_14[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[1]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1690),
    .D(_00848_),
    .Q_N(_14317_),
    .Q(\cpu.ex.r_14[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[2]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1691),
    .D(_00849_),
    .Q_N(_14316_),
    .Q(\cpu.ex.r_14[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[3]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1692),
    .D(_00850_),
    .Q_N(_14315_),
    .Q(\cpu.ex.r_14[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[4]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1693),
    .D(_00851_),
    .Q_N(_14314_),
    .Q(\cpu.ex.r_14[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[5]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1694),
    .D(_00852_),
    .Q_N(_14313_),
    .Q(\cpu.ex.r_14[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[6]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1695),
    .D(_00853_),
    .Q_N(_14312_),
    .Q(\cpu.ex.r_14[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[7]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1696),
    .D(_00854_),
    .Q_N(_14311_),
    .Q(\cpu.ex.r_14[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[8]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1697),
    .D(_00855_),
    .Q_N(_14310_),
    .Q(\cpu.ex.r_14[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[9]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1698),
    .D(_00856_),
    .Q_N(_14309_),
    .Q(\cpu.ex.r_14[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[0]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1699),
    .D(_00857_),
    .Q_N(_14308_),
    .Q(\cpu.ex.r_15[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[10]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1700),
    .D(_00858_),
    .Q_N(_00246_),
    .Q(\cpu.ex.r_15[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[11]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1701),
    .D(_00859_),
    .Q_N(_00247_),
    .Q(\cpu.ex.r_15[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[12]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1702),
    .D(_00860_),
    .Q_N(_00248_),
    .Q(\cpu.ex.r_15[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[13]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1703),
    .D(_00861_),
    .Q_N(_00249_),
    .Q(\cpu.ex.r_15[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[14]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1704),
    .D(_00862_),
    .Q_N(_00250_),
    .Q(\cpu.ex.r_15[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[15]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1705),
    .D(_00863_),
    .Q_N(_00251_),
    .Q(\cpu.ex.r_15[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[1]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1706),
    .D(_00864_),
    .Q_N(_00237_),
    .Q(\cpu.ex.r_15[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[2]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1707),
    .D(_00865_),
    .Q_N(_00238_),
    .Q(\cpu.ex.r_15[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[3]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1708),
    .D(_00866_),
    .Q_N(_00239_),
    .Q(\cpu.ex.r_15[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[4]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1709),
    .D(_00867_),
    .Q_N(_00240_),
    .Q(\cpu.ex.r_15[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[5]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1710),
    .D(_00868_),
    .Q_N(_00241_),
    .Q(\cpu.ex.r_15[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[6]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1711),
    .D(_00869_),
    .Q_N(_00242_),
    .Q(\cpu.ex.r_15[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[7]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1712),
    .D(_00870_),
    .Q_N(_00243_),
    .Q(\cpu.ex.r_15[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[8]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1713),
    .D(_00871_),
    .Q_N(_00244_),
    .Q(\cpu.ex.r_15[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[9]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1714),
    .D(_00872_),
    .Q_N(_00245_),
    .Q(\cpu.ex.r_15[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[0]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1715),
    .D(_00873_),
    .Q_N(_14307_),
    .Q(\cpu.ex.r_8[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[10]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1716),
    .D(_00874_),
    .Q_N(_14306_),
    .Q(\cpu.ex.r_8[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[11]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1717),
    .D(_00875_),
    .Q_N(_14305_),
    .Q(\cpu.ex.r_8[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[12]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1718),
    .D(_00876_),
    .Q_N(_14304_),
    .Q(\cpu.ex.r_8[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[13]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1719),
    .D(_00877_),
    .Q_N(_14303_),
    .Q(\cpu.ex.r_8[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[14]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1720),
    .D(_00878_),
    .Q_N(_14302_),
    .Q(\cpu.ex.r_8[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[15]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1721),
    .D(_00879_),
    .Q_N(_14301_),
    .Q(\cpu.ex.r_8[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[1]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1722),
    .D(_00880_),
    .Q_N(_14300_),
    .Q(\cpu.ex.r_8[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[2]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1723),
    .D(_00881_),
    .Q_N(_14299_),
    .Q(\cpu.ex.r_8[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[3]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1724),
    .D(_00882_),
    .Q_N(_14298_),
    .Q(\cpu.ex.r_8[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[4]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1725),
    .D(_00883_),
    .Q_N(_14297_),
    .Q(\cpu.ex.r_8[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[5]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1726),
    .D(_00884_),
    .Q_N(_14296_),
    .Q(\cpu.ex.r_8[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[6]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1727),
    .D(_00885_),
    .Q_N(_14295_),
    .Q(\cpu.ex.r_8[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[7]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1728),
    .D(_00886_),
    .Q_N(_14294_),
    .Q(\cpu.ex.r_8[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[8]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1729),
    .D(_00887_),
    .Q_N(_14293_),
    .Q(\cpu.ex.r_8[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[9]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1730),
    .D(_00888_),
    .Q_N(_14292_),
    .Q(\cpu.ex.r_8[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[0]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1731),
    .D(_00889_),
    .Q_N(_14291_),
    .Q(\cpu.ex.r_9[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[10]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1732),
    .D(_00890_),
    .Q_N(_14290_),
    .Q(\cpu.ex.r_9[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[11]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1733),
    .D(_00891_),
    .Q_N(_14289_),
    .Q(\cpu.ex.r_9[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[12]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1734),
    .D(_00892_),
    .Q_N(_14288_),
    .Q(\cpu.ex.r_9[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[13]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1735),
    .D(_00893_),
    .Q_N(_14287_),
    .Q(\cpu.ex.r_9[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[14]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1736),
    .D(_00894_),
    .Q_N(_14286_),
    .Q(\cpu.ex.r_9[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[15]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1737),
    .D(_00895_),
    .Q_N(_14285_),
    .Q(\cpu.ex.r_9[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[1]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1738),
    .D(_00896_),
    .Q_N(_14284_),
    .Q(\cpu.ex.r_9[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[2]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1739),
    .D(_00897_),
    .Q_N(_14283_),
    .Q(\cpu.ex.r_9[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[3]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1740),
    .D(_00898_),
    .Q_N(_14282_),
    .Q(\cpu.ex.r_9[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[4]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1741),
    .D(_00899_),
    .Q_N(_14281_),
    .Q(\cpu.ex.r_9[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[5]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1742),
    .D(_00900_),
    .Q_N(_14280_),
    .Q(\cpu.ex.r_9[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[6]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1743),
    .D(_00901_),
    .Q_N(_14279_),
    .Q(\cpu.ex.r_9[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[7]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1744),
    .D(_00902_),
    .Q_N(_14278_),
    .Q(\cpu.ex.r_9[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[8]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1745),
    .D(_00903_),
    .Q_N(_14277_),
    .Q(\cpu.ex.r_9[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[9]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1746),
    .D(_00904_),
    .Q_N(_14833_),
    .Q(\cpu.ex.r_9[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_branch_stall$_DFF_P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1747),
    .D(_00053_),
    .Q_N(_14276_),
    .Q(\cpu.ex.r_branch_stall ));
 sg13g2_dfrbp_1 \cpu.ex.r_d_flush_all$_SDFF_PP0_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1748),
    .D(_00905_),
    .Q_N(_14834_),
    .Q(\cpu.d_flush_all ));
 sg13g2_dfrbp_1 \cpu.ex.r_div_running$_DFF_P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1749),
    .D(\cpu.ex.c_div_running ),
    .Q_N(_14275_),
    .Q(\cpu.ex.r_div_running ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[0]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1750),
    .D(_00906_),
    .Q_N(_14274_),
    .Q(\cpu.ex.r_epc[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[10]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1751),
    .D(_00907_),
    .Q_N(_14273_),
    .Q(\cpu.ex.r_epc[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[11]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1752),
    .D(_00908_),
    .Q_N(_14272_),
    .Q(\cpu.ex.r_epc[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[12]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1753),
    .D(_00909_),
    .Q_N(_14271_),
    .Q(\cpu.ex.r_epc[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[13]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1754),
    .D(_00910_),
    .Q_N(_14270_),
    .Q(\cpu.ex.r_epc[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[14]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1755),
    .D(_00911_),
    .Q_N(_14269_),
    .Q(\cpu.ex.r_epc[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[1]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1756),
    .D(_00912_),
    .Q_N(_14268_),
    .Q(\cpu.ex.r_epc[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[2]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1757),
    .D(_00913_),
    .Q_N(_14267_),
    .Q(\cpu.ex.r_epc[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[3]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1758),
    .D(_00914_),
    .Q_N(_14266_),
    .Q(\cpu.ex.r_epc[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[4]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1759),
    .D(_00915_),
    .Q_N(_14265_),
    .Q(\cpu.ex.r_epc[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[5]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1760),
    .D(_00916_),
    .Q_N(_14264_),
    .Q(\cpu.ex.r_epc[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[6]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1761),
    .D(_00917_),
    .Q_N(_14263_),
    .Q(\cpu.ex.r_epc[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[7]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1762),
    .D(_00918_),
    .Q_N(_14262_),
    .Q(\cpu.ex.r_epc[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[8]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1763),
    .D(_00919_),
    .Q_N(_14261_),
    .Q(\cpu.ex.r_epc[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[9]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1764),
    .D(_00920_),
    .Q_N(_14260_),
    .Q(\cpu.ex.r_epc[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_fetch$_SDFF_PN1_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1765),
    .D(_00921_),
    .Q_N(_00173_),
    .Q(\cpu.ex.ifetch ));
 sg13g2_dfrbp_1 \cpu.ex.r_flush_write$_SDFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1766),
    .D(_00922_),
    .Q_N(_14259_),
    .Q(\cpu.dcache.flush_write ));
 sg13g2_dfrbp_1 \cpu.ex.r_i_flush_all$_SDFF_PP0_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1767),
    .D(_00923_),
    .Q_N(_14258_),
    .Q(\cpu.ex.i_flush_all ));
 sg13g2_dfrbp_1 \cpu.ex.r_ie$_SDFFE_PP0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1768),
    .D(_00924_),
    .Q_N(_14257_),
    .Q(\cpu.ex.r_ie ));
 sg13g2_dfrbp_1 \cpu.ex.r_io_access$_SDFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1769),
    .D(_00925_),
    .Q_N(_00181_),
    .Q(\cpu.ex.io_access ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[0]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1770),
    .D(_00926_),
    .Q_N(_14256_),
    .Q(\cpu.ex.r_lr[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[10]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1771),
    .D(_00927_),
    .Q_N(_14255_),
    .Q(\cpu.ex.r_lr[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[11]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1772),
    .D(_00928_),
    .Q_N(_14254_),
    .Q(\cpu.ex.r_lr[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[12]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1773),
    .D(_00929_),
    .Q_N(_14253_),
    .Q(\cpu.ex.r_lr[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[13]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1774),
    .D(_00930_),
    .Q_N(_14252_),
    .Q(\cpu.ex.r_lr[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[14]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1775),
    .D(_00931_),
    .Q_N(_14251_),
    .Q(\cpu.ex.r_lr[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[1]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1776),
    .D(_00932_),
    .Q_N(_14250_),
    .Q(\cpu.ex.r_lr[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[2]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1777),
    .D(_00933_),
    .Q_N(_14249_),
    .Q(\cpu.ex.r_lr[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[3]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1778),
    .D(_00934_),
    .Q_N(_14248_),
    .Q(\cpu.ex.r_lr[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[4]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1779),
    .D(_00935_),
    .Q_N(_14247_),
    .Q(\cpu.ex.r_lr[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[5]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1780),
    .D(_00936_),
    .Q_N(_14246_),
    .Q(\cpu.ex.r_lr[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[6]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1781),
    .D(_00937_),
    .Q_N(_14245_),
    .Q(\cpu.ex.r_lr[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[7]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1782),
    .D(_00938_),
    .Q_N(_14244_),
    .Q(\cpu.ex.r_lr[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[8]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1783),
    .D(_00939_),
    .Q_N(_14243_),
    .Q(\cpu.ex.r_lr[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[9]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1784),
    .D(_00940_),
    .Q_N(_14835_),
    .Q(\cpu.ex.r_lr[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[0]$_DFF_P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1785),
    .D(\cpu.ex.c_mult[0] ),
    .Q_N(_14836_),
    .Q(\cpu.ex.r_mult[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[10]$_DFF_P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1786),
    .D(\cpu.ex.c_mult[10] ),
    .Q_N(_14837_),
    .Q(\cpu.ex.r_mult[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[11]$_DFF_P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1787),
    .D(\cpu.ex.c_mult[11] ),
    .Q_N(_14838_),
    .Q(\cpu.ex.r_mult[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[12]$_DFF_P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1788),
    .D(\cpu.ex.c_mult[12] ),
    .Q_N(_14839_),
    .Q(\cpu.ex.r_mult[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[13]$_DFF_P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1789),
    .D(\cpu.ex.c_mult[13] ),
    .Q_N(_14840_),
    .Q(\cpu.ex.r_mult[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[14]$_DFF_P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1790),
    .D(\cpu.ex.c_mult[14] ),
    .Q_N(_00149_),
    .Q(\cpu.ex.r_mult[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[15]$_DFF_P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1791),
    .D(\cpu.ex.c_mult[15] ),
    .Q_N(_14242_),
    .Q(\cpu.ex.r_mult[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[16]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1792),
    .D(_00941_),
    .Q_N(_14241_),
    .Q(\cpu.ex.r_mult[16] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[17]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1793),
    .D(_00942_),
    .Q_N(_14240_),
    .Q(\cpu.ex.r_mult[17] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[18]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1794),
    .D(_00943_),
    .Q_N(_14239_),
    .Q(\cpu.ex.r_mult[18] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[19]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1795),
    .D(_00944_),
    .Q_N(_14841_),
    .Q(\cpu.ex.r_mult[19] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[1]$_DFF_P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1796),
    .D(\cpu.ex.c_mult[1] ),
    .Q_N(_14238_),
    .Q(\cpu.ex.r_mult[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[20]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1797),
    .D(_00945_),
    .Q_N(_14237_),
    .Q(\cpu.ex.r_mult[20] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[21]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1798),
    .D(_00946_),
    .Q_N(_14236_),
    .Q(\cpu.ex.r_mult[21] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[22]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1799),
    .D(_00947_),
    .Q_N(_14235_),
    .Q(\cpu.ex.r_mult[22] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[23]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1800),
    .D(_00948_),
    .Q_N(_14234_),
    .Q(\cpu.ex.r_mult[23] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[24]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1801),
    .D(_00949_),
    .Q_N(_14233_),
    .Q(\cpu.ex.r_mult[24] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[25]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1802),
    .D(_00950_),
    .Q_N(_14232_),
    .Q(\cpu.ex.r_mult[25] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[26]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1803),
    .D(_00951_),
    .Q_N(_14231_),
    .Q(\cpu.ex.r_mult[26] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[27]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1804),
    .D(_00952_),
    .Q_N(_14230_),
    .Q(\cpu.ex.r_mult[27] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[28]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1805),
    .D(_00953_),
    .Q_N(_14229_),
    .Q(\cpu.ex.r_mult[28] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[29]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1806),
    .D(_00954_),
    .Q_N(_14842_),
    .Q(\cpu.ex.r_mult[29] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[2]$_DFF_P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1807),
    .D(\cpu.ex.c_mult[2] ),
    .Q_N(_14228_),
    .Q(\cpu.ex.r_mult[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[30]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1808),
    .D(_00955_),
    .Q_N(_14227_),
    .Q(\cpu.ex.r_mult[30] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[31]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1809),
    .D(_00956_),
    .Q_N(_14843_),
    .Q(\cpu.ex.r_mult[31] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[3]$_DFF_P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1810),
    .D(\cpu.ex.c_mult[3] ),
    .Q_N(_14844_),
    .Q(\cpu.ex.r_mult[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[4]$_DFF_P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1811),
    .D(\cpu.ex.c_mult[4] ),
    .Q_N(_14845_),
    .Q(\cpu.ex.r_mult[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[5]$_DFF_P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1812),
    .D(\cpu.ex.c_mult[5] ),
    .Q_N(_14846_),
    .Q(\cpu.ex.r_mult[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[6]$_DFF_P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1813),
    .D(\cpu.ex.c_mult[6] ),
    .Q_N(_14847_),
    .Q(\cpu.ex.r_mult[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[7]$_DFF_P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1814),
    .D(\cpu.ex.c_mult[7] ),
    .Q_N(_14848_),
    .Q(\cpu.ex.r_mult[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[8]$_DFF_P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1815),
    .D(\cpu.ex.c_mult[8] ),
    .Q_N(_14849_),
    .Q(\cpu.ex.r_mult[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[9]$_DFF_P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1816),
    .D(\cpu.ex.c_mult[9] ),
    .Q_N(_14850_),
    .Q(\cpu.ex.r_mult[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[0]$_DFF_P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1817),
    .D(\cpu.ex.c_mult_off[0] ),
    .Q_N(_14851_),
    .Q(\cpu.ex.r_mult_off[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[1]$_DFF_P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1818),
    .D(\cpu.ex.c_mult_off[1] ),
    .Q_N(_14852_),
    .Q(\cpu.ex.r_mult_off[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[2]$_DFF_P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1819),
    .D(\cpu.ex.c_mult_off[2] ),
    .Q_N(_14853_),
    .Q(\cpu.ex.r_mult_off[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[3]$_DFF_P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1820),
    .D(\cpu.ex.c_mult_off[3] ),
    .Q_N(_14854_),
    .Q(\cpu.ex.r_mult_off[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_running$_DFF_P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1821),
    .D(\cpu.ex.c_mult_running ),
    .Q_N(_00183_),
    .Q(\cpu.ex.r_mult_running ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[0]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1822),
    .D(_00957_),
    .Q_N(_00184_),
    .Q(\cpu.ex.pc[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[10]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1823),
    .D(_00958_),
    .Q_N(_00271_),
    .Q(\cpu.ex.pc[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[11]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1824),
    .D(_00959_),
    .Q_N(_00270_),
    .Q(\cpu.ex.pc[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[12]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1825),
    .D(_00960_),
    .Q_N(_00180_),
    .Q(\cpu.ex.pc[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[13]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1826),
    .D(_00961_),
    .Q_N(_00179_),
    .Q(\cpu.ex.pc[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[14]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1827),
    .D(_00962_),
    .Q_N(_00178_),
    .Q(\cpu.ex.pc[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[1]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1828),
    .D(_00963_),
    .Q_N(_00269_),
    .Q(\cpu.ex.pc[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[2]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1829),
    .D(_00964_),
    .Q_N(_00175_),
    .Q(\cpu.ex.pc[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[3]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1830),
    .D(_00965_),
    .Q_N(_00174_),
    .Q(\cpu.ex.pc[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[4]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1831),
    .D(_00966_),
    .Q_N(_00276_),
    .Q(\cpu.ex.pc[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[5]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1832),
    .D(_00967_),
    .Q_N(_00275_),
    .Q(\cpu.ex.pc[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[6]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1833),
    .D(_00968_),
    .Q_N(_00274_),
    .Q(\cpu.ex.pc[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[7]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1834),
    .D(_00969_),
    .Q_N(_00268_),
    .Q(\cpu.ex.pc[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[8]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1835),
    .D(_00970_),
    .Q_N(_00273_),
    .Q(\cpu.ex.pc[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[9]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1836),
    .D(_00971_),
    .Q_N(_00272_),
    .Q(\cpu.ex.pc[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_prev_ie$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1837),
    .D(_00972_),
    .Q_N(_14226_),
    .Q(\cpu.ex.r_prev_ie ));
 sg13g2_dfrbp_1 \cpu.ex.r_read_stall$_SDFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1838),
    .D(_00973_),
    .Q_N(_00182_),
    .Q(\cpu.ex.r_read_stall ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[0]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1839),
    .D(_00974_),
    .Q_N(_14225_),
    .Q(\cpu.ex.r_sp[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[10]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1840),
    .D(_00975_),
    .Q_N(_14224_),
    .Q(\cpu.ex.r_sp[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[11]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1841),
    .D(_00976_),
    .Q_N(_14223_),
    .Q(\cpu.ex.r_sp[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[12]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1842),
    .D(_00977_),
    .Q_N(_14222_),
    .Q(\cpu.ex.r_sp[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[13]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1843),
    .D(_00978_),
    .Q_N(_14221_),
    .Q(\cpu.ex.r_sp[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[14]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1844),
    .D(_00979_),
    .Q_N(_14220_),
    .Q(\cpu.ex.r_sp[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[1]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1845),
    .D(_00980_),
    .Q_N(_14219_),
    .Q(\cpu.ex.r_sp[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[2]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1846),
    .D(_00981_),
    .Q_N(_14218_),
    .Q(\cpu.ex.r_sp[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[3]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1847),
    .D(_00982_),
    .Q_N(_14217_),
    .Q(\cpu.ex.r_sp[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[4]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1848),
    .D(_00983_),
    .Q_N(_14216_),
    .Q(\cpu.ex.r_sp[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[5]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1849),
    .D(_00984_),
    .Q_N(_14215_),
    .Q(\cpu.ex.r_sp[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[6]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1850),
    .D(_00985_),
    .Q_N(_14214_),
    .Q(\cpu.ex.r_sp[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[7]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1851),
    .D(_00986_),
    .Q_N(_14213_),
    .Q(\cpu.ex.r_sp[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[8]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1852),
    .D(_00987_),
    .Q_N(_14212_),
    .Q(\cpu.ex.r_sp[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[9]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1853),
    .D(_00988_),
    .Q_N(_14211_),
    .Q(\cpu.ex.r_sp[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1854),
    .D(_00989_),
    .Q_N(_14210_),
    .Q(\cpu.ex.r_stmp[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[10]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1855),
    .D(_00990_),
    .Q_N(_14209_),
    .Q(\cpu.ex.r_stmp[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[11]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1856),
    .D(_00991_),
    .Q_N(_14208_),
    .Q(\cpu.ex.r_stmp[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[12]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1857),
    .D(_00992_),
    .Q_N(_14207_),
    .Q(\cpu.ex.r_stmp[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[13]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1858),
    .D(_00993_),
    .Q_N(_14206_),
    .Q(\cpu.ex.r_stmp[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[14]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1859),
    .D(_00994_),
    .Q_N(_14205_),
    .Q(\cpu.ex.r_stmp[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[15]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1860),
    .D(_00995_),
    .Q_N(_14204_),
    .Q(\cpu.ex.r_stmp[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[1]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1861),
    .D(_00996_),
    .Q_N(_14203_),
    .Q(\cpu.ex.r_stmp[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[2]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1862),
    .D(_00997_),
    .Q_N(_14202_),
    .Q(\cpu.ex.r_stmp[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[3]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1863),
    .D(_00998_),
    .Q_N(_14201_),
    .Q(\cpu.ex.r_stmp[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[4]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1864),
    .D(_00999_),
    .Q_N(_14200_),
    .Q(\cpu.ex.r_stmp[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[5]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1865),
    .D(_01000_),
    .Q_N(_14199_),
    .Q(\cpu.ex.r_stmp[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[6]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1866),
    .D(_01001_),
    .Q_N(_14198_),
    .Q(\cpu.ex.r_stmp[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[7]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1867),
    .D(_01002_),
    .Q_N(_14197_),
    .Q(\cpu.ex.r_stmp[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[8]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1868),
    .D(_01003_),
    .Q_N(_14196_),
    .Q(\cpu.ex.r_stmp[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[9]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1869),
    .D(_01004_),
    .Q_N(_14195_),
    .Q(\cpu.ex.r_stmp[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[0]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1870),
    .D(_01005_),
    .Q_N(_00235_),
    .Q(\cpu.ex.mmu_reg_data[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[10]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1871),
    .D(_01006_),
    .Q_N(_00217_),
    .Q(\cpu.addr[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[11]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1872),
    .D(_01007_),
    .Q_N(_00219_),
    .Q(\cpu.addr[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[12]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1873),
    .D(_01008_),
    .Q_N(_14194_),
    .Q(\cpu.addr[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[13]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1874),
    .D(_01009_),
    .Q_N(_14193_),
    .Q(\cpu.addr[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[14]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1875),
    .D(_01010_),
    .Q_N(_14192_),
    .Q(\cpu.addr[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[15]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1876),
    .D(_01011_),
    .Q_N(_14191_),
    .Q(\cpu.addr[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[1]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1877),
    .D(_01012_),
    .Q_N(_00254_),
    .Q(\cpu.addr[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[2]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1878),
    .D(_01013_),
    .Q_N(_14190_),
    .Q(\cpu.addr[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[3]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1879),
    .D(_01014_),
    .Q_N(_00201_),
    .Q(\cpu.addr[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[4]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1880),
    .D(_01015_),
    .Q_N(_00206_),
    .Q(\cpu.addr[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[5]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1881),
    .D(_01016_),
    .Q_N(_00207_),
    .Q(\cpu.addr[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[6]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1882),
    .D(_01017_),
    .Q_N(_00209_),
    .Q(\cpu.addr[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[7]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1883),
    .D(_01018_),
    .Q_N(_00211_),
    .Q(\cpu.addr[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[8]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1884),
    .D(_01019_),
    .Q_N(_00213_),
    .Q(\cpu.addr[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[9]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1885),
    .D(_01020_),
    .Q_N(_00215_),
    .Q(\cpu.addr[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1886),
    .D(_01021_),
    .Q_N(_14189_),
    .Q(\cpu.ex.r_wb_addr[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1887),
    .D(_01022_),
    .Q_N(_14188_),
    .Q(\cpu.ex.r_wb_addr[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[2]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1888),
    .D(_01023_),
    .Q_N(_14187_),
    .Q(\cpu.ex.r_wb_addr[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[3]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1889),
    .D(_01024_),
    .Q_N(_14186_),
    .Q(\cpu.ex.r_wb_addr[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_swapsp$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1890),
    .D(_01025_),
    .Q_N(_14855_),
    .Q(\cpu.ex.r_wb_swapsp ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_valid$_DFF_P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1891),
    .D(_00054_),
    .Q_N(_00234_),
    .Q(\cpu.ex.r_wb_valid ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[0]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1892),
    .D(_01026_),
    .Q_N(_00202_),
    .Q(\cpu.dcache.wdata[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[10]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1893),
    .D(_01027_),
    .Q_N(_14185_),
    .Q(\cpu.dcache.wdata[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[11]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1894),
    .D(_01028_),
    .Q_N(_14184_),
    .Q(\cpu.dcache.wdata[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[12]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1895),
    .D(_01029_),
    .Q_N(_14183_),
    .Q(\cpu.dcache.wdata[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[13]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1896),
    .D(_01030_),
    .Q_N(_14182_),
    .Q(\cpu.dcache.wdata[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[14]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1897),
    .D(_01031_),
    .Q_N(_14181_),
    .Q(\cpu.dcache.wdata[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[15]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1898),
    .D(_01032_),
    .Q_N(_14180_),
    .Q(\cpu.dcache.wdata[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[1]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1899),
    .D(_01033_),
    .Q_N(_00162_),
    .Q(\cpu.dcache.wdata[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[2]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1900),
    .D(_01034_),
    .Q_N(_00163_),
    .Q(\cpu.dcache.wdata[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[3]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1901),
    .D(_01035_),
    .Q_N(_00266_),
    .Q(\cpu.dcache.wdata[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[4]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1902),
    .D(_01036_),
    .Q_N(_00164_),
    .Q(\cpu.dcache.wdata[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[5]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1903),
    .D(_01037_),
    .Q_N(_00165_),
    .Q(\cpu.dcache.wdata[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[6]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1904),
    .D(_01038_),
    .Q_N(_00166_),
    .Q(\cpu.dcache.wdata[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[7]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1905),
    .D(_01039_),
    .Q_N(_00260_),
    .Q(\cpu.dcache.wdata[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[8]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1906),
    .D(_01040_),
    .Q_N(_14179_),
    .Q(\cpu.dcache.wdata[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[9]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1907),
    .D(_01041_),
    .Q_N(_14178_),
    .Q(\cpu.dcache.wdata[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wmask[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1908),
    .D(_01042_),
    .Q_N(_14177_),
    .Q(\cpu.ex.r_wmask[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wmask[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1909),
    .D(_01043_),
    .Q_N(_14176_),
    .Q(\cpu.ex.r_wmask[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[0]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1910),
    .D(_01044_),
    .Q_N(_00267_),
    .Q(\cpu.ex.mmu_read[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[1]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1911),
    .D(_01045_),
    .Q_N(_14175_),
    .Q(\cpu.ex.mmu_read[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[2]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1912),
    .D(_01046_),
    .Q_N(_00172_),
    .Q(\cpu.ex.mmu_read[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[3]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1913),
    .D(_01047_),
    .Q_N(_14174_),
    .Q(\cpu.ex.mmu_read[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_ins$_SDFFE_PN0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1914),
    .D(_01048_),
    .Q_N(_00233_),
    .Q(\cpu.ex.mmu_read[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_sup$_SDFFE_PN0P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1915),
    .D(_01049_),
    .Q_N(_14173_),
    .Q(\cpu.ex.mmu_read[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_type$_SDFFE_PN0P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1916),
    .D(_01050_),
    .Q_N(_14172_),
    .Q(\cpu.ex.mmu_read[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1917),
    .D(_01051_),
    .Q_N(_14171_),
    .Q(\cpu.genblk1.mmu.r_valid_d[0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1918),
    .D(_01052_),
    .Q_N(_14170_),
    .Q(\cpu.genblk1.mmu.r_valid_d[10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1919),
    .D(_01053_),
    .Q_N(_14169_),
    .Q(\cpu.genblk1.mmu.r_valid_d[11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1920),
    .D(_01054_),
    .Q_N(_14168_),
    .Q(\cpu.genblk1.mmu.r_valid_d[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1921),
    .D(_01055_),
    .Q_N(_14167_),
    .Q(\cpu.genblk1.mmu.r_valid_d[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1922),
    .D(_01056_),
    .Q_N(_14166_),
    .Q(\cpu.genblk1.mmu.r_valid_d[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1923),
    .D(_01057_),
    .Q_N(_14165_),
    .Q(\cpu.genblk1.mmu.r_valid_d[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1924),
    .D(_01058_),
    .Q_N(_14164_),
    .Q(\cpu.genblk1.mmu.r_valid_d[16] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1925),
    .D(_01059_),
    .Q_N(_14163_),
    .Q(\cpu.genblk1.mmu.r_valid_d[17] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1926),
    .D(_01060_),
    .Q_N(_14162_),
    .Q(\cpu.genblk1.mmu.r_valid_d[18] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1927),
    .D(_01061_),
    .Q_N(_14161_),
    .Q(\cpu.genblk1.mmu.r_valid_d[19] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1928),
    .D(_01062_),
    .Q_N(_14160_),
    .Q(\cpu.genblk1.mmu.r_valid_d[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1929),
    .D(_01063_),
    .Q_N(_14159_),
    .Q(\cpu.genblk1.mmu.r_valid_d[20] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1930),
    .D(_01064_),
    .Q_N(_14158_),
    .Q(\cpu.genblk1.mmu.r_valid_d[21] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1931),
    .D(_01065_),
    .Q_N(_14157_),
    .Q(\cpu.genblk1.mmu.r_valid_d[22] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1932),
    .D(_01066_),
    .Q_N(_14156_),
    .Q(\cpu.genblk1.mmu.r_valid_d[23] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1933),
    .D(_01067_),
    .Q_N(_14155_),
    .Q(\cpu.genblk1.mmu.r_valid_d[24] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1934),
    .D(_01068_),
    .Q_N(_14154_),
    .Q(\cpu.genblk1.mmu.r_valid_d[25] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1935),
    .D(_01069_),
    .Q_N(_14153_),
    .Q(\cpu.genblk1.mmu.r_valid_d[26] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1936),
    .D(_01070_),
    .Q_N(_14152_),
    .Q(\cpu.genblk1.mmu.r_valid_d[27] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1937),
    .D(_01071_),
    .Q_N(_14151_),
    .Q(\cpu.genblk1.mmu.r_valid_d[28] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1938),
    .D(_01072_),
    .Q_N(_14150_),
    .Q(\cpu.genblk1.mmu.r_valid_d[29] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1939),
    .D(_01073_),
    .Q_N(_14149_),
    .Q(\cpu.genblk1.mmu.r_valid_d[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1940),
    .D(_01074_),
    .Q_N(_14148_),
    .Q(\cpu.genblk1.mmu.r_valid_d[30] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1941),
    .D(_01075_),
    .Q_N(_14147_),
    .Q(\cpu.genblk1.mmu.r_valid_d[31] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1942),
    .D(_01076_),
    .Q_N(_14146_),
    .Q(\cpu.genblk1.mmu.r_valid_d[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1943),
    .D(_01077_),
    .Q_N(_14145_),
    .Q(\cpu.genblk1.mmu.r_valid_d[4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1944),
    .D(_01078_),
    .Q_N(_14144_),
    .Q(\cpu.genblk1.mmu.r_valid_d[5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1945),
    .D(_01079_),
    .Q_N(_14143_),
    .Q(\cpu.genblk1.mmu.r_valid_d[6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1946),
    .D(_01080_),
    .Q_N(_14142_),
    .Q(\cpu.genblk1.mmu.r_valid_d[7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1947),
    .D(_01081_),
    .Q_N(_14141_),
    .Q(\cpu.genblk1.mmu.r_valid_d[8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1948),
    .D(_01082_),
    .Q_N(_14140_),
    .Q(\cpu.genblk1.mmu.r_valid_d[9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1949),
    .D(_01083_),
    .Q_N(_14139_),
    .Q(\cpu.genblk1.mmu.r_valid_i[0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1950),
    .D(_01084_),
    .Q_N(_14138_),
    .Q(\cpu.genblk1.mmu.r_valid_i[10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1951),
    .D(_01085_),
    .Q_N(_14137_),
    .Q(\cpu.genblk1.mmu.r_valid_i[11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1952),
    .D(_01086_),
    .Q_N(_14136_),
    .Q(\cpu.genblk1.mmu.r_valid_i[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1953),
    .D(_01087_),
    .Q_N(_14135_),
    .Q(\cpu.genblk1.mmu.r_valid_i[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1954),
    .D(_01088_),
    .Q_N(_14134_),
    .Q(\cpu.genblk1.mmu.r_valid_i[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1955),
    .D(_01089_),
    .Q_N(_14133_),
    .Q(\cpu.genblk1.mmu.r_valid_i[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1956),
    .D(_01090_),
    .Q_N(_14132_),
    .Q(\cpu.genblk1.mmu.r_valid_i[16] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1957),
    .D(_01091_),
    .Q_N(_14131_),
    .Q(\cpu.genblk1.mmu.r_valid_i[17] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1958),
    .D(_01092_),
    .Q_N(_14130_),
    .Q(\cpu.genblk1.mmu.r_valid_i[18] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1959),
    .D(_01093_),
    .Q_N(_14129_),
    .Q(\cpu.genblk1.mmu.r_valid_i[19] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1960),
    .D(_01094_),
    .Q_N(_14128_),
    .Q(\cpu.genblk1.mmu.r_valid_i[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1961),
    .D(_01095_),
    .Q_N(_14127_),
    .Q(\cpu.genblk1.mmu.r_valid_i[20] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1962),
    .D(_01096_),
    .Q_N(_14126_),
    .Q(\cpu.genblk1.mmu.r_valid_i[21] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1963),
    .D(_01097_),
    .Q_N(_14125_),
    .Q(\cpu.genblk1.mmu.r_valid_i[22] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1964),
    .D(_01098_),
    .Q_N(_14124_),
    .Q(\cpu.genblk1.mmu.r_valid_i[23] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1965),
    .D(_01099_),
    .Q_N(_14123_),
    .Q(\cpu.genblk1.mmu.r_valid_i[24] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1966),
    .D(_01100_),
    .Q_N(_14122_),
    .Q(\cpu.genblk1.mmu.r_valid_i[25] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1967),
    .D(_01101_),
    .Q_N(_14121_),
    .Q(\cpu.genblk1.mmu.r_valid_i[26] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1968),
    .D(_01102_),
    .Q_N(_14120_),
    .Q(\cpu.genblk1.mmu.r_valid_i[27] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1969),
    .D(_01103_),
    .Q_N(_14119_),
    .Q(\cpu.genblk1.mmu.r_valid_i[28] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1970),
    .D(_01104_),
    .Q_N(_14118_),
    .Q(\cpu.genblk1.mmu.r_valid_i[29] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1971),
    .D(_01105_),
    .Q_N(_14117_),
    .Q(\cpu.genblk1.mmu.r_valid_i[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1972),
    .D(_01106_),
    .Q_N(_14116_),
    .Q(\cpu.genblk1.mmu.r_valid_i[30] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1973),
    .D(_01107_),
    .Q_N(_14115_),
    .Q(\cpu.genblk1.mmu.r_valid_i[31] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1974),
    .D(_01108_),
    .Q_N(_14114_),
    .Q(\cpu.genblk1.mmu.r_valid_i[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1975),
    .D(_01109_),
    .Q_N(_14113_),
    .Q(\cpu.genblk1.mmu.r_valid_i[4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1976),
    .D(_01110_),
    .Q_N(_14112_),
    .Q(\cpu.genblk1.mmu.r_valid_i[5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1977),
    .D(_01111_),
    .Q_N(_14111_),
    .Q(\cpu.genblk1.mmu.r_valid_i[6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1978),
    .D(_01112_),
    .Q_N(_14110_),
    .Q(\cpu.genblk1.mmu.r_valid_i[7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1979),
    .D(_01113_),
    .Q_N(_14109_),
    .Q(\cpu.genblk1.mmu.r_valid_i[8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1980),
    .D(_01114_),
    .Q_N(_14108_),
    .Q(\cpu.genblk1.mmu.r_valid_i[9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1981),
    .D(_01115_),
    .Q_N(_14107_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1982),
    .D(_01116_),
    .Q_N(_14106_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1983),
    .D(_01117_),
    .Q_N(_14105_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1984),
    .D(_01118_),
    .Q_N(_14104_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1985),
    .D(_01119_),
    .Q_N(_14103_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1986),
    .D(_01120_),
    .Q_N(_14102_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1987),
    .D(_01121_),
    .Q_N(_14101_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1988),
    .D(_01122_),
    .Q_N(_14100_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1989),
    .D(_01123_),
    .Q_N(_14099_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1990),
    .D(_01124_),
    .Q_N(_14098_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1991),
    .D(_01125_),
    .Q_N(_14097_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1992),
    .D(_01126_),
    .Q_N(_14096_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][0]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1993),
    .D(_01127_),
    .Q_N(_14095_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][10]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1994),
    .D(_01128_),
    .Q_N(_14094_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][11]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1995),
    .D(_01129_),
    .Q_N(_14093_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][1]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1996),
    .D(_01130_),
    .Q_N(_14092_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][2]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1997),
    .D(_01131_),
    .Q_N(_14091_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][3]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1998),
    .D(_01132_),
    .Q_N(_14090_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][4]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1999),
    .D(_01133_),
    .Q_N(_14089_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][5]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2000),
    .D(_01134_),
    .Q_N(_14088_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][6]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2001),
    .D(_01135_),
    .Q_N(_14087_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][7]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2002),
    .D(_01136_),
    .Q_N(_14086_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][8]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2003),
    .D(_01137_),
    .Q_N(_14085_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][9]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2004),
    .D(_01138_),
    .Q_N(_14084_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][0]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2005),
    .D(_01139_),
    .Q_N(_14083_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][10]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2006),
    .D(_01140_),
    .Q_N(_14082_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][11]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2007),
    .D(_01141_),
    .Q_N(_14081_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][1]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2008),
    .D(_01142_),
    .Q_N(_14080_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][2]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2009),
    .D(_01143_),
    .Q_N(_14079_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][3]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2010),
    .D(_01144_),
    .Q_N(_14078_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][4]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2011),
    .D(_01145_),
    .Q_N(_14077_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][5]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2012),
    .D(_01146_),
    .Q_N(_14076_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][6]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2013),
    .D(_01147_),
    .Q_N(_14075_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][7]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2014),
    .D(_01148_),
    .Q_N(_14074_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][8]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2015),
    .D(_01149_),
    .Q_N(_14073_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][9]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2016),
    .D(_01150_),
    .Q_N(_14072_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][0]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2017),
    .D(_01151_),
    .Q_N(_14071_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][10]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2018),
    .D(_01152_),
    .Q_N(_14070_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][11]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2019),
    .D(_01153_),
    .Q_N(_14069_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][1]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2020),
    .D(_01154_),
    .Q_N(_14068_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][2]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2021),
    .D(_01155_),
    .Q_N(_14067_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][3]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2022),
    .D(_01156_),
    .Q_N(_14066_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][4]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2023),
    .D(_01157_),
    .Q_N(_14065_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][5]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2024),
    .D(_01158_),
    .Q_N(_14064_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][6]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2025),
    .D(_01159_),
    .Q_N(_14063_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][7]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2026),
    .D(_01160_),
    .Q_N(_14062_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][8]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2027),
    .D(_01161_),
    .Q_N(_14061_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][9]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2028),
    .D(_01162_),
    .Q_N(_14060_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][0]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2029),
    .D(_01163_),
    .Q_N(_14059_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][10]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2030),
    .D(_01164_),
    .Q_N(_14058_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][11]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2031),
    .D(_01165_),
    .Q_N(_14057_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][1]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2032),
    .D(_01166_),
    .Q_N(_14056_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][2]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2033),
    .D(_01167_),
    .Q_N(_14055_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][3]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2034),
    .D(_01168_),
    .Q_N(_14054_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][4]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2035),
    .D(_01169_),
    .Q_N(_14053_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][5]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2036),
    .D(_01170_),
    .Q_N(_14052_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][6]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2037),
    .D(_01171_),
    .Q_N(_14051_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][7]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2038),
    .D(_01172_),
    .Q_N(_14050_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][8]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2039),
    .D(_01173_),
    .Q_N(_14049_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][9]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2040),
    .D(_01174_),
    .Q_N(_14048_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][0]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2041),
    .D(_01175_),
    .Q_N(_14047_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][10]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2042),
    .D(_01176_),
    .Q_N(_14046_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][11]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2043),
    .D(_01177_),
    .Q_N(_14045_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][1]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2044),
    .D(_01178_),
    .Q_N(_14044_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][2]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2045),
    .D(_01179_),
    .Q_N(_14043_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][3]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2046),
    .D(_01180_),
    .Q_N(_14042_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][4]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2047),
    .D(_01181_),
    .Q_N(_14041_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][5]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2048),
    .D(_01182_),
    .Q_N(_14040_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][6]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2049),
    .D(_01183_),
    .Q_N(_14039_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][7]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2050),
    .D(_01184_),
    .Q_N(_14038_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][8]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2051),
    .D(_01185_),
    .Q_N(_14037_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][9]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2052),
    .D(_01186_),
    .Q_N(_14036_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][0]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2053),
    .D(_01187_),
    .Q_N(_14035_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][10]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2054),
    .D(_01188_),
    .Q_N(_14034_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][11]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2055),
    .D(_01189_),
    .Q_N(_14033_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][1]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2056),
    .D(_01190_),
    .Q_N(_14032_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][2]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2057),
    .D(_01191_),
    .Q_N(_14031_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][3]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2058),
    .D(_01192_),
    .Q_N(_14030_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][4]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2059),
    .D(_01193_),
    .Q_N(_14029_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][5]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2060),
    .D(_01194_),
    .Q_N(_14028_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][6]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2061),
    .D(_01195_),
    .Q_N(_14027_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][7]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2062),
    .D(_01196_),
    .Q_N(_14026_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][8]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2063),
    .D(_01197_),
    .Q_N(_14025_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][9]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2064),
    .D(_01198_),
    .Q_N(_14024_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][0]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2065),
    .D(_01199_),
    .Q_N(_14023_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][10]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2066),
    .D(_01200_),
    .Q_N(_14022_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][11]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2067),
    .D(_01201_),
    .Q_N(_14021_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][1]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2068),
    .D(_01202_),
    .Q_N(_14020_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][2]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2069),
    .D(_01203_),
    .Q_N(_14019_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][3]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2070),
    .D(_01204_),
    .Q_N(_14018_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][4]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2071),
    .D(_01205_),
    .Q_N(_14017_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][5]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2072),
    .D(_01206_),
    .Q_N(_14016_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][6]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2073),
    .D(_01207_),
    .Q_N(_14015_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][7]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2074),
    .D(_01208_),
    .Q_N(_14014_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][8]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2075),
    .D(_01209_),
    .Q_N(_14013_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][9]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2076),
    .D(_01210_),
    .Q_N(_14012_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][0]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2077),
    .D(_01211_),
    .Q_N(_14011_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][10]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2078),
    .D(_01212_),
    .Q_N(_14010_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][11]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2079),
    .D(_01213_),
    .Q_N(_14009_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][1]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2080),
    .D(_01214_),
    .Q_N(_14008_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][2]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2081),
    .D(_01215_),
    .Q_N(_14007_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][3]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2082),
    .D(_01216_),
    .Q_N(_14006_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][4]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2083),
    .D(_01217_),
    .Q_N(_14005_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][5]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2084),
    .D(_01218_),
    .Q_N(_14004_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][6]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2085),
    .D(_01219_),
    .Q_N(_14003_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][7]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2086),
    .D(_01220_),
    .Q_N(_14002_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][8]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2087),
    .D(_01221_),
    .Q_N(_14001_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][9]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2088),
    .D(_01222_),
    .Q_N(_14000_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][0]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2089),
    .D(_01223_),
    .Q_N(_13999_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][10]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2090),
    .D(_01224_),
    .Q_N(_13998_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][11]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2091),
    .D(_01225_),
    .Q_N(_13997_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][1]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2092),
    .D(_01226_),
    .Q_N(_13996_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][2]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2093),
    .D(_01227_),
    .Q_N(_13995_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][3]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2094),
    .D(_01228_),
    .Q_N(_13994_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][4]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2095),
    .D(_01229_),
    .Q_N(_13993_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][5]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2096),
    .D(_01230_),
    .Q_N(_13992_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][6]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2097),
    .D(_01231_),
    .Q_N(_13991_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][7]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2098),
    .D(_01232_),
    .Q_N(_13990_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][8]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2099),
    .D(_01233_),
    .Q_N(_13989_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][9]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2100),
    .D(_01234_),
    .Q_N(_13988_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][0]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2101),
    .D(_01235_),
    .Q_N(_13987_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][10]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2102),
    .D(_01236_),
    .Q_N(_13986_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][11]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2103),
    .D(_01237_),
    .Q_N(_13985_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][1]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2104),
    .D(_01238_),
    .Q_N(_13984_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][2]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2105),
    .D(_01239_),
    .Q_N(_13983_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][3]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2106),
    .D(_01240_),
    .Q_N(_13982_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][4]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2107),
    .D(_01241_),
    .Q_N(_13981_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][5]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2108),
    .D(_01242_),
    .Q_N(_13980_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][6]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2109),
    .D(_01243_),
    .Q_N(_13979_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][7]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2110),
    .D(_01244_),
    .Q_N(_13978_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][8]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2111),
    .D(_01245_),
    .Q_N(_13977_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][9]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2112),
    .D(_01246_),
    .Q_N(_13976_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2113),
    .D(_01247_),
    .Q_N(_13975_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2114),
    .D(_01248_),
    .Q_N(_13974_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2115),
    .D(_01249_),
    .Q_N(_13973_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2116),
    .D(_01250_),
    .Q_N(_13972_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2117),
    .D(_01251_),
    .Q_N(_13971_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2118),
    .D(_01252_),
    .Q_N(_13970_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2119),
    .D(_01253_),
    .Q_N(_13969_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2120),
    .D(_01254_),
    .Q_N(_13968_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2121),
    .D(_01255_),
    .Q_N(_13967_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2122),
    .D(_01256_),
    .Q_N(_13966_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2123),
    .D(_01257_),
    .Q_N(_13965_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2124),
    .D(_01258_),
    .Q_N(_13964_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][0]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2125),
    .D(_01259_),
    .Q_N(_13963_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][10]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2126),
    .D(_01260_),
    .Q_N(_13962_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][11]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2127),
    .D(_01261_),
    .Q_N(_13961_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][1]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2128),
    .D(_01262_),
    .Q_N(_13960_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][2]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2129),
    .D(_01263_),
    .Q_N(_13959_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][3]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2130),
    .D(_01264_),
    .Q_N(_13958_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][4]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2131),
    .D(_01265_),
    .Q_N(_13957_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][5]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2132),
    .D(_01266_),
    .Q_N(_13956_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][6]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2133),
    .D(_01267_),
    .Q_N(_13955_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][7]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2134),
    .D(_01268_),
    .Q_N(_13954_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][8]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2135),
    .D(_01269_),
    .Q_N(_13953_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][9]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2136),
    .D(_01270_),
    .Q_N(_13952_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][0]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2137),
    .D(_01271_),
    .Q_N(_13951_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][10]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2138),
    .D(_01272_),
    .Q_N(_13950_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][11]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2139),
    .D(_01273_),
    .Q_N(_13949_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][1]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2140),
    .D(_01274_),
    .Q_N(_13948_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][2]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2141),
    .D(_01275_),
    .Q_N(_13947_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][3]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2142),
    .D(_01276_),
    .Q_N(_13946_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][4]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2143),
    .D(_01277_),
    .Q_N(_13945_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][5]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2144),
    .D(_01278_),
    .Q_N(_13944_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][6]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2145),
    .D(_01279_),
    .Q_N(_13943_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][7]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2146),
    .D(_01280_),
    .Q_N(_13942_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][8]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2147),
    .D(_01281_),
    .Q_N(_13941_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][9]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2148),
    .D(_01282_),
    .Q_N(_13940_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][0]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2149),
    .D(_01283_),
    .Q_N(_13939_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][10]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2150),
    .D(_01284_),
    .Q_N(_13938_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][11]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2151),
    .D(_01285_),
    .Q_N(_13937_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][1]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2152),
    .D(_01286_),
    .Q_N(_13936_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][2]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2153),
    .D(_01287_),
    .Q_N(_13935_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][3]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2154),
    .D(_01288_),
    .Q_N(_13934_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][4]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2155),
    .D(_01289_),
    .Q_N(_13933_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][5]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2156),
    .D(_01290_),
    .Q_N(_13932_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][6]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2157),
    .D(_01291_),
    .Q_N(_13931_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][7]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2158),
    .D(_01292_),
    .Q_N(_13930_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][8]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2159),
    .D(_01293_),
    .Q_N(_13929_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][9]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2160),
    .D(_01294_),
    .Q_N(_13928_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][0]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2161),
    .D(_01295_),
    .Q_N(_13927_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][10]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2162),
    .D(_01296_),
    .Q_N(_13926_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][11]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2163),
    .D(_01297_),
    .Q_N(_13925_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][1]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2164),
    .D(_01298_),
    .Q_N(_13924_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][2]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2165),
    .D(_01299_),
    .Q_N(_13923_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][3]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2166),
    .D(_01300_),
    .Q_N(_13922_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][4]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2167),
    .D(_01301_),
    .Q_N(_13921_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][5]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2168),
    .D(_01302_),
    .Q_N(_13920_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][6]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2169),
    .D(_01303_),
    .Q_N(_13919_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][7]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2170),
    .D(_01304_),
    .Q_N(_13918_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][8]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2171),
    .D(_01305_),
    .Q_N(_13917_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][9]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2172),
    .D(_01306_),
    .Q_N(_13916_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][0]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2173),
    .D(_01307_),
    .Q_N(_13915_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][10]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2174),
    .D(_01308_),
    .Q_N(_13914_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][11]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2175),
    .D(_01309_),
    .Q_N(_13913_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][1]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2176),
    .D(_01310_),
    .Q_N(_13912_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][2]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2177),
    .D(_01311_),
    .Q_N(_13911_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][3]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2178),
    .D(_01312_),
    .Q_N(_13910_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][4]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2179),
    .D(_01313_),
    .Q_N(_13909_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][5]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2180),
    .D(_01314_),
    .Q_N(_13908_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][6]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2181),
    .D(_01315_),
    .Q_N(_13907_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][7]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2182),
    .D(_01316_),
    .Q_N(_13906_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][8]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2183),
    .D(_01317_),
    .Q_N(_13905_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][9]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2184),
    .D(_01318_),
    .Q_N(_13904_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][0]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2185),
    .D(_01319_),
    .Q_N(_13903_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][10]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2186),
    .D(_01320_),
    .Q_N(_13902_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][11]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2187),
    .D(_01321_),
    .Q_N(_13901_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][1]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2188),
    .D(_01322_),
    .Q_N(_13900_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][2]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2189),
    .D(_01323_),
    .Q_N(_13899_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][3]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2190),
    .D(_01324_),
    .Q_N(_13898_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][4]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2191),
    .D(_01325_),
    .Q_N(_13897_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][5]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2192),
    .D(_01326_),
    .Q_N(_13896_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][6]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2193),
    .D(_01327_),
    .Q_N(_13895_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][7]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2194),
    .D(_01328_),
    .Q_N(_13894_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][8]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2195),
    .D(_01329_),
    .Q_N(_13893_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][9]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2196),
    .D(_01330_),
    .Q_N(_13892_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][0]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2197),
    .D(_01331_),
    .Q_N(_13891_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][10]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2198),
    .D(_01332_),
    .Q_N(_13890_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][11]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2199),
    .D(_01333_),
    .Q_N(_13889_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][1]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2200),
    .D(_01334_),
    .Q_N(_13888_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][2]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2201),
    .D(_01335_),
    .Q_N(_13887_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][3]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2202),
    .D(_01336_),
    .Q_N(_13886_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][4]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2203),
    .D(_01337_),
    .Q_N(_13885_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][5]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2204),
    .D(_01338_),
    .Q_N(_13884_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][6]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2205),
    .D(_01339_),
    .Q_N(_13883_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][7]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2206),
    .D(_01340_),
    .Q_N(_13882_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][8]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2207),
    .D(_01341_),
    .Q_N(_13881_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][9]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2208),
    .D(_01342_),
    .Q_N(_13880_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][0]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2209),
    .D(_01343_),
    .Q_N(_13879_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][10]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2210),
    .D(_01344_),
    .Q_N(_13878_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][11]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2211),
    .D(_01345_),
    .Q_N(_13877_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][1]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2212),
    .D(_01346_),
    .Q_N(_13876_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][2]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2213),
    .D(_01347_),
    .Q_N(_13875_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][3]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2214),
    .D(_01348_),
    .Q_N(_13874_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][4]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2215),
    .D(_01349_),
    .Q_N(_13873_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][5]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2216),
    .D(_01350_),
    .Q_N(_13872_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][6]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2217),
    .D(_01351_),
    .Q_N(_13871_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][7]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2218),
    .D(_01352_),
    .Q_N(_13870_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][8]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2219),
    .D(_01353_),
    .Q_N(_13869_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][9]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2220),
    .D(_01354_),
    .Q_N(_13868_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][0]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2221),
    .D(_01355_),
    .Q_N(_13867_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][10]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2222),
    .D(_01356_),
    .Q_N(_13866_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][11]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2223),
    .D(_01357_),
    .Q_N(_13865_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][1]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2224),
    .D(_01358_),
    .Q_N(_13864_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][2]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2225),
    .D(_01359_),
    .Q_N(_13863_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][3]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2226),
    .D(_01360_),
    .Q_N(_13862_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][4]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2227),
    .D(_01361_),
    .Q_N(_13861_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][5]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2228),
    .D(_01362_),
    .Q_N(_13860_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][6]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2229),
    .D(_01363_),
    .Q_N(_13859_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][7]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2230),
    .D(_01364_),
    .Q_N(_13858_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][8]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2231),
    .D(_01365_),
    .Q_N(_13857_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][9]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2232),
    .D(_01366_),
    .Q_N(_13856_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][0]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2233),
    .D(_01367_),
    .Q_N(_13855_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][10]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2234),
    .D(_01368_),
    .Q_N(_13854_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][11]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2235),
    .D(_01369_),
    .Q_N(_13853_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][1]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2236),
    .D(_01370_),
    .Q_N(_13852_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][2]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2237),
    .D(_01371_),
    .Q_N(_13851_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][3]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2238),
    .D(_01372_),
    .Q_N(_13850_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][4]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2239),
    .D(_01373_),
    .Q_N(_13849_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][5]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2240),
    .D(_01374_),
    .Q_N(_13848_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][6]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2241),
    .D(_01375_),
    .Q_N(_13847_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][7]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2242),
    .D(_01376_),
    .Q_N(_13846_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][8]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2243),
    .D(_01377_),
    .Q_N(_13845_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][9]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2244),
    .D(_01378_),
    .Q_N(_13844_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2245),
    .D(_01379_),
    .Q_N(_13843_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2246),
    .D(_01380_),
    .Q_N(_13842_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2247),
    .D(_01381_),
    .Q_N(_13841_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2248),
    .D(_01382_),
    .Q_N(_13840_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2249),
    .D(_01383_),
    .Q_N(_13839_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2250),
    .D(_01384_),
    .Q_N(_13838_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2251),
    .D(_01385_),
    .Q_N(_13837_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2252),
    .D(_01386_),
    .Q_N(_13836_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2253),
    .D(_01387_),
    .Q_N(_13835_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2254),
    .D(_01388_),
    .Q_N(_13834_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2255),
    .D(_01389_),
    .Q_N(_13833_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2256),
    .D(_01390_),
    .Q_N(_13832_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][0]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2257),
    .D(_01391_),
    .Q_N(_13831_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][10]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2258),
    .D(_01392_),
    .Q_N(_13830_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][11]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2259),
    .D(_01393_),
    .Q_N(_13829_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][1]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2260),
    .D(_01394_),
    .Q_N(_13828_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][2]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2261),
    .D(_01395_),
    .Q_N(_13827_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][3]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2262),
    .D(_01396_),
    .Q_N(_13826_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][4]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2263),
    .D(_01397_),
    .Q_N(_13825_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][5]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2264),
    .D(_01398_),
    .Q_N(_13824_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][6]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2265),
    .D(_01399_),
    .Q_N(_13823_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][7]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2266),
    .D(_01400_),
    .Q_N(_13822_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][8]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2267),
    .D(_01401_),
    .Q_N(_13821_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][9]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2268),
    .D(_01402_),
    .Q_N(_13820_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][0]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2269),
    .D(_01403_),
    .Q_N(_13819_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][10]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2270),
    .D(_01404_),
    .Q_N(_13818_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][11]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2271),
    .D(_01405_),
    .Q_N(_13817_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][1]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2272),
    .D(_01406_),
    .Q_N(_13816_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][2]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2273),
    .D(_01407_),
    .Q_N(_13815_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][3]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2274),
    .D(_01408_),
    .Q_N(_13814_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][4]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2275),
    .D(_01409_),
    .Q_N(_13813_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][5]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2276),
    .D(_01410_),
    .Q_N(_13812_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][6]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2277),
    .D(_01411_),
    .Q_N(_13811_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][7]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2278),
    .D(_01412_),
    .Q_N(_13810_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][8]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2279),
    .D(_01413_),
    .Q_N(_13809_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][9]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2280),
    .D(_01414_),
    .Q_N(_13808_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2281),
    .D(_01415_),
    .Q_N(_13807_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2282),
    .D(_01416_),
    .Q_N(_13806_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2283),
    .D(_01417_),
    .Q_N(_13805_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2284),
    .D(_01418_),
    .Q_N(_13804_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2285),
    .D(_01419_),
    .Q_N(_13803_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2286),
    .D(_01420_),
    .Q_N(_13802_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2287),
    .D(_01421_),
    .Q_N(_13801_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2288),
    .D(_01422_),
    .Q_N(_13800_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2289),
    .D(_01423_),
    .Q_N(_13799_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2290),
    .D(_01424_),
    .Q_N(_13798_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2291),
    .D(_01425_),
    .Q_N(_13797_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2292),
    .D(_01426_),
    .Q_N(_13796_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2293),
    .D(_01427_),
    .Q_N(_13795_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2294),
    .D(_01428_),
    .Q_N(_13794_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2295),
    .D(_01429_),
    .Q_N(_13793_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2296),
    .D(_01430_),
    .Q_N(_13792_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2297),
    .D(_01431_),
    .Q_N(_13791_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2298),
    .D(_01432_),
    .Q_N(_13790_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2299),
    .D(_01433_),
    .Q_N(_13789_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2300),
    .D(_01434_),
    .Q_N(_13788_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2301),
    .D(_01435_),
    .Q_N(_13787_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2302),
    .D(_01436_),
    .Q_N(_13786_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2303),
    .D(_01437_),
    .Q_N(_13785_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2304),
    .D(_01438_),
    .Q_N(_13784_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2305),
    .D(_01439_),
    .Q_N(_13783_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2306),
    .D(_01440_),
    .Q_N(_13782_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2307),
    .D(_01441_),
    .Q_N(_13781_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2308),
    .D(_01442_),
    .Q_N(_13780_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2309),
    .D(_01443_),
    .Q_N(_13779_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2310),
    .D(_01444_),
    .Q_N(_13778_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2311),
    .D(_01445_),
    .Q_N(_13777_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2312),
    .D(_01446_),
    .Q_N(_13776_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2313),
    .D(_01447_),
    .Q_N(_13775_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2314),
    .D(_01448_),
    .Q_N(_13774_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2315),
    .D(_01449_),
    .Q_N(_13773_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2316),
    .D(_01450_),
    .Q_N(_13772_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2317),
    .D(_01451_),
    .Q_N(_13771_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2318),
    .D(_01452_),
    .Q_N(_13770_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2319),
    .D(_01453_),
    .Q_N(_13769_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2320),
    .D(_01454_),
    .Q_N(_13768_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2321),
    .D(_01455_),
    .Q_N(_13767_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2322),
    .D(_01456_),
    .Q_N(_13766_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2323),
    .D(_01457_),
    .Q_N(_13765_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2324),
    .D(_01458_),
    .Q_N(_13764_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2325),
    .D(_01459_),
    .Q_N(_13763_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2326),
    .D(_01460_),
    .Q_N(_13762_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2327),
    .D(_01461_),
    .Q_N(_13761_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2328),
    .D(_01462_),
    .Q_N(_13760_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2329),
    .D(_01463_),
    .Q_N(_13759_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2330),
    .D(_01464_),
    .Q_N(_13758_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2331),
    .D(_01465_),
    .Q_N(_13757_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2332),
    .D(_01466_),
    .Q_N(_13756_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2333),
    .D(_01467_),
    .Q_N(_13755_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2334),
    .D(_01468_),
    .Q_N(_13754_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2335),
    .D(_01469_),
    .Q_N(_13753_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2336),
    .D(_01470_),
    .Q_N(_13752_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2337),
    .D(_01471_),
    .Q_N(_13751_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2338),
    .D(_01472_),
    .Q_N(_13750_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2339),
    .D(_01473_),
    .Q_N(_13749_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2340),
    .D(_01474_),
    .Q_N(_13748_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][0]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2341),
    .D(_01475_),
    .Q_N(_13747_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][10]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2342),
    .D(_01476_),
    .Q_N(_13746_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][11]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2343),
    .D(_01477_),
    .Q_N(_13745_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][1]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2344),
    .D(_01478_),
    .Q_N(_13744_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][2]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2345),
    .D(_01479_),
    .Q_N(_13743_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][3]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2346),
    .D(_01480_),
    .Q_N(_13742_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][4]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2347),
    .D(_01481_),
    .Q_N(_13741_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][5]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2348),
    .D(_01482_),
    .Q_N(_13740_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][6]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2349),
    .D(_01483_),
    .Q_N(_13739_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][7]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2350),
    .D(_01484_),
    .Q_N(_13738_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][8]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2351),
    .D(_01485_),
    .Q_N(_13737_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][9]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2352),
    .D(_01486_),
    .Q_N(_13736_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][0]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2353),
    .D(_01487_),
    .Q_N(_13735_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][10]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2354),
    .D(_01488_),
    .Q_N(_13734_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][11]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2355),
    .D(_01489_),
    .Q_N(_13733_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][1]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2356),
    .D(_01490_),
    .Q_N(_13732_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][2]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2357),
    .D(_01491_),
    .Q_N(_13731_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][3]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2358),
    .D(_01492_),
    .Q_N(_13730_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][4]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2359),
    .D(_01493_),
    .Q_N(_13729_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][5]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2360),
    .D(_01494_),
    .Q_N(_13728_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][6]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2361),
    .D(_01495_),
    .Q_N(_13727_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][7]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2362),
    .D(_01496_),
    .Q_N(_13726_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][8]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2363),
    .D(_01497_),
    .Q_N(_13725_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][9]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2364),
    .D(_01498_),
    .Q_N(_13724_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2365),
    .D(_01499_),
    .Q_N(_13723_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2366),
    .D(_01500_),
    .Q_N(_13722_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2367),
    .D(_01501_),
    .Q_N(_13721_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2368),
    .D(_01502_),
    .Q_N(_13720_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2369),
    .D(_01503_),
    .Q_N(_13719_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2370),
    .D(_01504_),
    .Q_N(_13718_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2371),
    .D(_01505_),
    .Q_N(_13717_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2372),
    .D(_01506_),
    .Q_N(_13716_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2373),
    .D(_01507_),
    .Q_N(_13715_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2374),
    .D(_01508_),
    .Q_N(_13714_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2375),
    .D(_01509_),
    .Q_N(_13713_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2376),
    .D(_01510_),
    .Q_N(_13712_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][0]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2377),
    .D(_01511_),
    .Q_N(_13711_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][10]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2378),
    .D(_01512_),
    .Q_N(_13710_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][11]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2379),
    .D(_01513_),
    .Q_N(_13709_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][1]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2380),
    .D(_01514_),
    .Q_N(_13708_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][2]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2381),
    .D(_01515_),
    .Q_N(_13707_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][3]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2382),
    .D(_01516_),
    .Q_N(_13706_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][4]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2383),
    .D(_01517_),
    .Q_N(_13705_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][5]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2384),
    .D(_01518_),
    .Q_N(_13704_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][6]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2385),
    .D(_01519_),
    .Q_N(_13703_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][7]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2386),
    .D(_01520_),
    .Q_N(_13702_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][8]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2387),
    .D(_01521_),
    .Q_N(_13701_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][9]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2388),
    .D(_01522_),
    .Q_N(_13700_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][0]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2389),
    .D(_01523_),
    .Q_N(_13699_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][10]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2390),
    .D(_01524_),
    .Q_N(_13698_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][11]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2391),
    .D(_01525_),
    .Q_N(_13697_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][1]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2392),
    .D(_01526_),
    .Q_N(_13696_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][2]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2393),
    .D(_01527_),
    .Q_N(_13695_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][3]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2394),
    .D(_01528_),
    .Q_N(_13694_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][4]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2395),
    .D(_01529_),
    .Q_N(_13693_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][5]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2396),
    .D(_01530_),
    .Q_N(_13692_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][6]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2397),
    .D(_01531_),
    .Q_N(_13691_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][7]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2398),
    .D(_01532_),
    .Q_N(_13690_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][8]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2399),
    .D(_01533_),
    .Q_N(_13689_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][9]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2400),
    .D(_01534_),
    .Q_N(_13688_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][0]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2401),
    .D(_01535_),
    .Q_N(_13687_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][10]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2402),
    .D(_01536_),
    .Q_N(_13686_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][11]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2403),
    .D(_01537_),
    .Q_N(_13685_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][1]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2404),
    .D(_01538_),
    .Q_N(_13684_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][2]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2405),
    .D(_01539_),
    .Q_N(_13683_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][3]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2406),
    .D(_01540_),
    .Q_N(_13682_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][4]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2407),
    .D(_01541_),
    .Q_N(_13681_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][5]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2408),
    .D(_01542_),
    .Q_N(_13680_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][6]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2409),
    .D(_01543_),
    .Q_N(_13679_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][7]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2410),
    .D(_01544_),
    .Q_N(_13678_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][8]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2411),
    .D(_01545_),
    .Q_N(_13677_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][9]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2412),
    .D(_01546_),
    .Q_N(_13676_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][0]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2413),
    .D(_01547_),
    .Q_N(_13675_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][10]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2414),
    .D(_01548_),
    .Q_N(_13674_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][11]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2415),
    .D(_01549_),
    .Q_N(_13673_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][1]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2416),
    .D(_01550_),
    .Q_N(_13672_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][2]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2417),
    .D(_01551_),
    .Q_N(_13671_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][3]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2418),
    .D(_01552_),
    .Q_N(_13670_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][4]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2419),
    .D(_01553_),
    .Q_N(_13669_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][5]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2420),
    .D(_01554_),
    .Q_N(_13668_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][6]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2421),
    .D(_01555_),
    .Q_N(_13667_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][7]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2422),
    .D(_01556_),
    .Q_N(_13666_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][8]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2423),
    .D(_01557_),
    .Q_N(_13665_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][9]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2424),
    .D(_01558_),
    .Q_N(_13664_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][0]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2425),
    .D(_01559_),
    .Q_N(_13663_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][10]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2426),
    .D(_01560_),
    .Q_N(_13662_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][11]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2427),
    .D(_01561_),
    .Q_N(_13661_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][1]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2428),
    .D(_01562_),
    .Q_N(_13660_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][2]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2429),
    .D(_01563_),
    .Q_N(_13659_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][3]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2430),
    .D(_01564_),
    .Q_N(_13658_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][4]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2431),
    .D(_01565_),
    .Q_N(_13657_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][5]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2432),
    .D(_01566_),
    .Q_N(_13656_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][6]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2433),
    .D(_01567_),
    .Q_N(_13655_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][7]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2434),
    .D(_01568_),
    .Q_N(_13654_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][8]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2435),
    .D(_01569_),
    .Q_N(_13653_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][9]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2436),
    .D(_01570_),
    .Q_N(_13652_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][0]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2437),
    .D(_01571_),
    .Q_N(_13651_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][10]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2438),
    .D(_01572_),
    .Q_N(_13650_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][11]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2439),
    .D(_01573_),
    .Q_N(_13649_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][1]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2440),
    .D(_01574_),
    .Q_N(_13648_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][2]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2441),
    .D(_01575_),
    .Q_N(_13647_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][3]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2442),
    .D(_01576_),
    .Q_N(_13646_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][4]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2443),
    .D(_01577_),
    .Q_N(_13645_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][5]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2444),
    .D(_01578_),
    .Q_N(_13644_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][6]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2445),
    .D(_01579_),
    .Q_N(_13643_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][7]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2446),
    .D(_01580_),
    .Q_N(_13642_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][8]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2447),
    .D(_01581_),
    .Q_N(_13641_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][9]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2448),
    .D(_01582_),
    .Q_N(_13640_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][0]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2449),
    .D(_01583_),
    .Q_N(_13639_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][10]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2450),
    .D(_01584_),
    .Q_N(_13638_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][11]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2451),
    .D(_01585_),
    .Q_N(_13637_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][1]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2452),
    .D(_01586_),
    .Q_N(_13636_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][2]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2453),
    .D(_01587_),
    .Q_N(_13635_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][3]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2454),
    .D(_01588_),
    .Q_N(_13634_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][4]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2455),
    .D(_01589_),
    .Q_N(_13633_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][5]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2456),
    .D(_01590_),
    .Q_N(_13632_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][6]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2457),
    .D(_01591_),
    .Q_N(_13631_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][7]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2458),
    .D(_01592_),
    .Q_N(_13630_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][8]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2459),
    .D(_01593_),
    .Q_N(_13629_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][9]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2460),
    .D(_01594_),
    .Q_N(_13628_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][0]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2461),
    .D(_01595_),
    .Q_N(_13627_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][10]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2462),
    .D(_01596_),
    .Q_N(_13626_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][11]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2463),
    .D(_01597_),
    .Q_N(_13625_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][1]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2464),
    .D(_01598_),
    .Q_N(_13624_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][2]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2465),
    .D(_01599_),
    .Q_N(_13623_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][3]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2466),
    .D(_01600_),
    .Q_N(_13622_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][4]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2467),
    .D(_01601_),
    .Q_N(_13621_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][5]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2468),
    .D(_01602_),
    .Q_N(_13620_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][6]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2469),
    .D(_01603_),
    .Q_N(_13619_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][7]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2470),
    .D(_01604_),
    .Q_N(_13618_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][8]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2471),
    .D(_01605_),
    .Q_N(_13617_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][9]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2472),
    .D(_01606_),
    .Q_N(_13616_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][0]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2473),
    .D(_01607_),
    .Q_N(_13615_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][10]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2474),
    .D(_01608_),
    .Q_N(_13614_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][11]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2475),
    .D(_01609_),
    .Q_N(_13613_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][1]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2476),
    .D(_01610_),
    .Q_N(_13612_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][2]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2477),
    .D(_01611_),
    .Q_N(_13611_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][3]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2478),
    .D(_01612_),
    .Q_N(_13610_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][4]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2479),
    .D(_01613_),
    .Q_N(_13609_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][5]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2480),
    .D(_01614_),
    .Q_N(_13608_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][6]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2481),
    .D(_01615_),
    .Q_N(_13607_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][7]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2482),
    .D(_01616_),
    .Q_N(_13606_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][8]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2483),
    .D(_01617_),
    .Q_N(_13605_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][9]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2484),
    .D(_01618_),
    .Q_N(_13604_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][0]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2485),
    .D(_01619_),
    .Q_N(_13603_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][10]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2486),
    .D(_01620_),
    .Q_N(_13602_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][11]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2487),
    .D(_01621_),
    .Q_N(_13601_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][1]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2488),
    .D(_01622_),
    .Q_N(_13600_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][2]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2489),
    .D(_01623_),
    .Q_N(_13599_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][3]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2490),
    .D(_01624_),
    .Q_N(_13598_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][4]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2491),
    .D(_01625_),
    .Q_N(_13597_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][5]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2492),
    .D(_01626_),
    .Q_N(_13596_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][6]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2493),
    .D(_01627_),
    .Q_N(_13595_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][7]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2494),
    .D(_01628_),
    .Q_N(_13594_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][8]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2495),
    .D(_01629_),
    .Q_N(_13593_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][9]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2496),
    .D(_01630_),
    .Q_N(_13592_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2497),
    .D(_01631_),
    .Q_N(_13591_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2498),
    .D(_01632_),
    .Q_N(_13590_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2499),
    .D(_01633_),
    .Q_N(_13589_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2500),
    .D(_01634_),
    .Q_N(_13588_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2501),
    .D(_01635_),
    .Q_N(_13587_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2502),
    .D(_01636_),
    .Q_N(_13586_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2503),
    .D(_01637_),
    .Q_N(_13585_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2504),
    .D(_01638_),
    .Q_N(_13584_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2505),
    .D(_01639_),
    .Q_N(_13583_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2506),
    .D(_01640_),
    .Q_N(_13582_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2507),
    .D(_01641_),
    .Q_N(_13581_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2508),
    .D(_01642_),
    .Q_N(_13580_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][0]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2509),
    .D(_01643_),
    .Q_N(_13579_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][10]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2510),
    .D(_01644_),
    .Q_N(_13578_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][11]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2511),
    .D(_01645_),
    .Q_N(_13577_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][1]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2512),
    .D(_01646_),
    .Q_N(_13576_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][2]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2513),
    .D(_01647_),
    .Q_N(_13575_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][3]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2514),
    .D(_01648_),
    .Q_N(_13574_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][4]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2515),
    .D(_01649_),
    .Q_N(_13573_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][5]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2516),
    .D(_01650_),
    .Q_N(_13572_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][6]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2517),
    .D(_01651_),
    .Q_N(_13571_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][7]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2518),
    .D(_01652_),
    .Q_N(_13570_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][8]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2519),
    .D(_01653_),
    .Q_N(_13569_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][9]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2520),
    .D(_01654_),
    .Q_N(_13568_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][0]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2521),
    .D(_01655_),
    .Q_N(_13567_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][10]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2522),
    .D(_01656_),
    .Q_N(_13566_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][11]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2523),
    .D(_01657_),
    .Q_N(_13565_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][1]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2524),
    .D(_01658_),
    .Q_N(_13564_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][2]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2525),
    .D(_01659_),
    .Q_N(_13563_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][3]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2526),
    .D(_01660_),
    .Q_N(_13562_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][4]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2527),
    .D(_01661_),
    .Q_N(_13561_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][5]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2528),
    .D(_01662_),
    .Q_N(_13560_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][6]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2529),
    .D(_01663_),
    .Q_N(_13559_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][7]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2530),
    .D(_01664_),
    .Q_N(_13558_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][8]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2531),
    .D(_01665_),
    .Q_N(_13557_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][9]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2532),
    .D(_01666_),
    .Q_N(_13556_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][0]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2533),
    .D(_01667_),
    .Q_N(_13555_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][10]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2534),
    .D(_01668_),
    .Q_N(_13554_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][11]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2535),
    .D(_01669_),
    .Q_N(_13553_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][1]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2536),
    .D(_01670_),
    .Q_N(_13552_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][2]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2537),
    .D(_01671_),
    .Q_N(_13551_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][3]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2538),
    .D(_01672_),
    .Q_N(_13550_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][4]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2539),
    .D(_01673_),
    .Q_N(_13549_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][5]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2540),
    .D(_01674_),
    .Q_N(_13548_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][6]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2541),
    .D(_01675_),
    .Q_N(_13547_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][7]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2542),
    .D(_01676_),
    .Q_N(_13546_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][8]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2543),
    .D(_01677_),
    .Q_N(_13545_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][9]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2544),
    .D(_01678_),
    .Q_N(_13544_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][0]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2545),
    .D(_01679_),
    .Q_N(_13543_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][10]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2546),
    .D(_01680_),
    .Q_N(_13542_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][11]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2547),
    .D(_01681_),
    .Q_N(_13541_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][1]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2548),
    .D(_01682_),
    .Q_N(_13540_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][2]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2549),
    .D(_01683_),
    .Q_N(_13539_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][3]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2550),
    .D(_01684_),
    .Q_N(_13538_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][4]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2551),
    .D(_01685_),
    .Q_N(_13537_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][5]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2552),
    .D(_01686_),
    .Q_N(_13536_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][6]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2553),
    .D(_01687_),
    .Q_N(_13535_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][7]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2554),
    .D(_01688_),
    .Q_N(_13534_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][8]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2555),
    .D(_01689_),
    .Q_N(_13533_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][9]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2556),
    .D(_01690_),
    .Q_N(_13532_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][0]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2557),
    .D(_01691_),
    .Q_N(_13531_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][10]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2558),
    .D(_01692_),
    .Q_N(_13530_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][11]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2559),
    .D(_01693_),
    .Q_N(_13529_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][1]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2560),
    .D(_01694_),
    .Q_N(_13528_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][2]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2561),
    .D(_01695_),
    .Q_N(_13527_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][3]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2562),
    .D(_01696_),
    .Q_N(_13526_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][4]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2563),
    .D(_01697_),
    .Q_N(_13525_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][5]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2564),
    .D(_01698_),
    .Q_N(_13524_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][6]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2565),
    .D(_01699_),
    .Q_N(_13523_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][7]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2566),
    .D(_01700_),
    .Q_N(_13522_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][8]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2567),
    .D(_01701_),
    .Q_N(_13521_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][9]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2568),
    .D(_01702_),
    .Q_N(_13520_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][0]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2569),
    .D(_01703_),
    .Q_N(_13519_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][10]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2570),
    .D(_01704_),
    .Q_N(_13518_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][11]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2571),
    .D(_01705_),
    .Q_N(_13517_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][1]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2572),
    .D(_01706_),
    .Q_N(_13516_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][2]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2573),
    .D(_01707_),
    .Q_N(_13515_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][3]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2574),
    .D(_01708_),
    .Q_N(_13514_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][4]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2575),
    .D(_01709_),
    .Q_N(_13513_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][5]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2576),
    .D(_01710_),
    .Q_N(_13512_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][6]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2577),
    .D(_01711_),
    .Q_N(_13511_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][7]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2578),
    .D(_01712_),
    .Q_N(_13510_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][8]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2579),
    .D(_01713_),
    .Q_N(_13509_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][9]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2580),
    .D(_01714_),
    .Q_N(_13508_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][0]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2581),
    .D(_01715_),
    .Q_N(_13507_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][10]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2582),
    .D(_01716_),
    .Q_N(_13506_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][11]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2583),
    .D(_01717_),
    .Q_N(_13505_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][1]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2584),
    .D(_01718_),
    .Q_N(_13504_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][2]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2585),
    .D(_01719_),
    .Q_N(_13503_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][3]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2586),
    .D(_01720_),
    .Q_N(_13502_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][4]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2587),
    .D(_01721_),
    .Q_N(_13501_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][5]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2588),
    .D(_01722_),
    .Q_N(_13500_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][6]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2589),
    .D(_01723_),
    .Q_N(_13499_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][7]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2590),
    .D(_01724_),
    .Q_N(_13498_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][8]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2591),
    .D(_01725_),
    .Q_N(_13497_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][9]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2592),
    .D(_01726_),
    .Q_N(_13496_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][0]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2593),
    .D(_01727_),
    .Q_N(_13495_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][10]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2594),
    .D(_01728_),
    .Q_N(_13494_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][11]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2595),
    .D(_01729_),
    .Q_N(_13493_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][1]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2596),
    .D(_01730_),
    .Q_N(_13492_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][2]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2597),
    .D(_01731_),
    .Q_N(_13491_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][3]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2598),
    .D(_01732_),
    .Q_N(_13490_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][4]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2599),
    .D(_01733_),
    .Q_N(_13489_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][5]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2600),
    .D(_01734_),
    .Q_N(_13488_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][6]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2601),
    .D(_01735_),
    .Q_N(_13487_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][7]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2602),
    .D(_01736_),
    .Q_N(_13486_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][8]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2603),
    .D(_01737_),
    .Q_N(_13485_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][9]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2604),
    .D(_01738_),
    .Q_N(_13484_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][0]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2605),
    .D(_01739_),
    .Q_N(_13483_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][10]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2606),
    .D(_01740_),
    .Q_N(_13482_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][11]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2607),
    .D(_01741_),
    .Q_N(_13481_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][1]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2608),
    .D(_01742_),
    .Q_N(_13480_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][2]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2609),
    .D(_01743_),
    .Q_N(_13479_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][3]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2610),
    .D(_01744_),
    .Q_N(_13478_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][4]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2611),
    .D(_01745_),
    .Q_N(_13477_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][5]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2612),
    .D(_01746_),
    .Q_N(_13476_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][6]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2613),
    .D(_01747_),
    .Q_N(_13475_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][7]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2614),
    .D(_01748_),
    .Q_N(_13474_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][8]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2615),
    .D(_01749_),
    .Q_N(_13473_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][9]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2616),
    .D(_01750_),
    .Q_N(_13472_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][0]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2617),
    .D(_01751_),
    .Q_N(_13471_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][10]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2618),
    .D(_01752_),
    .Q_N(_13470_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][11]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2619),
    .D(_01753_),
    .Q_N(_13469_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][1]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2620),
    .D(_01754_),
    .Q_N(_13468_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][2]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2621),
    .D(_01755_),
    .Q_N(_13467_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][3]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2622),
    .D(_01756_),
    .Q_N(_13466_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][4]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2623),
    .D(_01757_),
    .Q_N(_13465_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][5]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2624),
    .D(_01758_),
    .Q_N(_13464_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][6]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2625),
    .D(_01759_),
    .Q_N(_13463_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][7]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2626),
    .D(_01760_),
    .Q_N(_13462_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][8]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2627),
    .D(_01761_),
    .Q_N(_13461_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][9]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2628),
    .D(_01762_),
    .Q_N(_13460_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2629),
    .D(_01763_),
    .Q_N(_13459_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2630),
    .D(_01764_),
    .Q_N(_13458_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2631),
    .D(_01765_),
    .Q_N(_13457_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2632),
    .D(_01766_),
    .Q_N(_13456_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2633),
    .D(_01767_),
    .Q_N(_13455_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2634),
    .D(_01768_),
    .Q_N(_13454_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2635),
    .D(_01769_),
    .Q_N(_13453_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2636),
    .D(_01770_),
    .Q_N(_13452_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2637),
    .D(_01771_),
    .Q_N(_13451_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2638),
    .D(_01772_),
    .Q_N(_13450_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2639),
    .D(_01773_),
    .Q_N(_13449_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2640),
    .D(_01774_),
    .Q_N(_13448_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][0]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2641),
    .D(_01775_),
    .Q_N(_13447_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][10]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2642),
    .D(_01776_),
    .Q_N(_13446_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][11]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2643),
    .D(_01777_),
    .Q_N(_13445_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][1]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2644),
    .D(_01778_),
    .Q_N(_13444_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][2]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2645),
    .D(_01779_),
    .Q_N(_13443_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][3]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2646),
    .D(_01780_),
    .Q_N(_13442_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][4]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2647),
    .D(_01781_),
    .Q_N(_13441_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][5]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2648),
    .D(_01782_),
    .Q_N(_13440_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][6]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2649),
    .D(_01783_),
    .Q_N(_13439_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][7]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2650),
    .D(_01784_),
    .Q_N(_13438_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][8]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2651),
    .D(_01785_),
    .Q_N(_13437_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][9]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2652),
    .D(_01786_),
    .Q_N(_13436_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][0]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2653),
    .D(_01787_),
    .Q_N(_13435_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][10]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2654),
    .D(_01788_),
    .Q_N(_13434_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][11]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2655),
    .D(_01789_),
    .Q_N(_13433_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][1]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2656),
    .D(_01790_),
    .Q_N(_13432_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][2]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2657),
    .D(_01791_),
    .Q_N(_13431_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][3]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2658),
    .D(_01792_),
    .Q_N(_13430_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][4]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2659),
    .D(_01793_),
    .Q_N(_13429_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][5]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2660),
    .D(_01794_),
    .Q_N(_13428_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][6]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2661),
    .D(_01795_),
    .Q_N(_13427_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][7]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2662),
    .D(_01796_),
    .Q_N(_13426_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][8]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2663),
    .D(_01797_),
    .Q_N(_13425_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][9]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2664),
    .D(_01798_),
    .Q_N(_13424_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2665),
    .D(_01799_),
    .Q_N(_13423_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2666),
    .D(_01800_),
    .Q_N(_13422_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2667),
    .D(_01801_),
    .Q_N(_13421_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2668),
    .D(_01802_),
    .Q_N(_13420_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2669),
    .D(_01803_),
    .Q_N(_13419_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2670),
    .D(_01804_),
    .Q_N(_13418_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2671),
    .D(_01805_),
    .Q_N(_13417_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2672),
    .D(_01806_),
    .Q_N(_13416_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2673),
    .D(_01807_),
    .Q_N(_13415_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2674),
    .D(_01808_),
    .Q_N(_13414_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2675),
    .D(_01809_),
    .Q_N(_13413_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2676),
    .D(_01810_),
    .Q_N(_13412_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2677),
    .D(_01811_),
    .Q_N(_13411_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2678),
    .D(_01812_),
    .Q_N(_13410_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2679),
    .D(_01813_),
    .Q_N(_13409_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2680),
    .D(_01814_),
    .Q_N(_13408_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2681),
    .D(_01815_),
    .Q_N(_13407_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2682),
    .D(_01816_),
    .Q_N(_13406_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2683),
    .D(_01817_),
    .Q_N(_13405_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2684),
    .D(_01818_),
    .Q_N(_13404_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2685),
    .D(_01819_),
    .Q_N(_13403_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2686),
    .D(_01820_),
    .Q_N(_13402_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2687),
    .D(_01821_),
    .Q_N(_13401_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2688),
    .D(_01822_),
    .Q_N(_13400_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2689),
    .D(_01823_),
    .Q_N(_13399_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2690),
    .D(_01824_),
    .Q_N(_13398_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2691),
    .D(_01825_),
    .Q_N(_13397_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2692),
    .D(_01826_),
    .Q_N(_13396_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2693),
    .D(_01827_),
    .Q_N(_13395_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2694),
    .D(_01828_),
    .Q_N(_13394_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2695),
    .D(_01829_),
    .Q_N(_13393_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2696),
    .D(_01830_),
    .Q_N(_13392_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2697),
    .D(_01831_),
    .Q_N(_13391_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2698),
    .D(_01832_),
    .Q_N(_13390_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2699),
    .D(_01833_),
    .Q_N(_13389_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2700),
    .D(_01834_),
    .Q_N(_13388_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2701),
    .D(_01835_),
    .Q_N(_13387_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2702),
    .D(_01836_),
    .Q_N(_13386_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2703),
    .D(_01837_),
    .Q_N(_13385_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2704),
    .D(_01838_),
    .Q_N(_13384_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2705),
    .D(_01839_),
    .Q_N(_13383_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2706),
    .D(_01840_),
    .Q_N(_13382_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2707),
    .D(_01841_),
    .Q_N(_13381_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2708),
    .D(_01842_),
    .Q_N(_13380_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2709),
    .D(_01843_),
    .Q_N(_13379_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2710),
    .D(_01844_),
    .Q_N(_13378_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2711),
    .D(_01845_),
    .Q_N(_13377_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2712),
    .D(_01846_),
    .Q_N(_13376_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2713),
    .D(_01847_),
    .Q_N(_13375_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2714),
    .D(_01848_),
    .Q_N(_13374_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2715),
    .D(_01849_),
    .Q_N(_13373_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2716),
    .D(_01850_),
    .Q_N(_13372_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2717),
    .D(_01851_),
    .Q_N(_13371_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2718),
    .D(_01852_),
    .Q_N(_13370_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2719),
    .D(_01853_),
    .Q_N(_13369_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2720),
    .D(_01854_),
    .Q_N(_13368_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2721),
    .D(_01855_),
    .Q_N(_13367_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2722),
    .D(_01856_),
    .Q_N(_13366_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2723),
    .D(_01857_),
    .Q_N(_13365_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2724),
    .D(_01858_),
    .Q_N(_13364_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][0]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2725),
    .D(_01859_),
    .Q_N(_13363_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][10]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2726),
    .D(_01860_),
    .Q_N(_13362_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][11]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2727),
    .D(_01861_),
    .Q_N(_13361_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][1]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2728),
    .D(_01862_),
    .Q_N(_13360_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][2]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2729),
    .D(_01863_),
    .Q_N(_13359_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][3]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2730),
    .D(_01864_),
    .Q_N(_13358_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][4]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2731),
    .D(_01865_),
    .Q_N(_13357_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][5]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2732),
    .D(_01866_),
    .Q_N(_13356_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][6]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2733),
    .D(_01867_),
    .Q_N(_13355_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][7]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2734),
    .D(_01868_),
    .Q_N(_13354_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][8]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2735),
    .D(_01869_),
    .Q_N(_13353_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][9]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2736),
    .D(_01870_),
    .Q_N(_13352_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][0]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2737),
    .D(_01871_),
    .Q_N(_13351_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][10]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2738),
    .D(_01872_),
    .Q_N(_13350_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][11]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2739),
    .D(_01873_),
    .Q_N(_13349_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][1]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2740),
    .D(_01874_),
    .Q_N(_13348_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][2]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2741),
    .D(_01875_),
    .Q_N(_13347_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][3]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2742),
    .D(_01876_),
    .Q_N(_13346_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][4]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2743),
    .D(_01877_),
    .Q_N(_13345_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][5]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2744),
    .D(_01878_),
    .Q_N(_13344_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][6]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2745),
    .D(_01879_),
    .Q_N(_13343_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][7]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2746),
    .D(_01880_),
    .Q_N(_13342_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][8]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2747),
    .D(_01881_),
    .Q_N(_13341_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][9]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2748),
    .D(_01882_),
    .Q_N(_13340_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[0]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2749),
    .D(_01883_),
    .Q_N(_13339_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[10]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2750),
    .D(_01884_),
    .Q_N(_13338_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[11]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2751),
    .D(_01885_),
    .Q_N(_13337_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[12]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2752),
    .D(_01886_),
    .Q_N(_13336_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[13]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2753),
    .D(_01887_),
    .Q_N(_13335_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[14]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2754),
    .D(_01888_),
    .Q_N(_13334_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[15]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2755),
    .D(_01889_),
    .Q_N(_13333_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[16]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2756),
    .D(_01890_),
    .Q_N(_13332_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[16] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[17]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2757),
    .D(_01891_),
    .Q_N(_13331_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[17] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[18]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2758),
    .D(_01892_),
    .Q_N(_13330_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[18] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[19]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2759),
    .D(_01893_),
    .Q_N(_13329_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[19] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[1]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2760),
    .D(_01894_),
    .Q_N(_13328_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[20]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2761),
    .D(_01895_),
    .Q_N(_13327_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[20] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[21]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2762),
    .D(_01896_),
    .Q_N(_13326_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[21] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[22]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2763),
    .D(_01897_),
    .Q_N(_13325_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[22] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[23]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2764),
    .D(_01898_),
    .Q_N(_13324_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[23] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[24]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2765),
    .D(_01899_),
    .Q_N(_13323_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[24] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[25]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2766),
    .D(_01900_),
    .Q_N(_13322_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[25] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[26]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2767),
    .D(_01901_),
    .Q_N(_13321_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[26] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[27]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2768),
    .D(_01902_),
    .Q_N(_13320_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[27] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[28]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2769),
    .D(_01903_),
    .Q_N(_13319_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[28] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[29]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2770),
    .D(_01904_),
    .Q_N(_13318_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[29] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[2]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2771),
    .D(_01905_),
    .Q_N(_13317_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[30]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2772),
    .D(_01906_),
    .Q_N(_13316_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[30] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[31]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2773),
    .D(_01907_),
    .Q_N(_13315_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[31] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[3]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2774),
    .D(_01908_),
    .Q_N(_13314_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[4]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2775),
    .D(_01909_),
    .Q_N(_13313_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[5]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2776),
    .D(_01910_),
    .Q_N(_13312_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[6]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2777),
    .D(_01911_),
    .Q_N(_13311_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[7]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2778),
    .D(_01912_),
    .Q_N(_13310_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[8]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2779),
    .D(_01913_),
    .Q_N(_13309_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[9]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2780),
    .D(_01914_),
    .Q_N(_13308_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[9] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net2781),
    .D(_01915_),
    .Q_N(_13307_),
    .Q(\cpu.gpio.r_enable_in[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net2782),
    .D(_01916_),
    .Q_N(_13306_),
    .Q(\cpu.gpio.r_enable_in[1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net2783),
    .D(_01917_),
    .Q_N(_13305_),
    .Q(\cpu.gpio.r_enable_in[2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net2784),
    .D(_01918_),
    .Q_N(_13304_),
    .Q(\cpu.gpio.r_enable_in[3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2785),
    .D(_01919_),
    .Q_N(_13303_),
    .Q(\cpu.gpio.r_enable_in[4] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net2786),
    .D(_01920_),
    .Q_N(_13302_),
    .Q(\cpu.gpio.r_enable_in[5] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net2787),
    .D(_01921_),
    .Q_N(_13301_),
    .Q(\cpu.gpio.r_enable_in[6] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net2788),
    .D(_01922_),
    .Q_N(_13300_),
    .Q(\cpu.gpio.r_enable_in[7] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net2789),
    .D(_01923_),
    .Q_N(_13299_),
    .Q(\cpu.gpio.r_enable_io[4] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net2790),
    .D(_01924_),
    .Q_N(_13298_),
    .Q(\cpu.gpio.r_enable_io[5] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net2791),
    .D(_01925_),
    .Q_N(_13297_),
    .Q(\cpu.gpio.r_enable_io[6] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net2792),
    .D(_01926_),
    .Q_N(_13296_),
    .Q(\cpu.gpio.r_enable_io[7] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net2793),
    .D(_01927_),
    .Q_N(_13295_),
    .Q(net7));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net2794),
    .D(_01928_),
    .Q_N(_13294_),
    .Q(net8));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2795),
    .D(_01929_),
    .Q_N(_13293_),
    .Q(net9));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net2796),
    .D(_01930_),
    .Q_N(_13292_),
    .Q(net10));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[0]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2797),
    .D(_01931_),
    .Q_N(_13291_),
    .Q(\cpu.gpio.genblk2[4].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[1]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2798),
    .D(_01932_),
    .Q_N(_13290_),
    .Q(\cpu.gpio.genblk2[5].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[2]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2799),
    .D(_01933_),
    .Q_N(_13289_),
    .Q(\cpu.gpio.genblk2[6].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[3]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2800),
    .D(_01934_),
    .Q_N(_13288_),
    .Q(\cpu.gpio.genblk2[7].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[0]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2801),
    .D(_01935_),
    .Q_N(_13287_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[1]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net2802),
    .D(_01936_),
    .Q_N(_13286_),
    .Q(\cpu.gpio.genblk1[4].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[2]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net2803),
    .D(_01937_),
    .Q_N(_13285_),
    .Q(\cpu.gpio.genblk1[5].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[3]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2804),
    .D(_01938_),
    .Q_N(_13284_),
    .Q(\cpu.gpio.genblk1[6].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[4]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net2805),
    .D(_01939_),
    .Q_N(_13283_),
    .Q(\cpu.gpio.genblk1[7].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2806),
    .D(_01940_),
    .Q_N(_13282_),
    .Q(\cpu.gpio.r_spi_miso_src[0][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2807),
    .D(_01941_),
    .Q_N(_00291_),
    .Q(\cpu.gpio.r_spi_miso_src[0][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2808),
    .D(_01942_),
    .Q_N(_00100_),
    .Q(\cpu.gpio.r_spi_miso_src[0][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2809),
    .D(_01943_),
    .Q_N(_00109_),
    .Q(\cpu.gpio.r_spi_miso_src[0][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2810),
    .D(_01944_),
    .Q_N(_13281_),
    .Q(\cpu.gpio.r_spi_miso_src[1][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2811),
    .D(_01945_),
    .Q_N(_00126_),
    .Q(\cpu.gpio.r_spi_miso_src[1][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2812),
    .D(_01946_),
    .Q_N(_00137_),
    .Q(\cpu.gpio.r_spi_miso_src[1][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2813),
    .D(_01947_),
    .Q_N(_00148_),
    .Q(\cpu.gpio.r_spi_miso_src[1][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2814),
    .D(_01948_),
    .Q_N(_13280_),
    .Q(\cpu.gpio.r_src_io[4][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2815),
    .D(_01949_),
    .Q_N(_13279_),
    .Q(\cpu.gpio.r_src_io[4][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2816),
    .D(_01950_),
    .Q_N(_00171_),
    .Q(\cpu.gpio.r_src_io[4][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2817),
    .D(_01951_),
    .Q_N(_13278_),
    .Q(\cpu.gpio.r_src_io[4][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2818),
    .D(_01952_),
    .Q_N(_13277_),
    .Q(\cpu.gpio.r_src_io[5][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2819),
    .D(_01953_),
    .Q_N(_13276_),
    .Q(\cpu.gpio.r_src_io[5][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2820),
    .D(_01954_),
    .Q_N(_00170_),
    .Q(\cpu.gpio.r_src_io[5][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2821),
    .D(_01955_),
    .Q_N(_13275_),
    .Q(\cpu.gpio.r_src_io[5][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2822),
    .D(_01956_),
    .Q_N(_13274_),
    .Q(\cpu.gpio.r_src_io[6][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2823),
    .D(_01957_),
    .Q_N(_00287_),
    .Q(\cpu.gpio.r_src_io[6][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2824),
    .D(_01958_),
    .Q_N(_00096_),
    .Q(\cpu.gpio.r_src_io[6][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net2825),
    .D(_01959_),
    .Q_N(_00106_),
    .Q(\cpu.gpio.r_src_io[6][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2826),
    .D(_01960_),
    .Q_N(_13273_),
    .Q(\cpu.gpio.r_src_io[7][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2827),
    .D(_01961_),
    .Q_N(_00122_),
    .Q(\cpu.gpio.r_src_io[7][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2828),
    .D(_01962_),
    .Q_N(_00133_),
    .Q(\cpu.gpio.r_src_io[7][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2829),
    .D(_01963_),
    .Q_N(_00144_),
    .Q(\cpu.gpio.r_src_io[7][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2830),
    .D(_01964_),
    .Q_N(_13272_),
    .Q(\cpu.gpio.r_src_o[3][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net2831),
    .D(_01965_),
    .Q_N(_00125_),
    .Q(\cpu.gpio.r_src_o[3][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2832),
    .D(_01966_),
    .Q_N(_00136_),
    .Q(\cpu.gpio.r_src_o[3][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2833),
    .D(_01967_),
    .Q_N(_00147_),
    .Q(\cpu.gpio.r_src_o[3][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net2834),
    .D(_01968_),
    .Q_N(_13271_),
    .Q(\cpu.gpio.r_src_o[4][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2835),
    .D(_01969_),
    .Q_N(_00289_),
    .Q(\cpu.gpio.r_src_o[4][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2836),
    .D(_01970_),
    .Q_N(_00098_),
    .Q(\cpu.gpio.r_src_o[4][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2837),
    .D(_01971_),
    .Q_N(_00108_),
    .Q(\cpu.gpio.r_src_o[4][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2838),
    .D(_01972_),
    .Q_N(_13270_),
    .Q(\cpu.gpio.r_src_o[5][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2839),
    .D(_01973_),
    .Q_N(_00124_),
    .Q(\cpu.gpio.r_src_o[5][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2840),
    .D(_01974_),
    .Q_N(_00135_),
    .Q(\cpu.gpio.r_src_o[5][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2841),
    .D(_01975_),
    .Q_N(_00146_),
    .Q(\cpu.gpio.r_src_o[5][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2842),
    .D(_01976_),
    .Q_N(_13269_),
    .Q(\cpu.gpio.r_src_o[6][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2843),
    .D(_01977_),
    .Q_N(_00288_),
    .Q(\cpu.gpio.r_src_o[6][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2844),
    .D(_01978_),
    .Q_N(_00097_),
    .Q(\cpu.gpio.r_src_o[6][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2845),
    .D(_01979_),
    .Q_N(_00107_),
    .Q(\cpu.gpio.r_src_o[6][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2846),
    .D(_01980_),
    .Q_N(_13268_),
    .Q(\cpu.gpio.r_src_o[7][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2847),
    .D(_01981_),
    .Q_N(_00123_),
    .Q(\cpu.gpio.r_src_o[7][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2848),
    .D(_01982_),
    .Q_N(_00134_),
    .Q(\cpu.gpio.r_src_o[7][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2849),
    .D(_01983_),
    .Q_N(_00145_),
    .Q(\cpu.gpio.r_src_o[7][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_uart_rx_src[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2850),
    .D(_01984_),
    .Q_N(_13267_),
    .Q(\cpu.gpio.r_uart_rx_src[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_uart_rx_src[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2851),
    .D(_01985_),
    .Q_N(_00290_),
    .Q(\cpu.gpio.r_uart_rx_src[1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_uart_rx_src[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net2852),
    .D(_01986_),
    .Q_N(_00099_),
    .Q(\cpu.gpio.r_uart_rx_src[2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2853),
    .D(_01987_),
    .Q_N(_13266_),
    .Q(\cpu.icache.r_data[0][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2854),
    .D(_01988_),
    .Q_N(_00185_),
    .Q(\cpu.icache.r_data[0][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2855),
    .D(_01989_),
    .Q_N(_00187_),
    .Q(\cpu.icache.r_data[0][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2856),
    .D(_01990_),
    .Q_N(_00197_),
    .Q(\cpu.icache.r_data[0][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2857),
    .D(_01991_),
    .Q_N(_13265_),
    .Q(\cpu.icache.r_data[0][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2858),
    .D(_01992_),
    .Q_N(_00189_),
    .Q(\cpu.icache.r_data[0][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2859),
    .D(_01993_),
    .Q_N(_00191_),
    .Q(\cpu.icache.r_data[0][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2860),
    .D(_01994_),
    .Q_N(_13264_),
    .Q(\cpu.icache.r_data[0][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2861),
    .D(_01995_),
    .Q_N(_13263_),
    .Q(\cpu.icache.r_data[0][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2862),
    .D(_01996_),
    .Q_N(_00157_),
    .Q(\cpu.icache.r_data[0][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][19]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2863),
    .D(_01997_),
    .Q_N(_00159_),
    .Q(\cpu.icache.r_data[0][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2864),
    .D(_01998_),
    .Q_N(_13262_),
    .Q(\cpu.icache.r_data[0][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][20]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2865),
    .D(_01999_),
    .Q_N(_00161_),
    .Q(\cpu.icache.r_data[0][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][21]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2866),
    .D(_02000_),
    .Q_N(_00194_),
    .Q(\cpu.icache.r_data[0][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][22]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2867),
    .D(_02001_),
    .Q_N(_00196_),
    .Q(\cpu.icache.r_data[0][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][23]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2868),
    .D(_02002_),
    .Q_N(_00151_),
    .Q(\cpu.icache.r_data[0][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][24]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2869),
    .D(_02003_),
    .Q_N(_00153_),
    .Q(\cpu.icache.r_data[0][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][25]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net2870),
    .D(_02004_),
    .Q_N(_00155_),
    .Q(\cpu.icache.r_data[0][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][26]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2871),
    .D(_02005_),
    .Q_N(_00186_),
    .Q(\cpu.icache.r_data[0][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][27]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2872),
    .D(_02006_),
    .Q_N(_00188_),
    .Q(\cpu.icache.r_data[0][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][28]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2873),
    .D(_02007_),
    .Q_N(_00198_),
    .Q(\cpu.icache.r_data[0][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][29]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2874),
    .D(_02008_),
    .Q_N(_13261_),
    .Q(\cpu.icache.r_data[0][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2875),
    .D(_02009_),
    .Q_N(_00156_),
    .Q(\cpu.icache.r_data[0][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][30]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2876),
    .D(_02010_),
    .Q_N(_00190_),
    .Q(\cpu.icache.r_data[0][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][31]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2877),
    .D(_02011_),
    .Q_N(_00192_),
    .Q(\cpu.icache.r_data[0][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2878),
    .D(_02012_),
    .Q_N(_00158_),
    .Q(\cpu.icache.r_data[0][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2879),
    .D(_02013_),
    .Q_N(_00160_),
    .Q(\cpu.icache.r_data[0][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2880),
    .D(_02014_),
    .Q_N(_00193_),
    .Q(\cpu.icache.r_data[0][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net2881),
    .D(_02015_),
    .Q_N(_00195_),
    .Q(\cpu.icache.r_data[0][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2882),
    .D(_02016_),
    .Q_N(_00150_),
    .Q(\cpu.icache.r_data[0][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2883),
    .D(_02017_),
    .Q_N(_00152_),
    .Q(\cpu.icache.r_data[0][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2884),
    .D(_02018_),
    .Q_N(_00154_),
    .Q(\cpu.icache.r_data[0][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2885),
    .D(_02019_),
    .Q_N(_13260_),
    .Q(\cpu.icache.r_data[1][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2886),
    .D(_02020_),
    .Q_N(_13259_),
    .Q(\cpu.icache.r_data[1][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2887),
    .D(_02021_),
    .Q_N(_13258_),
    .Q(\cpu.icache.r_data[1][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2888),
    .D(_02022_),
    .Q_N(_13257_),
    .Q(\cpu.icache.r_data[1][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2889),
    .D(_02023_),
    .Q_N(_13256_),
    .Q(\cpu.icache.r_data[1][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2890),
    .D(_02024_),
    .Q_N(_13255_),
    .Q(\cpu.icache.r_data[1][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2891),
    .D(_02025_),
    .Q_N(_13254_),
    .Q(\cpu.icache.r_data[1][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net2892),
    .D(_02026_),
    .Q_N(_13253_),
    .Q(\cpu.icache.r_data[1][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2893),
    .D(_02027_),
    .Q_N(_13252_),
    .Q(\cpu.icache.r_data[1][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2894),
    .D(_02028_),
    .Q_N(_13251_),
    .Q(\cpu.icache.r_data[1][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][19]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2895),
    .D(_02029_),
    .Q_N(_13250_),
    .Q(\cpu.icache.r_data[1][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2896),
    .D(_02030_),
    .Q_N(_13249_),
    .Q(\cpu.icache.r_data[1][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][20]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2897),
    .D(_02031_),
    .Q_N(_13248_),
    .Q(\cpu.icache.r_data[1][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][21]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2898),
    .D(_02032_),
    .Q_N(_13247_),
    .Q(\cpu.icache.r_data[1][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][22]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2899),
    .D(_02033_),
    .Q_N(_13246_),
    .Q(\cpu.icache.r_data[1][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][23]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2900),
    .D(_02034_),
    .Q_N(_13245_),
    .Q(\cpu.icache.r_data[1][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][24]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net2901),
    .D(_02035_),
    .Q_N(_13244_),
    .Q(\cpu.icache.r_data[1][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][25]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2902),
    .D(_02036_),
    .Q_N(_13243_),
    .Q(\cpu.icache.r_data[1][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][26]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net2903),
    .D(_02037_),
    .Q_N(_13242_),
    .Q(\cpu.icache.r_data[1][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][27]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net2904),
    .D(_02038_),
    .Q_N(_13241_),
    .Q(\cpu.icache.r_data[1][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][28]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2905),
    .D(_02039_),
    .Q_N(_13240_),
    .Q(\cpu.icache.r_data[1][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][29]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2906),
    .D(_02040_),
    .Q_N(_13239_),
    .Q(\cpu.icache.r_data[1][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2907),
    .D(_02041_),
    .Q_N(_13238_),
    .Q(\cpu.icache.r_data[1][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][30]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2908),
    .D(_02042_),
    .Q_N(_13237_),
    .Q(\cpu.icache.r_data[1][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][31]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2909),
    .D(_02043_),
    .Q_N(_13236_),
    .Q(\cpu.icache.r_data[1][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2910),
    .D(_02044_),
    .Q_N(_13235_),
    .Q(\cpu.icache.r_data[1][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2911),
    .D(_02045_),
    .Q_N(_13234_),
    .Q(\cpu.icache.r_data[1][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2912),
    .D(_02046_),
    .Q_N(_13233_),
    .Q(\cpu.icache.r_data[1][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2913),
    .D(_02047_),
    .Q_N(_13232_),
    .Q(\cpu.icache.r_data[1][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2914),
    .D(_02048_),
    .Q_N(_13231_),
    .Q(\cpu.icache.r_data[1][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2915),
    .D(_02049_),
    .Q_N(_13230_),
    .Q(\cpu.icache.r_data[1][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2916),
    .D(_02050_),
    .Q_N(_13229_),
    .Q(\cpu.icache.r_data[1][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2917),
    .D(_02051_),
    .Q_N(_13228_),
    .Q(\cpu.icache.r_data[2][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2918),
    .D(_02052_),
    .Q_N(_13227_),
    .Q(\cpu.icache.r_data[2][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2919),
    .D(_02053_),
    .Q_N(_13226_),
    .Q(\cpu.icache.r_data[2][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net2920),
    .D(_02054_),
    .Q_N(_13225_),
    .Q(\cpu.icache.r_data[2][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2921),
    .D(_02055_),
    .Q_N(_13224_),
    .Q(\cpu.icache.r_data[2][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2922),
    .D(_02056_),
    .Q_N(_13223_),
    .Q(\cpu.icache.r_data[2][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net2923),
    .D(_02057_),
    .Q_N(_13222_),
    .Q(\cpu.icache.r_data[2][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net2924),
    .D(_02058_),
    .Q_N(_13221_),
    .Q(\cpu.icache.r_data[2][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2925),
    .D(_02059_),
    .Q_N(_13220_),
    .Q(\cpu.icache.r_data[2][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net2926),
    .D(_02060_),
    .Q_N(_13219_),
    .Q(\cpu.icache.r_data[2][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][19]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2927),
    .D(_02061_),
    .Q_N(_13218_),
    .Q(\cpu.icache.r_data[2][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2928),
    .D(_02062_),
    .Q_N(_13217_),
    .Q(\cpu.icache.r_data[2][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][20]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2929),
    .D(_02063_),
    .Q_N(_13216_),
    .Q(\cpu.icache.r_data[2][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][21]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2930),
    .D(_02064_),
    .Q_N(_13215_),
    .Q(\cpu.icache.r_data[2][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][22]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2931),
    .D(_02065_),
    .Q_N(_13214_),
    .Q(\cpu.icache.r_data[2][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][23]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2932),
    .D(_02066_),
    .Q_N(_13213_),
    .Q(\cpu.icache.r_data[2][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][24]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net2933),
    .D(_02067_),
    .Q_N(_13212_),
    .Q(\cpu.icache.r_data[2][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][25]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2934),
    .D(_02068_),
    .Q_N(_13211_),
    .Q(\cpu.icache.r_data[2][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][26]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net2935),
    .D(_02069_),
    .Q_N(_13210_),
    .Q(\cpu.icache.r_data[2][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][27]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2936),
    .D(_02070_),
    .Q_N(_13209_),
    .Q(\cpu.icache.r_data[2][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][28]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2937),
    .D(_02071_),
    .Q_N(_13208_),
    .Q(\cpu.icache.r_data[2][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][29]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2938),
    .D(_02072_),
    .Q_N(_13207_),
    .Q(\cpu.icache.r_data[2][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2939),
    .D(_02073_),
    .Q_N(_13206_),
    .Q(\cpu.icache.r_data[2][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][30]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2940),
    .D(_02074_),
    .Q_N(_13205_),
    .Q(\cpu.icache.r_data[2][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][31]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2941),
    .D(_02075_),
    .Q_N(_13204_),
    .Q(\cpu.icache.r_data[2][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2942),
    .D(_02076_),
    .Q_N(_13203_),
    .Q(\cpu.icache.r_data[2][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2943),
    .D(_02077_),
    .Q_N(_13202_),
    .Q(\cpu.icache.r_data[2][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2944),
    .D(_02078_),
    .Q_N(_13201_),
    .Q(\cpu.icache.r_data[2][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2945),
    .D(_02079_),
    .Q_N(_13200_),
    .Q(\cpu.icache.r_data[2][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2946),
    .D(_02080_),
    .Q_N(_13199_),
    .Q(\cpu.icache.r_data[2][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net2947),
    .D(_02081_),
    .Q_N(_13198_),
    .Q(\cpu.icache.r_data[2][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2948),
    .D(_02082_),
    .Q_N(_13197_),
    .Q(\cpu.icache.r_data[2][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2949),
    .D(_02083_),
    .Q_N(_13196_),
    .Q(\cpu.icache.r_data[3][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2950),
    .D(_02084_),
    .Q_N(_13195_),
    .Q(\cpu.icache.r_data[3][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net2951),
    .D(_02085_),
    .Q_N(_13194_),
    .Q(\cpu.icache.r_data[3][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net2952),
    .D(_02086_),
    .Q_N(_13193_),
    .Q(\cpu.icache.r_data[3][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2953),
    .D(_02087_),
    .Q_N(_13192_),
    .Q(\cpu.icache.r_data[3][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2954),
    .D(_02088_),
    .Q_N(_13191_),
    .Q(\cpu.icache.r_data[3][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2955),
    .D(_02089_),
    .Q_N(_13190_),
    .Q(\cpu.icache.r_data[3][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2956),
    .D(_02090_),
    .Q_N(_13189_),
    .Q(\cpu.icache.r_data[3][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2957),
    .D(_02091_),
    .Q_N(_13188_),
    .Q(\cpu.icache.r_data[3][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net2958),
    .D(_02092_),
    .Q_N(_13187_),
    .Q(\cpu.icache.r_data[3][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][19]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2959),
    .D(_02093_),
    .Q_N(_13186_),
    .Q(\cpu.icache.r_data[3][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2960),
    .D(_02094_),
    .Q_N(_13185_),
    .Q(\cpu.icache.r_data[3][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][20]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2961),
    .D(_02095_),
    .Q_N(_13184_),
    .Q(\cpu.icache.r_data[3][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][21]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net2962),
    .D(_02096_),
    .Q_N(_13183_),
    .Q(\cpu.icache.r_data[3][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][22]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2963),
    .D(_02097_),
    .Q_N(_13182_),
    .Q(\cpu.icache.r_data[3][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][23]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net2964),
    .D(_02098_),
    .Q_N(_13181_),
    .Q(\cpu.icache.r_data[3][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][24]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2965),
    .D(_02099_),
    .Q_N(_13180_),
    .Q(\cpu.icache.r_data[3][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][25]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2966),
    .D(_02100_),
    .Q_N(_13179_),
    .Q(\cpu.icache.r_data[3][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][26]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2967),
    .D(_02101_),
    .Q_N(_13178_),
    .Q(\cpu.icache.r_data[3][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][27]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2968),
    .D(_02102_),
    .Q_N(_13177_),
    .Q(\cpu.icache.r_data[3][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][28]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2969),
    .D(_02103_),
    .Q_N(_13176_),
    .Q(\cpu.icache.r_data[3][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][29]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2970),
    .D(_02104_),
    .Q_N(_13175_),
    .Q(\cpu.icache.r_data[3][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2971),
    .D(_02105_),
    .Q_N(_13174_),
    .Q(\cpu.icache.r_data[3][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][30]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2972),
    .D(_02106_),
    .Q_N(_13173_),
    .Q(\cpu.icache.r_data[3][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][31]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net2973),
    .D(_02107_),
    .Q_N(_13172_),
    .Q(\cpu.icache.r_data[3][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2974),
    .D(_02108_),
    .Q_N(_13171_),
    .Q(\cpu.icache.r_data[3][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2975),
    .D(_02109_),
    .Q_N(_13170_),
    .Q(\cpu.icache.r_data[3][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2976),
    .D(_02110_),
    .Q_N(_13169_),
    .Q(\cpu.icache.r_data[3][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2977),
    .D(_02111_),
    .Q_N(_13168_),
    .Q(\cpu.icache.r_data[3][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2978),
    .D(_02112_),
    .Q_N(_13167_),
    .Q(\cpu.icache.r_data[3][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2979),
    .D(_02113_),
    .Q_N(_13166_),
    .Q(\cpu.icache.r_data[3][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2980),
    .D(_02114_),
    .Q_N(_13165_),
    .Q(\cpu.icache.r_data[3][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2981),
    .D(_02115_),
    .Q_N(_13164_),
    .Q(\cpu.icache.r_data[4][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2982),
    .D(_02116_),
    .Q_N(_13163_),
    .Q(\cpu.icache.r_data[4][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2983),
    .D(_02117_),
    .Q_N(_13162_),
    .Q(\cpu.icache.r_data[4][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2984),
    .D(_02118_),
    .Q_N(_13161_),
    .Q(\cpu.icache.r_data[4][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2985),
    .D(_02119_),
    .Q_N(_13160_),
    .Q(\cpu.icache.r_data[4][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2986),
    .D(_02120_),
    .Q_N(_13159_),
    .Q(\cpu.icache.r_data[4][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2987),
    .D(_02121_),
    .Q_N(_13158_),
    .Q(\cpu.icache.r_data[4][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2988),
    .D(_02122_),
    .Q_N(_13157_),
    .Q(\cpu.icache.r_data[4][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2989),
    .D(_02123_),
    .Q_N(_13156_),
    .Q(\cpu.icache.r_data[4][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2990),
    .D(_02124_),
    .Q_N(_13155_),
    .Q(\cpu.icache.r_data[4][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][19]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2991),
    .D(_02125_),
    .Q_N(_13154_),
    .Q(\cpu.icache.r_data[4][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2992),
    .D(_02126_),
    .Q_N(_13153_),
    .Q(\cpu.icache.r_data[4][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][20]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2993),
    .D(_02127_),
    .Q_N(_13152_),
    .Q(\cpu.icache.r_data[4][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][21]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2994),
    .D(_02128_),
    .Q_N(_13151_),
    .Q(\cpu.icache.r_data[4][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][22]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net2995),
    .D(_02129_),
    .Q_N(_13150_),
    .Q(\cpu.icache.r_data[4][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][23]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2996),
    .D(_02130_),
    .Q_N(_13149_),
    .Q(\cpu.icache.r_data[4][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][24]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net2997),
    .D(_02131_),
    .Q_N(_13148_),
    .Q(\cpu.icache.r_data[4][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][25]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2998),
    .D(_02132_),
    .Q_N(_13147_),
    .Q(\cpu.icache.r_data[4][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][26]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2999),
    .D(_02133_),
    .Q_N(_13146_),
    .Q(\cpu.icache.r_data[4][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][27]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3000),
    .D(_02134_),
    .Q_N(_13145_),
    .Q(\cpu.icache.r_data[4][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][28]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3001),
    .D(_02135_),
    .Q_N(_13144_),
    .Q(\cpu.icache.r_data[4][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][29]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3002),
    .D(_02136_),
    .Q_N(_13143_),
    .Q(\cpu.icache.r_data[4][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3003),
    .D(_02137_),
    .Q_N(_13142_),
    .Q(\cpu.icache.r_data[4][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][30]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3004),
    .D(_02138_),
    .Q_N(_13141_),
    .Q(\cpu.icache.r_data[4][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][31]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3005),
    .D(_02139_),
    .Q_N(_13140_),
    .Q(\cpu.icache.r_data[4][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3006),
    .D(_02140_),
    .Q_N(_13139_),
    .Q(\cpu.icache.r_data[4][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3007),
    .D(_02141_),
    .Q_N(_13138_),
    .Q(\cpu.icache.r_data[4][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3008),
    .D(_02142_),
    .Q_N(_13137_),
    .Q(\cpu.icache.r_data[4][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3009),
    .D(_02143_),
    .Q_N(_13136_),
    .Q(\cpu.icache.r_data[4][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3010),
    .D(_02144_),
    .Q_N(_13135_),
    .Q(\cpu.icache.r_data[4][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3011),
    .D(_02145_),
    .Q_N(_13134_),
    .Q(\cpu.icache.r_data[4][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3012),
    .D(_02146_),
    .Q_N(_13133_),
    .Q(\cpu.icache.r_data[4][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3013),
    .D(_02147_),
    .Q_N(_13132_),
    .Q(\cpu.icache.r_data[5][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3014),
    .D(_02148_),
    .Q_N(_13131_),
    .Q(\cpu.icache.r_data[5][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3015),
    .D(_02149_),
    .Q_N(_13130_),
    .Q(\cpu.icache.r_data[5][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3016),
    .D(_02150_),
    .Q_N(_13129_),
    .Q(\cpu.icache.r_data[5][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net3017),
    .D(_02151_),
    .Q_N(_13128_),
    .Q(\cpu.icache.r_data[5][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3018),
    .D(_02152_),
    .Q_N(_13127_),
    .Q(\cpu.icache.r_data[5][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3019),
    .D(_02153_),
    .Q_N(_13126_),
    .Q(\cpu.icache.r_data[5][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3020),
    .D(_02154_),
    .Q_N(_13125_),
    .Q(\cpu.icache.r_data[5][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3021),
    .D(_02155_),
    .Q_N(_13124_),
    .Q(\cpu.icache.r_data[5][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3022),
    .D(_02156_),
    .Q_N(_13123_),
    .Q(\cpu.icache.r_data[5][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][19]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3023),
    .D(_02157_),
    .Q_N(_13122_),
    .Q(\cpu.icache.r_data[5][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3024),
    .D(_02158_),
    .Q_N(_13121_),
    .Q(\cpu.icache.r_data[5][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][20]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3025),
    .D(_02159_),
    .Q_N(_13120_),
    .Q(\cpu.icache.r_data[5][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][21]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3026),
    .D(_02160_),
    .Q_N(_13119_),
    .Q(\cpu.icache.r_data[5][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][22]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3027),
    .D(_02161_),
    .Q_N(_13118_),
    .Q(\cpu.icache.r_data[5][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][23]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3028),
    .D(_02162_),
    .Q_N(_13117_),
    .Q(\cpu.icache.r_data[5][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][24]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3029),
    .D(_02163_),
    .Q_N(_13116_),
    .Q(\cpu.icache.r_data[5][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][25]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3030),
    .D(_02164_),
    .Q_N(_13115_),
    .Q(\cpu.icache.r_data[5][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][26]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3031),
    .D(_02165_),
    .Q_N(_13114_),
    .Q(\cpu.icache.r_data[5][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][27]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3032),
    .D(_02166_),
    .Q_N(_13113_),
    .Q(\cpu.icache.r_data[5][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][28]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3033),
    .D(_02167_),
    .Q_N(_13112_),
    .Q(\cpu.icache.r_data[5][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][29]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3034),
    .D(_02168_),
    .Q_N(_13111_),
    .Q(\cpu.icache.r_data[5][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3035),
    .D(_02169_),
    .Q_N(_13110_),
    .Q(\cpu.icache.r_data[5][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][30]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3036),
    .D(_02170_),
    .Q_N(_13109_),
    .Q(\cpu.icache.r_data[5][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][31]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3037),
    .D(_02171_),
    .Q_N(_13108_),
    .Q(\cpu.icache.r_data[5][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3038),
    .D(_02172_),
    .Q_N(_13107_),
    .Q(\cpu.icache.r_data[5][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3039),
    .D(_02173_),
    .Q_N(_13106_),
    .Q(\cpu.icache.r_data[5][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3040),
    .D(_02174_),
    .Q_N(_13105_),
    .Q(\cpu.icache.r_data[5][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3041),
    .D(_02175_),
    .Q_N(_13104_),
    .Q(\cpu.icache.r_data[5][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3042),
    .D(_02176_),
    .Q_N(_13103_),
    .Q(\cpu.icache.r_data[5][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3043),
    .D(_02177_),
    .Q_N(_13102_),
    .Q(\cpu.icache.r_data[5][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3044),
    .D(_02178_),
    .Q_N(_13101_),
    .Q(\cpu.icache.r_data[5][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3045),
    .D(_02179_),
    .Q_N(_13100_),
    .Q(\cpu.icache.r_data[6][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3046),
    .D(_02180_),
    .Q_N(_13099_),
    .Q(\cpu.icache.r_data[6][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3047),
    .D(_02181_),
    .Q_N(_13098_),
    .Q(\cpu.icache.r_data[6][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3048),
    .D(_02182_),
    .Q_N(_13097_),
    .Q(\cpu.icache.r_data[6][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net3049),
    .D(_02183_),
    .Q_N(_13096_),
    .Q(\cpu.icache.r_data[6][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3050),
    .D(_02184_),
    .Q_N(_13095_),
    .Q(\cpu.icache.r_data[6][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3051),
    .D(_02185_),
    .Q_N(_13094_),
    .Q(\cpu.icache.r_data[6][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3052),
    .D(_02186_),
    .Q_N(_13093_),
    .Q(\cpu.icache.r_data[6][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3053),
    .D(_02187_),
    .Q_N(_13092_),
    .Q(\cpu.icache.r_data[6][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3054),
    .D(_02188_),
    .Q_N(_13091_),
    .Q(\cpu.icache.r_data[6][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][19]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3055),
    .D(_02189_),
    .Q_N(_13090_),
    .Q(\cpu.icache.r_data[6][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3056),
    .D(_02190_),
    .Q_N(_13089_),
    .Q(\cpu.icache.r_data[6][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][20]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3057),
    .D(_02191_),
    .Q_N(_13088_),
    .Q(\cpu.icache.r_data[6][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][21]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3058),
    .D(_02192_),
    .Q_N(_13087_),
    .Q(\cpu.icache.r_data[6][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][22]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3059),
    .D(_02193_),
    .Q_N(_13086_),
    .Q(\cpu.icache.r_data[6][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][23]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3060),
    .D(_02194_),
    .Q_N(_13085_),
    .Q(\cpu.icache.r_data[6][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][24]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3061),
    .D(_02195_),
    .Q_N(_13084_),
    .Q(\cpu.icache.r_data[6][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][25]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3062),
    .D(_02196_),
    .Q_N(_13083_),
    .Q(\cpu.icache.r_data[6][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][26]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3063),
    .D(_02197_),
    .Q_N(_13082_),
    .Q(\cpu.icache.r_data[6][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][27]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3064),
    .D(_02198_),
    .Q_N(_13081_),
    .Q(\cpu.icache.r_data[6][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][28]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3065),
    .D(_02199_),
    .Q_N(_13080_),
    .Q(\cpu.icache.r_data[6][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][29]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3066),
    .D(_02200_),
    .Q_N(_13079_),
    .Q(\cpu.icache.r_data[6][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3067),
    .D(_02201_),
    .Q_N(_13078_),
    .Q(\cpu.icache.r_data[6][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][30]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3068),
    .D(_02202_),
    .Q_N(_13077_),
    .Q(\cpu.icache.r_data[6][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][31]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3069),
    .D(_02203_),
    .Q_N(_13076_),
    .Q(\cpu.icache.r_data[6][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3070),
    .D(_02204_),
    .Q_N(_13075_),
    .Q(\cpu.icache.r_data[6][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net3071),
    .D(_02205_),
    .Q_N(_13074_),
    .Q(\cpu.icache.r_data[6][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net3072),
    .D(_02206_),
    .Q_N(_13073_),
    .Q(\cpu.icache.r_data[6][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net3073),
    .D(_02207_),
    .Q_N(_13072_),
    .Q(\cpu.icache.r_data[6][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net3074),
    .D(_02208_),
    .Q_N(_13071_),
    .Q(\cpu.icache.r_data[6][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3075),
    .D(_02209_),
    .Q_N(_13070_),
    .Q(\cpu.icache.r_data[6][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3076),
    .D(_02210_),
    .Q_N(_13069_),
    .Q(\cpu.icache.r_data[6][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3077),
    .D(_02211_),
    .Q_N(_13068_),
    .Q(\cpu.icache.r_data[7][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3078),
    .D(_02212_),
    .Q_N(_13067_),
    .Q(\cpu.icache.r_data[7][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3079),
    .D(_02213_),
    .Q_N(_13066_),
    .Q(\cpu.icache.r_data[7][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3080),
    .D(_02214_),
    .Q_N(_13065_),
    .Q(\cpu.icache.r_data[7][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3081),
    .D(_02215_),
    .Q_N(_13064_),
    .Q(\cpu.icache.r_data[7][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3082),
    .D(_02216_),
    .Q_N(_13063_),
    .Q(\cpu.icache.r_data[7][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3083),
    .D(_02217_),
    .Q_N(_13062_),
    .Q(\cpu.icache.r_data[7][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3084),
    .D(_02218_),
    .Q_N(_13061_),
    .Q(\cpu.icache.r_data[7][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3085),
    .D(_02219_),
    .Q_N(_13060_),
    .Q(\cpu.icache.r_data[7][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3086),
    .D(_02220_),
    .Q_N(_13059_),
    .Q(\cpu.icache.r_data[7][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][19]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3087),
    .D(_02221_),
    .Q_N(_13058_),
    .Q(\cpu.icache.r_data[7][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3088),
    .D(_02222_),
    .Q_N(_13057_),
    .Q(\cpu.icache.r_data[7][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][20]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3089),
    .D(_02223_),
    .Q_N(_13056_),
    .Q(\cpu.icache.r_data[7][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][21]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3090),
    .D(_02224_),
    .Q_N(_13055_),
    .Q(\cpu.icache.r_data[7][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][22]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3091),
    .D(_02225_),
    .Q_N(_13054_),
    .Q(\cpu.icache.r_data[7][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][23]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3092),
    .D(_02226_),
    .Q_N(_13053_),
    .Q(\cpu.icache.r_data[7][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][24]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3093),
    .D(_02227_),
    .Q_N(_13052_),
    .Q(\cpu.icache.r_data[7][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][25]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3094),
    .D(_02228_),
    .Q_N(_13051_),
    .Q(\cpu.icache.r_data[7][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][26]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3095),
    .D(_02229_),
    .Q_N(_13050_),
    .Q(\cpu.icache.r_data[7][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][27]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3096),
    .D(_02230_),
    .Q_N(_13049_),
    .Q(\cpu.icache.r_data[7][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][28]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3097),
    .D(_02231_),
    .Q_N(_13048_),
    .Q(\cpu.icache.r_data[7][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][29]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3098),
    .D(_02232_),
    .Q_N(_13047_),
    .Q(\cpu.icache.r_data[7][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3099),
    .D(_02233_),
    .Q_N(_13046_),
    .Q(\cpu.icache.r_data[7][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][30]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3100),
    .D(_02234_),
    .Q_N(_13045_),
    .Q(\cpu.icache.r_data[7][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][31]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3101),
    .D(_02235_),
    .Q_N(_13044_),
    .Q(\cpu.icache.r_data[7][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3102),
    .D(_02236_),
    .Q_N(_13043_),
    .Q(\cpu.icache.r_data[7][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3103),
    .D(_02237_),
    .Q_N(_13042_),
    .Q(\cpu.icache.r_data[7][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3104),
    .D(_02238_),
    .Q_N(_13041_),
    .Q(\cpu.icache.r_data[7][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3105),
    .D(_02239_),
    .Q_N(_13040_),
    .Q(\cpu.icache.r_data[7][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3106),
    .D(_02240_),
    .Q_N(_13039_),
    .Q(\cpu.icache.r_data[7][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3107),
    .D(_02241_),
    .Q_N(_13038_),
    .Q(\cpu.icache.r_data[7][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3108),
    .D(_02242_),
    .Q_N(_13037_),
    .Q(\cpu.icache.r_data[7][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_offset[0]$_SDFF_PN0_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3109),
    .D(_02243_),
    .Q_N(_00293_),
    .Q(\cpu.icache.r_offset[0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_offset[1]$_SDFF_PN0_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3110),
    .D(_02244_),
    .Q_N(_13036_),
    .Q(\cpu.icache.r_offset[1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_offset[2]$_SDFF_PN0_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3111),
    .D(_02245_),
    .Q_N(_00232_),
    .Q(\cpu.icache.r_offset[2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net3112),
    .D(_02246_),
    .Q_N(_13035_),
    .Q(\cpu.icache.r_tag[0][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net3113),
    .D(_02247_),
    .Q_N(_13034_),
    .Q(\cpu.icache.r_tag[0][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net3114),
    .D(_02248_),
    .Q_N(_13033_),
    .Q(\cpu.icache.r_tag[0][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net3115),
    .D(_02249_),
    .Q_N(_13032_),
    .Q(\cpu.icache.r_tag[0][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net3116),
    .D(_02250_),
    .Q_N(_13031_),
    .Q(\cpu.icache.r_tag[0][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net3117),
    .D(_02251_),
    .Q_N(_13030_),
    .Q(\cpu.icache.r_tag[0][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3118),
    .D(_02252_),
    .Q_N(_13029_),
    .Q(\cpu.icache.r_tag[0][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net3119),
    .D(_02253_),
    .Q_N(_13028_),
    .Q(\cpu.icache.r_tag[0][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net3120),
    .D(_02254_),
    .Q_N(_13027_),
    .Q(\cpu.icache.r_tag[0][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net3121),
    .D(_02255_),
    .Q_N(_13026_),
    .Q(\cpu.icache.r_tag[0][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net3122),
    .D(_02256_),
    .Q_N(_13025_),
    .Q(\cpu.icache.r_tag[0][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net3123),
    .D(_02257_),
    .Q_N(_13024_),
    .Q(\cpu.icache.r_tag[0][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net3124),
    .D(_02258_),
    .Q_N(_13023_),
    .Q(\cpu.icache.r_tag[0][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net3125),
    .D(_02259_),
    .Q_N(_13022_),
    .Q(\cpu.icache.r_tag[0][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net3126),
    .D(_02260_),
    .Q_N(_13021_),
    .Q(\cpu.icache.r_tag[0][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net3127),
    .D(_02261_),
    .Q_N(_13020_),
    .Q(\cpu.icache.r_tag[0][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net3128),
    .D(_02262_),
    .Q_N(_13019_),
    .Q(\cpu.icache.r_tag[0][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net3129),
    .D(_02263_),
    .Q_N(_13018_),
    .Q(\cpu.icache.r_tag[0][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net3130),
    .D(_02264_),
    .Q_N(_13017_),
    .Q(\cpu.icache.r_tag[0][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net3131),
    .D(_02265_),
    .Q_N(_13016_),
    .Q(\cpu.icache.r_tag[1][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net3132),
    .D(_02266_),
    .Q_N(_13015_),
    .Q(\cpu.icache.r_tag[1][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net3133),
    .D(_02267_),
    .Q_N(_13014_),
    .Q(\cpu.icache.r_tag[1][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net3134),
    .D(_02268_),
    .Q_N(_13013_),
    .Q(\cpu.icache.r_tag[1][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net3135),
    .D(_02269_),
    .Q_N(_13012_),
    .Q(\cpu.icache.r_tag[1][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3136),
    .D(_02270_),
    .Q_N(_13011_),
    .Q(\cpu.icache.r_tag[1][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3137),
    .D(_02271_),
    .Q_N(_13010_),
    .Q(\cpu.icache.r_tag[1][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3138),
    .D(_02272_),
    .Q_N(_13009_),
    .Q(\cpu.icache.r_tag[1][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net3139),
    .D(_02273_),
    .Q_N(_13008_),
    .Q(\cpu.icache.r_tag[1][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3140),
    .D(_02274_),
    .Q_N(_13007_),
    .Q(\cpu.icache.r_tag[1][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net3141),
    .D(_02275_),
    .Q_N(_13006_),
    .Q(\cpu.icache.r_tag[1][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net3142),
    .D(_02276_),
    .Q_N(_13005_),
    .Q(\cpu.icache.r_tag[1][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net3143),
    .D(_02277_),
    .Q_N(_13004_),
    .Q(\cpu.icache.r_tag[1][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net3144),
    .D(_02278_),
    .Q_N(_13003_),
    .Q(\cpu.icache.r_tag[1][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net3145),
    .D(_02279_),
    .Q_N(_13002_),
    .Q(\cpu.icache.r_tag[1][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net3146),
    .D(_02280_),
    .Q_N(_13001_),
    .Q(\cpu.icache.r_tag[1][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net3147),
    .D(_02281_),
    .Q_N(_13000_),
    .Q(\cpu.icache.r_tag[1][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net3148),
    .D(_02282_),
    .Q_N(_12999_),
    .Q(\cpu.icache.r_tag[1][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net3149),
    .D(_02283_),
    .Q_N(_12998_),
    .Q(\cpu.icache.r_tag[1][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net3150),
    .D(_02284_),
    .Q_N(_12997_),
    .Q(\cpu.icache.r_tag[2][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net3151),
    .D(_02285_),
    .Q_N(_12996_),
    .Q(\cpu.icache.r_tag[2][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net3152),
    .D(_02286_),
    .Q_N(_12995_),
    .Q(\cpu.icache.r_tag[2][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net3153),
    .D(_02287_),
    .Q_N(_12994_),
    .Q(\cpu.icache.r_tag[2][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net3154),
    .D(_02288_),
    .Q_N(_12993_),
    .Q(\cpu.icache.r_tag[2][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3155),
    .D(_02289_),
    .Q_N(_12992_),
    .Q(\cpu.icache.r_tag[2][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3156),
    .D(_02290_),
    .Q_N(_12991_),
    .Q(\cpu.icache.r_tag[2][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3157),
    .D(_02291_),
    .Q_N(_12990_),
    .Q(\cpu.icache.r_tag[2][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net3158),
    .D(_02292_),
    .Q_N(_12989_),
    .Q(\cpu.icache.r_tag[2][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net3159),
    .D(_02293_),
    .Q_N(_12988_),
    .Q(\cpu.icache.r_tag[2][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net3160),
    .D(_02294_),
    .Q_N(_12987_),
    .Q(\cpu.icache.r_tag[2][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net3161),
    .D(_02295_),
    .Q_N(_12986_),
    .Q(\cpu.icache.r_tag[2][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net3162),
    .D(_02296_),
    .Q_N(_12985_),
    .Q(\cpu.icache.r_tag[2][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net3163),
    .D(_02297_),
    .Q_N(_12984_),
    .Q(\cpu.icache.r_tag[2][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net3164),
    .D(_02298_),
    .Q_N(_12983_),
    .Q(\cpu.icache.r_tag[2][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net3165),
    .D(_02299_),
    .Q_N(_12982_),
    .Q(\cpu.icache.r_tag[2][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net3166),
    .D(_02300_),
    .Q_N(_12981_),
    .Q(\cpu.icache.r_tag[2][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net3167),
    .D(_02301_),
    .Q_N(_12980_),
    .Q(\cpu.icache.r_tag[2][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net3168),
    .D(_02302_),
    .Q_N(_12979_),
    .Q(\cpu.icache.r_tag[2][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net3169),
    .D(_02303_),
    .Q_N(_12978_),
    .Q(\cpu.icache.r_tag[3][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net3170),
    .D(_02304_),
    .Q_N(_12977_),
    .Q(\cpu.icache.r_tag[3][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3171),
    .D(_02305_),
    .Q_N(_12976_),
    .Q(\cpu.icache.r_tag[3][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net3172),
    .D(_02306_),
    .Q_N(_12975_),
    .Q(\cpu.icache.r_tag[3][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net3173),
    .D(_02307_),
    .Q_N(_12974_),
    .Q(\cpu.icache.r_tag[3][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3174),
    .D(_02308_),
    .Q_N(_12973_),
    .Q(\cpu.icache.r_tag[3][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3175),
    .D(_02309_),
    .Q_N(_12972_),
    .Q(\cpu.icache.r_tag[3][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net3176),
    .D(_02310_),
    .Q_N(_12971_),
    .Q(\cpu.icache.r_tag[3][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net3177),
    .D(_02311_),
    .Q_N(_12970_),
    .Q(\cpu.icache.r_tag[3][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net3178),
    .D(_02312_),
    .Q_N(_12969_),
    .Q(\cpu.icache.r_tag[3][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net3179),
    .D(_02313_),
    .Q_N(_12968_),
    .Q(\cpu.icache.r_tag[3][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net3180),
    .D(_02314_),
    .Q_N(_12967_),
    .Q(\cpu.icache.r_tag[3][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net3181),
    .D(_02315_),
    .Q_N(_12966_),
    .Q(\cpu.icache.r_tag[3][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net3182),
    .D(_02316_),
    .Q_N(_12965_),
    .Q(\cpu.icache.r_tag[3][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net3183),
    .D(_02317_),
    .Q_N(_12964_),
    .Q(\cpu.icache.r_tag[3][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net3184),
    .D(_02318_),
    .Q_N(_12963_),
    .Q(\cpu.icache.r_tag[3][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net3185),
    .D(_02319_),
    .Q_N(_12962_),
    .Q(\cpu.icache.r_tag[3][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net3186),
    .D(_02320_),
    .Q_N(_12961_),
    .Q(\cpu.icache.r_tag[3][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net3187),
    .D(_02321_),
    .Q_N(_12960_),
    .Q(\cpu.icache.r_tag[3][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net3188),
    .D(_02322_),
    .Q_N(_12959_),
    .Q(\cpu.icache.r_tag[4][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net3189),
    .D(_02323_),
    .Q_N(_12958_),
    .Q(\cpu.icache.r_tag[4][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net3190),
    .D(_02324_),
    .Q_N(_12957_),
    .Q(\cpu.icache.r_tag[4][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net3191),
    .D(_02325_),
    .Q_N(_12956_),
    .Q(\cpu.icache.r_tag[4][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net3192),
    .D(_02326_),
    .Q_N(_12955_),
    .Q(\cpu.icache.r_tag[4][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3193),
    .D(_02327_),
    .Q_N(_12954_),
    .Q(\cpu.icache.r_tag[4][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3194),
    .D(_02328_),
    .Q_N(_12953_),
    .Q(\cpu.icache.r_tag[4][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3195),
    .D(_02329_),
    .Q_N(_12952_),
    .Q(\cpu.icache.r_tag[4][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net3196),
    .D(_02330_),
    .Q_N(_12951_),
    .Q(\cpu.icache.r_tag[4][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3197),
    .D(_02331_),
    .Q_N(_12950_),
    .Q(\cpu.icache.r_tag[4][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net3198),
    .D(_02332_),
    .Q_N(_12949_),
    .Q(\cpu.icache.r_tag[4][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net3199),
    .D(_02333_),
    .Q_N(_12948_),
    .Q(\cpu.icache.r_tag[4][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net3200),
    .D(_02334_),
    .Q_N(_12947_),
    .Q(\cpu.icache.r_tag[4][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net3201),
    .D(_02335_),
    .Q_N(_12946_),
    .Q(\cpu.icache.r_tag[4][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net3202),
    .D(_02336_),
    .Q_N(_12945_),
    .Q(\cpu.icache.r_tag[4][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net3203),
    .D(_02337_),
    .Q_N(_12944_),
    .Q(\cpu.icache.r_tag[4][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net3204),
    .D(_02338_),
    .Q_N(_12943_),
    .Q(\cpu.icache.r_tag[4][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net3205),
    .D(_02339_),
    .Q_N(_12942_),
    .Q(\cpu.icache.r_tag[4][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net3206),
    .D(_02340_),
    .Q_N(_12941_),
    .Q(\cpu.icache.r_tag[4][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net3207),
    .D(_02341_),
    .Q_N(_12940_),
    .Q(\cpu.icache.r_tag[5][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net3208),
    .D(_02342_),
    .Q_N(_12939_),
    .Q(\cpu.icache.r_tag[5][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3209),
    .D(_02343_),
    .Q_N(_12938_),
    .Q(\cpu.icache.r_tag[5][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net3210),
    .D(_02344_),
    .Q_N(_12937_),
    .Q(\cpu.icache.r_tag[5][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3211),
    .D(_02345_),
    .Q_N(_12936_),
    .Q(\cpu.icache.r_tag[5][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3212),
    .D(_02346_),
    .Q_N(_12935_),
    .Q(\cpu.icache.r_tag[5][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3213),
    .D(_02347_),
    .Q_N(_12934_),
    .Q(\cpu.icache.r_tag[5][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net3214),
    .D(_02348_),
    .Q_N(_12933_),
    .Q(\cpu.icache.r_tag[5][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net3215),
    .D(_02349_),
    .Q_N(_12932_),
    .Q(\cpu.icache.r_tag[5][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net3216),
    .D(_02350_),
    .Q_N(_12931_),
    .Q(\cpu.icache.r_tag[5][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net3217),
    .D(_02351_),
    .Q_N(_12930_),
    .Q(\cpu.icache.r_tag[5][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net3218),
    .D(_02352_),
    .Q_N(_12929_),
    .Q(\cpu.icache.r_tag[5][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net3219),
    .D(_02353_),
    .Q_N(_12928_),
    .Q(\cpu.icache.r_tag[5][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net3220),
    .D(_02354_),
    .Q_N(_12927_),
    .Q(\cpu.icache.r_tag[5][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net3221),
    .D(_02355_),
    .Q_N(_12926_),
    .Q(\cpu.icache.r_tag[5][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net3222),
    .D(_02356_),
    .Q_N(_12925_),
    .Q(\cpu.icache.r_tag[5][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net3223),
    .D(_02357_),
    .Q_N(_12924_),
    .Q(\cpu.icache.r_tag[5][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net3224),
    .D(_02358_),
    .Q_N(_12923_),
    .Q(\cpu.icache.r_tag[5][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net3225),
    .D(_02359_),
    .Q_N(_12922_),
    .Q(\cpu.icache.r_tag[5][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net3226),
    .D(_02360_),
    .Q_N(_12921_),
    .Q(\cpu.icache.r_tag[6][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net3227),
    .D(_02361_),
    .Q_N(_12920_),
    .Q(\cpu.icache.r_tag[6][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net3228),
    .D(_02362_),
    .Q_N(_12919_),
    .Q(\cpu.icache.r_tag[6][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3229),
    .D(_02363_),
    .Q_N(_12918_),
    .Q(\cpu.icache.r_tag[6][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net3230),
    .D(_02364_),
    .Q_N(_12917_),
    .Q(\cpu.icache.r_tag[6][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3231),
    .D(_02365_),
    .Q_N(_12916_),
    .Q(\cpu.icache.r_tag[6][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3232),
    .D(_02366_),
    .Q_N(_12915_),
    .Q(\cpu.icache.r_tag[6][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net3233),
    .D(_02367_),
    .Q_N(_12914_),
    .Q(\cpu.icache.r_tag[6][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net3234),
    .D(_02368_),
    .Q_N(_12913_),
    .Q(\cpu.icache.r_tag[6][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net3235),
    .D(_02369_),
    .Q_N(_12912_),
    .Q(\cpu.icache.r_tag[6][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net3236),
    .D(_02370_),
    .Q_N(_12911_),
    .Q(\cpu.icache.r_tag[6][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net3237),
    .D(_02371_),
    .Q_N(_12910_),
    .Q(\cpu.icache.r_tag[6][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net3238),
    .D(_02372_),
    .Q_N(_12909_),
    .Q(\cpu.icache.r_tag[6][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net3239),
    .D(_02373_),
    .Q_N(_12908_),
    .Q(\cpu.icache.r_tag[6][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net3240),
    .D(_02374_),
    .Q_N(_12907_),
    .Q(\cpu.icache.r_tag[6][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net3241),
    .D(_02375_),
    .Q_N(_12906_),
    .Q(\cpu.icache.r_tag[6][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net3242),
    .D(_02376_),
    .Q_N(_12905_),
    .Q(\cpu.icache.r_tag[6][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net3243),
    .D(_02377_),
    .Q_N(_12904_),
    .Q(\cpu.icache.r_tag[6][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net3244),
    .D(_02378_),
    .Q_N(_12903_),
    .Q(\cpu.icache.r_tag[6][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net3245),
    .D(_02379_),
    .Q_N(_12902_),
    .Q(\cpu.icache.r_tag[7][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net3246),
    .D(_02380_),
    .Q_N(_12901_),
    .Q(\cpu.icache.r_tag[7][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3247),
    .D(_02381_),
    .Q_N(_12900_),
    .Q(\cpu.icache.r_tag[7][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net3248),
    .D(_02382_),
    .Q_N(_12899_),
    .Q(\cpu.icache.r_tag[7][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3249),
    .D(_02383_),
    .Q_N(_12898_),
    .Q(\cpu.icache.r_tag[7][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3250),
    .D(_02384_),
    .Q_N(_12897_),
    .Q(\cpu.icache.r_tag[7][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3251),
    .D(_02385_),
    .Q_N(_12896_),
    .Q(\cpu.icache.r_tag[7][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3252),
    .D(_02386_),
    .Q_N(_12895_),
    .Q(\cpu.icache.r_tag[7][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net3253),
    .D(_02387_),
    .Q_N(_12894_),
    .Q(\cpu.icache.r_tag[7][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net3254),
    .D(_02388_),
    .Q_N(_12893_),
    .Q(\cpu.icache.r_tag[7][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net3255),
    .D(_02389_),
    .Q_N(_12892_),
    .Q(\cpu.icache.r_tag[7][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net3256),
    .D(_02390_),
    .Q_N(_12891_),
    .Q(\cpu.icache.r_tag[7][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net3257),
    .D(_02391_),
    .Q_N(_12890_),
    .Q(\cpu.icache.r_tag[7][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net3258),
    .D(_02392_),
    .Q_N(_12889_),
    .Q(\cpu.icache.r_tag[7][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net3259),
    .D(_02393_),
    .Q_N(_12888_),
    .Q(\cpu.icache.r_tag[7][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net3260),
    .D(_02394_),
    .Q_N(_12887_),
    .Q(\cpu.icache.r_tag[7][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net3261),
    .D(_02395_),
    .Q_N(_12886_),
    .Q(\cpu.icache.r_tag[7][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net3262),
    .D(_02396_),
    .Q_N(_12885_),
    .Q(\cpu.icache.r_tag[7][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net3263),
    .D(_02397_),
    .Q_N(_12884_),
    .Q(\cpu.icache.r_tag[7][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3264),
    .D(_02398_),
    .Q_N(_12883_),
    .Q(\cpu.icache.r_valid[0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3265),
    .D(_02399_),
    .Q_N(_12882_),
    .Q(\cpu.icache.r_valid[1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3266),
    .D(_02400_),
    .Q_N(_12881_),
    .Q(\cpu.icache.r_valid[2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3267),
    .D(_02401_),
    .Q_N(_12880_),
    .Q(\cpu.icache.r_valid[3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3268),
    .D(_02402_),
    .Q_N(_12879_),
    .Q(\cpu.icache.r_valid[4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3269),
    .D(_02403_),
    .Q_N(_12878_),
    .Q(\cpu.icache.r_valid[5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3270),
    .D(_02404_),
    .Q_N(_12877_),
    .Q(\cpu.icache.r_valid[6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3271),
    .D(_02405_),
    .Q_N(_12876_),
    .Q(\cpu.icache.r_valid[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3272),
    .D(_02406_),
    .Q_N(_12875_),
    .Q(\cpu.intr.r_clock ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[0]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3273),
    .D(_02407_),
    .Q_N(_12874_),
    .Q(\cpu.intr.r_clock_cmp[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[10]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3274),
    .D(_02408_),
    .Q_N(_12873_),
    .Q(\cpu.intr.r_clock_cmp[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[11]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3275),
    .D(_02409_),
    .Q_N(_12872_),
    .Q(\cpu.intr.r_clock_cmp[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[12]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3276),
    .D(_02410_),
    .Q_N(_12871_),
    .Q(\cpu.intr.r_clock_cmp[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[13]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3277),
    .D(_02411_),
    .Q_N(_12870_),
    .Q(\cpu.intr.r_clock_cmp[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[14]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3278),
    .D(_02412_),
    .Q_N(_12869_),
    .Q(\cpu.intr.r_clock_cmp[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[15]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3279),
    .D(_02413_),
    .Q_N(_12868_),
    .Q(\cpu.intr.r_clock_cmp[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[16]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3280),
    .D(_02414_),
    .Q_N(_12867_),
    .Q(\cpu.intr.r_clock_cmp[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[17]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3281),
    .D(_02415_),
    .Q_N(_12866_),
    .Q(\cpu.intr.r_clock_cmp[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[18]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3282),
    .D(_02416_),
    .Q_N(_12865_),
    .Q(\cpu.intr.r_clock_cmp[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[19]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3283),
    .D(_02417_),
    .Q_N(_12864_),
    .Q(\cpu.intr.r_clock_cmp[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[1]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3284),
    .D(_02418_),
    .Q_N(_12863_),
    .Q(\cpu.intr.r_clock_cmp[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[20]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3285),
    .D(_02419_),
    .Q_N(_12862_),
    .Q(\cpu.intr.r_clock_cmp[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[21]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3286),
    .D(_02420_),
    .Q_N(_12861_),
    .Q(\cpu.intr.r_clock_cmp[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[22]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3287),
    .D(_02421_),
    .Q_N(_12860_),
    .Q(\cpu.intr.r_clock_cmp[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[23]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3288),
    .D(_02422_),
    .Q_N(_12859_),
    .Q(\cpu.intr.r_clock_cmp[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[24]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3289),
    .D(_02423_),
    .Q_N(_12858_),
    .Q(\cpu.intr.r_clock_cmp[24] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[25]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3290),
    .D(_02424_),
    .Q_N(_12857_),
    .Q(\cpu.intr.r_clock_cmp[25] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[26]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3291),
    .D(_02425_),
    .Q_N(_12856_),
    .Q(\cpu.intr.r_clock_cmp[26] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[27]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3292),
    .D(_02426_),
    .Q_N(_12855_),
    .Q(\cpu.intr.r_clock_cmp[27] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[28]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3293),
    .D(_02427_),
    .Q_N(_12854_),
    .Q(\cpu.intr.r_clock_cmp[28] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[29]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3294),
    .D(_02428_),
    .Q_N(_12853_),
    .Q(\cpu.intr.r_clock_cmp[29] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[2]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3295),
    .D(_02429_),
    .Q_N(_12852_),
    .Q(\cpu.intr.r_clock_cmp[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[30]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3296),
    .D(_02430_),
    .Q_N(_12851_),
    .Q(\cpu.intr.r_clock_cmp[30] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[31]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3297),
    .D(_02431_),
    .Q_N(_12850_),
    .Q(\cpu.intr.r_clock_cmp[31] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[3]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3298),
    .D(_02432_),
    .Q_N(_12849_),
    .Q(\cpu.intr.r_clock_cmp[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[4]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3299),
    .D(_02433_),
    .Q_N(_12848_),
    .Q(\cpu.intr.r_clock_cmp[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[5]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3300),
    .D(_02434_),
    .Q_N(_12847_),
    .Q(\cpu.intr.r_clock_cmp[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[6]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3301),
    .D(_02435_),
    .Q_N(_12846_),
    .Q(\cpu.intr.r_clock_cmp[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[7]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3302),
    .D(_02436_),
    .Q_N(_12845_),
    .Q(\cpu.intr.r_clock_cmp[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[8]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3303),
    .D(_02437_),
    .Q_N(_12844_),
    .Q(\cpu.intr.r_clock_cmp[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[9]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3304),
    .D(_02438_),
    .Q_N(_14856_),
    .Q(\cpu.intr.r_clock_cmp[9] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[0]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3305),
    .D(_00036_),
    .Q_N(_00265_),
    .Q(\cpu.intr.r_clock_count[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[10]$_DFF_P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3306),
    .D(_00037_),
    .Q_N(_14857_),
    .Q(\cpu.intr.r_clock_count[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[11]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3307),
    .D(_00038_),
    .Q_N(_14858_),
    .Q(\cpu.intr.r_clock_count[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[12]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3308),
    .D(_00039_),
    .Q_N(_14859_),
    .Q(\cpu.intr.r_clock_count[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[13]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3309),
    .D(_00040_),
    .Q_N(_14860_),
    .Q(\cpu.intr.r_clock_count[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[14]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3310),
    .D(_00041_),
    .Q_N(_14861_),
    .Q(\cpu.intr.r_clock_count[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[15]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net3311),
    .D(_00042_),
    .Q_N(_12843_),
    .Q(\cpu.intr.r_clock_count[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[16]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3312),
    .D(_02439_),
    .Q_N(_12842_),
    .Q(\cpu.intr.r_clock_count[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[17]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3313),
    .D(_02440_),
    .Q_N(_12841_),
    .Q(\cpu.intr.r_clock_count[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[18]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3314),
    .D(_02441_),
    .Q_N(_12840_),
    .Q(\cpu.intr.r_clock_count[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[19]$_DFFE_PN_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3315),
    .D(_02442_),
    .Q_N(_14862_),
    .Q(\cpu.intr.r_clock_count[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[1]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3316),
    .D(_00043_),
    .Q_N(_12839_),
    .Q(\cpu.intr.r_clock_count[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[20]$_DFFE_PN_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3317),
    .D(_02443_),
    .Q_N(_12838_),
    .Q(\cpu.intr.r_clock_count[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[21]$_DFFE_PN_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3318),
    .D(_02444_),
    .Q_N(_12837_),
    .Q(\cpu.intr.r_clock_count[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[22]$_DFFE_PN_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3319),
    .D(_02445_),
    .Q_N(_12836_),
    .Q(\cpu.intr.r_clock_count[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[23]$_DFFE_PN_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net3320),
    .D(_02446_),
    .Q_N(_12835_),
    .Q(\cpu.intr.r_clock_count[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[24]$_DFFE_PN_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3321),
    .D(_02447_),
    .Q_N(_12834_),
    .Q(\cpu.intr.r_clock_count[24] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[25]$_DFFE_PN_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3322),
    .D(_02448_),
    .Q_N(_12833_),
    .Q(\cpu.intr.r_clock_count[25] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[26]$_DFFE_PN_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3323),
    .D(_02449_),
    .Q_N(_12832_),
    .Q(\cpu.intr.r_clock_count[26] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[27]$_DFFE_PN_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3324),
    .D(_02450_),
    .Q_N(_12831_),
    .Q(\cpu.intr.r_clock_count[27] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[28]$_DFFE_PN_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3325),
    .D(_02451_),
    .Q_N(_12830_),
    .Q(\cpu.intr.r_clock_count[28] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[29]$_DFFE_PN_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3326),
    .D(_02452_),
    .Q_N(_14863_),
    .Q(\cpu.intr.r_clock_count[29] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[2]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3327),
    .D(_00044_),
    .Q_N(_12829_),
    .Q(\cpu.intr.r_clock_count[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[30]$_DFFE_PN_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net3328),
    .D(_02453_),
    .Q_N(_12828_),
    .Q(\cpu.intr.r_clock_count[30] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[31]$_DFFE_PN_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3329),
    .D(_02454_),
    .Q_N(_14864_),
    .Q(\cpu.intr.r_clock_count[31] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[3]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3330),
    .D(_00045_),
    .Q_N(_14865_),
    .Q(\cpu.intr.r_clock_count[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[4]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3331),
    .D(_00046_),
    .Q_N(_14866_),
    .Q(\cpu.intr.r_clock_count[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[5]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3332),
    .D(_00047_),
    .Q_N(_14867_),
    .Q(\cpu.intr.r_clock_count[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[6]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3333),
    .D(_00048_),
    .Q_N(_14868_),
    .Q(\cpu.intr.r_clock_count[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[7]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3334),
    .D(_00049_),
    .Q_N(_14869_),
    .Q(\cpu.intr.r_clock_count[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[8]$_DFF_P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3335),
    .D(_00050_),
    .Q_N(_14870_),
    .Q(\cpu.intr.r_clock_count[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[9]$_DFF_P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3336),
    .D(_00051_),
    .Q_N(_12827_),
    .Q(\cpu.intr.r_clock_count[9] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3337),
    .D(_02455_),
    .Q_N(_12826_),
    .Q(\cpu.intr.r_enable[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3338),
    .D(_02456_),
    .Q_N(_12825_),
    .Q(\cpu.intr.r_enable[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3339),
    .D(_02457_),
    .Q_N(_12824_),
    .Q(\cpu.intr.r_enable[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3340),
    .D(_02458_),
    .Q_N(_12823_),
    .Q(\cpu.intr.r_enable[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3341),
    .D(_02459_),
    .Q_N(_12822_),
    .Q(\cpu.intr.r_enable[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3342),
    .D(_02460_),
    .Q_N(_12821_),
    .Q(\cpu.intr.r_enable[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3343),
    .D(_02461_),
    .Q_N(_14871_),
    .Q(\cpu.intr.r_timer ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[0]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3344),
    .D(_00055_),
    .Q_N(_00264_),
    .Q(\cpu.intr.r_timer_count[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[10]$_DFF_P_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net3345),
    .D(_00056_),
    .Q_N(_14872_),
    .Q(\cpu.intr.r_timer_count[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[11]$_DFF_P_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net3346),
    .D(_00057_),
    .Q_N(_14873_),
    .Q(\cpu.intr.r_timer_count[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[12]$_DFF_P_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net3347),
    .D(_00058_),
    .Q_N(_14874_),
    .Q(\cpu.intr.r_timer_count[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[13]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3348),
    .D(_00059_),
    .Q_N(_14875_),
    .Q(\cpu.intr.r_timer_count[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[14]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3349),
    .D(_00060_),
    .Q_N(_14876_),
    .Q(\cpu.intr.r_timer_count[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[15]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3350),
    .D(_00061_),
    .Q_N(_14877_),
    .Q(\cpu.intr.r_timer_count[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[16]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3351),
    .D(_00062_),
    .Q_N(_14878_),
    .Q(\cpu.intr.r_timer_count[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[17]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3352),
    .D(_00063_),
    .Q_N(_14879_),
    .Q(\cpu.intr.r_timer_count[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[18]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3353),
    .D(_00064_),
    .Q_N(_14880_),
    .Q(\cpu.intr.r_timer_count[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[19]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3354),
    .D(_00065_),
    .Q_N(_14881_),
    .Q(\cpu.intr.r_timer_count[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[1]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3355),
    .D(_00066_),
    .Q_N(_14882_),
    .Q(\cpu.intr.r_timer_count[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[20]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3356),
    .D(_00067_),
    .Q_N(_14883_),
    .Q(\cpu.intr.r_timer_count[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[21]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3357),
    .D(_00068_),
    .Q_N(_14884_),
    .Q(\cpu.intr.r_timer_count[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[22]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3358),
    .D(_00069_),
    .Q_N(_14885_),
    .Q(\cpu.intr.r_timer_count[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[23]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3359),
    .D(_00070_),
    .Q_N(_14886_),
    .Q(\cpu.intr.r_timer_count[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[2]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3360),
    .D(_00071_),
    .Q_N(_14887_),
    .Q(\cpu.intr.r_timer_count[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[3]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3361),
    .D(_00072_),
    .Q_N(_14888_),
    .Q(\cpu.intr.r_timer_count[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[4]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3362),
    .D(_00073_),
    .Q_N(_14889_),
    .Q(\cpu.intr.r_timer_count[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[5]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3363),
    .D(_00074_),
    .Q_N(_14890_),
    .Q(\cpu.intr.r_timer_count[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[6]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3364),
    .D(_00075_),
    .Q_N(_14891_),
    .Q(\cpu.intr.r_timer_count[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[7]$_DFF_P_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net3365),
    .D(_00076_),
    .Q_N(_14892_),
    .Q(\cpu.intr.r_timer_count[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[8]$_DFF_P_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net3366),
    .D(_00077_),
    .Q_N(_14893_),
    .Q(\cpu.intr.r_timer_count[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[9]$_DFF_P_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net3367),
    .D(_00078_),
    .Q_N(_12820_),
    .Q(\cpu.intr.r_timer_count[9] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[0]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3368),
    .D(_02462_),
    .Q_N(_12819_),
    .Q(\cpu.intr.r_timer_reload[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[10]$_DFFE_PP_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net3369),
    .D(_02463_),
    .Q_N(_12818_),
    .Q(\cpu.intr.r_timer_reload[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[11]$_DFFE_PP_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net3370),
    .D(_02464_),
    .Q_N(_12817_),
    .Q(\cpu.intr.r_timer_reload[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[12]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3371),
    .D(_02465_),
    .Q_N(_12816_),
    .Q(\cpu.intr.r_timer_reload[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[13]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3372),
    .D(_02466_),
    .Q_N(_12815_),
    .Q(\cpu.intr.r_timer_reload[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[14]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3373),
    .D(_02467_),
    .Q_N(_12814_),
    .Q(\cpu.intr.r_timer_reload[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[15]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3374),
    .D(_02468_),
    .Q_N(_12813_),
    .Q(\cpu.intr.r_timer_reload[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[16]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3375),
    .D(_02469_),
    .Q_N(_12812_),
    .Q(\cpu.intr.r_timer_reload[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[17]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3376),
    .D(_02470_),
    .Q_N(_12811_),
    .Q(\cpu.intr.r_timer_reload[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[18]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3377),
    .D(_02471_),
    .Q_N(_12810_),
    .Q(\cpu.intr.r_timer_reload[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[19]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3378),
    .D(_02472_),
    .Q_N(_12809_),
    .Q(\cpu.intr.r_timer_reload[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[1]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3379),
    .D(_02473_),
    .Q_N(_12808_),
    .Q(\cpu.intr.r_timer_reload[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[20]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3380),
    .D(_02474_),
    .Q_N(_12807_),
    .Q(\cpu.intr.r_timer_reload[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[21]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3381),
    .D(_02475_),
    .Q_N(_12806_),
    .Q(\cpu.intr.r_timer_reload[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[22]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3382),
    .D(_02476_),
    .Q_N(_12805_),
    .Q(\cpu.intr.r_timer_reload[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[23]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3383),
    .D(_02477_),
    .Q_N(_12804_),
    .Q(\cpu.intr.r_timer_reload[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[2]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3384),
    .D(_02478_),
    .Q_N(_12803_),
    .Q(\cpu.intr.r_timer_reload[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[3]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3385),
    .D(_02479_),
    .Q_N(_12802_),
    .Q(\cpu.intr.r_timer_reload[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[4]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3386),
    .D(_02480_),
    .Q_N(_12801_),
    .Q(\cpu.intr.r_timer_reload[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[5]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3387),
    .D(_02481_),
    .Q_N(_12800_),
    .Q(\cpu.intr.r_timer_reload[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[6]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3388),
    .D(_02482_),
    .Q_N(_12799_),
    .Q(\cpu.intr.r_timer_reload[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[7]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3389),
    .D(_02483_),
    .Q_N(_12798_),
    .Q(\cpu.intr.r_timer_reload[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[8]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3390),
    .D(_02484_),
    .Q_N(_12797_),
    .Q(\cpu.intr.r_timer_reload[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[9]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3391),
    .D(_02485_),
    .Q_N(_12796_),
    .Q(\cpu.intr.r_timer_reload[9] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[0]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3392),
    .D(_02486_),
    .Q_N(_00167_),
    .Q(\cpu.qspi.r_count[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[1]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3393),
    .D(_02487_),
    .Q_N(_12795_),
    .Q(\cpu.qspi.r_count[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[2]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3394),
    .D(_02488_),
    .Q_N(_00168_),
    .Q(\cpu.qspi.r_count[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[3]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3395),
    .D(_02489_),
    .Q_N(_12794_),
    .Q(\cpu.qspi.r_count[3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[4]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3396),
    .D(_02490_),
    .Q_N(_00230_),
    .Q(\cpu.qspi.r_count[4] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_cs[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3397),
    .D(_02491_),
    .Q_N(_12793_),
    .Q(net19));
 sg13g2_dfrbp_1 \cpu.qspi.r_cs[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3398),
    .D(_02492_),
    .Q_N(_12792_),
    .Q(net20));
 sg13g2_dfrbp_1 \cpu.qspi.r_cs[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3399),
    .D(_02493_),
    .Q_N(_12791_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[11] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_ind$_SDFFE_PN0N_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3400),
    .D(_02494_),
    .Q_N(_12790_),
    .Q(\cpu.qspi.r_ind ));
 sg13g2_dfrbp_1 \cpu.qspi.r_mask[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3401),
    .D(_02495_),
    .Q_N(_12789_),
    .Q(\cpu.qspi.r_mask[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_mask[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3402),
    .D(_02496_),
    .Q_N(_12788_),
    .Q(\cpu.qspi.r_mask[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_mask[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3403),
    .D(_02497_),
    .Q_N(_12787_),
    .Q(\cpu.qspi.r_mask[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_quad[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3404),
    .D(_02498_),
    .Q_N(_12786_),
    .Q(\cpu.qspi.r_quad[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_quad[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3405),
    .D(_02499_),
    .Q_N(_12785_),
    .Q(\cpu.qspi.r_quad[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_quad[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3406),
    .D(_02500_),
    .Q_N(_12784_),
    .Q(\cpu.qspi.r_quad[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3407),
    .D(_02501_),
    .Q_N(_12783_),
    .Q(\cpu.qspi.r_read_delay[0][0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3408),
    .D(_02502_),
    .Q_N(_12782_),
    .Q(\cpu.qspi.r_read_delay[0][1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][2]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3409),
    .D(_02503_),
    .Q_N(_12781_),
    .Q(\cpu.qspi.r_read_delay[0][2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3410),
    .D(_02504_),
    .Q_N(_12780_),
    .Q(\cpu.qspi.r_read_delay[0][3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3411),
    .D(_02505_),
    .Q_N(_12779_),
    .Q(\cpu.qspi.r_read_delay[1][0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3412),
    .D(_02506_),
    .Q_N(_12778_),
    .Q(\cpu.qspi.r_read_delay[1][1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][2]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3413),
    .D(_02507_),
    .Q_N(_12777_),
    .Q(\cpu.qspi.r_read_delay[1][2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3414),
    .D(_02508_),
    .Q_N(_12776_),
    .Q(\cpu.qspi.r_read_delay[1][3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3415),
    .D(_02509_),
    .Q_N(_12775_),
    .Q(\cpu.qspi.r_read_delay[2][0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net3416),
    .D(_02510_),
    .Q_N(_12774_),
    .Q(\cpu.qspi.r_read_delay[2][1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][2]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3417),
    .D(_02511_),
    .Q_N(_12773_),
    .Q(\cpu.qspi.r_read_delay[2][2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3418),
    .D(_02512_),
    .Q_N(_12772_),
    .Q(\cpu.qspi.r_read_delay[2][3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_rom_mode[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3419),
    .D(_02513_),
    .Q_N(_12771_),
    .Q(\cpu.qspi.r_rom_mode[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_rom_mode[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3420),
    .D(_02514_),
    .Q_N(_14894_),
    .Q(\cpu.qspi.r_rom_mode[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_rstrobe_d$_DFF_P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3421),
    .D(\cpu.qspi.c_rstrobe_d ),
    .Q_N(_14895_),
    .Q(\cpu.d_rstrobe_d ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[0]$_DFF_P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3422),
    .D(_00021_),
    .Q_N(_00257_),
    .Q(\cpu.qspi.r_state[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[10]$_DFF_P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net3423),
    .D(_00008_),
    .Q_N(_14896_),
    .Q(\cpu.qspi.r_state[10] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[11]$_DFF_P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net3424),
    .D(_00022_),
    .Q_N(_14897_),
    .Q(\cpu.qspi.r_state[11] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[12]$_DFF_P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3425),
    .D(_00023_),
    .Q_N(_14898_),
    .Q(\cpu.qspi.r_state[12] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[13]$_DFF_P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net3426),
    .D(_00009_),
    .Q_N(_14899_),
    .Q(\cpu.qspi.r_state[13] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[14]$_DFF_P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3427),
    .D(_00024_),
    .Q_N(_14900_),
    .Q(\cpu.qspi.r_state[14] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[15]$_DFF_P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net3428),
    .D(_00010_),
    .Q_N(_14901_),
    .Q(\cpu.qspi.r_state[15] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[16]$_DFF_P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net3429),
    .D(_00025_),
    .Q_N(_14902_),
    .Q(\cpu.qspi.r_state[16] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[17]$_DFF_P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3430),
    .D(_00026_),
    .Q_N(_14903_),
    .Q(\cpu.qspi.r_state[17] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[1]$_DFF_P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3431),
    .D(_00001_),
    .Q_N(_14904_),
    .Q(\cpu.qspi.r_state[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[2]$_DFF_P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3432),
    .D(_00027_),
    .Q_N(_14905_),
    .Q(\cpu.qspi.r_state[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[3]$_DFF_P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net3433),
    .D(_00002_),
    .Q_N(_14906_),
    .Q(\cpu.qspi.r_state[3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[4]$_DFF_P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3434),
    .D(_00028_),
    .Q_N(_14907_),
    .Q(\cpu.qspi.r_state[4] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[5]$_DFF_P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3435),
    .D(_00003_),
    .Q_N(_14908_),
    .Q(\cpu.qspi.r_state[5] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[6]$_DFF_P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net3436),
    .D(_00004_),
    .Q_N(_14909_),
    .Q(\cpu.qspi.r_state[6] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[7]$_DFF_P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3437),
    .D(_00005_),
    .Q_N(_14910_),
    .Q(\cpu.qspi.r_state[7] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[8]$_DFF_P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net3438),
    .D(_00006_),
    .Q_N(_00169_),
    .Q(\cpu.qspi.r_state[8] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[9]$_DFF_P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3439),
    .D(_00007_),
    .Q_N(_12770_),
    .Q(\cpu.qspi.r_state[9] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_oe[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3440),
    .D(_02515_),
    .Q_N(_12769_),
    .Q(net3));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_oe[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3441),
    .D(_02516_),
    .Q_N(_12768_),
    .Q(net6));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3442),
    .D(_02517_),
    .Q_N(_12767_),
    .Q(net11));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3443),
    .D(_02518_),
    .Q_N(_12766_),
    .Q(net12));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3444),
    .D(_02519_),
    .Q_N(_12765_),
    .Q(net13));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3445),
    .D(_02520_),
    .Q_N(_14911_),
    .Q(net14));
 sg13g2_dfrbp_1 \cpu.qspi.r_wstrobe_d$_DFF_P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net3446),
    .D(\cpu.qspi.c_wstrobe_d ),
    .Q_N(_14912_),
    .Q(\cpu.d_wstrobe_d ));
 sg13g2_dfrbp_1 \cpu.qspi.r_wstrobe_i$_DFF_P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3447),
    .D(\cpu.qspi.c_wstrobe_i ),
    .Q_N(_00231_),
    .Q(\cpu.i_wstrobe_d ));
 sg13g2_dfrbp_1 \cpu.r_clk_invert$_DFFE_PN_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net3448),
    .D(_02521_),
    .Q_N(_12764_),
    .Q(\cpu.r_clk_invert ));
 sg13g2_dfrbp_1 \cpu.spi.r_bits[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3449),
    .D(_02522_),
    .Q_N(_12763_),
    .Q(\cpu.spi.r_bits[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_bits[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3450),
    .D(_02523_),
    .Q_N(_12762_),
    .Q(\cpu.spi.r_bits[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_bits[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3451),
    .D(_02524_),
    .Q_N(_12761_),
    .Q(\cpu.spi.r_bits[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3452),
    .D(_02525_),
    .Q_N(_00281_),
    .Q(\cpu.spi.r_clk_count[0][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3453),
    .D(_02526_),
    .Q_N(_00286_),
    .Q(\cpu.spi.r_clk_count[0][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3454),
    .D(_02527_),
    .Q_N(_00095_),
    .Q(\cpu.spi.r_clk_count[0][2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3455),
    .D(_02528_),
    .Q_N(_00105_),
    .Q(\cpu.spi.r_clk_count[0][3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3456),
    .D(_02529_),
    .Q_N(_00115_),
    .Q(\cpu.spi.r_clk_count[0][4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3457),
    .D(_02530_),
    .Q_N(_00121_),
    .Q(\cpu.spi.r_clk_count[0][5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3458),
    .D(_02531_),
    .Q_N(_00132_),
    .Q(\cpu.spi.r_clk_count[0][6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3459),
    .D(_02532_),
    .Q_N(_00143_),
    .Q(\cpu.spi.r_clk_count[0][7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3460),
    .D(_02533_),
    .Q_N(_00280_),
    .Q(\cpu.spi.r_clk_count[1][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3461),
    .D(_02534_),
    .Q_N(_00285_),
    .Q(\cpu.spi.r_clk_count[1][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3462),
    .D(_02535_),
    .Q_N(_00094_),
    .Q(\cpu.spi.r_clk_count[1][2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3463),
    .D(_02536_),
    .Q_N(_00104_),
    .Q(\cpu.spi.r_clk_count[1][3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3464),
    .D(_02537_),
    .Q_N(_00114_),
    .Q(\cpu.spi.r_clk_count[1][4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3465),
    .D(_02538_),
    .Q_N(_00120_),
    .Q(\cpu.spi.r_clk_count[1][5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3466),
    .D(_02539_),
    .Q_N(_00131_),
    .Q(\cpu.spi.r_clk_count[1][6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3467),
    .D(_02540_),
    .Q_N(_00142_),
    .Q(\cpu.spi.r_clk_count[1][7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3468),
    .D(_02541_),
    .Q_N(_12760_),
    .Q(\cpu.spi.r_clk_count[2][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3469),
    .D(_02542_),
    .Q_N(_12759_),
    .Q(\cpu.spi.r_clk_count[2][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3470),
    .D(_02543_),
    .Q_N(_12758_),
    .Q(\cpu.spi.r_clk_count[2][2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3471),
    .D(_02544_),
    .Q_N(_12757_),
    .Q(\cpu.spi.r_clk_count[2][3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3472),
    .D(_02545_),
    .Q_N(_12756_),
    .Q(\cpu.spi.r_clk_count[2][4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3473),
    .D(_02546_),
    .Q_N(_12755_),
    .Q(\cpu.spi.r_clk_count[2][5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3474),
    .D(_02547_),
    .Q_N(_12754_),
    .Q(\cpu.spi.r_clk_count[2][6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3475),
    .D(_02548_),
    .Q_N(_12753_),
    .Q(\cpu.spi.r_clk_count[2][7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[0]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3476),
    .D(_02549_),
    .Q_N(_12752_),
    .Q(\cpu.spi.r_count[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[1]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3477),
    .D(_02550_),
    .Q_N(_12751_),
    .Q(\cpu.spi.r_count[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[2]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3478),
    .D(_02551_),
    .Q_N(_12750_),
    .Q(\cpu.spi.r_count[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[3]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3479),
    .D(_02552_),
    .Q_N(_12749_),
    .Q(\cpu.spi.r_count[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[4]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3480),
    .D(_02553_),
    .Q_N(_12748_),
    .Q(\cpu.spi.r_count[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[5]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3481),
    .D(_02554_),
    .Q_N(_12747_),
    .Q(\cpu.spi.r_count[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[6]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3482),
    .D(_02555_),
    .Q_N(_12746_),
    .Q(\cpu.spi.r_count[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[7]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3483),
    .D(_02556_),
    .Q_N(_12745_),
    .Q(\cpu.spi.r_count[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_cs[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3484),
    .D(_02557_),
    .Q_N(_12744_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_cs[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3485),
    .D(_02558_),
    .Q_N(_12743_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_cs[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3486),
    .D(_02559_),
    .Q_N(_12742_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[8] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[0]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3487),
    .D(_02560_),
    .Q_N(_12741_),
    .Q(\cpu.spi.r_in[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[1]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3488),
    .D(_02561_),
    .Q_N(_12740_),
    .Q(\cpu.spi.r_in[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[2]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3489),
    .D(_02562_),
    .Q_N(_12739_),
    .Q(\cpu.spi.r_in[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[3]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3490),
    .D(_02563_),
    .Q_N(_12738_),
    .Q(\cpu.spi.r_in[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[4]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3491),
    .D(_02564_),
    .Q_N(_12737_),
    .Q(\cpu.spi.r_in[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[5]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3492),
    .D(_02565_),
    .Q_N(_12736_),
    .Q(\cpu.spi.r_in[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[6]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3493),
    .D(_02566_),
    .Q_N(_12735_),
    .Q(\cpu.spi.r_in[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[7]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3494),
    .D(_02567_),
    .Q_N(_00200_),
    .Q(\cpu.spi.r_in[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_interrupt$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3495),
    .D(_02568_),
    .Q_N(_12734_),
    .Q(\cpu.intr.spi_intr ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3496),
    .D(_02569_),
    .Q_N(_00203_),
    .Q(\cpu.spi.r_mode[0][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3497),
    .D(_02570_),
    .Q_N(_12733_),
    .Q(\cpu.spi.r_mode[0][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3498),
    .D(_02571_),
    .Q_N(_12732_),
    .Q(\cpu.spi.r_mode[1][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3499),
    .D(_02572_),
    .Q_N(_12731_),
    .Q(\cpu.spi.r_mode[1][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3500),
    .D(_02573_),
    .Q_N(_12730_),
    .Q(\cpu.spi.r_mode[2][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3501),
    .D(_02574_),
    .Q_N(_12729_),
    .Q(\cpu.spi.r_mode[2][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3502),
    .D(_02575_),
    .Q_N(_12728_),
    .Q(\cpu.spi.r_out[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3503),
    .D(_02576_),
    .Q_N(_12727_),
    .Q(\cpu.spi.r_out[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3504),
    .D(_02577_),
    .Q_N(_12726_),
    .Q(\cpu.spi.r_out[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net3505),
    .D(_02578_),
    .Q_N(_12725_),
    .Q(\cpu.spi.r_out[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[4]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3506),
    .D(_02579_),
    .Q_N(_12724_),
    .Q(\cpu.spi.r_out[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[5]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3507),
    .D(_02580_),
    .Q_N(_12723_),
    .Q(\cpu.spi.r_out[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[6]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3508),
    .D(_02581_),
    .Q_N(_12722_),
    .Q(\cpu.spi.r_out[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[7]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3509),
    .D(_02582_),
    .Q_N(_12721_),
    .Q(\cpu.spi.r_out[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_ready$_SDFFE_PN1P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3510),
    .D(_02583_),
    .Q_N(_12720_),
    .Q(\cpu.spi.r_ready ));
 sg13g2_dfrbp_1 \cpu.spi.r_searching$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3511),
    .D(_02584_),
    .Q_N(_00199_),
    .Q(\cpu.spi.r_searching ));
 sg13g2_dfrbp_1 \cpu.spi.r_sel[0]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3512),
    .D(_02585_),
    .Q_N(_12719_),
    .Q(\cpu.spi.r_sel[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_sel[1]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3513),
    .D(_02586_),
    .Q_N(_12718_),
    .Q(\cpu.spi.r_sel[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_src[0]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3514),
    .D(_02587_),
    .Q_N(_00261_),
    .Q(\cpu.spi.r_src[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_src[1]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3515),
    .D(_02588_),
    .Q_N(_00262_),
    .Q(\cpu.spi.r_src[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_src[2]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3516),
    .D(_02589_),
    .Q_N(_14913_),
    .Q(\cpu.spi.r_src[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[0]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3517),
    .D(_00029_),
    .Q_N(_14914_),
    .Q(\cpu.spi.r_state[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[1]$_DFF_P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3518),
    .D(_00030_),
    .Q_N(_00204_),
    .Q(\cpu.spi.r_state[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[2]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3519),
    .D(_00031_),
    .Q_N(_14915_),
    .Q(\cpu.spi.r_state[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[3]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3520),
    .D(_00032_),
    .Q_N(_14916_),
    .Q(\cpu.spi.r_state[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[4]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3521),
    .D(_00033_),
    .Q_N(_00256_),
    .Q(\cpu.spi.r_state[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[5]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3522),
    .D(_00034_),
    .Q_N(_14917_),
    .Q(\cpu.spi.r_state[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[6]$_DFF_P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3523),
    .D(_00035_),
    .Q_N(_00205_),
    .Q(\cpu.spi.r_state[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[0]$_DFFE_PP_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net3524),
    .D(_02590_),
    .Q_N(_12717_),
    .Q(\cpu.spi.r_timeout[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[1]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3525),
    .D(_02591_),
    .Q_N(_12716_),
    .Q(\cpu.spi.r_timeout[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[2]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3526),
    .D(_02592_),
    .Q_N(_12715_),
    .Q(\cpu.spi.r_timeout[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[3]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3527),
    .D(_02593_),
    .Q_N(_12714_),
    .Q(\cpu.spi.r_timeout[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[4]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3528),
    .D(_02594_),
    .Q_N(_12713_),
    .Q(\cpu.spi.r_timeout[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[5]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3529),
    .D(_02595_),
    .Q_N(_12712_),
    .Q(\cpu.spi.r_timeout[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[6]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3530),
    .D(_02596_),
    .Q_N(_12711_),
    .Q(\cpu.spi.r_timeout[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[7]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3531),
    .D(_02597_),
    .Q_N(_12710_),
    .Q(\cpu.spi.r_timeout[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[0]$_DFFE_PP_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net3532),
    .D(_02598_),
    .Q_N(_00263_),
    .Q(\cpu.spi.r_timeout_count[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[1]$_DFFE_PP_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net3533),
    .D(_02599_),
    .Q_N(_12709_),
    .Q(\cpu.spi.r_timeout_count[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[2]$_DFFE_PP_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net3534),
    .D(_02600_),
    .Q_N(_12708_),
    .Q(\cpu.spi.r_timeout_count[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[3]$_DFFE_PP_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net3535),
    .D(_02601_),
    .Q_N(_12707_),
    .Q(\cpu.spi.r_timeout_count[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[4]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3536),
    .D(_02602_),
    .Q_N(_12706_),
    .Q(\cpu.spi.r_timeout_count[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[5]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3537),
    .D(_02603_),
    .Q_N(_12705_),
    .Q(\cpu.spi.r_timeout_count[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[6]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3538),
    .D(_02604_),
    .Q_N(_12704_),
    .Q(\cpu.spi.r_timeout_count[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[7]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3539),
    .D(_02605_),
    .Q_N(_14918_),
    .Q(\cpu.spi.r_timeout_count[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[0]$_DFF_P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net3540),
    .D(_00079_),
    .Q_N(_00258_),
    .Q(\cpu.uart.r_div[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[10]$_DFF_P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3541),
    .D(_00080_),
    .Q_N(_14919_),
    .Q(\cpu.uart.r_div[10] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[11]$_DFF_P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3542),
    .D(_00081_),
    .Q_N(_14920_),
    .Q(\cpu.uart.r_div[11] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[1]$_DFF_P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net3543),
    .D(_00082_),
    .Q_N(_14921_),
    .Q(\cpu.uart.r_div[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[2]$_DFF_P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net3544),
    .D(_00083_),
    .Q_N(_14922_),
    .Q(\cpu.uart.r_div[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[3]$_DFF_P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net3545),
    .D(_00084_),
    .Q_N(_14923_),
    .Q(\cpu.uart.r_div[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[4]$_DFF_P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net3546),
    .D(_00085_),
    .Q_N(_14924_),
    .Q(\cpu.uart.r_div[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[5]$_DFF_P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net3547),
    .D(_00086_),
    .Q_N(_14925_),
    .Q(\cpu.uart.r_div[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[6]$_DFF_P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net3548),
    .D(_00087_),
    .Q_N(_14926_),
    .Q(\cpu.uart.r_div[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[7]$_DFF_P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net3549),
    .D(_00088_),
    .Q_N(_14927_),
    .Q(\cpu.uart.r_div[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[8]$_DFF_P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net3550),
    .D(_00089_),
    .Q_N(_14928_),
    .Q(\cpu.uart.r_div[8] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[9]$_DFF_P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net3551),
    .D(_00090_),
    .Q_N(_12703_),
    .Q(\cpu.uart.r_div[9] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net3552),
    .D(_02606_),
    .Q_N(_12702_),
    .Q(\cpu.uart.r_div_value[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3553),
    .D(_02607_),
    .Q_N(_12701_),
    .Q(\cpu.uart.r_div_value[10] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3554),
    .D(_02608_),
    .Q_N(_12700_),
    .Q(\cpu.uart.r_div_value[11] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3555),
    .D(_02609_),
    .Q_N(_12699_),
    .Q(\cpu.uart.r_div_value[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3556),
    .D(_02610_),
    .Q_N(_12698_),
    .Q(\cpu.uart.r_div_value[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3557),
    .D(_02611_),
    .Q_N(_12697_),
    .Q(\cpu.uart.r_div_value[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3558),
    .D(_02612_),
    .Q_N(_12696_),
    .Q(\cpu.uart.r_div_value[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3559),
    .D(_02613_),
    .Q_N(_12695_),
    .Q(\cpu.uart.r_div_value[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3560),
    .D(_02614_),
    .Q_N(_12694_),
    .Q(\cpu.uart.r_div_value[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3561),
    .D(_02615_),
    .Q_N(_12693_),
    .Q(\cpu.uart.r_div_value[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3562),
    .D(_02616_),
    .Q_N(_12692_),
    .Q(\cpu.uart.r_div_value[8] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3563),
    .D(_02617_),
    .Q_N(_12691_),
    .Q(\cpu.uart.r_div_value[9] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[0]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3564),
    .D(_02618_),
    .Q_N(_12690_),
    .Q(\cpu.uart.r_ib[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[1]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3565),
    .D(_02619_),
    .Q_N(_12689_),
    .Q(\cpu.uart.r_ib[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[2]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3566),
    .D(_02620_),
    .Q_N(_12688_),
    .Q(\cpu.uart.r_ib[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[3]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3567),
    .D(_02621_),
    .Q_N(_12687_),
    .Q(\cpu.uart.r_ib[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[4]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3568),
    .D(_02622_),
    .Q_N(_12686_),
    .Q(\cpu.uart.r_ib[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[5]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3569),
    .D(_02623_),
    .Q_N(_12685_),
    .Q(\cpu.uart.r_ib[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[6]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3570),
    .D(_02624_),
    .Q_N(_12684_),
    .Q(\cpu.uart.r_ib[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[0]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3571),
    .D(_02625_),
    .Q_N(_12683_),
    .Q(\cpu.uart.r_in[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[1]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3572),
    .D(_02626_),
    .Q_N(_12682_),
    .Q(\cpu.uart.r_in[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[2]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3573),
    .D(_02627_),
    .Q_N(_12681_),
    .Q(\cpu.uart.r_in[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[3]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3574),
    .D(_02628_),
    .Q_N(_12680_),
    .Q(\cpu.uart.r_in[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[4]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3575),
    .D(_02629_),
    .Q_N(_12679_),
    .Q(\cpu.uart.r_in[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[5]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3576),
    .D(_02630_),
    .Q_N(_12678_),
    .Q(\cpu.uart.r_in[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[6]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3577),
    .D(_02631_),
    .Q_N(_12677_),
    .Q(\cpu.uart.r_in[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[7]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3578),
    .D(_02632_),
    .Q_N(_12676_),
    .Q(\cpu.uart.r_in[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3579),
    .D(_02633_),
    .Q_N(_12675_),
    .Q(\cpu.uart.r_out[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3580),
    .D(_02634_),
    .Q_N(_12674_),
    .Q(\cpu.uart.r_out[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3581),
    .D(_02635_),
    .Q_N(_12673_),
    .Q(\cpu.uart.r_out[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3582),
    .D(_02636_),
    .Q_N(_12672_),
    .Q(\cpu.uart.r_out[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[4]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3583),
    .D(_02637_),
    .Q_N(_12671_),
    .Q(\cpu.uart.r_out[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[5]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3584),
    .D(_02638_),
    .Q_N(_12670_),
    .Q(\cpu.uart.r_out[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[6]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3585),
    .D(_02639_),
    .Q_N(_12669_),
    .Q(\cpu.uart.r_out[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[7]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3586),
    .D(_02640_),
    .Q_N(_14929_),
    .Q(\cpu.uart.r_out[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_r$_DFF_P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3587),
    .D(\cpu.gpio.uart_rx ),
    .Q_N(_12668_),
    .Q(\cpu.uart.r_r ));
 sg13g2_dfrbp_1 \cpu.uart.r_r_int$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3588),
    .D(_02641_),
    .Q_N(_12667_),
    .Q(\cpu.uart.r_r_int ));
 sg13g2_dfrbp_1 \cpu.uart.r_r_invert$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3589),
    .D(_02642_),
    .Q_N(_12666_),
    .Q(\cpu.uart.r_r_invert ));
 sg13g2_dfrbp_1 \cpu.uart.r_rcnt[0]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net3590),
    .D(_02643_),
    .Q_N(_12665_),
    .Q(\cpu.uart.r_rcnt[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rcnt[1]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net3591),
    .D(_02644_),
    .Q_N(_12664_),
    .Q(\cpu.uart.r_rcnt[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net3592),
    .D(_02645_),
    .Q_N(_12663_),
    .Q(\cpu.uart.r_rstate[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net3593),
    .D(_02646_),
    .Q_N(_12662_),
    .Q(\cpu.uart.r_rstate[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net3594),
    .D(_02647_),
    .Q_N(_12661_),
    .Q(\cpu.uart.r_rstate[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net3595),
    .D(_02648_),
    .Q_N(_12660_),
    .Q(\cpu.uart.r_rstate[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_x$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3596),
    .D(_02649_),
    .Q_N(_12659_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_x_int$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3597),
    .D(_02650_),
    .Q_N(_12658_),
    .Q(\cpu.uart.r_x_int ));
 sg13g2_dfrbp_1 \cpu.uart.r_x_invert$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3598),
    .D(_02651_),
    .Q_N(_00259_),
    .Q(\cpu.uart.r_x_invert ));
 sg13g2_dfrbp_1 \cpu.uart.r_xcnt[0]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3599),
    .D(_02652_),
    .Q_N(_12657_),
    .Q(\cpu.uart.r_xcnt[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xcnt[1]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3600),
    .D(_02653_),
    .Q_N(_12656_),
    .Q(\cpu.uart.r_xcnt[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3601),
    .D(_02654_),
    .Q_N(_12655_),
    .Q(\cpu.uart.r_xstate[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3602),
    .D(_02655_),
    .Q_N(_12654_),
    .Q(\cpu.uart.r_xstate[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3603),
    .D(_02656_),
    .Q_N(_12653_),
    .Q(\cpu.uart.r_xstate[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3604),
    .D(_02657_),
    .Q_N(_14930_),
    .Q(\cpu.uart.r_xstate[3] ));
 sg13g2_dfrbp_1 \r_reset$_DFF_P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3605),
    .D(_00000_),
    .Q_N(_12652_),
    .Q(r_reset));
 sg13g2_buf_1 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_1 input2 (.A(rst_n),
    .X(net2));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uio_oe[0]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uio_oe[1]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uio_oe[2]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_oe[3]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_oe[4]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_oe[5]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_oe[6]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_oe[7]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[0]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[1]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[2]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[3]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_out[4]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_out[5]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_out[6]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_out[7]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[0]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[1]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[2]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[3]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[4]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[5]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[6]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout27 (.A(_11539_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_06614_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_03722_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_04309_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_06894_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_04141_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_03009_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_02983_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_02957_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_02949_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_02893_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_02861_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_02836_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_02827_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_02771_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_02738_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_02711_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_02703_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_12617_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_12591_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_12583_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_12528_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_12501_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_12476_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_12468_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_12407_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_12375_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_12350_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_12342_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_12284_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_12253_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_12226_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_12217_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_12093_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_12028_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_12004_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_09834_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_09823_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_09822_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_07119_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_07070_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_05004_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_12649_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_12155_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_11661_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_11583_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_11564_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_07206_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_06255_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_06240_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_04143_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_11582_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_11563_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_11471_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_06565_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_06564_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_04254_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_09934_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_07491_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_07304_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_07107_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_06859_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_06591_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_06590_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_06573_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_06572_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_05742_),
    .X(net93));
 sg13g2_buf_4 fanout94 (.X(net94),
    .A(_05147_));
 sg13g2_buf_2 fanout95 (.A(_04130_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_04090_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_03428_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_09958_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_09933_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_09926_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_09919_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_09865_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_09109_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_08927_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_08926_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_07956_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_07755_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_07654_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_05745_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_05228_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_04810_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_04089_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_04068_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_04023_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_03357_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_03167_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_03139_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_11236_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_11100_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_08943_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_08925_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_08883_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_08688_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_07542_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_07501_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_07500_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_07168_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_06702_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_06695_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_06561_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_04217_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_04102_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_04093_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_04088_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_04072_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_04054_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_04016_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_03449_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_03319_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_03153_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_03150_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_11846_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_11795_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_11518_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_11263_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_11235_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_11073_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_09879_),
    .X(net148));
 sg13g2_buf_4 fanout149 (.X(net149),
    .A(_08960_));
 sg13g2_buf_2 fanout150 (.A(_08804_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_08765_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_08687_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_07709_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_07685_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_07674_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_07658_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_07657_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_07484_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_07297_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_04290_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_04234_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_04229_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_04191_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_04078_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_04065_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_04060_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_04057_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_04055_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_04051_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_04046_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_04040_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_04037_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_04031_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_03257_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_03160_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_03154_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_03146_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_11485_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_11451_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_11435_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_11033_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_10996_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_10913_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_09747_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_08941_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_08905_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_08686_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_07647_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_04232_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_04216_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_04062_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_04050_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_03432_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_03276_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_03169_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_03163_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_03159_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_11652_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_11445_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_11385_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_11277_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_11213_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_11177_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_10967_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_10820_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_10817_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_10769_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_09746_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_09726_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_08912_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_08902_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_08783_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_04074_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_04005_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_03350_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_03252_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_03213_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_03158_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_03156_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_03144_),
    .X(net220));
 sg13g2_buf_4 fanout221 (.X(net221),
    .A(_03121_));
 sg13g2_buf_4 fanout222 (.X(net222),
    .A(_03120_));
 sg13g2_buf_2 fanout223 (.A(_11665_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_11284_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_11256_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_11244_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_10826_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_10800_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_10611_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_10541_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_09710_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_08937_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_08929_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_08878_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_06469_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_06365_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_03753_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_03377_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_03290_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_12530_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_11586_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_11584_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_11560_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_11543_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_11467_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_11295_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_11293_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_10877_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_10812_),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(_10676_),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(_10126_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(_09744_),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_08939_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_08928_),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(_06528_),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(_06526_),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(_06525_),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(_06470_),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(_06455_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_06453_),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(_06452_),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(_06364_),
    .X(net262));
 sg13g2_buf_4 fanout263 (.X(net263),
    .A(_06221_));
 sg13g2_buf_4 fanout264 (.X(net264),
    .A(_06196_));
 sg13g2_buf_4 fanout265 (.X(net265),
    .A(_06171_));
 sg13g2_buf_4 fanout266 (.X(net266),
    .A(_06166_));
 sg13g2_buf_4 fanout267 (.X(net267),
    .A(_06138_));
 sg13g2_buf_4 fanout268 (.X(net268),
    .A(_06118_));
 sg13g2_buf_4 fanout269 (.X(net269),
    .A(_06113_));
 sg13g2_buf_4 fanout270 (.X(net270),
    .A(_06107_));
 sg13g2_buf_4 fanout271 (.X(net271),
    .A(_06087_));
 sg13g2_buf_4 fanout272 (.X(net272),
    .A(_06058_));
 sg13g2_buf_4 fanout273 (.X(net273),
    .A(_06051_));
 sg13g2_buf_4 fanout274 (.X(net274),
    .A(_06034_));
 sg13g2_buf_4 fanout275 (.X(net275),
    .A(_06025_));
 sg13g2_buf_4 fanout276 (.X(net276),
    .A(_06002_));
 sg13g2_buf_4 fanout277 (.X(net277),
    .A(_05985_));
 sg13g2_buf_4 fanout278 (.X(net278),
    .A(_05979_));
 sg13g2_buf_4 fanout279 (.X(net279),
    .A(_05958_));
 sg13g2_buf_4 fanout280 (.X(net280),
    .A(_05943_));
 sg13g2_buf_4 fanout281 (.X(net281),
    .A(_05939_));
 sg13g2_buf_4 fanout282 (.X(net282),
    .A(_05934_));
 sg13g2_buf_4 fanout283 (.X(net283),
    .A(_05911_));
 sg13g2_buf_4 fanout284 (.X(net284),
    .A(_05890_));
 sg13g2_buf_4 fanout285 (.X(net285),
    .A(_05883_));
 sg13g2_buf_4 fanout286 (.X(net286),
    .A(_05859_));
 sg13g2_buf_2 fanout287 (.A(_05459_),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(_05016_),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(_04924_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(_04439_),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(_04098_),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(_03752_),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(_03721_),
    .X(net293));
 sg13g2_buf_4 fanout294 (.X(net294),
    .A(_03112_));
 sg13g2_buf_4 fanout295 (.X(net295),
    .A(_03110_));
 sg13g2_buf_2 fanout296 (.A(_11565_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_11542_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(_11466_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(_11405_),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(_11400_),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(_11399_),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(_11274_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(_10339_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_09095_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(_08737_),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(_06436_),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_06434_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(_06433_),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(_06413_),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_06304_),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(_06226_),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(_06225_),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(_06224_),
    .X(net313));
 sg13g2_buf_4 fanout314 (.X(net314),
    .A(_06216_));
 sg13g2_buf_4 fanout315 (.X(net315),
    .A(_06211_));
 sg13g2_buf_4 fanout316 (.X(net316),
    .A(_06206_));
 sg13g2_buf_4 fanout317 (.X(net317),
    .A(_06201_));
 sg13g2_buf_4 fanout318 (.X(net318),
    .A(_06191_));
 sg13g2_buf_4 fanout319 (.X(net319),
    .A(_06186_));
 sg13g2_buf_4 fanout320 (.X(net320),
    .A(_06181_));
 sg13g2_buf_4 fanout321 (.X(net321),
    .A(_06176_));
 sg13g2_buf_4 fanout322 (.X(net322),
    .A(_06156_));
 sg13g2_buf_4 fanout323 (.X(net323),
    .A(_06150_));
 sg13g2_buf_4 fanout324 (.X(net324),
    .A(_06133_));
 sg13g2_buf_4 fanout325 (.X(net325),
    .A(_06128_));
 sg13g2_buf_4 fanout326 (.X(net326),
    .A(_06123_));
 sg13g2_buf_4 fanout327 (.X(net327),
    .A(_06102_));
 sg13g2_buf_4 fanout328 (.X(net328),
    .A(_06093_));
 sg13g2_buf_4 fanout329 (.X(net329),
    .A(_06075_));
 sg13g2_buf_4 fanout330 (.X(net330),
    .A(_06069_));
 sg13g2_buf_4 fanout331 (.X(net331),
    .A(_06063_));
 sg13g2_buf_4 fanout332 (.X(net332),
    .A(_06045_));
 sg13g2_buf_4 fanout333 (.X(net333),
    .A(_06040_));
 sg13g2_buf_4 fanout334 (.X(net334),
    .A(_06022_));
 sg13g2_buf_4 fanout335 (.X(net335),
    .A(_06019_));
 sg13g2_buf_4 fanout336 (.X(net336),
    .A(_06014_));
 sg13g2_buf_4 fanout337 (.X(net337),
    .A(_06007_));
 sg13g2_buf_4 fanout338 (.X(net338),
    .A(_05998_));
 sg13g2_buf_4 fanout339 (.X(net339),
    .A(_05995_));
 sg13g2_buf_4 fanout340 (.X(net340),
    .A(_05992_));
 sg13g2_buf_4 fanout341 (.X(net341),
    .A(_05988_));
 sg13g2_buf_4 fanout342 (.X(net342),
    .A(_05970_));
 sg13g2_buf_4 fanout343 (.X(net343),
    .A(_05964_));
 sg13g2_buf_4 fanout344 (.X(net344),
    .A(_05955_));
 sg13g2_buf_4 fanout345 (.X(net345),
    .A(_05949_));
 sg13g2_buf_4 fanout346 (.X(net346),
    .A(_05946_));
 sg13g2_buf_4 fanout347 (.X(net347),
    .A(_05928_));
 sg13g2_buf_4 fanout348 (.X(net348),
    .A(_05919_));
 sg13g2_buf_4 fanout349 (.X(net349),
    .A(_05906_));
 sg13g2_buf_4 fanout350 (.X(net350),
    .A(_05898_));
 sg13g2_buf_4 fanout351 (.X(net351),
    .A(_05894_));
 sg13g2_buf_4 fanout352 (.X(net352),
    .A(_05876_));
 sg13g2_buf_4 fanout353 (.X(net353),
    .A(_05871_));
 sg13g2_buf_2 fanout354 (.A(_04973_),
    .X(net354));
 sg13g2_buf_2 fanout355 (.A(_04902_),
    .X(net355));
 sg13g2_buf_2 fanout356 (.A(_04898_),
    .X(net356));
 sg13g2_buf_2 fanout357 (.A(_04890_),
    .X(net357));
 sg13g2_buf_2 fanout358 (.A(_03769_),
    .X(net358));
 sg13g2_buf_2 fanout359 (.A(_03663_),
    .X(net359));
 sg13g2_buf_4 fanout360 (.X(net360),
    .A(_03126_));
 sg13g2_buf_4 fanout361 (.X(net361),
    .A(_03125_));
 sg13g2_buf_4 fanout362 (.X(net362),
    .A(_03119_));
 sg13g2_buf_4 fanout363 (.X(net363),
    .A(_03118_));
 sg13g2_buf_4 fanout364 (.X(net364),
    .A(_03091_));
 sg13g2_buf_4 fanout365 (.X(net365),
    .A(_03090_));
 sg13g2_buf_2 fanout366 (.A(_12463_),
    .X(net366));
 sg13g2_buf_2 fanout367 (.A(_12286_),
    .X(net367));
 sg13g2_buf_2 fanout368 (.A(_12171_),
    .X(net368));
 sg13g2_buf_2 fanout369 (.A(_12161_),
    .X(net369));
 sg13g2_buf_2 fanout370 (.A(_11369_),
    .X(net370));
 sg13g2_buf_2 fanout371 (.A(_10463_),
    .X(net371));
 sg13g2_buf_2 fanout372 (.A(_10431_),
    .X(net372));
 sg13g2_buf_2 fanout373 (.A(_10264_),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(_10211_),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(_09687_),
    .X(net375));
 sg13g2_buf_2 fanout376 (.A(_09502_),
    .X(net376));
 sg13g2_buf_2 fanout377 (.A(_09486_),
    .X(net377));
 sg13g2_buf_2 fanout378 (.A(_09113_),
    .X(net378));
 sg13g2_buf_2 fanout379 (.A(_09094_),
    .X(net379));
 sg13g2_buf_2 fanout380 (.A(_08515_),
    .X(net380));
 sg13g2_buf_2 fanout381 (.A(_08494_),
    .X(net381));
 sg13g2_buf_2 fanout382 (.A(_08473_),
    .X(net382));
 sg13g2_buf_2 fanout383 (.A(_08447_),
    .X(net383));
 sg13g2_buf_2 fanout384 (.A(_08422_),
    .X(net384));
 sg13g2_buf_2 fanout385 (.A(_08400_),
    .X(net385));
 sg13g2_buf_2 fanout386 (.A(_08356_),
    .X(net386));
 sg13g2_buf_2 fanout387 (.A(_08259_),
    .X(net387));
 sg13g2_buf_2 fanout388 (.A(_06547_),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(_06545_),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(_06544_),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(_06509_),
    .X(net391));
 sg13g2_buf_2 fanout392 (.A(_06507_),
    .X(net392));
 sg13g2_buf_2 fanout393 (.A(_06506_),
    .X(net393));
 sg13g2_buf_2 fanout394 (.A(_06490_),
    .X(net394));
 sg13g2_buf_2 fanout395 (.A(_06488_),
    .X(net395));
 sg13g2_buf_2 fanout396 (.A(_06487_),
    .X(net396));
 sg13g2_buf_2 fanout397 (.A(_06414_),
    .X(net397));
 sg13g2_buf_2 fanout398 (.A(_06303_),
    .X(net398));
 sg13g2_buf_2 fanout399 (.A(_05974_),
    .X(net399));
 sg13g2_buf_2 fanout400 (.A(_05923_),
    .X(net400));
 sg13g2_buf_2 fanout401 (.A(_05848_),
    .X(net401));
 sg13g2_buf_2 fanout402 (.A(_05340_),
    .X(net402));
 sg13g2_buf_2 fanout403 (.A(_05024_),
    .X(net403));
 sg13g2_buf_2 fanout404 (.A(_04893_),
    .X(net404));
 sg13g2_buf_2 fanout405 (.A(_04889_),
    .X(net405));
 sg13g2_buf_2 fanout406 (.A(_04784_),
    .X(net406));
 sg13g2_buf_4 fanout407 (.X(net407),
    .A(_04781_));
 sg13g2_buf_2 fanout408 (.A(_03658_),
    .X(net408));
 sg13g2_buf_2 fanout409 (.A(_03655_),
    .X(net409));
 sg13g2_buf_2 fanout410 (.A(_03653_),
    .X(net410));
 sg13g2_buf_4 fanout411 (.X(net411),
    .A(_03124_));
 sg13g2_buf_4 fanout412 (.X(net412),
    .A(_03122_));
 sg13g2_buf_2 fanout413 (.A(_03070_),
    .X(net413));
 sg13g2_buf_2 fanout414 (.A(_02773_),
    .X(net414));
 sg13g2_buf_2 fanout415 (.A(_12409_),
    .X(net415));
 sg13g2_buf_2 fanout416 (.A(_12185_),
    .X(net416));
 sg13g2_buf_2 fanout417 (.A(_12181_),
    .X(net417));
 sg13g2_buf_2 fanout418 (.A(_12175_),
    .X(net418));
 sg13g2_buf_2 fanout419 (.A(_12164_),
    .X(net419));
 sg13g2_buf_2 fanout420 (.A(_12149_),
    .X(net420));
 sg13g2_buf_2 fanout421 (.A(_12043_),
    .X(net421));
 sg13g2_buf_2 fanout422 (.A(_11641_),
    .X(net422));
 sg13g2_buf_2 fanout423 (.A(_09966_),
    .X(net423));
 sg13g2_buf_2 fanout424 (.A(_09638_),
    .X(net424));
 sg13g2_buf_2 fanout425 (.A(_09607_),
    .X(net425));
 sg13g2_buf_2 fanout426 (.A(_09446_),
    .X(net426));
 sg13g2_buf_2 fanout427 (.A(_09399_),
    .X(net427));
 sg13g2_buf_2 fanout428 (.A(_09362_),
    .X(net428));
 sg13g2_buf_2 fanout429 (.A(_09329_),
    .X(net429));
 sg13g2_buf_2 fanout430 (.A(_09294_),
    .X(net430));
 sg13g2_buf_2 fanout431 (.A(_09252_),
    .X(net431));
 sg13g2_buf_2 fanout432 (.A(_09208_),
    .X(net432));
 sg13g2_buf_4 fanout433 (.X(net433),
    .A(_08889_));
 sg13g2_buf_2 fanout434 (.A(_08689_),
    .X(net434));
 sg13g2_buf_2 fanout435 (.A(_08601_),
    .X(net435));
 sg13g2_buf_2 fanout436 (.A(_08577_),
    .X(net436));
 sg13g2_buf_2 fanout437 (.A(_08557_),
    .X(net437));
 sg13g2_buf_2 fanout438 (.A(_08285_),
    .X(net438));
 sg13g2_buf_2 fanout439 (.A(_06869_),
    .X(net439));
 sg13g2_buf_2 fanout440 (.A(_06162_),
    .X(net440));
 sg13g2_buf_2 fanout441 (.A(_06161_),
    .X(net441));
 sg13g2_buf_2 fanout442 (.A(_06099_),
    .X(net442));
 sg13g2_buf_2 fanout443 (.A(_06098_),
    .X(net443));
 sg13g2_buf_2 fanout444 (.A(_05027_),
    .X(net444));
 sg13g2_buf_2 fanout445 (.A(_03712_),
    .X(net445));
 sg13g2_buf_2 fanout446 (.A(_03711_),
    .X(net446));
 sg13g2_buf_2 fanout447 (.A(_03697_),
    .X(net447));
 sg13g2_buf_4 fanout448 (.X(net448),
    .A(_03657_));
 sg13g2_buf_2 fanout449 (.A(_03645_),
    .X(net449));
 sg13g2_buf_2 fanout450 (.A(_03643_),
    .X(net450));
 sg13g2_buf_4 fanout451 (.X(net451),
    .A(_03130_));
 sg13g2_buf_4 fanout452 (.X(net452),
    .A(_03127_));
 sg13g2_buf_2 fanout453 (.A(_03081_),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(_03073_),
    .X(net454));
 sg13g2_buf_2 fanout455 (.A(_03069_),
    .X(net455));
 sg13g2_buf_4 fanout456 (.X(net456),
    .A(_12461_));
 sg13g2_buf_2 fanout457 (.A(_12212_),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(_11465_),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(_11043_),
    .X(net459));
 sg13g2_buf_2 fanout460 (.A(_10119_),
    .X(net460));
 sg13g2_buf_2 fanout461 (.A(_09965_),
    .X(net461));
 sg13g2_buf_2 fanout462 (.A(_09923_),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(_09916_),
    .X(net463));
 sg13g2_buf_4 fanout464 (.X(net464),
    .A(_09106_));
 sg13g2_buf_2 fanout465 (.A(_08784_),
    .X(net465));
 sg13g2_buf_4 fanout466 (.X(net466),
    .A(_08770_));
 sg13g2_buf_2 fanout467 (.A(_08716_),
    .X(net467));
 sg13g2_buf_2 fanout468 (.A(_08700_),
    .X(net468));
 sg13g2_buf_2 fanout469 (.A(_08535_),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(_08357_),
    .X(net470));
 sg13g2_buf_2 fanout471 (.A(_08298_),
    .X(net471));
 sg13g2_buf_2 fanout472 (.A(_07566_),
    .X(net472));
 sg13g2_buf_2 fanout473 (.A(_07535_),
    .X(net473));
 sg13g2_buf_2 fanout474 (.A(_07404_),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(_06153_),
    .X(net475));
 sg13g2_buf_2 fanout476 (.A(_06090_),
    .X(net476));
 sg13g2_buf_2 fanout477 (.A(_06066_),
    .X(net477));
 sg13g2_buf_2 fanout478 (.A(_06037_),
    .X(net478));
 sg13g2_buf_2 fanout479 (.A(_05960_),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(_05959_),
    .X(net480));
 sg13g2_buf_2 fanout481 (.A(_05908_),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(_05907_),
    .X(net482));
 sg13g2_buf_2 fanout483 (.A(_05891_),
    .X(net483));
 sg13g2_buf_2 fanout484 (.A(_05863_),
    .X(net484));
 sg13g2_buf_2 fanout485 (.A(_05048_),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(_05033_),
    .X(net486));
 sg13g2_buf_2 fanout487 (.A(_05030_),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(_05023_),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(_04862_),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(_04855_),
    .X(net490));
 sg13g2_buf_4 fanout491 (.X(net491),
    .A(_04788_));
 sg13g2_buf_2 fanout492 (.A(_04774_),
    .X(net492));
 sg13g2_buf_4 fanout493 (.X(net493),
    .A(_04768_));
 sg13g2_buf_2 fanout494 (.A(_03763_),
    .X(net494));
 sg13g2_buf_2 fanout495 (.A(_03718_),
    .X(net495));
 sg13g2_buf_2 fanout496 (.A(_03696_),
    .X(net496));
 sg13g2_buf_4 fanout497 (.X(net497),
    .A(_03695_));
 sg13g2_buf_4 fanout498 (.X(net498),
    .A(_03691_));
 sg13g2_buf_4 fanout499 (.X(net499),
    .A(_03681_));
 sg13g2_buf_4 fanout500 (.X(net500),
    .A(_03662_));
 sg13g2_buf_2 fanout501 (.A(_03656_),
    .X(net501));
 sg13g2_buf_2 fanout502 (.A(_03652_),
    .X(net502));
 sg13g2_buf_2 fanout503 (.A(_03644_),
    .X(net503));
 sg13g2_buf_2 fanout504 (.A(_03642_),
    .X(net504));
 sg13g2_buf_4 fanout505 (.X(net505),
    .A(_03641_));
 sg13g2_buf_4 fanout506 (.X(net506),
    .A(_03131_));
 sg13g2_buf_4 fanout507 (.X(net507),
    .A(_03128_));
 sg13g2_buf_2 fanout508 (.A(_03109_),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(_03084_),
    .X(net509));
 sg13g2_buf_2 fanout510 (.A(_03080_),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(_03076_),
    .X(net511));
 sg13g2_buf_2 fanout512 (.A(_03072_),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(_03068_),
    .X(net513));
 sg13g2_buf_2 fanout514 (.A(_03011_),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(_02895_),
    .X(net515));
 sg13g2_buf_2 fanout516 (.A(_02698_),
    .X(net516));
 sg13g2_buf_4 fanout517 (.X(net517),
    .A(_12460_));
 sg13g2_buf_2 fanout518 (.A(_12337_),
    .X(net518));
 sg13g2_buf_2 fanout519 (.A(_12008_),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(_11948_),
    .X(net520));
 sg13g2_buf_2 fanout521 (.A(_11546_),
    .X(net521));
 sg13g2_buf_2 fanout522 (.A(_11541_),
    .X(net522));
 sg13g2_buf_2 fanout523 (.A(_11418_),
    .X(net523));
 sg13g2_buf_2 fanout524 (.A(_11049_),
    .X(net524));
 sg13g2_buf_2 fanout525 (.A(_10792_),
    .X(net525));
 sg13g2_buf_2 fanout526 (.A(_10533_),
    .X(net526));
 sg13g2_buf_2 fanout527 (.A(_10357_),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(_09922_),
    .X(net528));
 sg13g2_buf_2 fanout529 (.A(_09915_),
    .X(net529));
 sg13g2_buf_2 fanout530 (.A(_09780_),
    .X(net530));
 sg13g2_buf_2 fanout531 (.A(_09330_),
    .X(net531));
 sg13g2_buf_4 fanout532 (.X(net532),
    .A(_09105_));
 sg13g2_buf_2 fanout533 (.A(_08785_),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(_08698_),
    .X(net534));
 sg13g2_buf_2 fanout535 (.A(_08697_),
    .X(net535));
 sg13g2_buf_4 fanout536 (.X(net536),
    .A(_08374_));
 sg13g2_buf_2 fanout537 (.A(_08358_),
    .X(net537));
 sg13g2_buf_2 fanout538 (.A(_08321_),
    .X(net538));
 sg13g2_buf_2 fanout539 (.A(_08306_),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(_08300_),
    .X(net540));
 sg13g2_buf_2 fanout541 (.A(_08297_),
    .X(net541));
 sg13g2_buf_2 fanout542 (.A(_07854_),
    .X(net542));
 sg13g2_buf_2 fanout543 (.A(_07763_),
    .X(net543));
 sg13g2_buf_2 fanout544 (.A(_07740_),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(_07729_),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(_07706_),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(_07682_),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(_07641_),
    .X(net548));
 sg13g2_buf_2 fanout549 (.A(_07609_),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(_07570_),
    .X(net550));
 sg13g2_buf_2 fanout551 (.A(_07551_),
    .X(net551));
 sg13g2_buf_2 fanout552 (.A(_07534_),
    .X(net552));
 sg13g2_buf_2 fanout553 (.A(_07504_),
    .X(net553));
 sg13g2_buf_2 fanout554 (.A(_07210_),
    .X(net554));
 sg13g2_buf_2 fanout555 (.A(_07072_),
    .X(net555));
 sg13g2_buf_2 fanout556 (.A(_06674_),
    .X(net556));
 sg13g2_buf_2 fanout557 (.A(_06159_),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(_06158_),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(_06096_),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(_06095_),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(_05950_),
    .X(net561));
 sg13g2_buf_2 fanout562 (.A(_05895_),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(_05014_),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(_04849_),
    .X(net564));
 sg13g2_buf_2 fanout565 (.A(_04769_),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(_03717_),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(_03714_),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(_03713_),
    .X(net568));
 sg13g2_buf_4 fanout569 (.X(net569),
    .A(_03703_));
 sg13g2_buf_2 fanout570 (.A(_03688_),
    .X(net570));
 sg13g2_buf_4 fanout571 (.X(net571),
    .A(_03687_));
 sg13g2_buf_2 fanout572 (.A(_03680_),
    .X(net572));
 sg13g2_buf_4 fanout573 (.X(net573),
    .A(_03674_));
 sg13g2_buf_4 fanout574 (.X(net574),
    .A(_03668_));
 sg13g2_buf_4 fanout575 (.X(net575),
    .A(_03651_));
 sg13g2_buf_2 fanout576 (.A(_03649_),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(_03647_),
    .X(net577));
 sg13g2_buf_4 fanout578 (.X(net578),
    .A(_03640_));
 sg13g2_buf_4 fanout579 (.X(net579),
    .A(_03108_));
 sg13g2_buf_2 fanout580 (.A(_03083_),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(_03079_),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(_03075_),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(_12578_),
    .X(net583));
 sg13g2_buf_2 fanout584 (.A(_12040_),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(_11947_),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(_11568_),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(_11545_),
    .X(net587));
 sg13g2_buf_2 fanout588 (.A(_11249_),
    .X(net588));
 sg13g2_buf_2 fanout589 (.A(_11023_),
    .X(net589));
 sg13g2_buf_2 fanout590 (.A(_10973_),
    .X(net590));
 sg13g2_buf_2 fanout591 (.A(_10897_),
    .X(net591));
 sg13g2_buf_2 fanout592 (.A(_10625_),
    .X(net592));
 sg13g2_buf_2 fanout593 (.A(_10507_),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(_10213_),
    .X(net594));
 sg13g2_buf_2 fanout595 (.A(_10052_),
    .X(net595));
 sg13g2_buf_2 fanout596 (.A(_10047_),
    .X(net596));
 sg13g2_buf_2 fanout597 (.A(_10029_),
    .X(net597));
 sg13g2_buf_2 fanout598 (.A(_09963_),
    .X(net598));
 sg13g2_buf_2 fanout599 (.A(_09779_),
    .X(net599));
 sg13g2_buf_2 fanout600 (.A(_09675_),
    .X(net600));
 sg13g2_buf_2 fanout601 (.A(_09483_),
    .X(net601));
 sg13g2_buf_2 fanout602 (.A(_09449_),
    .X(net602));
 sg13g2_buf_2 fanout603 (.A(_09447_),
    .X(net603));
 sg13g2_buf_2 fanout604 (.A(_09300_),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(_09259_),
    .X(net605));
 sg13g2_buf_2 fanout606 (.A(_09137_),
    .X(net606));
 sg13g2_buf_4 fanout607 (.X(net607),
    .A(_09130_));
 sg13g2_buf_4 fanout608 (.X(net608),
    .A(_09104_));
 sg13g2_buf_2 fanout609 (.A(_09037_),
    .X(net609));
 sg13g2_buf_2 fanout610 (.A(_08888_),
    .X(net610));
 sg13g2_buf_2 fanout611 (.A(_08712_),
    .X(net611));
 sg13g2_buf_2 fanout612 (.A(_08710_),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(_08402_),
    .X(net613));
 sg13g2_buf_2 fanout614 (.A(_08373_),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(_08367_),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(_08339_),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(_08320_),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(_08315_),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(_08305_),
    .X(net619));
 sg13g2_buf_2 fanout620 (.A(_08299_),
    .X(net620));
 sg13g2_buf_2 fanout621 (.A(_08296_),
    .X(net621));
 sg13g2_buf_2 fanout622 (.A(_07450_),
    .X(net622));
 sg13g2_buf_2 fanout623 (.A(_06866_),
    .X(net623));
 sg13g2_buf_2 fanout624 (.A(_06140_),
    .X(net624));
 sg13g2_buf_2 fanout625 (.A(_06077_),
    .X(net625));
 sg13g2_buf_2 fanout626 (.A(_05971_),
    .X(net626));
 sg13g2_buf_2 fanout627 (.A(_05965_),
    .X(net627));
 sg13g2_buf_2 fanout628 (.A(_05920_),
    .X(net628));
 sg13g2_buf_2 fanout629 (.A(_05912_),
    .X(net629));
 sg13g2_buf_2 fanout630 (.A(_05013_),
    .X(net630));
 sg13g2_buf_2 fanout631 (.A(_04852_),
    .X(net631));
 sg13g2_buf_2 fanout632 (.A(_04270_),
    .X(net632));
 sg13g2_buf_2 fanout633 (.A(_03709_),
    .X(net633));
 sg13g2_buf_2 fanout634 (.A(_03708_),
    .X(net634));
 sg13g2_buf_2 fanout635 (.A(_03705_),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(_03673_),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(_03650_),
    .X(net637));
 sg13g2_buf_2 fanout638 (.A(_03648_),
    .X(net638));
 sg13g2_buf_2 fanout639 (.A(_03646_),
    .X(net639));
 sg13g2_buf_4 fanout640 (.X(net640),
    .A(_03107_));
 sg13g2_buf_2 fanout641 (.A(_03089_),
    .X(net641));
 sg13g2_buf_2 fanout642 (.A(_02822_),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(_11995_),
    .X(net643));
 sg13g2_buf_4 fanout644 (.X(net644),
    .A(_11988_));
 sg13g2_buf_2 fanout645 (.A(_11942_),
    .X(net645));
 sg13g2_buf_2 fanout646 (.A(_11939_),
    .X(net646));
 sg13g2_buf_2 fanout647 (.A(_11904_),
    .X(net647));
 sg13g2_buf_2 fanout648 (.A(_11884_),
    .X(net648));
 sg13g2_buf_2 fanout649 (.A(_11507_),
    .X(net649));
 sg13g2_buf_2 fanout650 (.A(_11473_),
    .X(net650));
 sg13g2_buf_2 fanout651 (.A(_11267_),
    .X(net651));
 sg13g2_buf_2 fanout652 (.A(_11248_),
    .X(net652));
 sg13g2_buf_2 fanout653 (.A(_10624_),
    .X(net653));
 sg13g2_buf_2 fanout654 (.A(_10620_),
    .X(net654));
 sg13g2_buf_2 fanout655 (.A(_10601_),
    .X(net655));
 sg13g2_buf_2 fanout656 (.A(_10549_),
    .X(net656));
 sg13g2_buf_2 fanout657 (.A(_10519_),
    .X(net657));
 sg13g2_buf_2 fanout658 (.A(_10516_),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(_10506_),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(_10248_),
    .X(net660));
 sg13g2_buf_2 fanout661 (.A(_10245_),
    .X(net661));
 sg13g2_buf_2 fanout662 (.A(_10229_),
    .X(net662));
 sg13g2_buf_2 fanout663 (.A(_10163_),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(_10099_),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(_10096_),
    .X(net665));
 sg13g2_buf_2 fanout666 (.A(_10084_),
    .X(net666));
 sg13g2_buf_2 fanout667 (.A(_10077_),
    .X(net667));
 sg13g2_buf_2 fanout668 (.A(_10063_),
    .X(net668));
 sg13g2_buf_2 fanout669 (.A(_10059_),
    .X(net669));
 sg13g2_buf_2 fanout670 (.A(_10056_),
    .X(net670));
 sg13g2_buf_2 fanout671 (.A(_10051_),
    .X(net671));
 sg13g2_buf_2 fanout672 (.A(_09876_),
    .X(net672));
 sg13g2_buf_2 fanout673 (.A(_09875_),
    .X(net673));
 sg13g2_buf_2 fanout674 (.A(_09784_),
    .X(net674));
 sg13g2_buf_2 fanout675 (.A(_09778_),
    .X(net675));
 sg13g2_buf_2 fanout676 (.A(_09582_),
    .X(net676));
 sg13g2_buf_2 fanout677 (.A(_09420_),
    .X(net677));
 sg13g2_buf_4 fanout678 (.X(net678),
    .A(_09402_));
 sg13g2_buf_4 fanout679 (.X(net679),
    .A(_09401_));
 sg13g2_buf_2 fanout680 (.A(_09297_),
    .X(net680));
 sg13g2_buf_2 fanout681 (.A(_09255_),
    .X(net681));
 sg13g2_buf_2 fanout682 (.A(_09198_),
    .X(net682));
 sg13g2_buf_2 fanout683 (.A(_09157_),
    .X(net683));
 sg13g2_buf_4 fanout684 (.X(net684),
    .A(_09124_));
 sg13g2_buf_2 fanout685 (.A(_09103_),
    .X(net685));
 sg13g2_buf_4 fanout686 (.X(net686),
    .A(_09036_));
 sg13g2_buf_2 fanout687 (.A(_08965_),
    .X(net687));
 sg13g2_buf_2 fanout688 (.A(_08766_),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(_08739_),
    .X(net689));
 sg13g2_buf_2 fanout690 (.A(_08701_),
    .X(net690));
 sg13g2_buf_2 fanout691 (.A(_08695_),
    .X(net691));
 sg13g2_buf_4 fanout692 (.X(net692),
    .A(_08693_));
 sg13g2_buf_4 fanout693 (.X(net693),
    .A(_08433_));
 sg13g2_buf_4 fanout694 (.X(net694),
    .A(_08393_));
 sg13g2_buf_4 fanout695 (.X(net695),
    .A(_08383_));
 sg13g2_buf_2 fanout696 (.A(_08361_),
    .X(net696));
 sg13g2_buf_4 fanout697 (.X(net697),
    .A(_08338_));
 sg13g2_buf_2 fanout698 (.A(_08314_),
    .X(net698));
 sg13g2_buf_2 fanout699 (.A(_08310_),
    .X(net699));
 sg13g2_buf_2 fanout700 (.A(_06694_),
    .X(net700));
 sg13g2_buf_2 fanout701 (.A(_06693_),
    .X(net701));
 sg13g2_buf_2 fanout702 (.A(_06144_),
    .X(net702));
 sg13g2_buf_2 fanout703 (.A(_06143_),
    .X(net703));
 sg13g2_buf_2 fanout704 (.A(_06142_),
    .X(net704));
 sg13g2_buf_2 fanout705 (.A(_06081_),
    .X(net705));
 sg13g2_buf_2 fanout706 (.A(_06080_),
    .X(net706));
 sg13g2_buf_2 fanout707 (.A(_06079_),
    .X(net707));
 sg13g2_buf_2 fanout708 (.A(_05865_),
    .X(net708));
 sg13g2_buf_2 fanout709 (.A(_03135_),
    .X(net709));
 sg13g2_buf_2 fanout710 (.A(_03134_),
    .X(net710));
 sg13g2_buf_2 fanout711 (.A(_03133_),
    .X(net711));
 sg13g2_buf_1 fanout712 (.A(_03114_),
    .X(net712));
 sg13g2_buf_1 fanout713 (.A(_03113_),
    .X(net713));
 sg13g2_buf_2 fanout714 (.A(_03111_),
    .X(net714));
 sg13g2_buf_2 fanout715 (.A(_03100_),
    .X(net715));
 sg13g2_buf_2 fanout716 (.A(_03098_),
    .X(net716));
 sg13g2_buf_2 fanout717 (.A(_03095_),
    .X(net717));
 sg13g2_buf_2 fanout718 (.A(_03088_),
    .X(net718));
 sg13g2_buf_2 fanout719 (.A(_02766_),
    .X(net719));
 sg13g2_buf_2 fanout720 (.A(_02755_),
    .X(net720));
 sg13g2_buf_2 fanout721 (.A(_02749_),
    .X(net721));
 sg13g2_buf_2 fanout722 (.A(_12140_),
    .X(net722));
 sg13g2_buf_2 fanout723 (.A(_12121_),
    .X(net723));
 sg13g2_buf_2 fanout724 (.A(_12112_),
    .X(net724));
 sg13g2_buf_2 fanout725 (.A(_12106_),
    .X(net725));
 sg13g2_buf_2 fanout726 (.A(_11959_),
    .X(net726));
 sg13g2_buf_2 fanout727 (.A(_11946_),
    .X(net727));
 sg13g2_buf_2 fanout728 (.A(_11930_),
    .X(net728));
 sg13g2_buf_2 fanout729 (.A(_11900_),
    .X(net729));
 sg13g2_buf_2 fanout730 (.A(_11323_),
    .X(net730));
 sg13g2_buf_2 fanout731 (.A(_11186_),
    .X(net731));
 sg13g2_buf_2 fanout732 (.A(_11042_),
    .X(net732));
 sg13g2_buf_2 fanout733 (.A(_10771_),
    .X(net733));
 sg13g2_buf_2 fanout734 (.A(_10511_),
    .X(net734));
 sg13g2_buf_2 fanout735 (.A(_10508_),
    .X(net735));
 sg13g2_buf_2 fanout736 (.A(_10433_),
    .X(net736));
 sg13g2_buf_2 fanout737 (.A(_10391_),
    .X(net737));
 sg13g2_buf_2 fanout738 (.A(_10306_),
    .X(net738));
 sg13g2_buf_2 fanout739 (.A(_10301_),
    .X(net739));
 sg13g2_buf_2 fanout740 (.A(_10272_),
    .X(net740));
 sg13g2_buf_2 fanout741 (.A(_10266_),
    .X(net741));
 sg13g2_buf_2 fanout742 (.A(_10214_),
    .X(net742));
 sg13g2_buf_2 fanout743 (.A(_10199_),
    .X(net743));
 sg13g2_buf_2 fanout744 (.A(_10194_),
    .X(net744));
 sg13g2_buf_2 fanout745 (.A(_10178_),
    .X(net745));
 sg13g2_buf_2 fanout746 (.A(_10158_),
    .X(net746));
 sg13g2_buf_2 fanout747 (.A(_10147_),
    .X(net747));
 sg13g2_buf_2 fanout748 (.A(_10088_),
    .X(net748));
 sg13g2_buf_2 fanout749 (.A(_10078_),
    .X(net749));
 sg13g2_buf_2 fanout750 (.A(_10066_),
    .X(net750));
 sg13g2_buf_2 fanout751 (.A(_10055_),
    .X(net751));
 sg13g2_buf_2 fanout752 (.A(_10050_),
    .X(net752));
 sg13g2_buf_2 fanout753 (.A(_09884_),
    .X(net753));
 sg13g2_buf_2 fanout754 (.A(_09874_),
    .X(net754));
 sg13g2_buf_2 fanout755 (.A(_09777_),
    .X(net755));
 sg13g2_buf_8 fanout756 (.A(_09476_),
    .X(net756));
 sg13g2_buf_4 fanout757 (.X(net757),
    .A(_09474_));
 sg13g2_buf_2 fanout758 (.A(_09462_),
    .X(net758));
 sg13g2_buf_4 fanout759 (.X(net759),
    .A(_09432_));
 sg13g2_buf_8 fanout760 (.A(_09431_),
    .X(net760));
 sg13g2_buf_4 fanout761 (.X(net761),
    .A(_09412_));
 sg13g2_buf_8 fanout762 (.A(_09411_),
    .X(net762));
 sg13g2_buf_2 fanout763 (.A(_09382_),
    .X(net763));
 sg13g2_buf_8 fanout764 (.A(_09322_),
    .X(net764));
 sg13g2_buf_4 fanout765 (.X(net765),
    .A(_09320_));
 sg13g2_buf_4 fanout766 (.X(net766),
    .A(_09280_));
 sg13g2_buf_8 fanout767 (.A(_09279_),
    .X(net767));
 sg13g2_buf_2 fanout768 (.A(_09269_),
    .X(net768));
 sg13g2_buf_2 fanout769 (.A(_09265_),
    .X(net769));
 sg13g2_buf_4 fanout770 (.X(net770),
    .A(_09236_));
 sg13g2_buf_4 fanout771 (.X(net771),
    .A(_09235_));
 sg13g2_buf_2 fanout772 (.A(_09230_),
    .X(net772));
 sg13g2_buf_4 fanout773 (.X(net773),
    .A(_09191_));
 sg13g2_buf_4 fanout774 (.X(net774),
    .A(_09187_));
 sg13g2_buf_8 fanout775 (.A(_09185_),
    .X(net775));
 sg13g2_buf_2 fanout776 (.A(_09183_),
    .X(net776));
 sg13g2_buf_2 fanout777 (.A(_09174_),
    .X(net777));
 sg13g2_buf_4 fanout778 (.X(net778),
    .A(_09123_));
 sg13g2_buf_2 fanout779 (.A(_09118_),
    .X(net779));
 sg13g2_buf_2 fanout780 (.A(_09102_),
    .X(net780));
 sg13g2_buf_4 fanout781 (.X(net781),
    .A(_09052_));
 sg13g2_buf_2 fanout782 (.A(_09035_),
    .X(net782));
 sg13g2_buf_2 fanout783 (.A(_08964_),
    .X(net783));
 sg13g2_buf_2 fanout784 (.A(_08707_),
    .X(net784));
 sg13g2_buf_2 fanout785 (.A(_08691_),
    .X(net785));
 sg13g2_buf_4 fanout786 (.X(net786),
    .A(_08545_));
 sg13g2_buf_8 fanout787 (.A(_08464_),
    .X(net787));
 sg13g2_buf_4 fanout788 (.X(net788),
    .A(_08424_));
 sg13g2_buf_4 fanout789 (.X(net789),
    .A(_08397_));
 sg13g2_buf_4 fanout790 (.X(net790),
    .A(_08389_));
 sg13g2_buf_4 fanout791 (.X(net791),
    .A(_08349_));
 sg13g2_buf_2 fanout792 (.A(_08337_),
    .X(net792));
 sg13g2_buf_2 fanout793 (.A(_08332_),
    .X(net793));
 sg13g2_buf_4 fanout794 (.X(net794),
    .A(_08325_));
 sg13g2_buf_2 fanout795 (.A(_08309_),
    .X(net795));
 sg13g2_buf_8 fanout796 (.A(_08272_),
    .X(net796));
 sg13g2_buf_4 fanout797 (.X(net797),
    .A(_08269_));
 sg13g2_buf_4 fanout798 (.X(net798),
    .A(_08265_));
 sg13g2_buf_2 fanout799 (.A(_07071_),
    .X(net799));
 sg13g2_buf_2 fanout800 (.A(_06872_),
    .X(net800));
 sg13g2_buf_2 fanout801 (.A(_06763_),
    .X(net801));
 sg13g2_buf_2 fanout802 (.A(_06362_),
    .X(net802));
 sg13g2_buf_2 fanout803 (.A(_06361_),
    .X(net803));
 sg13g2_buf_2 fanout804 (.A(_06348_),
    .X(net804));
 sg13g2_buf_2 fanout805 (.A(_06324_),
    .X(net805));
 sg13g2_buf_2 fanout806 (.A(_06323_),
    .X(net806));
 sg13g2_buf_2 fanout807 (.A(_06318_),
    .X(net807));
 sg13g2_buf_2 fanout808 (.A(_06316_),
    .X(net808));
 sg13g2_buf_2 fanout809 (.A(_06283_),
    .X(net809));
 sg13g2_buf_2 fanout810 (.A(_06276_),
    .X(net810));
 sg13g2_buf_2 fanout811 (.A(_06147_),
    .X(net811));
 sg13g2_buf_2 fanout812 (.A(_06146_),
    .X(net812));
 sg13g2_buf_2 fanout813 (.A(_06145_),
    .X(net813));
 sg13g2_buf_2 fanout814 (.A(_06084_),
    .X(net814));
 sg13g2_buf_2 fanout815 (.A(_06083_),
    .X(net815));
 sg13g2_buf_2 fanout816 (.A(_06082_),
    .X(net816));
 sg13g2_buf_2 fanout817 (.A(_05989_),
    .X(net817));
 sg13g2_buf_2 fanout818 (.A(_05980_),
    .X(net818));
 sg13g2_buf_2 fanout819 (.A(_05972_),
    .X(net819));
 sg13g2_buf_2 fanout820 (.A(_05940_),
    .X(net820));
 sg13g2_buf_2 fanout821 (.A(_05929_),
    .X(net821));
 sg13g2_buf_2 fanout822 (.A(_05921_),
    .X(net822));
 sg13g2_buf_2 fanout823 (.A(_05877_),
    .X(net823));
 sg13g2_buf_2 fanout824 (.A(_05862_),
    .X(net824));
 sg13g2_buf_2 fanout825 (.A(_05861_),
    .X(net825));
 sg13g2_buf_2 fanout826 (.A(_05860_),
    .X(net826));
 sg13g2_buf_2 fanout827 (.A(_05828_),
    .X(net827));
 sg13g2_buf_2 fanout828 (.A(_05826_),
    .X(net828));
 sg13g2_buf_2 fanout829 (.A(_05780_),
    .X(net829));
 sg13g2_buf_2 fanout830 (.A(_05369_),
    .X(net830));
 sg13g2_buf_2 fanout831 (.A(_05151_),
    .X(net831));
 sg13g2_buf_2 fanout832 (.A(_05018_),
    .X(net832));
 sg13g2_buf_2 fanout833 (.A(_04770_),
    .X(net833));
 sg13g2_buf_2 fanout834 (.A(_04083_),
    .X(net834));
 sg13g2_buf_2 fanout835 (.A(_03633_),
    .X(net835));
 sg13g2_buf_2 fanout836 (.A(_03138_),
    .X(net836));
 sg13g2_buf_2 fanout837 (.A(_03137_),
    .X(net837));
 sg13g2_buf_2 fanout838 (.A(_03136_),
    .X(net838));
 sg13g2_buf_2 fanout839 (.A(_03117_),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(_03116_),
    .X(net840));
 sg13g2_buf_2 fanout841 (.A(_03115_),
    .X(net841));
 sg13g2_buf_2 fanout842 (.A(_03106_),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(_03104_),
    .X(net843));
 sg13g2_buf_2 fanout844 (.A(_03102_),
    .X(net844));
 sg13g2_buf_2 fanout845 (.A(_03099_),
    .X(net845));
 sg13g2_buf_2 fanout846 (.A(_03097_),
    .X(net846));
 sg13g2_buf_2 fanout847 (.A(_03094_),
    .X(net847));
 sg13g2_buf_2 fanout848 (.A(_03087_),
    .X(net848));
 sg13g2_buf_2 fanout849 (.A(_12522_),
    .X(net849));
 sg13g2_buf_2 fanout850 (.A(_12391_),
    .X(net850));
 sg13g2_buf_2 fanout851 (.A(_12222_),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(_12139_),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(_12120_),
    .X(net853));
 sg13g2_buf_2 fanout854 (.A(_12111_),
    .X(net854));
 sg13g2_buf_2 fanout855 (.A(_12104_),
    .X(net855));
 sg13g2_buf_2 fanout856 (.A(_11965_),
    .X(net856));
 sg13g2_buf_2 fanout857 (.A(_11938_),
    .X(net857));
 sg13g2_buf_2 fanout858 (.A(_11929_),
    .X(net858));
 sg13g2_buf_2 fanout859 (.A(_11914_),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(_10795_),
    .X(net860));
 sg13g2_buf_2 fanout861 (.A(_10452_),
    .X(net861));
 sg13g2_buf_2 fanout862 (.A(_10235_),
    .X(net862));
 sg13g2_buf_2 fanout863 (.A(_10224_),
    .X(net863));
 sg13g2_buf_2 fanout864 (.A(_10187_),
    .X(net864));
 sg13g2_buf_2 fanout865 (.A(_10177_),
    .X(net865));
 sg13g2_buf_2 fanout866 (.A(_10176_),
    .X(net866));
 sg13g2_buf_2 fanout867 (.A(_10173_),
    .X(net867));
 sg13g2_buf_2 fanout868 (.A(_10169_),
    .X(net868));
 sg13g2_buf_2 fanout869 (.A(_10168_),
    .X(net869));
 sg13g2_buf_2 fanout870 (.A(_10101_),
    .X(net870));
 sg13g2_buf_2 fanout871 (.A(_10069_),
    .X(net871));
 sg13g2_buf_2 fanout872 (.A(_10065_),
    .X(net872));
 sg13g2_buf_2 fanout873 (.A(_10054_),
    .X(net873));
 sg13g2_buf_2 fanout874 (.A(_10049_),
    .X(net874));
 sg13g2_buf_2 fanout875 (.A(_09957_),
    .X(net875));
 sg13g2_buf_2 fanout876 (.A(_09937_),
    .X(net876));
 sg13g2_buf_2 fanout877 (.A(_09927_),
    .X(net877));
 sg13g2_buf_2 fanout878 (.A(_09883_),
    .X(net878));
 sg13g2_buf_2 fanout879 (.A(_09873_),
    .X(net879));
 sg13g2_buf_2 fanout880 (.A(_09861_),
    .X(net880));
 sg13g2_buf_2 fanout881 (.A(_09776_),
    .X(net881));
 sg13g2_buf_2 fanout882 (.A(_09686_),
    .X(net882));
 sg13g2_buf_2 fanout883 (.A(_09544_),
    .X(net883));
 sg13g2_buf_4 fanout884 (.X(net884),
    .A(_09385_));
 sg13g2_buf_2 fanout885 (.A(_09381_),
    .X(net885));
 sg13g2_buf_4 fanout886 (.X(net886),
    .A(_09313_));
 sg13g2_buf_2 fanout887 (.A(_09306_),
    .X(net887));
 sg13g2_buf_4 fanout888 (.X(net888),
    .A(_09242_));
 sg13g2_buf_8 fanout889 (.A(_09241_),
    .X(net889));
 sg13g2_buf_2 fanout890 (.A(_09224_),
    .X(net890));
 sg13g2_buf_2 fanout891 (.A(_09217_),
    .X(net891));
 sg13g2_buf_4 fanout892 (.X(net892),
    .A(_09202_));
 sg13g2_buf_8 fanout893 (.A(_09201_),
    .X(net893));
 sg13g2_buf_8 fanout894 (.A(_09190_),
    .X(net894));
 sg13g2_buf_2 fanout895 (.A(_09173_),
    .X(net895));
 sg13g2_buf_2 fanout896 (.A(_09166_),
    .X(net896));
 sg13g2_buf_2 fanout897 (.A(_09122_),
    .X(net897));
 sg13g2_buf_2 fanout898 (.A(_09101_),
    .X(net898));
 sg13g2_buf_2 fanout899 (.A(_09099_),
    .X(net899));
 sg13g2_buf_2 fanout900 (.A(_09034_),
    .X(net900));
 sg13g2_buf_2 fanout901 (.A(_08963_),
    .X(net901));
 sg13g2_buf_2 fanout902 (.A(_08706_),
    .X(net902));
 sg13g2_buf_4 fanout903 (.X(net903),
    .A(_08605_));
 sg13g2_buf_8 fanout904 (.A(_08551_),
    .X(net904));
 sg13g2_buf_4 fanout905 (.X(net905),
    .A(_08463_));
 sg13g2_buf_2 fanout906 (.A(_08438_),
    .X(net906));
 sg13g2_buf_8 fanout907 (.A(_08432_),
    .X(net907));
 sg13g2_buf_2 fanout908 (.A(_08425_),
    .X(net908));
 sg13g2_buf_8 fanout909 (.A(_08386_),
    .X(net909));
 sg13g2_buf_8 fanout910 (.A(_08382_),
    .X(net910));
 sg13g2_buf_8 fanout911 (.A(_08342_),
    .X(net911));
 sg13g2_buf_2 fanout912 (.A(_08331_),
    .X(net912));
 sg13g2_buf_2 fanout913 (.A(_08328_),
    .X(net913));
 sg13g2_buf_2 fanout914 (.A(_08324_),
    .X(net914));
 sg13g2_buf_2 fanout915 (.A(_08302_),
    .X(net915));
 sg13g2_buf_4 fanout916 (.X(net916),
    .A(_08281_));
 sg13g2_buf_4 fanout917 (.X(net917),
    .A(_08274_));
 sg13g2_buf_8 fanout918 (.A(_08268_),
    .X(net918));
 sg13g2_buf_8 fanout919 (.A(_08263_),
    .X(net919));
 sg13g2_buf_2 fanout920 (.A(_08261_),
    .X(net920));
 sg13g2_buf_2 fanout921 (.A(_07239_),
    .X(net921));
 sg13g2_buf_2 fanout922 (.A(_07173_),
    .X(net922));
 sg13g2_buf_2 fanout923 (.A(_07171_),
    .X(net923));
 sg13g2_buf_2 fanout924 (.A(_07156_),
    .X(net924));
 sg13g2_buf_2 fanout925 (.A(_06708_),
    .X(net925));
 sg13g2_buf_2 fanout926 (.A(_06387_),
    .X(net926));
 sg13g2_buf_2 fanout927 (.A(_06386_),
    .X(net927));
 sg13g2_buf_2 fanout928 (.A(_06385_),
    .X(net928));
 sg13g2_buf_2 fanout929 (.A(_06383_),
    .X(net929));
 sg13g2_buf_2 fanout930 (.A(_06359_),
    .X(net930));
 sg13g2_buf_2 fanout931 (.A(_06357_),
    .X(net931));
 sg13g2_buf_2 fanout932 (.A(_06347_),
    .X(net932));
 sg13g2_buf_2 fanout933 (.A(_06346_),
    .X(net933));
 sg13g2_buf_2 fanout934 (.A(_06344_),
    .X(net934));
 sg13g2_buf_2 fanout935 (.A(_06327_),
    .X(net935));
 sg13g2_buf_2 fanout936 (.A(_06322_),
    .X(net936));
 sg13g2_buf_2 fanout937 (.A(_06319_),
    .X(net937));
 sg13g2_buf_2 fanout938 (.A(_06311_),
    .X(net938));
 sg13g2_buf_2 fanout939 (.A(_06289_),
    .X(net939));
 sg13g2_buf_2 fanout940 (.A(_06264_),
    .X(net940));
 sg13g2_buf_2 fanout941 (.A(_05982_),
    .X(net941));
 sg13g2_buf_2 fanout942 (.A(_05981_),
    .X(net942));
 sg13g2_buf_2 fanout943 (.A(_05973_),
    .X(net943));
 sg13g2_buf_2 fanout944 (.A(_05951_),
    .X(net944));
 sg13g2_buf_2 fanout945 (.A(_05931_),
    .X(net945));
 sg13g2_buf_2 fanout946 (.A(_05930_),
    .X(net946));
 sg13g2_buf_2 fanout947 (.A(_05922_),
    .X(net947));
 sg13g2_buf_2 fanout948 (.A(_05913_),
    .X(net948));
 sg13g2_buf_2 fanout949 (.A(_05824_),
    .X(net949));
 sg13g2_buf_2 fanout950 (.A(_05816_),
    .X(net950));
 sg13g2_buf_2 fanout951 (.A(_05811_),
    .X(net951));
 sg13g2_buf_2 fanout952 (.A(_04954_),
    .X(net952));
 sg13g2_buf_2 fanout953 (.A(_04771_),
    .X(net953));
 sg13g2_buf_2 fanout954 (.A(_04762_),
    .X(net954));
 sg13g2_buf_2 fanout955 (.A(_04693_),
    .X(net955));
 sg13g2_buf_2 fanout956 (.A(_04656_),
    .X(net956));
 sg13g2_buf_2 fanout957 (.A(_04561_),
    .X(net957));
 sg13g2_buf_2 fanout958 (.A(_04245_),
    .X(net958));
 sg13g2_buf_2 fanout959 (.A(_04244_),
    .X(net959));
 sg13g2_buf_2 fanout960 (.A(_03632_),
    .X(net960));
 sg13g2_buf_2 fanout961 (.A(_03598_),
    .X(net961));
 sg13g2_buf_2 fanout962 (.A(_03105_),
    .X(net962));
 sg13g2_buf_2 fanout963 (.A(_03103_),
    .X(net963));
 sg13g2_buf_2 fanout964 (.A(_03101_),
    .X(net964));
 sg13g2_buf_4 fanout965 (.X(net965),
    .A(_03096_));
 sg13g2_buf_2 fanout966 (.A(_03093_),
    .X(net966));
 sg13g2_buf_2 fanout967 (.A(_03057_),
    .X(net967));
 sg13g2_buf_2 fanout968 (.A(_02963_),
    .X(net968));
 sg13g2_buf_2 fanout969 (.A(_02918_),
    .X(net969));
 sg13g2_buf_2 fanout970 (.A(_02832_),
    .X(net970));
 sg13g2_buf_2 fanout971 (.A(_02712_),
    .X(net971));
 sg13g2_buf_2 fanout972 (.A(_02659_),
    .X(net972));
 sg13g2_buf_2 fanout973 (.A(_12611_),
    .X(net973));
 sg13g2_buf_2 fanout974 (.A(_12569_),
    .X(net974));
 sg13g2_buf_2 fanout975 (.A(_12534_),
    .X(net975));
 sg13g2_buf_2 fanout976 (.A(_12453_),
    .X(net976));
 sg13g2_buf_2 fanout977 (.A(_12447_),
    .X(net977));
 sg13g2_buf_2 fanout978 (.A(_12381_),
    .X(net978));
 sg13g2_buf_2 fanout979 (.A(_12312_),
    .X(net979));
 sg13g2_buf_2 fanout980 (.A(_12244_),
    .X(net980));
 sg13g2_buf_2 fanout981 (.A(_12235_),
    .X(net981));
 sg13g2_buf_2 fanout982 (.A(_12208_),
    .X(net982));
 sg13g2_buf_2 fanout983 (.A(_12202_),
    .X(net983));
 sg13g2_buf_2 fanout984 (.A(_12197_),
    .X(net984));
 sg13g2_buf_2 fanout985 (.A(_12136_),
    .X(net985));
 sg13g2_buf_2 fanout986 (.A(_12132_),
    .X(net986));
 sg13g2_buf_2 fanout987 (.A(_12094_),
    .X(net987));
 sg13g2_buf_4 fanout988 (.X(net988),
    .A(_12067_));
 sg13g2_buf_4 fanout989 (.X(net989),
    .A(_12047_));
 sg13g2_buf_4 fanout990 (.X(net990),
    .A(_12031_));
 sg13g2_buf_2 fanout991 (.A(_12011_),
    .X(net991));
 sg13g2_buf_4 fanout992 (.X(net992),
    .A(_12007_));
 sg13g2_buf_2 fanout993 (.A(_11985_),
    .X(net993));
 sg13g2_buf_2 fanout994 (.A(_11937_),
    .X(net994));
 sg13g2_buf_2 fanout995 (.A(_11918_),
    .X(net995));
 sg13g2_buf_2 fanout996 (.A(_11913_),
    .X(net996));
 sg13g2_buf_2 fanout997 (.A(_11472_),
    .X(net997));
 sg13g2_buf_2 fanout998 (.A(_11431_),
    .X(net998));
 sg13g2_buf_2 fanout999 (.A(_11409_),
    .X(net999));
 sg13g2_buf_2 fanout1000 (.A(_11395_),
    .X(net1000));
 sg13g2_buf_2 fanout1001 (.A(_11275_),
    .X(net1001));
 sg13g2_buf_2 fanout1002 (.A(_11270_),
    .X(net1002));
 sg13g2_buf_2 fanout1003 (.A(_11269_),
    .X(net1003));
 sg13g2_buf_2 fanout1004 (.A(_11243_),
    .X(net1004));
 sg13g2_buf_2 fanout1005 (.A(_10642_),
    .X(net1005));
 sg13g2_buf_2 fanout1006 (.A(_10424_),
    .X(net1006));
 sg13g2_buf_2 fanout1007 (.A(_10165_),
    .X(net1007));
 sg13g2_buf_2 fanout1008 (.A(_10156_),
    .X(net1008));
 sg13g2_buf_2 fanout1009 (.A(_10144_),
    .X(net1009));
 sg13g2_buf_2 fanout1010 (.A(_10139_),
    .X(net1010));
 sg13g2_buf_2 fanout1011 (.A(_10060_),
    .X(net1011));
 sg13g2_buf_2 fanout1012 (.A(_10053_),
    .X(net1012));
 sg13g2_buf_2 fanout1013 (.A(_10043_),
    .X(net1013));
 sg13g2_buf_2 fanout1014 (.A(_10036_),
    .X(net1014));
 sg13g2_buf_2 fanout1015 (.A(_10025_),
    .X(net1015));
 sg13g2_buf_2 fanout1016 (.A(_09942_),
    .X(net1016));
 sg13g2_buf_2 fanout1017 (.A(_09936_),
    .X(net1017));
 sg13g2_buf_2 fanout1018 (.A(_09929_),
    .X(net1018));
 sg13g2_buf_2 fanout1019 (.A(_09911_),
    .X(net1019));
 sg13g2_buf_2 fanout1020 (.A(_09908_),
    .X(net1020));
 sg13g2_buf_2 fanout1021 (.A(_09902_),
    .X(net1021));
 sg13g2_buf_2 fanout1022 (.A(_09896_),
    .X(net1022));
 sg13g2_buf_2 fanout1023 (.A(_09871_),
    .X(net1023));
 sg13g2_buf_2 fanout1024 (.A(_09860_),
    .X(net1024));
 sg13g2_buf_2 fanout1025 (.A(_09775_),
    .X(net1025));
 sg13g2_buf_2 fanout1026 (.A(_09732_),
    .X(net1026));
 sg13g2_buf_2 fanout1027 (.A(_09719_),
    .X(net1027));
 sg13g2_buf_2 fanout1028 (.A(_09274_),
    .X(net1028));
 sg13g2_buf_2 fanout1029 (.A(_09218_),
    .X(net1029));
 sg13g2_buf_2 fanout1030 (.A(_09164_),
    .X(net1030));
 sg13g2_buf_2 fanout1031 (.A(_09144_),
    .X(net1031));
 sg13g2_buf_2 fanout1032 (.A(_09100_),
    .X(net1032));
 sg13g2_buf_2 fanout1033 (.A(_09098_),
    .X(net1033));
 sg13g2_buf_2 fanout1034 (.A(_09058_),
    .X(net1034));
 sg13g2_buf_2 fanout1035 (.A(_09050_),
    .X(net1035));
 sg13g2_buf_2 fanout1036 (.A(_09033_),
    .X(net1036));
 sg13g2_buf_4 fanout1037 (.X(net1037),
    .A(_09025_));
 sg13g2_buf_2 fanout1038 (.A(_09021_),
    .X(net1038));
 sg13g2_buf_2 fanout1039 (.A(_08962_),
    .X(net1039));
 sg13g2_buf_2 fanout1040 (.A(_08959_),
    .X(net1040));
 sg13g2_buf_2 fanout1041 (.A(_08933_),
    .X(net1041));
 sg13g2_buf_2 fanout1042 (.A(_08911_),
    .X(net1042));
 sg13g2_buf_2 fanout1043 (.A(_08882_),
    .X(net1043));
 sg13g2_buf_2 fanout1044 (.A(_08709_),
    .X(net1044));
 sg13g2_buf_2 fanout1045 (.A(_08705_),
    .X(net1045));
 sg13g2_buf_2 fanout1046 (.A(_08667_),
    .X(net1046));
 sg13g2_buf_2 fanout1047 (.A(_08648_),
    .X(net1047));
 sg13g2_buf_4 fanout1048 (.X(net1048),
    .A(_08462_));
 sg13g2_buf_2 fanout1049 (.A(_08381_),
    .X(net1049));
 sg13g2_buf_2 fanout1050 (.A(_08362_),
    .X(net1050));
 sg13g2_buf_2 fanout1051 (.A(_08330_),
    .X(net1051));
 sg13g2_buf_2 fanout1052 (.A(_08323_),
    .X(net1052));
 sg13g2_buf_4 fanout1053 (.X(net1053),
    .A(_08287_));
 sg13g2_buf_4 fanout1054 (.X(net1054),
    .A(_08273_));
 sg13g2_buf_4 fanout1055 (.X(net1055),
    .A(_08237_));
 sg13g2_buf_2 fanout1056 (.A(_08184_),
    .X(net1056));
 sg13g2_buf_2 fanout1057 (.A(_08169_),
    .X(net1057));
 sg13g2_buf_4 fanout1058 (.X(net1058),
    .A(_08161_));
 sg13g2_buf_2 fanout1059 (.A(_08154_),
    .X(net1059));
 sg13g2_buf_8 fanout1060 (.A(_08150_),
    .X(net1060));
 sg13g2_buf_4 fanout1061 (.X(net1061),
    .A(_08143_));
 sg13g2_buf_4 fanout1062 (.X(net1062),
    .A(_08138_));
 sg13g2_buf_2 fanout1063 (.A(_08122_),
    .X(net1063));
 sg13g2_buf_2 fanout1064 (.A(_07937_),
    .X(net1064));
 sg13g2_buf_2 fanout1065 (.A(_07935_),
    .X(net1065));
 sg13g2_buf_2 fanout1066 (.A(_07919_),
    .X(net1066));
 sg13g2_buf_2 fanout1067 (.A(_07871_),
    .X(net1067));
 sg13g2_buf_2 fanout1068 (.A(_07260_),
    .X(net1068));
 sg13g2_buf_2 fanout1069 (.A(_07175_),
    .X(net1069));
 sg13g2_buf_2 fanout1070 (.A(_07169_),
    .X(net1070));
 sg13g2_buf_2 fanout1071 (.A(_07157_),
    .X(net1071));
 sg13g2_buf_2 fanout1072 (.A(_05803_),
    .X(net1072));
 sg13g2_buf_2 fanout1073 (.A(_05629_),
    .X(net1073));
 sg13g2_buf_2 fanout1074 (.A(_02875_),
    .X(net1074));
 sg13g2_buf_2 fanout1075 (.A(_02862_),
    .X(net1075));
 sg13g2_buf_2 fanout1076 (.A(_02726_),
    .X(net1076));
 sg13g2_buf_2 fanout1077 (.A(_12560_),
    .X(net1077));
 sg13g2_buf_2 fanout1078 (.A(_12262_),
    .X(net1078));
 sg13g2_buf_2 fanout1079 (.A(_12122_),
    .X(net1079));
 sg13g2_buf_2 fanout1080 (.A(_12113_),
    .X(net1080));
 sg13g2_buf_2 fanout1081 (.A(_12107_),
    .X(net1081));
 sg13g2_buf_2 fanout1082 (.A(_12066_),
    .X(net1082));
 sg13g2_buf_2 fanout1083 (.A(_12046_),
    .X(net1083));
 sg13g2_buf_2 fanout1084 (.A(_12030_),
    .X(net1084));
 sg13g2_buf_2 fanout1085 (.A(_12012_),
    .X(net1085));
 sg13g2_buf_2 fanout1086 (.A(_12009_),
    .X(net1086));
 sg13g2_buf_2 fanout1087 (.A(_12006_),
    .X(net1087));
 sg13g2_buf_2 fanout1088 (.A(_11981_),
    .X(net1088));
 sg13g2_buf_2 fanout1089 (.A(_11964_),
    .X(net1089));
 sg13g2_buf_2 fanout1090 (.A(_11962_),
    .X(net1090));
 sg13g2_buf_2 fanout1091 (.A(_11956_),
    .X(net1091));
 sg13g2_buf_2 fanout1092 (.A(_11763_),
    .X(net1092));
 sg13g2_buf_2 fanout1093 (.A(_11698_),
    .X(net1093));
 sg13g2_buf_2 fanout1094 (.A(_11680_),
    .X(net1094));
 sg13g2_buf_2 fanout1095 (.A(_10963_),
    .X(net1095));
 sg13g2_buf_2 fanout1096 (.A(_10725_),
    .X(net1096));
 sg13g2_buf_2 fanout1097 (.A(_10627_),
    .X(net1097));
 sg13g2_buf_2 fanout1098 (.A(_10141_),
    .X(net1098));
 sg13g2_buf_2 fanout1099 (.A(_10138_),
    .X(net1099));
 sg13g2_buf_2 fanout1100 (.A(_10134_),
    .X(net1100));
 sg13g2_buf_2 fanout1101 (.A(_10129_),
    .X(net1101));
 sg13g2_buf_2 fanout1102 (.A(_10023_),
    .X(net1102));
 sg13g2_buf_2 fanout1103 (.A(_10019_),
    .X(net1103));
 sg13g2_buf_2 fanout1104 (.A(_09910_),
    .X(net1104));
 sg13g2_buf_2 fanout1105 (.A(_09895_),
    .X(net1105));
 sg13g2_buf_2 fanout1106 (.A(_09890_),
    .X(net1106));
 sg13g2_buf_2 fanout1107 (.A(_09721_),
    .X(net1107));
 sg13g2_buf_2 fanout1108 (.A(_09209_),
    .X(net1108));
 sg13g2_buf_2 fanout1109 (.A(_09139_),
    .X(net1109));
 sg13g2_buf_2 fanout1110 (.A(_09111_),
    .X(net1110));
 sg13g2_buf_2 fanout1111 (.A(_09038_),
    .X(net1111));
 sg13g2_buf_2 fanout1112 (.A(_09032_),
    .X(net1112));
 sg13g2_buf_2 fanout1113 (.A(_08958_),
    .X(net1113));
 sg13g2_buf_2 fanout1114 (.A(_08881_),
    .X(net1114));
 sg13g2_buf_2 fanout1115 (.A(_08290_),
    .X(net1115));
 sg13g2_buf_2 fanout1116 (.A(_08286_),
    .X(net1116));
 sg13g2_buf_2 fanout1117 (.A(_08225_),
    .X(net1117));
 sg13g2_buf_2 fanout1118 (.A(_08189_),
    .X(net1118));
 sg13g2_buf_2 fanout1119 (.A(_08186_),
    .X(net1119));
 sg13g2_buf_4 fanout1120 (.X(net1120),
    .A(_08142_));
 sg13g2_buf_2 fanout1121 (.A(_08140_),
    .X(net1121));
 sg13g2_buf_2 fanout1122 (.A(_08124_),
    .X(net1122));
 sg13g2_buf_2 fanout1123 (.A(_08121_),
    .X(net1123));
 sg13g2_tiehi _27418__1124 (.L_HI(net1124));
 sg13g2_tiehi _27419__1125 (.L_HI(net1125));
 sg13g2_tiehi _27420__1126 (.L_HI(net1126));
 sg13g2_tiehi _27421__1127 (.L_HI(net1127));
 sg13g2_tiehi _27422__1128 (.L_HI(net1128));
 sg13g2_tiehi \cpu.dcache.r_data[0][0]$_DFFE_PP__1129  (.L_HI(net1129));
 sg13g2_tiehi \cpu.dcache.r_data[0][10]$_DFFE_PP__1130  (.L_HI(net1130));
 sg13g2_tiehi \cpu.dcache.r_data[0][11]$_DFFE_PP__1131  (.L_HI(net1131));
 sg13g2_tiehi \cpu.dcache.r_data[0][12]$_DFFE_PP__1132  (.L_HI(net1132));
 sg13g2_tiehi \cpu.dcache.r_data[0][13]$_DFFE_PP__1133  (.L_HI(net1133));
 sg13g2_tiehi \cpu.dcache.r_data[0][14]$_DFFE_PP__1134  (.L_HI(net1134));
 sg13g2_tiehi \cpu.dcache.r_data[0][15]$_DFFE_PP__1135  (.L_HI(net1135));
 sg13g2_tiehi \cpu.dcache.r_data[0][16]$_DFFE_PP__1136  (.L_HI(net1136));
 sg13g2_tiehi \cpu.dcache.r_data[0][17]$_DFFE_PP__1137  (.L_HI(net1137));
 sg13g2_tiehi \cpu.dcache.r_data[0][18]$_DFFE_PP__1138  (.L_HI(net1138));
 sg13g2_tiehi \cpu.dcache.r_data[0][19]$_DFFE_PP__1139  (.L_HI(net1139));
 sg13g2_tiehi \cpu.dcache.r_data[0][1]$_DFFE_PP__1140  (.L_HI(net1140));
 sg13g2_tiehi \cpu.dcache.r_data[0][20]$_DFFE_PP__1141  (.L_HI(net1141));
 sg13g2_tiehi \cpu.dcache.r_data[0][21]$_DFFE_PP__1142  (.L_HI(net1142));
 sg13g2_tiehi \cpu.dcache.r_data[0][22]$_DFFE_PP__1143  (.L_HI(net1143));
 sg13g2_tiehi \cpu.dcache.r_data[0][23]$_DFFE_PP__1144  (.L_HI(net1144));
 sg13g2_tiehi \cpu.dcache.r_data[0][24]$_DFFE_PP__1145  (.L_HI(net1145));
 sg13g2_tiehi \cpu.dcache.r_data[0][25]$_DFFE_PP__1146  (.L_HI(net1146));
 sg13g2_tiehi \cpu.dcache.r_data[0][26]$_DFFE_PP__1147  (.L_HI(net1147));
 sg13g2_tiehi \cpu.dcache.r_data[0][27]$_DFFE_PP__1148  (.L_HI(net1148));
 sg13g2_tiehi \cpu.dcache.r_data[0][28]$_DFFE_PP__1149  (.L_HI(net1149));
 sg13g2_tiehi \cpu.dcache.r_data[0][29]$_DFFE_PP__1150  (.L_HI(net1150));
 sg13g2_tiehi \cpu.dcache.r_data[0][2]$_DFFE_PP__1151  (.L_HI(net1151));
 sg13g2_tiehi \cpu.dcache.r_data[0][30]$_DFFE_PP__1152  (.L_HI(net1152));
 sg13g2_tiehi \cpu.dcache.r_data[0][31]$_DFFE_PP__1153  (.L_HI(net1153));
 sg13g2_tiehi \cpu.dcache.r_data[0][3]$_DFFE_PP__1154  (.L_HI(net1154));
 sg13g2_tiehi \cpu.dcache.r_data[0][4]$_DFFE_PP__1155  (.L_HI(net1155));
 sg13g2_tiehi \cpu.dcache.r_data[0][5]$_DFFE_PP__1156  (.L_HI(net1156));
 sg13g2_tiehi \cpu.dcache.r_data[0][6]$_DFFE_PP__1157  (.L_HI(net1157));
 sg13g2_tiehi \cpu.dcache.r_data[0][7]$_DFFE_PP__1158  (.L_HI(net1158));
 sg13g2_tiehi \cpu.dcache.r_data[0][8]$_DFFE_PP__1159  (.L_HI(net1159));
 sg13g2_tiehi \cpu.dcache.r_data[0][9]$_DFFE_PP__1160  (.L_HI(net1160));
 sg13g2_tiehi \cpu.dcache.r_data[1][0]$_DFFE_PP__1161  (.L_HI(net1161));
 sg13g2_tiehi \cpu.dcache.r_data[1][10]$_DFFE_PP__1162  (.L_HI(net1162));
 sg13g2_tiehi \cpu.dcache.r_data[1][11]$_DFFE_PP__1163  (.L_HI(net1163));
 sg13g2_tiehi \cpu.dcache.r_data[1][12]$_DFFE_PP__1164  (.L_HI(net1164));
 sg13g2_tiehi \cpu.dcache.r_data[1][13]$_DFFE_PP__1165  (.L_HI(net1165));
 sg13g2_tiehi \cpu.dcache.r_data[1][14]$_DFFE_PP__1166  (.L_HI(net1166));
 sg13g2_tiehi \cpu.dcache.r_data[1][15]$_DFFE_PP__1167  (.L_HI(net1167));
 sg13g2_tiehi \cpu.dcache.r_data[1][16]$_DFFE_PP__1168  (.L_HI(net1168));
 sg13g2_tiehi \cpu.dcache.r_data[1][17]$_DFFE_PP__1169  (.L_HI(net1169));
 sg13g2_tiehi \cpu.dcache.r_data[1][18]$_DFFE_PP__1170  (.L_HI(net1170));
 sg13g2_tiehi \cpu.dcache.r_data[1][19]$_DFFE_PP__1171  (.L_HI(net1171));
 sg13g2_tiehi \cpu.dcache.r_data[1][1]$_DFFE_PP__1172  (.L_HI(net1172));
 sg13g2_tiehi \cpu.dcache.r_data[1][20]$_DFFE_PP__1173  (.L_HI(net1173));
 sg13g2_tiehi \cpu.dcache.r_data[1][21]$_DFFE_PP__1174  (.L_HI(net1174));
 sg13g2_tiehi \cpu.dcache.r_data[1][22]$_DFFE_PP__1175  (.L_HI(net1175));
 sg13g2_tiehi \cpu.dcache.r_data[1][23]$_DFFE_PP__1176  (.L_HI(net1176));
 sg13g2_tiehi \cpu.dcache.r_data[1][24]$_DFFE_PP__1177  (.L_HI(net1177));
 sg13g2_tiehi \cpu.dcache.r_data[1][25]$_DFFE_PP__1178  (.L_HI(net1178));
 sg13g2_tiehi \cpu.dcache.r_data[1][26]$_DFFE_PP__1179  (.L_HI(net1179));
 sg13g2_tiehi \cpu.dcache.r_data[1][27]$_DFFE_PP__1180  (.L_HI(net1180));
 sg13g2_tiehi \cpu.dcache.r_data[1][28]$_DFFE_PP__1181  (.L_HI(net1181));
 sg13g2_tiehi \cpu.dcache.r_data[1][29]$_DFFE_PP__1182  (.L_HI(net1182));
 sg13g2_tiehi \cpu.dcache.r_data[1][2]$_DFFE_PP__1183  (.L_HI(net1183));
 sg13g2_tiehi \cpu.dcache.r_data[1][30]$_DFFE_PP__1184  (.L_HI(net1184));
 sg13g2_tiehi \cpu.dcache.r_data[1][31]$_DFFE_PP__1185  (.L_HI(net1185));
 sg13g2_tiehi \cpu.dcache.r_data[1][3]$_DFFE_PP__1186  (.L_HI(net1186));
 sg13g2_tiehi \cpu.dcache.r_data[1][4]$_DFFE_PP__1187  (.L_HI(net1187));
 sg13g2_tiehi \cpu.dcache.r_data[1][5]$_DFFE_PP__1188  (.L_HI(net1188));
 sg13g2_tiehi \cpu.dcache.r_data[1][6]$_DFFE_PP__1189  (.L_HI(net1189));
 sg13g2_tiehi \cpu.dcache.r_data[1][7]$_DFFE_PP__1190  (.L_HI(net1190));
 sg13g2_tiehi \cpu.dcache.r_data[1][8]$_DFFE_PP__1191  (.L_HI(net1191));
 sg13g2_tiehi \cpu.dcache.r_data[1][9]$_DFFE_PP__1192  (.L_HI(net1192));
 sg13g2_tiehi \cpu.dcache.r_data[2][0]$_DFFE_PP__1193  (.L_HI(net1193));
 sg13g2_tiehi \cpu.dcache.r_data[2][10]$_DFFE_PP__1194  (.L_HI(net1194));
 sg13g2_tiehi \cpu.dcache.r_data[2][11]$_DFFE_PP__1195  (.L_HI(net1195));
 sg13g2_tiehi \cpu.dcache.r_data[2][12]$_DFFE_PP__1196  (.L_HI(net1196));
 sg13g2_tiehi \cpu.dcache.r_data[2][13]$_DFFE_PP__1197  (.L_HI(net1197));
 sg13g2_tiehi \cpu.dcache.r_data[2][14]$_DFFE_PP__1198  (.L_HI(net1198));
 sg13g2_tiehi \cpu.dcache.r_data[2][15]$_DFFE_PP__1199  (.L_HI(net1199));
 sg13g2_tiehi \cpu.dcache.r_data[2][16]$_DFFE_PP__1200  (.L_HI(net1200));
 sg13g2_tiehi \cpu.dcache.r_data[2][17]$_DFFE_PP__1201  (.L_HI(net1201));
 sg13g2_tiehi \cpu.dcache.r_data[2][18]$_DFFE_PP__1202  (.L_HI(net1202));
 sg13g2_tiehi \cpu.dcache.r_data[2][19]$_DFFE_PP__1203  (.L_HI(net1203));
 sg13g2_tiehi \cpu.dcache.r_data[2][1]$_DFFE_PP__1204  (.L_HI(net1204));
 sg13g2_tiehi \cpu.dcache.r_data[2][20]$_DFFE_PP__1205  (.L_HI(net1205));
 sg13g2_tiehi \cpu.dcache.r_data[2][21]$_DFFE_PP__1206  (.L_HI(net1206));
 sg13g2_tiehi \cpu.dcache.r_data[2][22]$_DFFE_PP__1207  (.L_HI(net1207));
 sg13g2_tiehi \cpu.dcache.r_data[2][23]$_DFFE_PP__1208  (.L_HI(net1208));
 sg13g2_tiehi \cpu.dcache.r_data[2][24]$_DFFE_PP__1209  (.L_HI(net1209));
 sg13g2_tiehi \cpu.dcache.r_data[2][25]$_DFFE_PP__1210  (.L_HI(net1210));
 sg13g2_tiehi \cpu.dcache.r_data[2][26]$_DFFE_PP__1211  (.L_HI(net1211));
 sg13g2_tiehi \cpu.dcache.r_data[2][27]$_DFFE_PP__1212  (.L_HI(net1212));
 sg13g2_tiehi \cpu.dcache.r_data[2][28]$_DFFE_PP__1213  (.L_HI(net1213));
 sg13g2_tiehi \cpu.dcache.r_data[2][29]$_DFFE_PP__1214  (.L_HI(net1214));
 sg13g2_tiehi \cpu.dcache.r_data[2][2]$_DFFE_PP__1215  (.L_HI(net1215));
 sg13g2_tiehi \cpu.dcache.r_data[2][30]$_DFFE_PP__1216  (.L_HI(net1216));
 sg13g2_tiehi \cpu.dcache.r_data[2][31]$_DFFE_PP__1217  (.L_HI(net1217));
 sg13g2_tiehi \cpu.dcache.r_data[2][3]$_DFFE_PP__1218  (.L_HI(net1218));
 sg13g2_tiehi \cpu.dcache.r_data[2][4]$_DFFE_PP__1219  (.L_HI(net1219));
 sg13g2_tiehi \cpu.dcache.r_data[2][5]$_DFFE_PP__1220  (.L_HI(net1220));
 sg13g2_tiehi \cpu.dcache.r_data[2][6]$_DFFE_PP__1221  (.L_HI(net1221));
 sg13g2_tiehi \cpu.dcache.r_data[2][7]$_DFFE_PP__1222  (.L_HI(net1222));
 sg13g2_tiehi \cpu.dcache.r_data[2][8]$_DFFE_PP__1223  (.L_HI(net1223));
 sg13g2_tiehi \cpu.dcache.r_data[2][9]$_DFFE_PP__1224  (.L_HI(net1224));
 sg13g2_tiehi \cpu.dcache.r_data[3][0]$_DFFE_PP__1225  (.L_HI(net1225));
 sg13g2_tiehi \cpu.dcache.r_data[3][10]$_DFFE_PP__1226  (.L_HI(net1226));
 sg13g2_tiehi \cpu.dcache.r_data[3][11]$_DFFE_PP__1227  (.L_HI(net1227));
 sg13g2_tiehi \cpu.dcache.r_data[3][12]$_DFFE_PP__1228  (.L_HI(net1228));
 sg13g2_tiehi \cpu.dcache.r_data[3][13]$_DFFE_PP__1229  (.L_HI(net1229));
 sg13g2_tiehi \cpu.dcache.r_data[3][14]$_DFFE_PP__1230  (.L_HI(net1230));
 sg13g2_tiehi \cpu.dcache.r_data[3][15]$_DFFE_PP__1231  (.L_HI(net1231));
 sg13g2_tiehi \cpu.dcache.r_data[3][16]$_DFFE_PP__1232  (.L_HI(net1232));
 sg13g2_tiehi \cpu.dcache.r_data[3][17]$_DFFE_PP__1233  (.L_HI(net1233));
 sg13g2_tiehi \cpu.dcache.r_data[3][18]$_DFFE_PP__1234  (.L_HI(net1234));
 sg13g2_tiehi \cpu.dcache.r_data[3][19]$_DFFE_PP__1235  (.L_HI(net1235));
 sg13g2_tiehi \cpu.dcache.r_data[3][1]$_DFFE_PP__1236  (.L_HI(net1236));
 sg13g2_tiehi \cpu.dcache.r_data[3][20]$_DFFE_PP__1237  (.L_HI(net1237));
 sg13g2_tiehi \cpu.dcache.r_data[3][21]$_DFFE_PP__1238  (.L_HI(net1238));
 sg13g2_tiehi \cpu.dcache.r_data[3][22]$_DFFE_PP__1239  (.L_HI(net1239));
 sg13g2_tiehi \cpu.dcache.r_data[3][23]$_DFFE_PP__1240  (.L_HI(net1240));
 sg13g2_tiehi \cpu.dcache.r_data[3][24]$_DFFE_PP__1241  (.L_HI(net1241));
 sg13g2_tiehi \cpu.dcache.r_data[3][25]$_DFFE_PP__1242  (.L_HI(net1242));
 sg13g2_tiehi \cpu.dcache.r_data[3][26]$_DFFE_PP__1243  (.L_HI(net1243));
 sg13g2_tiehi \cpu.dcache.r_data[3][27]$_DFFE_PP__1244  (.L_HI(net1244));
 sg13g2_tiehi \cpu.dcache.r_data[3][28]$_DFFE_PP__1245  (.L_HI(net1245));
 sg13g2_tiehi \cpu.dcache.r_data[3][29]$_DFFE_PP__1246  (.L_HI(net1246));
 sg13g2_tiehi \cpu.dcache.r_data[3][2]$_DFFE_PP__1247  (.L_HI(net1247));
 sg13g2_tiehi \cpu.dcache.r_data[3][30]$_DFFE_PP__1248  (.L_HI(net1248));
 sg13g2_tiehi \cpu.dcache.r_data[3][31]$_DFFE_PP__1249  (.L_HI(net1249));
 sg13g2_tiehi \cpu.dcache.r_data[3][3]$_DFFE_PP__1250  (.L_HI(net1250));
 sg13g2_tiehi \cpu.dcache.r_data[3][4]$_DFFE_PP__1251  (.L_HI(net1251));
 sg13g2_tiehi \cpu.dcache.r_data[3][5]$_DFFE_PP__1252  (.L_HI(net1252));
 sg13g2_tiehi \cpu.dcache.r_data[3][6]$_DFFE_PP__1253  (.L_HI(net1253));
 sg13g2_tiehi \cpu.dcache.r_data[3][7]$_DFFE_PP__1254  (.L_HI(net1254));
 sg13g2_tiehi \cpu.dcache.r_data[3][8]$_DFFE_PP__1255  (.L_HI(net1255));
 sg13g2_tiehi \cpu.dcache.r_data[3][9]$_DFFE_PP__1256  (.L_HI(net1256));
 sg13g2_tiehi \cpu.dcache.r_data[4][0]$_DFFE_PP__1257  (.L_HI(net1257));
 sg13g2_tiehi \cpu.dcache.r_data[4][10]$_DFFE_PP__1258  (.L_HI(net1258));
 sg13g2_tiehi \cpu.dcache.r_data[4][11]$_DFFE_PP__1259  (.L_HI(net1259));
 sg13g2_tiehi \cpu.dcache.r_data[4][12]$_DFFE_PP__1260  (.L_HI(net1260));
 sg13g2_tiehi \cpu.dcache.r_data[4][13]$_DFFE_PP__1261  (.L_HI(net1261));
 sg13g2_tiehi \cpu.dcache.r_data[4][14]$_DFFE_PP__1262  (.L_HI(net1262));
 sg13g2_tiehi \cpu.dcache.r_data[4][15]$_DFFE_PP__1263  (.L_HI(net1263));
 sg13g2_tiehi \cpu.dcache.r_data[4][16]$_DFFE_PP__1264  (.L_HI(net1264));
 sg13g2_tiehi \cpu.dcache.r_data[4][17]$_DFFE_PP__1265  (.L_HI(net1265));
 sg13g2_tiehi \cpu.dcache.r_data[4][18]$_DFFE_PP__1266  (.L_HI(net1266));
 sg13g2_tiehi \cpu.dcache.r_data[4][19]$_DFFE_PP__1267  (.L_HI(net1267));
 sg13g2_tiehi \cpu.dcache.r_data[4][1]$_DFFE_PP__1268  (.L_HI(net1268));
 sg13g2_tiehi \cpu.dcache.r_data[4][20]$_DFFE_PP__1269  (.L_HI(net1269));
 sg13g2_tiehi \cpu.dcache.r_data[4][21]$_DFFE_PP__1270  (.L_HI(net1270));
 sg13g2_tiehi \cpu.dcache.r_data[4][22]$_DFFE_PP__1271  (.L_HI(net1271));
 sg13g2_tiehi \cpu.dcache.r_data[4][23]$_DFFE_PP__1272  (.L_HI(net1272));
 sg13g2_tiehi \cpu.dcache.r_data[4][24]$_DFFE_PP__1273  (.L_HI(net1273));
 sg13g2_tiehi \cpu.dcache.r_data[4][25]$_DFFE_PP__1274  (.L_HI(net1274));
 sg13g2_tiehi \cpu.dcache.r_data[4][26]$_DFFE_PP__1275  (.L_HI(net1275));
 sg13g2_tiehi \cpu.dcache.r_data[4][27]$_DFFE_PP__1276  (.L_HI(net1276));
 sg13g2_tiehi \cpu.dcache.r_data[4][28]$_DFFE_PP__1277  (.L_HI(net1277));
 sg13g2_tiehi \cpu.dcache.r_data[4][29]$_DFFE_PP__1278  (.L_HI(net1278));
 sg13g2_tiehi \cpu.dcache.r_data[4][2]$_DFFE_PP__1279  (.L_HI(net1279));
 sg13g2_tiehi \cpu.dcache.r_data[4][30]$_DFFE_PP__1280  (.L_HI(net1280));
 sg13g2_tiehi \cpu.dcache.r_data[4][31]$_DFFE_PP__1281  (.L_HI(net1281));
 sg13g2_tiehi \cpu.dcache.r_data[4][3]$_DFFE_PP__1282  (.L_HI(net1282));
 sg13g2_tiehi \cpu.dcache.r_data[4][4]$_DFFE_PP__1283  (.L_HI(net1283));
 sg13g2_tiehi \cpu.dcache.r_data[4][5]$_DFFE_PP__1284  (.L_HI(net1284));
 sg13g2_tiehi \cpu.dcache.r_data[4][6]$_DFFE_PP__1285  (.L_HI(net1285));
 sg13g2_tiehi \cpu.dcache.r_data[4][7]$_DFFE_PP__1286  (.L_HI(net1286));
 sg13g2_tiehi \cpu.dcache.r_data[4][8]$_DFFE_PP__1287  (.L_HI(net1287));
 sg13g2_tiehi \cpu.dcache.r_data[4][9]$_DFFE_PP__1288  (.L_HI(net1288));
 sg13g2_tiehi \cpu.dcache.r_data[5][0]$_DFFE_PP__1289  (.L_HI(net1289));
 sg13g2_tiehi \cpu.dcache.r_data[5][10]$_DFFE_PP__1290  (.L_HI(net1290));
 sg13g2_tiehi \cpu.dcache.r_data[5][11]$_DFFE_PP__1291  (.L_HI(net1291));
 sg13g2_tiehi \cpu.dcache.r_data[5][12]$_DFFE_PP__1292  (.L_HI(net1292));
 sg13g2_tiehi \cpu.dcache.r_data[5][13]$_DFFE_PP__1293  (.L_HI(net1293));
 sg13g2_tiehi \cpu.dcache.r_data[5][14]$_DFFE_PP__1294  (.L_HI(net1294));
 sg13g2_tiehi \cpu.dcache.r_data[5][15]$_DFFE_PP__1295  (.L_HI(net1295));
 sg13g2_tiehi \cpu.dcache.r_data[5][16]$_DFFE_PP__1296  (.L_HI(net1296));
 sg13g2_tiehi \cpu.dcache.r_data[5][17]$_DFFE_PP__1297  (.L_HI(net1297));
 sg13g2_tiehi \cpu.dcache.r_data[5][18]$_DFFE_PP__1298  (.L_HI(net1298));
 sg13g2_tiehi \cpu.dcache.r_data[5][19]$_DFFE_PP__1299  (.L_HI(net1299));
 sg13g2_tiehi \cpu.dcache.r_data[5][1]$_DFFE_PP__1300  (.L_HI(net1300));
 sg13g2_tiehi \cpu.dcache.r_data[5][20]$_DFFE_PP__1301  (.L_HI(net1301));
 sg13g2_tiehi \cpu.dcache.r_data[5][21]$_DFFE_PP__1302  (.L_HI(net1302));
 sg13g2_tiehi \cpu.dcache.r_data[5][22]$_DFFE_PP__1303  (.L_HI(net1303));
 sg13g2_tiehi \cpu.dcache.r_data[5][23]$_DFFE_PP__1304  (.L_HI(net1304));
 sg13g2_tiehi \cpu.dcache.r_data[5][24]$_DFFE_PP__1305  (.L_HI(net1305));
 sg13g2_tiehi \cpu.dcache.r_data[5][25]$_DFFE_PP__1306  (.L_HI(net1306));
 sg13g2_tiehi \cpu.dcache.r_data[5][26]$_DFFE_PP__1307  (.L_HI(net1307));
 sg13g2_tiehi \cpu.dcache.r_data[5][27]$_DFFE_PP__1308  (.L_HI(net1308));
 sg13g2_tiehi \cpu.dcache.r_data[5][28]$_DFFE_PP__1309  (.L_HI(net1309));
 sg13g2_tiehi \cpu.dcache.r_data[5][29]$_DFFE_PP__1310  (.L_HI(net1310));
 sg13g2_tiehi \cpu.dcache.r_data[5][2]$_DFFE_PP__1311  (.L_HI(net1311));
 sg13g2_tiehi \cpu.dcache.r_data[5][30]$_DFFE_PP__1312  (.L_HI(net1312));
 sg13g2_tiehi \cpu.dcache.r_data[5][31]$_DFFE_PP__1313  (.L_HI(net1313));
 sg13g2_tiehi \cpu.dcache.r_data[5][3]$_DFFE_PP__1314  (.L_HI(net1314));
 sg13g2_tiehi \cpu.dcache.r_data[5][4]$_DFFE_PP__1315  (.L_HI(net1315));
 sg13g2_tiehi \cpu.dcache.r_data[5][5]$_DFFE_PP__1316  (.L_HI(net1316));
 sg13g2_tiehi \cpu.dcache.r_data[5][6]$_DFFE_PP__1317  (.L_HI(net1317));
 sg13g2_tiehi \cpu.dcache.r_data[5][7]$_DFFE_PP__1318  (.L_HI(net1318));
 sg13g2_tiehi \cpu.dcache.r_data[5][8]$_DFFE_PP__1319  (.L_HI(net1319));
 sg13g2_tiehi \cpu.dcache.r_data[5][9]$_DFFE_PP__1320  (.L_HI(net1320));
 sg13g2_tiehi \cpu.dcache.r_data[6][0]$_DFFE_PP__1321  (.L_HI(net1321));
 sg13g2_tiehi \cpu.dcache.r_data[6][10]$_DFFE_PP__1322  (.L_HI(net1322));
 sg13g2_tiehi \cpu.dcache.r_data[6][11]$_DFFE_PP__1323  (.L_HI(net1323));
 sg13g2_tiehi \cpu.dcache.r_data[6][12]$_DFFE_PP__1324  (.L_HI(net1324));
 sg13g2_tiehi \cpu.dcache.r_data[6][13]$_DFFE_PP__1325  (.L_HI(net1325));
 sg13g2_tiehi \cpu.dcache.r_data[6][14]$_DFFE_PP__1326  (.L_HI(net1326));
 sg13g2_tiehi \cpu.dcache.r_data[6][15]$_DFFE_PP__1327  (.L_HI(net1327));
 sg13g2_tiehi \cpu.dcache.r_data[6][16]$_DFFE_PP__1328  (.L_HI(net1328));
 sg13g2_tiehi \cpu.dcache.r_data[6][17]$_DFFE_PP__1329  (.L_HI(net1329));
 sg13g2_tiehi \cpu.dcache.r_data[6][18]$_DFFE_PP__1330  (.L_HI(net1330));
 sg13g2_tiehi \cpu.dcache.r_data[6][19]$_DFFE_PP__1331  (.L_HI(net1331));
 sg13g2_tiehi \cpu.dcache.r_data[6][1]$_DFFE_PP__1332  (.L_HI(net1332));
 sg13g2_tiehi \cpu.dcache.r_data[6][20]$_DFFE_PP__1333  (.L_HI(net1333));
 sg13g2_tiehi \cpu.dcache.r_data[6][21]$_DFFE_PP__1334  (.L_HI(net1334));
 sg13g2_tiehi \cpu.dcache.r_data[6][22]$_DFFE_PP__1335  (.L_HI(net1335));
 sg13g2_tiehi \cpu.dcache.r_data[6][23]$_DFFE_PP__1336  (.L_HI(net1336));
 sg13g2_tiehi \cpu.dcache.r_data[6][24]$_DFFE_PP__1337  (.L_HI(net1337));
 sg13g2_tiehi \cpu.dcache.r_data[6][25]$_DFFE_PP__1338  (.L_HI(net1338));
 sg13g2_tiehi \cpu.dcache.r_data[6][26]$_DFFE_PP__1339  (.L_HI(net1339));
 sg13g2_tiehi \cpu.dcache.r_data[6][27]$_DFFE_PP__1340  (.L_HI(net1340));
 sg13g2_tiehi \cpu.dcache.r_data[6][28]$_DFFE_PP__1341  (.L_HI(net1341));
 sg13g2_tiehi \cpu.dcache.r_data[6][29]$_DFFE_PP__1342  (.L_HI(net1342));
 sg13g2_tiehi \cpu.dcache.r_data[6][2]$_DFFE_PP__1343  (.L_HI(net1343));
 sg13g2_tiehi \cpu.dcache.r_data[6][30]$_DFFE_PP__1344  (.L_HI(net1344));
 sg13g2_tiehi \cpu.dcache.r_data[6][31]$_DFFE_PP__1345  (.L_HI(net1345));
 sg13g2_tiehi \cpu.dcache.r_data[6][3]$_DFFE_PP__1346  (.L_HI(net1346));
 sg13g2_tiehi \cpu.dcache.r_data[6][4]$_DFFE_PP__1347  (.L_HI(net1347));
 sg13g2_tiehi \cpu.dcache.r_data[6][5]$_DFFE_PP__1348  (.L_HI(net1348));
 sg13g2_tiehi \cpu.dcache.r_data[6][6]$_DFFE_PP__1349  (.L_HI(net1349));
 sg13g2_tiehi \cpu.dcache.r_data[6][7]$_DFFE_PP__1350  (.L_HI(net1350));
 sg13g2_tiehi \cpu.dcache.r_data[6][8]$_DFFE_PP__1351  (.L_HI(net1351));
 sg13g2_tiehi \cpu.dcache.r_data[6][9]$_DFFE_PP__1352  (.L_HI(net1352));
 sg13g2_tiehi \cpu.dcache.r_data[7][0]$_DFFE_PP__1353  (.L_HI(net1353));
 sg13g2_tiehi \cpu.dcache.r_data[7][10]$_DFFE_PP__1354  (.L_HI(net1354));
 sg13g2_tiehi \cpu.dcache.r_data[7][11]$_DFFE_PP__1355  (.L_HI(net1355));
 sg13g2_tiehi \cpu.dcache.r_data[7][12]$_DFFE_PP__1356  (.L_HI(net1356));
 sg13g2_tiehi \cpu.dcache.r_data[7][13]$_DFFE_PP__1357  (.L_HI(net1357));
 sg13g2_tiehi \cpu.dcache.r_data[7][14]$_DFFE_PP__1358  (.L_HI(net1358));
 sg13g2_tiehi \cpu.dcache.r_data[7][15]$_DFFE_PP__1359  (.L_HI(net1359));
 sg13g2_tiehi \cpu.dcache.r_data[7][16]$_DFFE_PP__1360  (.L_HI(net1360));
 sg13g2_tiehi \cpu.dcache.r_data[7][17]$_DFFE_PP__1361  (.L_HI(net1361));
 sg13g2_tiehi \cpu.dcache.r_data[7][18]$_DFFE_PP__1362  (.L_HI(net1362));
 sg13g2_tiehi \cpu.dcache.r_data[7][19]$_DFFE_PP__1363  (.L_HI(net1363));
 sg13g2_tiehi \cpu.dcache.r_data[7][1]$_DFFE_PP__1364  (.L_HI(net1364));
 sg13g2_tiehi \cpu.dcache.r_data[7][20]$_DFFE_PP__1365  (.L_HI(net1365));
 sg13g2_tiehi \cpu.dcache.r_data[7][21]$_DFFE_PP__1366  (.L_HI(net1366));
 sg13g2_tiehi \cpu.dcache.r_data[7][22]$_DFFE_PP__1367  (.L_HI(net1367));
 sg13g2_tiehi \cpu.dcache.r_data[7][23]$_DFFE_PP__1368  (.L_HI(net1368));
 sg13g2_tiehi \cpu.dcache.r_data[7][24]$_DFFE_PP__1369  (.L_HI(net1369));
 sg13g2_tiehi \cpu.dcache.r_data[7][25]$_DFFE_PP__1370  (.L_HI(net1370));
 sg13g2_tiehi \cpu.dcache.r_data[7][26]$_DFFE_PP__1371  (.L_HI(net1371));
 sg13g2_tiehi \cpu.dcache.r_data[7][27]$_DFFE_PP__1372  (.L_HI(net1372));
 sg13g2_tiehi \cpu.dcache.r_data[7][28]$_DFFE_PP__1373  (.L_HI(net1373));
 sg13g2_tiehi \cpu.dcache.r_data[7][29]$_DFFE_PP__1374  (.L_HI(net1374));
 sg13g2_tiehi \cpu.dcache.r_data[7][2]$_DFFE_PP__1375  (.L_HI(net1375));
 sg13g2_tiehi \cpu.dcache.r_data[7][30]$_DFFE_PP__1376  (.L_HI(net1376));
 sg13g2_tiehi \cpu.dcache.r_data[7][31]$_DFFE_PP__1377  (.L_HI(net1377));
 sg13g2_tiehi \cpu.dcache.r_data[7][3]$_DFFE_PP__1378  (.L_HI(net1378));
 sg13g2_tiehi \cpu.dcache.r_data[7][4]$_DFFE_PP__1379  (.L_HI(net1379));
 sg13g2_tiehi \cpu.dcache.r_data[7][5]$_DFFE_PP__1380  (.L_HI(net1380));
 sg13g2_tiehi \cpu.dcache.r_data[7][6]$_DFFE_PP__1381  (.L_HI(net1381));
 sg13g2_tiehi \cpu.dcache.r_data[7][7]$_DFFE_PP__1382  (.L_HI(net1382));
 sg13g2_tiehi \cpu.dcache.r_data[7][8]$_DFFE_PP__1383  (.L_HI(net1383));
 sg13g2_tiehi \cpu.dcache.r_data[7][9]$_DFFE_PP__1384  (.L_HI(net1384));
 sg13g2_tiehi \cpu.dcache.r_dirty[0]$_SDFFCE_PP1P__1385  (.L_HI(net1385));
 sg13g2_tiehi \cpu.dcache.r_dirty[1]$_SDFFCE_PP1P__1386  (.L_HI(net1386));
 sg13g2_tiehi \cpu.dcache.r_dirty[2]$_SDFFCE_PP1P__1387  (.L_HI(net1387));
 sg13g2_tiehi \cpu.dcache.r_dirty[3]$_SDFFCE_PP1P__1388  (.L_HI(net1388));
 sg13g2_tiehi \cpu.dcache.r_dirty[4]$_SDFFCE_PP1P__1389  (.L_HI(net1389));
 sg13g2_tiehi \cpu.dcache.r_dirty[5]$_SDFFCE_PP1P__1390  (.L_HI(net1390));
 sg13g2_tiehi \cpu.dcache.r_dirty[6]$_SDFFCE_PP1P__1391  (.L_HI(net1391));
 sg13g2_tiehi \cpu.dcache.r_dirty[7]$_SDFFCE_PP1P__1392  (.L_HI(net1392));
 sg13g2_tiehi \cpu.dcache.r_offset[0]$_SDFF_PN0__1393  (.L_HI(net1393));
 sg13g2_tiehi \cpu.dcache.r_offset[1]$_SDFF_PN0__1394  (.L_HI(net1394));
 sg13g2_tiehi \cpu.dcache.r_offset[2]$_SDFF_PN0__1395  (.L_HI(net1395));
 sg13g2_tiehi \cpu.dcache.r_tag[0][0]$_DFFE_PP__1396  (.L_HI(net1396));
 sg13g2_tiehi \cpu.dcache.r_tag[0][10]$_DFFE_PP__1397  (.L_HI(net1397));
 sg13g2_tiehi \cpu.dcache.r_tag[0][11]$_DFFE_PP__1398  (.L_HI(net1398));
 sg13g2_tiehi \cpu.dcache.r_tag[0][12]$_DFFE_PP__1399  (.L_HI(net1399));
 sg13g2_tiehi \cpu.dcache.r_tag[0][13]$_DFFE_PP__1400  (.L_HI(net1400));
 sg13g2_tiehi \cpu.dcache.r_tag[0][14]$_DFFE_PP__1401  (.L_HI(net1401));
 sg13g2_tiehi \cpu.dcache.r_tag[0][15]$_DFFE_PP__1402  (.L_HI(net1402));
 sg13g2_tiehi \cpu.dcache.r_tag[0][16]$_DFFE_PP__1403  (.L_HI(net1403));
 sg13g2_tiehi \cpu.dcache.r_tag[0][17]$_DFFE_PP__1404  (.L_HI(net1404));
 sg13g2_tiehi \cpu.dcache.r_tag[0][18]$_DFFE_PP__1405  (.L_HI(net1405));
 sg13g2_tiehi \cpu.dcache.r_tag[0][1]$_DFFE_PP__1406  (.L_HI(net1406));
 sg13g2_tiehi \cpu.dcache.r_tag[0][2]$_DFFE_PP__1407  (.L_HI(net1407));
 sg13g2_tiehi \cpu.dcache.r_tag[0][3]$_DFFE_PP__1408  (.L_HI(net1408));
 sg13g2_tiehi \cpu.dcache.r_tag[0][4]$_DFFE_PP__1409  (.L_HI(net1409));
 sg13g2_tiehi \cpu.dcache.r_tag[0][5]$_DFFE_PP__1410  (.L_HI(net1410));
 sg13g2_tiehi \cpu.dcache.r_tag[0][6]$_DFFE_PP__1411  (.L_HI(net1411));
 sg13g2_tiehi \cpu.dcache.r_tag[0][7]$_DFFE_PP__1412  (.L_HI(net1412));
 sg13g2_tiehi \cpu.dcache.r_tag[0][8]$_DFFE_PP__1413  (.L_HI(net1413));
 sg13g2_tiehi \cpu.dcache.r_tag[0][9]$_DFFE_PP__1414  (.L_HI(net1414));
 sg13g2_tiehi \cpu.dcache.r_tag[1][0]$_DFFE_PP__1415  (.L_HI(net1415));
 sg13g2_tiehi \cpu.dcache.r_tag[1][10]$_DFFE_PP__1416  (.L_HI(net1416));
 sg13g2_tiehi \cpu.dcache.r_tag[1][11]$_DFFE_PP__1417  (.L_HI(net1417));
 sg13g2_tiehi \cpu.dcache.r_tag[1][12]$_DFFE_PP__1418  (.L_HI(net1418));
 sg13g2_tiehi \cpu.dcache.r_tag[1][13]$_DFFE_PP__1419  (.L_HI(net1419));
 sg13g2_tiehi \cpu.dcache.r_tag[1][14]$_DFFE_PP__1420  (.L_HI(net1420));
 sg13g2_tiehi \cpu.dcache.r_tag[1][15]$_DFFE_PP__1421  (.L_HI(net1421));
 sg13g2_tiehi \cpu.dcache.r_tag[1][16]$_DFFE_PP__1422  (.L_HI(net1422));
 sg13g2_tiehi \cpu.dcache.r_tag[1][17]$_DFFE_PP__1423  (.L_HI(net1423));
 sg13g2_tiehi \cpu.dcache.r_tag[1][18]$_DFFE_PP__1424  (.L_HI(net1424));
 sg13g2_tiehi \cpu.dcache.r_tag[1][1]$_DFFE_PP__1425  (.L_HI(net1425));
 sg13g2_tiehi \cpu.dcache.r_tag[1][2]$_DFFE_PP__1426  (.L_HI(net1426));
 sg13g2_tiehi \cpu.dcache.r_tag[1][3]$_DFFE_PP__1427  (.L_HI(net1427));
 sg13g2_tiehi \cpu.dcache.r_tag[1][4]$_DFFE_PP__1428  (.L_HI(net1428));
 sg13g2_tiehi \cpu.dcache.r_tag[1][5]$_DFFE_PP__1429  (.L_HI(net1429));
 sg13g2_tiehi \cpu.dcache.r_tag[1][6]$_DFFE_PP__1430  (.L_HI(net1430));
 sg13g2_tiehi \cpu.dcache.r_tag[1][7]$_DFFE_PP__1431  (.L_HI(net1431));
 sg13g2_tiehi \cpu.dcache.r_tag[1][8]$_DFFE_PP__1432  (.L_HI(net1432));
 sg13g2_tiehi \cpu.dcache.r_tag[1][9]$_DFFE_PP__1433  (.L_HI(net1433));
 sg13g2_tiehi \cpu.dcache.r_tag[2][0]$_DFFE_PP__1434  (.L_HI(net1434));
 sg13g2_tiehi \cpu.dcache.r_tag[2][10]$_DFFE_PP__1435  (.L_HI(net1435));
 sg13g2_tiehi \cpu.dcache.r_tag[2][11]$_DFFE_PP__1436  (.L_HI(net1436));
 sg13g2_tiehi \cpu.dcache.r_tag[2][12]$_DFFE_PP__1437  (.L_HI(net1437));
 sg13g2_tiehi \cpu.dcache.r_tag[2][13]$_DFFE_PP__1438  (.L_HI(net1438));
 sg13g2_tiehi \cpu.dcache.r_tag[2][14]$_DFFE_PP__1439  (.L_HI(net1439));
 sg13g2_tiehi \cpu.dcache.r_tag[2][15]$_DFFE_PP__1440  (.L_HI(net1440));
 sg13g2_tiehi \cpu.dcache.r_tag[2][16]$_DFFE_PP__1441  (.L_HI(net1441));
 sg13g2_tiehi \cpu.dcache.r_tag[2][17]$_DFFE_PP__1442  (.L_HI(net1442));
 sg13g2_tiehi \cpu.dcache.r_tag[2][18]$_DFFE_PP__1443  (.L_HI(net1443));
 sg13g2_tiehi \cpu.dcache.r_tag[2][1]$_DFFE_PP__1444  (.L_HI(net1444));
 sg13g2_tiehi \cpu.dcache.r_tag[2][2]$_DFFE_PP__1445  (.L_HI(net1445));
 sg13g2_tiehi \cpu.dcache.r_tag[2][3]$_DFFE_PP__1446  (.L_HI(net1446));
 sg13g2_tiehi \cpu.dcache.r_tag[2][4]$_DFFE_PP__1447  (.L_HI(net1447));
 sg13g2_tiehi \cpu.dcache.r_tag[2][5]$_DFFE_PP__1448  (.L_HI(net1448));
 sg13g2_tiehi \cpu.dcache.r_tag[2][6]$_DFFE_PP__1449  (.L_HI(net1449));
 sg13g2_tiehi \cpu.dcache.r_tag[2][7]$_DFFE_PP__1450  (.L_HI(net1450));
 sg13g2_tiehi \cpu.dcache.r_tag[2][8]$_DFFE_PP__1451  (.L_HI(net1451));
 sg13g2_tiehi \cpu.dcache.r_tag[2][9]$_DFFE_PP__1452  (.L_HI(net1452));
 sg13g2_tiehi \cpu.dcache.r_tag[3][0]$_DFFE_PP__1453  (.L_HI(net1453));
 sg13g2_tiehi \cpu.dcache.r_tag[3][10]$_DFFE_PP__1454  (.L_HI(net1454));
 sg13g2_tiehi \cpu.dcache.r_tag[3][11]$_DFFE_PP__1455  (.L_HI(net1455));
 sg13g2_tiehi \cpu.dcache.r_tag[3][12]$_DFFE_PP__1456  (.L_HI(net1456));
 sg13g2_tiehi \cpu.dcache.r_tag[3][13]$_DFFE_PP__1457  (.L_HI(net1457));
 sg13g2_tiehi \cpu.dcache.r_tag[3][14]$_DFFE_PP__1458  (.L_HI(net1458));
 sg13g2_tiehi \cpu.dcache.r_tag[3][15]$_DFFE_PP__1459  (.L_HI(net1459));
 sg13g2_tiehi \cpu.dcache.r_tag[3][16]$_DFFE_PP__1460  (.L_HI(net1460));
 sg13g2_tiehi \cpu.dcache.r_tag[3][17]$_DFFE_PP__1461  (.L_HI(net1461));
 sg13g2_tiehi \cpu.dcache.r_tag[3][18]$_DFFE_PP__1462  (.L_HI(net1462));
 sg13g2_tiehi \cpu.dcache.r_tag[3][1]$_DFFE_PP__1463  (.L_HI(net1463));
 sg13g2_tiehi \cpu.dcache.r_tag[3][2]$_DFFE_PP__1464  (.L_HI(net1464));
 sg13g2_tiehi \cpu.dcache.r_tag[3][3]$_DFFE_PP__1465  (.L_HI(net1465));
 sg13g2_tiehi \cpu.dcache.r_tag[3][4]$_DFFE_PP__1466  (.L_HI(net1466));
 sg13g2_tiehi \cpu.dcache.r_tag[3][5]$_DFFE_PP__1467  (.L_HI(net1467));
 sg13g2_tiehi \cpu.dcache.r_tag[3][6]$_DFFE_PP__1468  (.L_HI(net1468));
 sg13g2_tiehi \cpu.dcache.r_tag[3][7]$_DFFE_PP__1469  (.L_HI(net1469));
 sg13g2_tiehi \cpu.dcache.r_tag[3][8]$_DFFE_PP__1470  (.L_HI(net1470));
 sg13g2_tiehi \cpu.dcache.r_tag[3][9]$_DFFE_PP__1471  (.L_HI(net1471));
 sg13g2_tiehi \cpu.dcache.r_tag[4][0]$_DFFE_PP__1472  (.L_HI(net1472));
 sg13g2_tiehi \cpu.dcache.r_tag[4][10]$_DFFE_PP__1473  (.L_HI(net1473));
 sg13g2_tiehi \cpu.dcache.r_tag[4][11]$_DFFE_PP__1474  (.L_HI(net1474));
 sg13g2_tiehi \cpu.dcache.r_tag[4][12]$_DFFE_PP__1475  (.L_HI(net1475));
 sg13g2_tiehi \cpu.dcache.r_tag[4][13]$_DFFE_PP__1476  (.L_HI(net1476));
 sg13g2_tiehi \cpu.dcache.r_tag[4][14]$_DFFE_PP__1477  (.L_HI(net1477));
 sg13g2_tiehi \cpu.dcache.r_tag[4][15]$_DFFE_PP__1478  (.L_HI(net1478));
 sg13g2_tiehi \cpu.dcache.r_tag[4][16]$_DFFE_PP__1479  (.L_HI(net1479));
 sg13g2_tiehi \cpu.dcache.r_tag[4][17]$_DFFE_PP__1480  (.L_HI(net1480));
 sg13g2_tiehi \cpu.dcache.r_tag[4][18]$_DFFE_PP__1481  (.L_HI(net1481));
 sg13g2_tiehi \cpu.dcache.r_tag[4][1]$_DFFE_PP__1482  (.L_HI(net1482));
 sg13g2_tiehi \cpu.dcache.r_tag[4][2]$_DFFE_PP__1483  (.L_HI(net1483));
 sg13g2_tiehi \cpu.dcache.r_tag[4][3]$_DFFE_PP__1484  (.L_HI(net1484));
 sg13g2_tiehi \cpu.dcache.r_tag[4][4]$_DFFE_PP__1485  (.L_HI(net1485));
 sg13g2_tiehi \cpu.dcache.r_tag[4][5]$_DFFE_PP__1486  (.L_HI(net1486));
 sg13g2_tiehi \cpu.dcache.r_tag[4][6]$_DFFE_PP__1487  (.L_HI(net1487));
 sg13g2_tiehi \cpu.dcache.r_tag[4][7]$_DFFE_PP__1488  (.L_HI(net1488));
 sg13g2_tiehi \cpu.dcache.r_tag[4][8]$_DFFE_PP__1489  (.L_HI(net1489));
 sg13g2_tiehi \cpu.dcache.r_tag[4][9]$_DFFE_PP__1490  (.L_HI(net1490));
 sg13g2_tiehi \cpu.dcache.r_tag[5][0]$_DFFE_PP__1491  (.L_HI(net1491));
 sg13g2_tiehi \cpu.dcache.r_tag[5][10]$_DFFE_PP__1492  (.L_HI(net1492));
 sg13g2_tiehi \cpu.dcache.r_tag[5][11]$_DFFE_PP__1493  (.L_HI(net1493));
 sg13g2_tiehi \cpu.dcache.r_tag[5][12]$_DFFE_PP__1494  (.L_HI(net1494));
 sg13g2_tiehi \cpu.dcache.r_tag[5][13]$_DFFE_PP__1495  (.L_HI(net1495));
 sg13g2_tiehi \cpu.dcache.r_tag[5][14]$_DFFE_PP__1496  (.L_HI(net1496));
 sg13g2_tiehi \cpu.dcache.r_tag[5][15]$_DFFE_PP__1497  (.L_HI(net1497));
 sg13g2_tiehi \cpu.dcache.r_tag[5][16]$_DFFE_PP__1498  (.L_HI(net1498));
 sg13g2_tiehi \cpu.dcache.r_tag[5][17]$_DFFE_PP__1499  (.L_HI(net1499));
 sg13g2_tiehi \cpu.dcache.r_tag[5][18]$_DFFE_PP__1500  (.L_HI(net1500));
 sg13g2_tiehi \cpu.dcache.r_tag[5][1]$_DFFE_PP__1501  (.L_HI(net1501));
 sg13g2_tiehi \cpu.dcache.r_tag[5][2]$_DFFE_PP__1502  (.L_HI(net1502));
 sg13g2_tiehi \cpu.dcache.r_tag[5][3]$_DFFE_PP__1503  (.L_HI(net1503));
 sg13g2_tiehi \cpu.dcache.r_tag[5][4]$_DFFE_PP__1504  (.L_HI(net1504));
 sg13g2_tiehi \cpu.dcache.r_tag[5][5]$_DFFE_PP__1505  (.L_HI(net1505));
 sg13g2_tiehi \cpu.dcache.r_tag[5][6]$_DFFE_PP__1506  (.L_HI(net1506));
 sg13g2_tiehi \cpu.dcache.r_tag[5][7]$_DFFE_PP__1507  (.L_HI(net1507));
 sg13g2_tiehi \cpu.dcache.r_tag[5][8]$_DFFE_PP__1508  (.L_HI(net1508));
 sg13g2_tiehi \cpu.dcache.r_tag[5][9]$_DFFE_PP__1509  (.L_HI(net1509));
 sg13g2_tiehi \cpu.dcache.r_tag[6][0]$_DFFE_PP__1510  (.L_HI(net1510));
 sg13g2_tiehi \cpu.dcache.r_tag[6][10]$_DFFE_PP__1511  (.L_HI(net1511));
 sg13g2_tiehi \cpu.dcache.r_tag[6][11]$_DFFE_PP__1512  (.L_HI(net1512));
 sg13g2_tiehi \cpu.dcache.r_tag[6][12]$_DFFE_PP__1513  (.L_HI(net1513));
 sg13g2_tiehi \cpu.dcache.r_tag[6][13]$_DFFE_PP__1514  (.L_HI(net1514));
 sg13g2_tiehi \cpu.dcache.r_tag[6][14]$_DFFE_PP__1515  (.L_HI(net1515));
 sg13g2_tiehi \cpu.dcache.r_tag[6][15]$_DFFE_PP__1516  (.L_HI(net1516));
 sg13g2_tiehi \cpu.dcache.r_tag[6][16]$_DFFE_PP__1517  (.L_HI(net1517));
 sg13g2_tiehi \cpu.dcache.r_tag[6][17]$_DFFE_PP__1518  (.L_HI(net1518));
 sg13g2_tiehi \cpu.dcache.r_tag[6][18]$_DFFE_PP__1519  (.L_HI(net1519));
 sg13g2_tiehi \cpu.dcache.r_tag[6][1]$_DFFE_PP__1520  (.L_HI(net1520));
 sg13g2_tiehi \cpu.dcache.r_tag[6][2]$_DFFE_PP__1521  (.L_HI(net1521));
 sg13g2_tiehi \cpu.dcache.r_tag[6][3]$_DFFE_PP__1522  (.L_HI(net1522));
 sg13g2_tiehi \cpu.dcache.r_tag[6][4]$_DFFE_PP__1523  (.L_HI(net1523));
 sg13g2_tiehi \cpu.dcache.r_tag[6][5]$_DFFE_PP__1524  (.L_HI(net1524));
 sg13g2_tiehi \cpu.dcache.r_tag[6][6]$_DFFE_PP__1525  (.L_HI(net1525));
 sg13g2_tiehi \cpu.dcache.r_tag[6][7]$_DFFE_PP__1526  (.L_HI(net1526));
 sg13g2_tiehi \cpu.dcache.r_tag[6][8]$_DFFE_PP__1527  (.L_HI(net1527));
 sg13g2_tiehi \cpu.dcache.r_tag[6][9]$_DFFE_PP__1528  (.L_HI(net1528));
 sg13g2_tiehi \cpu.dcache.r_tag[7][0]$_DFFE_PP__1529  (.L_HI(net1529));
 sg13g2_tiehi \cpu.dcache.r_tag[7][10]$_DFFE_PP__1530  (.L_HI(net1530));
 sg13g2_tiehi \cpu.dcache.r_tag[7][11]$_DFFE_PP__1531  (.L_HI(net1531));
 sg13g2_tiehi \cpu.dcache.r_tag[7][12]$_DFFE_PP__1532  (.L_HI(net1532));
 sg13g2_tiehi \cpu.dcache.r_tag[7][13]$_DFFE_PP__1533  (.L_HI(net1533));
 sg13g2_tiehi \cpu.dcache.r_tag[7][14]$_DFFE_PP__1534  (.L_HI(net1534));
 sg13g2_tiehi \cpu.dcache.r_tag[7][15]$_DFFE_PP__1535  (.L_HI(net1535));
 sg13g2_tiehi \cpu.dcache.r_tag[7][16]$_DFFE_PP__1536  (.L_HI(net1536));
 sg13g2_tiehi \cpu.dcache.r_tag[7][17]$_DFFE_PP__1537  (.L_HI(net1537));
 sg13g2_tiehi \cpu.dcache.r_tag[7][18]$_DFFE_PP__1538  (.L_HI(net1538));
 sg13g2_tiehi \cpu.dcache.r_tag[7][1]$_DFFE_PP__1539  (.L_HI(net1539));
 sg13g2_tiehi \cpu.dcache.r_tag[7][2]$_DFFE_PP__1540  (.L_HI(net1540));
 sg13g2_tiehi \cpu.dcache.r_tag[7][3]$_DFFE_PP__1541  (.L_HI(net1541));
 sg13g2_tiehi \cpu.dcache.r_tag[7][4]$_DFFE_PP__1542  (.L_HI(net1542));
 sg13g2_tiehi \cpu.dcache.r_tag[7][5]$_DFFE_PP__1543  (.L_HI(net1543));
 sg13g2_tiehi \cpu.dcache.r_tag[7][6]$_DFFE_PP__1544  (.L_HI(net1544));
 sg13g2_tiehi \cpu.dcache.r_tag[7][7]$_DFFE_PP__1545  (.L_HI(net1545));
 sg13g2_tiehi \cpu.dcache.r_tag[7][8]$_DFFE_PP__1546  (.L_HI(net1546));
 sg13g2_tiehi \cpu.dcache.r_tag[7][9]$_DFFE_PP__1547  (.L_HI(net1547));
 sg13g2_tiehi \cpu.dcache.r_valid[0]$_SDFFE_PP0P__1548  (.L_HI(net1548));
 sg13g2_tiehi \cpu.dcache.r_valid[1]$_SDFFE_PP0P__1549  (.L_HI(net1549));
 sg13g2_tiehi \cpu.dcache.r_valid[2]$_SDFFE_PP0P__1550  (.L_HI(net1550));
 sg13g2_tiehi \cpu.dcache.r_valid[3]$_SDFFE_PP0P__1551  (.L_HI(net1551));
 sg13g2_tiehi \cpu.dcache.r_valid[4]$_SDFFE_PP0P__1552  (.L_HI(net1552));
 sg13g2_tiehi \cpu.dcache.r_valid[5]$_SDFFE_PP0P__1553  (.L_HI(net1553));
 sg13g2_tiehi \cpu.dcache.r_valid[6]$_SDFFE_PP0P__1554  (.L_HI(net1554));
 sg13g2_tiehi \cpu.dcache.r_valid[7]$_SDFFE_PP0P__1555  (.L_HI(net1555));
 sg13g2_tiehi \cpu.dec.r_br$_DFFE_PP__1556  (.L_HI(net1556));
 sg13g2_tiehi \cpu.dec.r_cond[0]$_DFFE_PP__1557  (.L_HI(net1557));
 sg13g2_tiehi \cpu.dec.r_cond[1]$_DFFE_PP__1558  (.L_HI(net1558));
 sg13g2_tiehi \cpu.dec.r_cond[2]$_DFFE_PP__1559  (.L_HI(net1559));
 sg13g2_tiehi \cpu.dec.r_div$_DFFE_PP__1560  (.L_HI(net1560));
 sg13g2_tiehi \cpu.dec.r_flush_all$_DFFE_PP__1561  (.L_HI(net1561));
 sg13g2_tiehi \cpu.dec.r_flush_write$_DFFE_PP__1562  (.L_HI(net1562));
 sg13g2_tiehi \cpu.dec.r_imm[0]$_DFFE_PP__1563  (.L_HI(net1563));
 sg13g2_tiehi \cpu.dec.r_imm[10]$_DFFE_PP__1564  (.L_HI(net1564));
 sg13g2_tiehi \cpu.dec.r_imm[11]$_DFFE_PP__1565  (.L_HI(net1565));
 sg13g2_tiehi \cpu.dec.r_imm[12]$_DFFE_PP__1566  (.L_HI(net1566));
 sg13g2_tiehi \cpu.dec.r_imm[13]$_DFFE_PP__1567  (.L_HI(net1567));
 sg13g2_tiehi \cpu.dec.r_imm[14]$_DFFE_PP__1568  (.L_HI(net1568));
 sg13g2_tiehi \cpu.dec.r_imm[15]$_DFFE_PP__1569  (.L_HI(net1569));
 sg13g2_tiehi \cpu.dec.r_imm[1]$_DFFE_PP__1570  (.L_HI(net1570));
 sg13g2_tiehi \cpu.dec.r_imm[2]$_DFFE_PP__1571  (.L_HI(net1571));
 sg13g2_tiehi \cpu.dec.r_imm[3]$_DFFE_PP__1572  (.L_HI(net1572));
 sg13g2_tiehi \cpu.dec.r_imm[4]$_DFFE_PP__1573  (.L_HI(net1573));
 sg13g2_tiehi \cpu.dec.r_imm[5]$_DFFE_PP__1574  (.L_HI(net1574));
 sg13g2_tiehi \cpu.dec.r_imm[6]$_DFFE_PP__1575  (.L_HI(net1575));
 sg13g2_tiehi \cpu.dec.r_imm[7]$_DFFE_PP__1576  (.L_HI(net1576));
 sg13g2_tiehi \cpu.dec.r_imm[8]$_DFFE_PP__1577  (.L_HI(net1577));
 sg13g2_tiehi \cpu.dec.r_imm[9]$_DFFE_PP__1578  (.L_HI(net1578));
 sg13g2_tiehi \cpu.dec.r_inv_mmu$_DFFE_PP__1579  (.L_HI(net1579));
 sg13g2_tiehi \cpu.dec.r_io$_DFFE_PP__1580  (.L_HI(net1580));
 sg13g2_tiehi \cpu.dec.r_jmp$_SDFFCE_PP0P__1581  (.L_HI(net1581));
 sg13g2_tiehi \cpu.dec.r_load$_DFFE_PP__1582  (.L_HI(net1582));
 sg13g2_tiehi \cpu.dec.r_mult$_DFFE_PP__1583  (.L_HI(net1583));
 sg13g2_tiehi \cpu.dec.r_needs_rs2$_DFFE_PP__1584  (.L_HI(net1584));
 sg13g2_tiehi \cpu.dec.r_op[10]$_DFF_P__1585  (.L_HI(net1585));
 sg13g2_tiehi \cpu.dec.r_op[1]$_DFF_P__1586  (.L_HI(net1586));
 sg13g2_tiehi \cpu.dec.r_op[2]$_DFF_P__1587  (.L_HI(net1587));
 sg13g2_tiehi \cpu.dec.r_op[3]$_DFF_P__1588  (.L_HI(net1588));
 sg13g2_tiehi \cpu.dec.r_op[4]$_DFF_P__1589  (.L_HI(net1589));
 sg13g2_tiehi \cpu.dec.r_op[5]$_DFF_P__1590  (.L_HI(net1590));
 sg13g2_tiehi \cpu.dec.r_op[6]$_DFF_P__1591  (.L_HI(net1591));
 sg13g2_tiehi \cpu.dec.r_op[7]$_DFF_P__1592  (.L_HI(net1592));
 sg13g2_tiehi \cpu.dec.r_op[8]$_DFF_P__1593  (.L_HI(net1593));
 sg13g2_tiehi \cpu.dec.r_op[9]$_DFF_P__1594  (.L_HI(net1594));
 sg13g2_tiehi \cpu.dec.r_rd[0]$_DFFE_PP__1595  (.L_HI(net1595));
 sg13g2_tiehi \cpu.dec.r_rd[1]$_DFFE_PP__1596  (.L_HI(net1596));
 sg13g2_tiehi \cpu.dec.r_rd[2]$_DFFE_PP__1597  (.L_HI(net1597));
 sg13g2_tiehi \cpu.dec.r_rd[3]$_DFFE_PP__1598  (.L_HI(net1598));
 sg13g2_tiehi \cpu.dec.r_ready$_DFF_P__1599  (.L_HI(net1599));
 sg13g2_tiehi \cpu.dec.r_rs1[0]$_DFFE_PP__1600  (.L_HI(net1600));
 sg13g2_tiehi \cpu.dec.r_rs1[1]$_DFFE_PP__1601  (.L_HI(net1601));
 sg13g2_tiehi \cpu.dec.r_rs1[2]$_DFFE_PP__1602  (.L_HI(net1602));
 sg13g2_tiehi \cpu.dec.r_rs1[3]$_DFFE_PP__1603  (.L_HI(net1603));
 sg13g2_tiehi \cpu.dec.r_rs2[0]$_DFFE_PP__1604  (.L_HI(net1604));
 sg13g2_tiehi \cpu.dec.r_rs2[1]$_DFFE_PP__1605  (.L_HI(net1605));
 sg13g2_tiehi \cpu.dec.r_rs2[2]$_DFFE_PP__1606  (.L_HI(net1606));
 sg13g2_tiehi \cpu.dec.r_rs2[3]$_DFFE_PP__1607  (.L_HI(net1607));
 sg13g2_tiehi \cpu.dec.r_rs2_pc$_DFFE_PP__1608  (.L_HI(net1608));
 sg13g2_tiehi \cpu.dec.r_set_cc$_SDFFCE_PP0P__1609  (.L_HI(net1609));
 sg13g2_tiehi \cpu.dec.r_store$_DFFE_PP__1610  (.L_HI(net1610));
 sg13g2_tiehi \cpu.dec.r_swapsp$_DFFE_PP__1611  (.L_HI(net1611));
 sg13g2_tiehi \cpu.dec.r_sys_call$_DFFE_PP__1612  (.L_HI(net1612));
 sg13g2_tiehi \cpu.dec.r_trap$_DFFE_PP__1613  (.L_HI(net1613));
 sg13g2_tiehi \cpu.ex.genblk3.r_mmu_d_proxy$_SDFFE_PP0P__1614  (.L_HI(net1614));
 sg13g2_tiehi \cpu.ex.genblk3.r_mmu_enable$_SDFFE_PN0P__1615  (.L_HI(net1615));
 sg13g2_tiehi \cpu.ex.genblk3.r_prev_supmode$_SDFFE_PN1P__1616  (.L_HI(net1616));
 sg13g2_tiehi \cpu.ex.genblk3.r_supmode$_DFF_P__1617  (.L_HI(net1617));
 sg13g2_tiehi \cpu.ex.genblk3.r_user_io$_SDFFE_PN0P__1618  (.L_HI(net1618));
 sg13g2_tiehi \cpu.ex.r_10[0]$_DFFE_PP__1619  (.L_HI(net1619));
 sg13g2_tiehi \cpu.ex.r_10[10]$_DFFE_PP__1620  (.L_HI(net1620));
 sg13g2_tiehi \cpu.ex.r_10[11]$_DFFE_PP__1621  (.L_HI(net1621));
 sg13g2_tiehi \cpu.ex.r_10[12]$_DFFE_PP__1622  (.L_HI(net1622));
 sg13g2_tiehi \cpu.ex.r_10[13]$_DFFE_PP__1623  (.L_HI(net1623));
 sg13g2_tiehi \cpu.ex.r_10[14]$_DFFE_PP__1624  (.L_HI(net1624));
 sg13g2_tiehi \cpu.ex.r_10[15]$_DFFE_PP__1625  (.L_HI(net1625));
 sg13g2_tiehi \cpu.ex.r_10[1]$_DFFE_PP__1626  (.L_HI(net1626));
 sg13g2_tiehi \cpu.ex.r_10[2]$_DFFE_PP__1627  (.L_HI(net1627));
 sg13g2_tiehi \cpu.ex.r_10[3]$_DFFE_PP__1628  (.L_HI(net1628));
 sg13g2_tiehi \cpu.ex.r_10[4]$_DFFE_PP__1629  (.L_HI(net1629));
 sg13g2_tiehi \cpu.ex.r_10[5]$_DFFE_PP__1630  (.L_HI(net1630));
 sg13g2_tiehi \cpu.ex.r_10[6]$_DFFE_PP__1631  (.L_HI(net1631));
 sg13g2_tiehi \cpu.ex.r_10[7]$_DFFE_PP__1632  (.L_HI(net1632));
 sg13g2_tiehi \cpu.ex.r_10[8]$_DFFE_PP__1633  (.L_HI(net1633));
 sg13g2_tiehi \cpu.ex.r_10[9]$_DFFE_PP__1634  (.L_HI(net1634));
 sg13g2_tiehi \cpu.ex.r_11[0]$_DFFE_PP__1635  (.L_HI(net1635));
 sg13g2_tiehi \cpu.ex.r_11[10]$_DFFE_PP__1636  (.L_HI(net1636));
 sg13g2_tiehi \cpu.ex.r_11[11]$_DFFE_PP__1637  (.L_HI(net1637));
 sg13g2_tiehi \cpu.ex.r_11[12]$_DFFE_PP__1638  (.L_HI(net1638));
 sg13g2_tiehi \cpu.ex.r_11[13]$_DFFE_PP__1639  (.L_HI(net1639));
 sg13g2_tiehi \cpu.ex.r_11[14]$_DFFE_PP__1640  (.L_HI(net1640));
 sg13g2_tiehi \cpu.ex.r_11[15]$_DFFE_PP__1641  (.L_HI(net1641));
 sg13g2_tiehi \cpu.ex.r_11[1]$_DFFE_PP__1642  (.L_HI(net1642));
 sg13g2_tiehi \cpu.ex.r_11[2]$_DFFE_PP__1643  (.L_HI(net1643));
 sg13g2_tiehi \cpu.ex.r_11[3]$_DFFE_PP__1644  (.L_HI(net1644));
 sg13g2_tiehi \cpu.ex.r_11[4]$_DFFE_PP__1645  (.L_HI(net1645));
 sg13g2_tiehi \cpu.ex.r_11[5]$_DFFE_PP__1646  (.L_HI(net1646));
 sg13g2_tiehi \cpu.ex.r_11[6]$_DFFE_PP__1647  (.L_HI(net1647));
 sg13g2_tiehi \cpu.ex.r_11[7]$_DFFE_PP__1648  (.L_HI(net1648));
 sg13g2_tiehi \cpu.ex.r_11[8]$_DFFE_PP__1649  (.L_HI(net1649));
 sg13g2_tiehi \cpu.ex.r_11[9]$_DFFE_PP__1650  (.L_HI(net1650));
 sg13g2_tiehi \cpu.ex.r_12[0]$_DFFE_PP__1651  (.L_HI(net1651));
 sg13g2_tiehi \cpu.ex.r_12[10]$_DFFE_PP__1652  (.L_HI(net1652));
 sg13g2_tiehi \cpu.ex.r_12[11]$_DFFE_PP__1653  (.L_HI(net1653));
 sg13g2_tiehi \cpu.ex.r_12[12]$_DFFE_PP__1654  (.L_HI(net1654));
 sg13g2_tiehi \cpu.ex.r_12[13]$_DFFE_PP__1655  (.L_HI(net1655));
 sg13g2_tiehi \cpu.ex.r_12[14]$_DFFE_PP__1656  (.L_HI(net1656));
 sg13g2_tiehi \cpu.ex.r_12[15]$_DFFE_PP__1657  (.L_HI(net1657));
 sg13g2_tiehi \cpu.ex.r_12[1]$_DFFE_PP__1658  (.L_HI(net1658));
 sg13g2_tiehi \cpu.ex.r_12[2]$_DFFE_PP__1659  (.L_HI(net1659));
 sg13g2_tiehi \cpu.ex.r_12[3]$_DFFE_PP__1660  (.L_HI(net1660));
 sg13g2_tiehi \cpu.ex.r_12[4]$_DFFE_PP__1661  (.L_HI(net1661));
 sg13g2_tiehi \cpu.ex.r_12[5]$_DFFE_PP__1662  (.L_HI(net1662));
 sg13g2_tiehi \cpu.ex.r_12[6]$_DFFE_PP__1663  (.L_HI(net1663));
 sg13g2_tiehi \cpu.ex.r_12[7]$_DFFE_PP__1664  (.L_HI(net1664));
 sg13g2_tiehi \cpu.ex.r_12[8]$_DFFE_PP__1665  (.L_HI(net1665));
 sg13g2_tiehi \cpu.ex.r_12[9]$_DFFE_PP__1666  (.L_HI(net1666));
 sg13g2_tiehi \cpu.ex.r_13[0]$_DFFE_PP__1667  (.L_HI(net1667));
 sg13g2_tiehi \cpu.ex.r_13[10]$_DFFE_PP__1668  (.L_HI(net1668));
 sg13g2_tiehi \cpu.ex.r_13[11]$_DFFE_PP__1669  (.L_HI(net1669));
 sg13g2_tiehi \cpu.ex.r_13[12]$_DFFE_PP__1670  (.L_HI(net1670));
 sg13g2_tiehi \cpu.ex.r_13[13]$_DFFE_PP__1671  (.L_HI(net1671));
 sg13g2_tiehi \cpu.ex.r_13[14]$_DFFE_PP__1672  (.L_HI(net1672));
 sg13g2_tiehi \cpu.ex.r_13[15]$_DFFE_PP__1673  (.L_HI(net1673));
 sg13g2_tiehi \cpu.ex.r_13[1]$_DFFE_PP__1674  (.L_HI(net1674));
 sg13g2_tiehi \cpu.ex.r_13[2]$_DFFE_PP__1675  (.L_HI(net1675));
 sg13g2_tiehi \cpu.ex.r_13[3]$_DFFE_PP__1676  (.L_HI(net1676));
 sg13g2_tiehi \cpu.ex.r_13[4]$_DFFE_PP__1677  (.L_HI(net1677));
 sg13g2_tiehi \cpu.ex.r_13[5]$_DFFE_PP__1678  (.L_HI(net1678));
 sg13g2_tiehi \cpu.ex.r_13[6]$_DFFE_PP__1679  (.L_HI(net1679));
 sg13g2_tiehi \cpu.ex.r_13[7]$_DFFE_PP__1680  (.L_HI(net1680));
 sg13g2_tiehi \cpu.ex.r_13[8]$_DFFE_PP__1681  (.L_HI(net1681));
 sg13g2_tiehi \cpu.ex.r_13[9]$_DFFE_PP__1682  (.L_HI(net1682));
 sg13g2_tiehi \cpu.ex.r_14[0]$_DFFE_PP__1683  (.L_HI(net1683));
 sg13g2_tiehi \cpu.ex.r_14[10]$_DFFE_PP__1684  (.L_HI(net1684));
 sg13g2_tiehi \cpu.ex.r_14[11]$_DFFE_PP__1685  (.L_HI(net1685));
 sg13g2_tiehi \cpu.ex.r_14[12]$_DFFE_PP__1686  (.L_HI(net1686));
 sg13g2_tiehi \cpu.ex.r_14[13]$_DFFE_PP__1687  (.L_HI(net1687));
 sg13g2_tiehi \cpu.ex.r_14[14]$_DFFE_PP__1688  (.L_HI(net1688));
 sg13g2_tiehi \cpu.ex.r_14[15]$_DFFE_PP__1689  (.L_HI(net1689));
 sg13g2_tiehi \cpu.ex.r_14[1]$_DFFE_PP__1690  (.L_HI(net1690));
 sg13g2_tiehi \cpu.ex.r_14[2]$_DFFE_PP__1691  (.L_HI(net1691));
 sg13g2_tiehi \cpu.ex.r_14[3]$_DFFE_PP__1692  (.L_HI(net1692));
 sg13g2_tiehi \cpu.ex.r_14[4]$_DFFE_PP__1693  (.L_HI(net1693));
 sg13g2_tiehi \cpu.ex.r_14[5]$_DFFE_PP__1694  (.L_HI(net1694));
 sg13g2_tiehi \cpu.ex.r_14[6]$_DFFE_PP__1695  (.L_HI(net1695));
 sg13g2_tiehi \cpu.ex.r_14[7]$_DFFE_PP__1696  (.L_HI(net1696));
 sg13g2_tiehi \cpu.ex.r_14[8]$_DFFE_PP__1697  (.L_HI(net1697));
 sg13g2_tiehi \cpu.ex.r_14[9]$_DFFE_PP__1698  (.L_HI(net1698));
 sg13g2_tiehi \cpu.ex.r_15[0]$_DFFE_PP__1699  (.L_HI(net1699));
 sg13g2_tiehi \cpu.ex.r_15[10]$_DFFE_PP__1700  (.L_HI(net1700));
 sg13g2_tiehi \cpu.ex.r_15[11]$_DFFE_PP__1701  (.L_HI(net1701));
 sg13g2_tiehi \cpu.ex.r_15[12]$_DFFE_PP__1702  (.L_HI(net1702));
 sg13g2_tiehi \cpu.ex.r_15[13]$_DFFE_PP__1703  (.L_HI(net1703));
 sg13g2_tiehi \cpu.ex.r_15[14]$_DFFE_PP__1704  (.L_HI(net1704));
 sg13g2_tiehi \cpu.ex.r_15[15]$_DFFE_PP__1705  (.L_HI(net1705));
 sg13g2_tiehi \cpu.ex.r_15[1]$_DFFE_PP__1706  (.L_HI(net1706));
 sg13g2_tiehi \cpu.ex.r_15[2]$_DFFE_PP__1707  (.L_HI(net1707));
 sg13g2_tiehi \cpu.ex.r_15[3]$_DFFE_PP__1708  (.L_HI(net1708));
 sg13g2_tiehi \cpu.ex.r_15[4]$_DFFE_PP__1709  (.L_HI(net1709));
 sg13g2_tiehi \cpu.ex.r_15[5]$_DFFE_PP__1710  (.L_HI(net1710));
 sg13g2_tiehi \cpu.ex.r_15[6]$_DFFE_PP__1711  (.L_HI(net1711));
 sg13g2_tiehi \cpu.ex.r_15[7]$_DFFE_PP__1712  (.L_HI(net1712));
 sg13g2_tiehi \cpu.ex.r_15[8]$_DFFE_PP__1713  (.L_HI(net1713));
 sg13g2_tiehi \cpu.ex.r_15[9]$_DFFE_PP__1714  (.L_HI(net1714));
 sg13g2_tiehi \cpu.ex.r_8[0]$_DFFE_PP__1715  (.L_HI(net1715));
 sg13g2_tiehi \cpu.ex.r_8[10]$_DFFE_PP__1716  (.L_HI(net1716));
 sg13g2_tiehi \cpu.ex.r_8[11]$_DFFE_PP__1717  (.L_HI(net1717));
 sg13g2_tiehi \cpu.ex.r_8[12]$_DFFE_PP__1718  (.L_HI(net1718));
 sg13g2_tiehi \cpu.ex.r_8[13]$_DFFE_PP__1719  (.L_HI(net1719));
 sg13g2_tiehi \cpu.ex.r_8[14]$_DFFE_PP__1720  (.L_HI(net1720));
 sg13g2_tiehi \cpu.ex.r_8[15]$_DFFE_PP__1721  (.L_HI(net1721));
 sg13g2_tiehi \cpu.ex.r_8[1]$_DFFE_PP__1722  (.L_HI(net1722));
 sg13g2_tiehi \cpu.ex.r_8[2]$_DFFE_PP__1723  (.L_HI(net1723));
 sg13g2_tiehi \cpu.ex.r_8[3]$_DFFE_PP__1724  (.L_HI(net1724));
 sg13g2_tiehi \cpu.ex.r_8[4]$_DFFE_PP__1725  (.L_HI(net1725));
 sg13g2_tiehi \cpu.ex.r_8[5]$_DFFE_PP__1726  (.L_HI(net1726));
 sg13g2_tiehi \cpu.ex.r_8[6]$_DFFE_PP__1727  (.L_HI(net1727));
 sg13g2_tiehi \cpu.ex.r_8[7]$_DFFE_PP__1728  (.L_HI(net1728));
 sg13g2_tiehi \cpu.ex.r_8[8]$_DFFE_PP__1729  (.L_HI(net1729));
 sg13g2_tiehi \cpu.ex.r_8[9]$_DFFE_PP__1730  (.L_HI(net1730));
 sg13g2_tiehi \cpu.ex.r_9[0]$_DFFE_PP__1731  (.L_HI(net1731));
 sg13g2_tiehi \cpu.ex.r_9[10]$_DFFE_PP__1732  (.L_HI(net1732));
 sg13g2_tiehi \cpu.ex.r_9[11]$_DFFE_PP__1733  (.L_HI(net1733));
 sg13g2_tiehi \cpu.ex.r_9[12]$_DFFE_PP__1734  (.L_HI(net1734));
 sg13g2_tiehi \cpu.ex.r_9[13]$_DFFE_PP__1735  (.L_HI(net1735));
 sg13g2_tiehi \cpu.ex.r_9[14]$_DFFE_PP__1736  (.L_HI(net1736));
 sg13g2_tiehi \cpu.ex.r_9[15]$_DFFE_PP__1737  (.L_HI(net1737));
 sg13g2_tiehi \cpu.ex.r_9[1]$_DFFE_PP__1738  (.L_HI(net1738));
 sg13g2_tiehi \cpu.ex.r_9[2]$_DFFE_PP__1739  (.L_HI(net1739));
 sg13g2_tiehi \cpu.ex.r_9[3]$_DFFE_PP__1740  (.L_HI(net1740));
 sg13g2_tiehi \cpu.ex.r_9[4]$_DFFE_PP__1741  (.L_HI(net1741));
 sg13g2_tiehi \cpu.ex.r_9[5]$_DFFE_PP__1742  (.L_HI(net1742));
 sg13g2_tiehi \cpu.ex.r_9[6]$_DFFE_PP__1743  (.L_HI(net1743));
 sg13g2_tiehi \cpu.ex.r_9[7]$_DFFE_PP__1744  (.L_HI(net1744));
 sg13g2_tiehi \cpu.ex.r_9[8]$_DFFE_PP__1745  (.L_HI(net1745));
 sg13g2_tiehi \cpu.ex.r_9[9]$_DFFE_PP__1746  (.L_HI(net1746));
 sg13g2_tiehi \cpu.ex.r_branch_stall$_DFF_P__1747  (.L_HI(net1747));
 sg13g2_tiehi \cpu.ex.r_d_flush_all$_SDFF_PP0__1748  (.L_HI(net1748));
 sg13g2_tiehi \cpu.ex.r_div_running$_DFF_P__1749  (.L_HI(net1749));
 sg13g2_tiehi \cpu.ex.r_epc[0]$_DFFE_PP__1750  (.L_HI(net1750));
 sg13g2_tiehi \cpu.ex.r_epc[10]$_DFFE_PP__1751  (.L_HI(net1751));
 sg13g2_tiehi \cpu.ex.r_epc[11]$_DFFE_PP__1752  (.L_HI(net1752));
 sg13g2_tiehi \cpu.ex.r_epc[12]$_DFFE_PP__1753  (.L_HI(net1753));
 sg13g2_tiehi \cpu.ex.r_epc[13]$_DFFE_PP__1754  (.L_HI(net1754));
 sg13g2_tiehi \cpu.ex.r_epc[14]$_DFFE_PP__1755  (.L_HI(net1755));
 sg13g2_tiehi \cpu.ex.r_epc[1]$_DFFE_PP__1756  (.L_HI(net1756));
 sg13g2_tiehi \cpu.ex.r_epc[2]$_DFFE_PP__1757  (.L_HI(net1757));
 sg13g2_tiehi \cpu.ex.r_epc[3]$_DFFE_PP__1758  (.L_HI(net1758));
 sg13g2_tiehi \cpu.ex.r_epc[4]$_DFFE_PP__1759  (.L_HI(net1759));
 sg13g2_tiehi \cpu.ex.r_epc[5]$_DFFE_PP__1760  (.L_HI(net1760));
 sg13g2_tiehi \cpu.ex.r_epc[6]$_DFFE_PP__1761  (.L_HI(net1761));
 sg13g2_tiehi \cpu.ex.r_epc[7]$_DFFE_PP__1762  (.L_HI(net1762));
 sg13g2_tiehi \cpu.ex.r_epc[8]$_DFFE_PP__1763  (.L_HI(net1763));
 sg13g2_tiehi \cpu.ex.r_epc[9]$_DFFE_PP__1764  (.L_HI(net1764));
 sg13g2_tiehi \cpu.ex.r_fetch$_SDFF_PN1__1765  (.L_HI(net1765));
 sg13g2_tiehi \cpu.ex.r_flush_write$_SDFFE_PN0P__1766  (.L_HI(net1766));
 sg13g2_tiehi \cpu.ex.r_i_flush_all$_SDFF_PP0__1767  (.L_HI(net1767));
 sg13g2_tiehi \cpu.ex.r_ie$_SDFFE_PP0P__1768  (.L_HI(net1768));
 sg13g2_tiehi \cpu.ex.r_io_access$_SDFFE_PN0P__1769  (.L_HI(net1769));
 sg13g2_tiehi \cpu.ex.r_lr[0]$_DFFE_PP__1770  (.L_HI(net1770));
 sg13g2_tiehi \cpu.ex.r_lr[10]$_DFFE_PP__1771  (.L_HI(net1771));
 sg13g2_tiehi \cpu.ex.r_lr[11]$_DFFE_PP__1772  (.L_HI(net1772));
 sg13g2_tiehi \cpu.ex.r_lr[12]$_DFFE_PP__1773  (.L_HI(net1773));
 sg13g2_tiehi \cpu.ex.r_lr[13]$_DFFE_PP__1774  (.L_HI(net1774));
 sg13g2_tiehi \cpu.ex.r_lr[14]$_DFFE_PP__1775  (.L_HI(net1775));
 sg13g2_tiehi \cpu.ex.r_lr[1]$_DFFE_PP__1776  (.L_HI(net1776));
 sg13g2_tiehi \cpu.ex.r_lr[2]$_DFFE_PP__1777  (.L_HI(net1777));
 sg13g2_tiehi \cpu.ex.r_lr[3]$_DFFE_PP__1778  (.L_HI(net1778));
 sg13g2_tiehi \cpu.ex.r_lr[4]$_DFFE_PP__1779  (.L_HI(net1779));
 sg13g2_tiehi \cpu.ex.r_lr[5]$_DFFE_PP__1780  (.L_HI(net1780));
 sg13g2_tiehi \cpu.ex.r_lr[6]$_DFFE_PP__1781  (.L_HI(net1781));
 sg13g2_tiehi \cpu.ex.r_lr[7]$_DFFE_PP__1782  (.L_HI(net1782));
 sg13g2_tiehi \cpu.ex.r_lr[8]$_DFFE_PP__1783  (.L_HI(net1783));
 sg13g2_tiehi \cpu.ex.r_lr[9]$_DFFE_PP__1784  (.L_HI(net1784));
 sg13g2_tiehi \cpu.ex.r_mult[0]$_DFF_P__1785  (.L_HI(net1785));
 sg13g2_tiehi \cpu.ex.r_mult[10]$_DFF_P__1786  (.L_HI(net1786));
 sg13g2_tiehi \cpu.ex.r_mult[11]$_DFF_P__1787  (.L_HI(net1787));
 sg13g2_tiehi \cpu.ex.r_mult[12]$_DFF_P__1788  (.L_HI(net1788));
 sg13g2_tiehi \cpu.ex.r_mult[13]$_DFF_P__1789  (.L_HI(net1789));
 sg13g2_tiehi \cpu.ex.r_mult[14]$_DFF_P__1790  (.L_HI(net1790));
 sg13g2_tiehi \cpu.ex.r_mult[15]$_DFF_P__1791  (.L_HI(net1791));
 sg13g2_tiehi \cpu.ex.r_mult[16]$_DFFE_PP__1792  (.L_HI(net1792));
 sg13g2_tiehi \cpu.ex.r_mult[17]$_DFFE_PP__1793  (.L_HI(net1793));
 sg13g2_tiehi \cpu.ex.r_mult[18]$_DFFE_PP__1794  (.L_HI(net1794));
 sg13g2_tiehi \cpu.ex.r_mult[19]$_DFFE_PP__1795  (.L_HI(net1795));
 sg13g2_tiehi \cpu.ex.r_mult[1]$_DFF_P__1796  (.L_HI(net1796));
 sg13g2_tiehi \cpu.ex.r_mult[20]$_DFFE_PP__1797  (.L_HI(net1797));
 sg13g2_tiehi \cpu.ex.r_mult[21]$_DFFE_PP__1798  (.L_HI(net1798));
 sg13g2_tiehi \cpu.ex.r_mult[22]$_DFFE_PP__1799  (.L_HI(net1799));
 sg13g2_tiehi \cpu.ex.r_mult[23]$_DFFE_PP__1800  (.L_HI(net1800));
 sg13g2_tiehi \cpu.ex.r_mult[24]$_DFFE_PP__1801  (.L_HI(net1801));
 sg13g2_tiehi \cpu.ex.r_mult[25]$_DFFE_PP__1802  (.L_HI(net1802));
 sg13g2_tiehi \cpu.ex.r_mult[26]$_DFFE_PP__1803  (.L_HI(net1803));
 sg13g2_tiehi \cpu.ex.r_mult[27]$_DFFE_PP__1804  (.L_HI(net1804));
 sg13g2_tiehi \cpu.ex.r_mult[28]$_DFFE_PP__1805  (.L_HI(net1805));
 sg13g2_tiehi \cpu.ex.r_mult[29]$_DFFE_PP__1806  (.L_HI(net1806));
 sg13g2_tiehi \cpu.ex.r_mult[2]$_DFF_P__1807  (.L_HI(net1807));
 sg13g2_tiehi \cpu.ex.r_mult[30]$_DFFE_PP__1808  (.L_HI(net1808));
 sg13g2_tiehi \cpu.ex.r_mult[31]$_DFFE_PP__1809  (.L_HI(net1809));
 sg13g2_tiehi \cpu.ex.r_mult[3]$_DFF_P__1810  (.L_HI(net1810));
 sg13g2_tiehi \cpu.ex.r_mult[4]$_DFF_P__1811  (.L_HI(net1811));
 sg13g2_tiehi \cpu.ex.r_mult[5]$_DFF_P__1812  (.L_HI(net1812));
 sg13g2_tiehi \cpu.ex.r_mult[6]$_DFF_P__1813  (.L_HI(net1813));
 sg13g2_tiehi \cpu.ex.r_mult[7]$_DFF_P__1814  (.L_HI(net1814));
 sg13g2_tiehi \cpu.ex.r_mult[8]$_DFF_P__1815  (.L_HI(net1815));
 sg13g2_tiehi \cpu.ex.r_mult[9]$_DFF_P__1816  (.L_HI(net1816));
 sg13g2_tiehi \cpu.ex.r_mult_off[0]$_DFF_P__1817  (.L_HI(net1817));
 sg13g2_tiehi \cpu.ex.r_mult_off[1]$_DFF_P__1818  (.L_HI(net1818));
 sg13g2_tiehi \cpu.ex.r_mult_off[2]$_DFF_P__1819  (.L_HI(net1819));
 sg13g2_tiehi \cpu.ex.r_mult_off[3]$_DFF_P__1820  (.L_HI(net1820));
 sg13g2_tiehi \cpu.ex.r_mult_running$_DFF_P__1821  (.L_HI(net1821));
 sg13g2_tiehi \cpu.ex.r_pc[0]$_DFFE_PP__1822  (.L_HI(net1822));
 sg13g2_tiehi \cpu.ex.r_pc[10]$_DFFE_PP__1823  (.L_HI(net1823));
 sg13g2_tiehi \cpu.ex.r_pc[11]$_DFFE_PP__1824  (.L_HI(net1824));
 sg13g2_tiehi \cpu.ex.r_pc[12]$_DFFE_PP__1825  (.L_HI(net1825));
 sg13g2_tiehi \cpu.ex.r_pc[13]$_DFFE_PP__1826  (.L_HI(net1826));
 sg13g2_tiehi \cpu.ex.r_pc[14]$_DFFE_PP__1827  (.L_HI(net1827));
 sg13g2_tiehi \cpu.ex.r_pc[1]$_DFFE_PP__1828  (.L_HI(net1828));
 sg13g2_tiehi \cpu.ex.r_pc[2]$_DFFE_PP__1829  (.L_HI(net1829));
 sg13g2_tiehi \cpu.ex.r_pc[3]$_DFFE_PP__1830  (.L_HI(net1830));
 sg13g2_tiehi \cpu.ex.r_pc[4]$_DFFE_PP__1831  (.L_HI(net1831));
 sg13g2_tiehi \cpu.ex.r_pc[5]$_DFFE_PP__1832  (.L_HI(net1832));
 sg13g2_tiehi \cpu.ex.r_pc[6]$_DFFE_PP__1833  (.L_HI(net1833));
 sg13g2_tiehi \cpu.ex.r_pc[7]$_DFFE_PP__1834  (.L_HI(net1834));
 sg13g2_tiehi \cpu.ex.r_pc[8]$_DFFE_PP__1835  (.L_HI(net1835));
 sg13g2_tiehi \cpu.ex.r_pc[9]$_DFFE_PP__1836  (.L_HI(net1836));
 sg13g2_tiehi \cpu.ex.r_prev_ie$_SDFFE_PN0P__1837  (.L_HI(net1837));
 sg13g2_tiehi \cpu.ex.r_read_stall$_SDFFE_PN0P__1838  (.L_HI(net1838));
 sg13g2_tiehi \cpu.ex.r_sp[0]$_DFFE_PP__1839  (.L_HI(net1839));
 sg13g2_tiehi \cpu.ex.r_sp[10]$_DFFE_PP__1840  (.L_HI(net1840));
 sg13g2_tiehi \cpu.ex.r_sp[11]$_DFFE_PP__1841  (.L_HI(net1841));
 sg13g2_tiehi \cpu.ex.r_sp[12]$_DFFE_PP__1842  (.L_HI(net1842));
 sg13g2_tiehi \cpu.ex.r_sp[13]$_DFFE_PP__1843  (.L_HI(net1843));
 sg13g2_tiehi \cpu.ex.r_sp[14]$_DFFE_PP__1844  (.L_HI(net1844));
 sg13g2_tiehi \cpu.ex.r_sp[1]$_DFFE_PP__1845  (.L_HI(net1845));
 sg13g2_tiehi \cpu.ex.r_sp[2]$_DFFE_PP__1846  (.L_HI(net1846));
 sg13g2_tiehi \cpu.ex.r_sp[3]$_DFFE_PP__1847  (.L_HI(net1847));
 sg13g2_tiehi \cpu.ex.r_sp[4]$_DFFE_PP__1848  (.L_HI(net1848));
 sg13g2_tiehi \cpu.ex.r_sp[5]$_DFFE_PP__1849  (.L_HI(net1849));
 sg13g2_tiehi \cpu.ex.r_sp[6]$_DFFE_PP__1850  (.L_HI(net1850));
 sg13g2_tiehi \cpu.ex.r_sp[7]$_DFFE_PP__1851  (.L_HI(net1851));
 sg13g2_tiehi \cpu.ex.r_sp[8]$_DFFE_PP__1852  (.L_HI(net1852));
 sg13g2_tiehi \cpu.ex.r_sp[9]$_DFFE_PP__1853  (.L_HI(net1853));
 sg13g2_tiehi \cpu.ex.r_stmp[0]$_SDFFCE_PN0P__1854  (.L_HI(net1854));
 sg13g2_tiehi \cpu.ex.r_stmp[10]$_DFFE_PP__1855  (.L_HI(net1855));
 sg13g2_tiehi \cpu.ex.r_stmp[11]$_DFFE_PP__1856  (.L_HI(net1856));
 sg13g2_tiehi \cpu.ex.r_stmp[12]$_DFFE_PP__1857  (.L_HI(net1857));
 sg13g2_tiehi \cpu.ex.r_stmp[13]$_DFFE_PP__1858  (.L_HI(net1858));
 sg13g2_tiehi \cpu.ex.r_stmp[14]$_DFFE_PP__1859  (.L_HI(net1859));
 sg13g2_tiehi \cpu.ex.r_stmp[15]$_DFFE_PP__1860  (.L_HI(net1860));
 sg13g2_tiehi \cpu.ex.r_stmp[1]$_DFFE_PP__1861  (.L_HI(net1861));
 sg13g2_tiehi \cpu.ex.r_stmp[2]$_DFFE_PP__1862  (.L_HI(net1862));
 sg13g2_tiehi \cpu.ex.r_stmp[3]$_DFFE_PP__1863  (.L_HI(net1863));
 sg13g2_tiehi \cpu.ex.r_stmp[4]$_DFFE_PP__1864  (.L_HI(net1864));
 sg13g2_tiehi \cpu.ex.r_stmp[5]$_DFFE_PP__1865  (.L_HI(net1865));
 sg13g2_tiehi \cpu.ex.r_stmp[6]$_DFFE_PP__1866  (.L_HI(net1866));
 sg13g2_tiehi \cpu.ex.r_stmp[7]$_DFFE_PP__1867  (.L_HI(net1867));
 sg13g2_tiehi \cpu.ex.r_stmp[8]$_DFFE_PP__1868  (.L_HI(net1868));
 sg13g2_tiehi \cpu.ex.r_stmp[9]$_DFFE_PP__1869  (.L_HI(net1869));
 sg13g2_tiehi \cpu.ex.r_wb[0]$_DFFE_PP__1870  (.L_HI(net1870));
 sg13g2_tiehi \cpu.ex.r_wb[10]$_DFFE_PP__1871  (.L_HI(net1871));
 sg13g2_tiehi \cpu.ex.r_wb[11]$_DFFE_PP__1872  (.L_HI(net1872));
 sg13g2_tiehi \cpu.ex.r_wb[12]$_DFFE_PP__1873  (.L_HI(net1873));
 sg13g2_tiehi \cpu.ex.r_wb[13]$_DFFE_PP__1874  (.L_HI(net1874));
 sg13g2_tiehi \cpu.ex.r_wb[14]$_DFFE_PP__1875  (.L_HI(net1875));
 sg13g2_tiehi \cpu.ex.r_wb[15]$_DFFE_PP__1876  (.L_HI(net1876));
 sg13g2_tiehi \cpu.ex.r_wb[1]$_DFFE_PP__1877  (.L_HI(net1877));
 sg13g2_tiehi \cpu.ex.r_wb[2]$_DFFE_PP__1878  (.L_HI(net1878));
 sg13g2_tiehi \cpu.ex.r_wb[3]$_DFFE_PP__1879  (.L_HI(net1879));
 sg13g2_tiehi \cpu.ex.r_wb[4]$_DFFE_PP__1880  (.L_HI(net1880));
 sg13g2_tiehi \cpu.ex.r_wb[5]$_DFFE_PP__1881  (.L_HI(net1881));
 sg13g2_tiehi \cpu.ex.r_wb[6]$_DFFE_PP__1882  (.L_HI(net1882));
 sg13g2_tiehi \cpu.ex.r_wb[7]$_DFFE_PP__1883  (.L_HI(net1883));
 sg13g2_tiehi \cpu.ex.r_wb[8]$_DFFE_PP__1884  (.L_HI(net1884));
 sg13g2_tiehi \cpu.ex.r_wb[9]$_DFFE_PP__1885  (.L_HI(net1885));
 sg13g2_tiehi \cpu.ex.r_wb_addr[0]$_SDFFCE_PN0P__1886  (.L_HI(net1886));
 sg13g2_tiehi \cpu.ex.r_wb_addr[1]$_SDFFCE_PN0P__1887  (.L_HI(net1887));
 sg13g2_tiehi \cpu.ex.r_wb_addr[2]$_SDFFCE_PP0P__1888  (.L_HI(net1888));
 sg13g2_tiehi \cpu.ex.r_wb_addr[3]$_SDFFCE_PP0P__1889  (.L_HI(net1889));
 sg13g2_tiehi \cpu.ex.r_wb_swapsp$_DFFE_PP__1890  (.L_HI(net1890));
 sg13g2_tiehi \cpu.ex.r_wb_valid$_DFF_P__1891  (.L_HI(net1891));
 sg13g2_tiehi \cpu.ex.r_wdata[0]$_DFFE_PP__1892  (.L_HI(net1892));
 sg13g2_tiehi \cpu.ex.r_wdata[10]$_DFFE_PP__1893  (.L_HI(net1893));
 sg13g2_tiehi \cpu.ex.r_wdata[11]$_DFFE_PP__1894  (.L_HI(net1894));
 sg13g2_tiehi \cpu.ex.r_wdata[12]$_DFFE_PP__1895  (.L_HI(net1895));
 sg13g2_tiehi \cpu.ex.r_wdata[13]$_DFFE_PP__1896  (.L_HI(net1896));
 sg13g2_tiehi \cpu.ex.r_wdata[14]$_DFFE_PP__1897  (.L_HI(net1897));
 sg13g2_tiehi \cpu.ex.r_wdata[15]$_DFFE_PP__1898  (.L_HI(net1898));
 sg13g2_tiehi \cpu.ex.r_wdata[1]$_DFFE_PP__1899  (.L_HI(net1899));
 sg13g2_tiehi \cpu.ex.r_wdata[2]$_DFFE_PP__1900  (.L_HI(net1900));
 sg13g2_tiehi \cpu.ex.r_wdata[3]$_DFFE_PP__1901  (.L_HI(net1901));
 sg13g2_tiehi \cpu.ex.r_wdata[4]$_DFFE_PP__1902  (.L_HI(net1902));
 sg13g2_tiehi \cpu.ex.r_wdata[5]$_DFFE_PP__1903  (.L_HI(net1903));
 sg13g2_tiehi \cpu.ex.r_wdata[6]$_DFFE_PP__1904  (.L_HI(net1904));
 sg13g2_tiehi \cpu.ex.r_wdata[7]$_DFFE_PP__1905  (.L_HI(net1905));
 sg13g2_tiehi \cpu.ex.r_wdata[8]$_DFFE_PP__1906  (.L_HI(net1906));
 sg13g2_tiehi \cpu.ex.r_wdata[9]$_DFFE_PP__1907  (.L_HI(net1907));
 sg13g2_tiehi \cpu.ex.r_wmask[0]$_SDFFE_PP0P__1908  (.L_HI(net1908));
 sg13g2_tiehi \cpu.ex.r_wmask[1]$_SDFFE_PP0P__1909  (.L_HI(net1909));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[0]$_DFFE_PP__1910  (.L_HI(net1910));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[1]$_DFFE_PP__1911  (.L_HI(net1911));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[2]$_DFFE_PP__1912  (.L_HI(net1912));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[3]$_DFFE_PP__1913  (.L_HI(net1913));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_ins$_SDFFE_PN0P__1914  (.L_HI(net1914));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_sup$_SDFFE_PN0P__1915  (.L_HI(net1915));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_type$_SDFFE_PN0P__1916  (.L_HI(net1916));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[0]$_SDFFE_PN0P__1917  (.L_HI(net1917));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[10]$_SDFFE_PN0P__1918  (.L_HI(net1918));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[11]$_SDFFE_PN0P__1919  (.L_HI(net1919));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[12]$_SDFFE_PN0P__1920  (.L_HI(net1920));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[13]$_SDFFE_PN0P__1921  (.L_HI(net1921));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[14]$_SDFFE_PN0P__1922  (.L_HI(net1922));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[15]$_SDFFE_PN0P__1923  (.L_HI(net1923));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[16]$_SDFFE_PN0P__1924  (.L_HI(net1924));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[17]$_SDFFE_PN0P__1925  (.L_HI(net1925));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[18]$_SDFFE_PN0P__1926  (.L_HI(net1926));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[19]$_SDFFE_PN0P__1927  (.L_HI(net1927));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[1]$_SDFFE_PN0P__1928  (.L_HI(net1928));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[20]$_SDFFE_PN0P__1929  (.L_HI(net1929));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[21]$_SDFFE_PN0P__1930  (.L_HI(net1930));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[22]$_SDFFE_PN0P__1931  (.L_HI(net1931));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[23]$_SDFFE_PN0P__1932  (.L_HI(net1932));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[24]$_SDFFE_PN0P__1933  (.L_HI(net1933));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[25]$_SDFFE_PN0P__1934  (.L_HI(net1934));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[26]$_SDFFE_PN0P__1935  (.L_HI(net1935));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[27]$_SDFFE_PN0P__1936  (.L_HI(net1936));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[28]$_SDFFE_PN0P__1937  (.L_HI(net1937));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[29]$_SDFFE_PN0P__1938  (.L_HI(net1938));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[2]$_SDFFE_PN0P__1939  (.L_HI(net1939));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[30]$_SDFFE_PN0P__1940  (.L_HI(net1940));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[31]$_SDFFE_PN0P__1941  (.L_HI(net1941));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[3]$_SDFFE_PN0P__1942  (.L_HI(net1942));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[4]$_SDFFE_PN0P__1943  (.L_HI(net1943));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[5]$_SDFFE_PN0P__1944  (.L_HI(net1944));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[6]$_SDFFE_PN0P__1945  (.L_HI(net1945));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[7]$_SDFFE_PN0P__1946  (.L_HI(net1946));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[8]$_SDFFE_PN0P__1947  (.L_HI(net1947));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[9]$_SDFFE_PN0P__1948  (.L_HI(net1948));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[0]$_SDFFE_PN0P__1949  (.L_HI(net1949));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[10]$_SDFFE_PN0P__1950  (.L_HI(net1950));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[11]$_SDFFE_PN0P__1951  (.L_HI(net1951));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[12]$_SDFFE_PN0P__1952  (.L_HI(net1952));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[13]$_SDFFE_PN0P__1953  (.L_HI(net1953));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[14]$_SDFFE_PN0P__1954  (.L_HI(net1954));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[15]$_SDFFE_PN0P__1955  (.L_HI(net1955));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[16]$_SDFFE_PN0P__1956  (.L_HI(net1956));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[17]$_SDFFE_PN0P__1957  (.L_HI(net1957));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[18]$_SDFFE_PN0P__1958  (.L_HI(net1958));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[19]$_SDFFE_PN0P__1959  (.L_HI(net1959));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[1]$_SDFFE_PN0P__1960  (.L_HI(net1960));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[20]$_SDFFE_PN0P__1961  (.L_HI(net1961));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[21]$_SDFFE_PN0P__1962  (.L_HI(net1962));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[22]$_SDFFE_PN0P__1963  (.L_HI(net1963));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[23]$_SDFFE_PN0P__1964  (.L_HI(net1964));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[24]$_SDFFE_PN0P__1965  (.L_HI(net1965));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[25]$_SDFFE_PN0P__1966  (.L_HI(net1966));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[26]$_SDFFE_PN0P__1967  (.L_HI(net1967));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[27]$_SDFFE_PN0P__1968  (.L_HI(net1968));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[28]$_SDFFE_PN0P__1969  (.L_HI(net1969));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[29]$_SDFFE_PN0P__1970  (.L_HI(net1970));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[2]$_SDFFE_PN0P__1971  (.L_HI(net1971));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[30]$_SDFFE_PN0P__1972  (.L_HI(net1972));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[31]$_SDFFE_PN0P__1973  (.L_HI(net1973));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[3]$_SDFFE_PN0P__1974  (.L_HI(net1974));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[4]$_SDFFE_PN0P__1975  (.L_HI(net1975));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[5]$_SDFFE_PN0P__1976  (.L_HI(net1976));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[6]$_SDFFE_PN0P__1977  (.L_HI(net1977));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[7]$_SDFFE_PN0P__1978  (.L_HI(net1978));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[8]$_SDFFE_PN0P__1979  (.L_HI(net1979));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[9]$_SDFFE_PN0P__1980  (.L_HI(net1980));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][0]$_DFFE_PP__1981  (.L_HI(net1981));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][10]$_DFFE_PP__1982  (.L_HI(net1982));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][11]$_DFFE_PP__1983  (.L_HI(net1983));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][1]$_DFFE_PP__1984  (.L_HI(net1984));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][2]$_DFFE_PP__1985  (.L_HI(net1985));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][3]$_DFFE_PP__1986  (.L_HI(net1986));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][4]$_DFFE_PP__1987  (.L_HI(net1987));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][5]$_DFFE_PP__1988  (.L_HI(net1988));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][6]$_DFFE_PP__1989  (.L_HI(net1989));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][7]$_DFFE_PP__1990  (.L_HI(net1990));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][8]$_DFFE_PP__1991  (.L_HI(net1991));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][9]$_DFFE_PP__1992  (.L_HI(net1992));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][0]$_DFFE_PP__1993  (.L_HI(net1993));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][10]$_DFFE_PP__1994  (.L_HI(net1994));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][11]$_DFFE_PP__1995  (.L_HI(net1995));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][1]$_DFFE_PP__1996  (.L_HI(net1996));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][2]$_DFFE_PP__1997  (.L_HI(net1997));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][3]$_DFFE_PP__1998  (.L_HI(net1998));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][4]$_DFFE_PP__1999  (.L_HI(net1999));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][5]$_DFFE_PP__2000  (.L_HI(net2000));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][6]$_DFFE_PP__2001  (.L_HI(net2001));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][7]$_DFFE_PP__2002  (.L_HI(net2002));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][8]$_DFFE_PP__2003  (.L_HI(net2003));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][9]$_DFFE_PP__2004  (.L_HI(net2004));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][0]$_DFFE_PP__2005  (.L_HI(net2005));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][10]$_DFFE_PP__2006  (.L_HI(net2006));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][11]$_DFFE_PP__2007  (.L_HI(net2007));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][1]$_DFFE_PP__2008  (.L_HI(net2008));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][2]$_DFFE_PP__2009  (.L_HI(net2009));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][3]$_DFFE_PP__2010  (.L_HI(net2010));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][4]$_DFFE_PP__2011  (.L_HI(net2011));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][5]$_DFFE_PP__2012  (.L_HI(net2012));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][6]$_DFFE_PP__2013  (.L_HI(net2013));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][7]$_DFFE_PP__2014  (.L_HI(net2014));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][8]$_DFFE_PP__2015  (.L_HI(net2015));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][9]$_DFFE_PP__2016  (.L_HI(net2016));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][0]$_DFFE_PP__2017  (.L_HI(net2017));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][10]$_DFFE_PP__2018  (.L_HI(net2018));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][11]$_DFFE_PP__2019  (.L_HI(net2019));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][1]$_DFFE_PP__2020  (.L_HI(net2020));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][2]$_DFFE_PP__2021  (.L_HI(net2021));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][3]$_DFFE_PP__2022  (.L_HI(net2022));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][4]$_DFFE_PP__2023  (.L_HI(net2023));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][5]$_DFFE_PP__2024  (.L_HI(net2024));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][6]$_DFFE_PP__2025  (.L_HI(net2025));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][7]$_DFFE_PP__2026  (.L_HI(net2026));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][8]$_DFFE_PP__2027  (.L_HI(net2027));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][9]$_DFFE_PP__2028  (.L_HI(net2028));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][0]$_DFFE_PP__2029  (.L_HI(net2029));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][10]$_DFFE_PP__2030  (.L_HI(net2030));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][11]$_DFFE_PP__2031  (.L_HI(net2031));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][1]$_DFFE_PP__2032  (.L_HI(net2032));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][2]$_DFFE_PP__2033  (.L_HI(net2033));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][3]$_DFFE_PP__2034  (.L_HI(net2034));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][4]$_DFFE_PP__2035  (.L_HI(net2035));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][5]$_DFFE_PP__2036  (.L_HI(net2036));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][6]$_DFFE_PP__2037  (.L_HI(net2037));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][7]$_DFFE_PP__2038  (.L_HI(net2038));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][8]$_DFFE_PP__2039  (.L_HI(net2039));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][9]$_DFFE_PP__2040  (.L_HI(net2040));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][0]$_DFFE_PP__2041  (.L_HI(net2041));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][10]$_DFFE_PP__2042  (.L_HI(net2042));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][11]$_DFFE_PP__2043  (.L_HI(net2043));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][1]$_DFFE_PP__2044  (.L_HI(net2044));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][2]$_DFFE_PP__2045  (.L_HI(net2045));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][3]$_DFFE_PP__2046  (.L_HI(net2046));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][4]$_DFFE_PP__2047  (.L_HI(net2047));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][5]$_DFFE_PP__2048  (.L_HI(net2048));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][6]$_DFFE_PP__2049  (.L_HI(net2049));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][7]$_DFFE_PP__2050  (.L_HI(net2050));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][8]$_DFFE_PP__2051  (.L_HI(net2051));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][9]$_DFFE_PP__2052  (.L_HI(net2052));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][0]$_DFFE_PP__2053  (.L_HI(net2053));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][10]$_DFFE_PP__2054  (.L_HI(net2054));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][11]$_DFFE_PP__2055  (.L_HI(net2055));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][1]$_DFFE_PP__2056  (.L_HI(net2056));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][2]$_DFFE_PP__2057  (.L_HI(net2057));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][3]$_DFFE_PP__2058  (.L_HI(net2058));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][4]$_DFFE_PP__2059  (.L_HI(net2059));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][5]$_DFFE_PP__2060  (.L_HI(net2060));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][6]$_DFFE_PP__2061  (.L_HI(net2061));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][7]$_DFFE_PP__2062  (.L_HI(net2062));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][8]$_DFFE_PP__2063  (.L_HI(net2063));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][9]$_DFFE_PP__2064  (.L_HI(net2064));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][0]$_DFFE_PP__2065  (.L_HI(net2065));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][10]$_DFFE_PP__2066  (.L_HI(net2066));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][11]$_DFFE_PP__2067  (.L_HI(net2067));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][1]$_DFFE_PP__2068  (.L_HI(net2068));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][2]$_DFFE_PP__2069  (.L_HI(net2069));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][3]$_DFFE_PP__2070  (.L_HI(net2070));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][4]$_DFFE_PP__2071  (.L_HI(net2071));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][5]$_DFFE_PP__2072  (.L_HI(net2072));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][6]$_DFFE_PP__2073  (.L_HI(net2073));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][7]$_DFFE_PP__2074  (.L_HI(net2074));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][8]$_DFFE_PP__2075  (.L_HI(net2075));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][9]$_DFFE_PP__2076  (.L_HI(net2076));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][0]$_DFFE_PP__2077  (.L_HI(net2077));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][10]$_DFFE_PP__2078  (.L_HI(net2078));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][11]$_DFFE_PP__2079  (.L_HI(net2079));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][1]$_DFFE_PP__2080  (.L_HI(net2080));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][2]$_DFFE_PP__2081  (.L_HI(net2081));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][3]$_DFFE_PP__2082  (.L_HI(net2082));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][4]$_DFFE_PP__2083  (.L_HI(net2083));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][5]$_DFFE_PP__2084  (.L_HI(net2084));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][6]$_DFFE_PP__2085  (.L_HI(net2085));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][7]$_DFFE_PP__2086  (.L_HI(net2086));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][8]$_DFFE_PP__2087  (.L_HI(net2087));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][9]$_DFFE_PP__2088  (.L_HI(net2088));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][0]$_DFFE_PP__2089  (.L_HI(net2089));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][10]$_DFFE_PP__2090  (.L_HI(net2090));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][11]$_DFFE_PP__2091  (.L_HI(net2091));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][1]$_DFFE_PP__2092  (.L_HI(net2092));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][2]$_DFFE_PP__2093  (.L_HI(net2093));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][3]$_DFFE_PP__2094  (.L_HI(net2094));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][4]$_DFFE_PP__2095  (.L_HI(net2095));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][5]$_DFFE_PP__2096  (.L_HI(net2096));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][6]$_DFFE_PP__2097  (.L_HI(net2097));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][7]$_DFFE_PP__2098  (.L_HI(net2098));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][8]$_DFFE_PP__2099  (.L_HI(net2099));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][9]$_DFFE_PP__2100  (.L_HI(net2100));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][0]$_DFFE_PP__2101  (.L_HI(net2101));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][10]$_DFFE_PP__2102  (.L_HI(net2102));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][11]$_DFFE_PP__2103  (.L_HI(net2103));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][1]$_DFFE_PP__2104  (.L_HI(net2104));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][2]$_DFFE_PP__2105  (.L_HI(net2105));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][3]$_DFFE_PP__2106  (.L_HI(net2106));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][4]$_DFFE_PP__2107  (.L_HI(net2107));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][5]$_DFFE_PP__2108  (.L_HI(net2108));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][6]$_DFFE_PP__2109  (.L_HI(net2109));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][7]$_DFFE_PP__2110  (.L_HI(net2110));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][8]$_DFFE_PP__2111  (.L_HI(net2111));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][9]$_DFFE_PP__2112  (.L_HI(net2112));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][0]$_DFFE_PP__2113  (.L_HI(net2113));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][10]$_DFFE_PP__2114  (.L_HI(net2114));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][11]$_DFFE_PP__2115  (.L_HI(net2115));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][1]$_DFFE_PP__2116  (.L_HI(net2116));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][2]$_DFFE_PP__2117  (.L_HI(net2117));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][3]$_DFFE_PP__2118  (.L_HI(net2118));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][4]$_DFFE_PP__2119  (.L_HI(net2119));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][5]$_DFFE_PP__2120  (.L_HI(net2120));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][6]$_DFFE_PP__2121  (.L_HI(net2121));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][7]$_DFFE_PP__2122  (.L_HI(net2122));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][8]$_DFFE_PP__2123  (.L_HI(net2123));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][9]$_DFFE_PP__2124  (.L_HI(net2124));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][0]$_DFFE_PP__2125  (.L_HI(net2125));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][10]$_DFFE_PP__2126  (.L_HI(net2126));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][11]$_DFFE_PP__2127  (.L_HI(net2127));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][1]$_DFFE_PP__2128  (.L_HI(net2128));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][2]$_DFFE_PP__2129  (.L_HI(net2129));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][3]$_DFFE_PP__2130  (.L_HI(net2130));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][4]$_DFFE_PP__2131  (.L_HI(net2131));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][5]$_DFFE_PP__2132  (.L_HI(net2132));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][6]$_DFFE_PP__2133  (.L_HI(net2133));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][7]$_DFFE_PP__2134  (.L_HI(net2134));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][8]$_DFFE_PP__2135  (.L_HI(net2135));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][9]$_DFFE_PP__2136  (.L_HI(net2136));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][0]$_DFFE_PP__2137  (.L_HI(net2137));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][10]$_DFFE_PP__2138  (.L_HI(net2138));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][11]$_DFFE_PP__2139  (.L_HI(net2139));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][1]$_DFFE_PP__2140  (.L_HI(net2140));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][2]$_DFFE_PP__2141  (.L_HI(net2141));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][3]$_DFFE_PP__2142  (.L_HI(net2142));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][4]$_DFFE_PP__2143  (.L_HI(net2143));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][5]$_DFFE_PP__2144  (.L_HI(net2144));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][6]$_DFFE_PP__2145  (.L_HI(net2145));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][7]$_DFFE_PP__2146  (.L_HI(net2146));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][8]$_DFFE_PP__2147  (.L_HI(net2147));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][9]$_DFFE_PP__2148  (.L_HI(net2148));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][0]$_DFFE_PP__2149  (.L_HI(net2149));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][10]$_DFFE_PP__2150  (.L_HI(net2150));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][11]$_DFFE_PP__2151  (.L_HI(net2151));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][1]$_DFFE_PP__2152  (.L_HI(net2152));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][2]$_DFFE_PP__2153  (.L_HI(net2153));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][3]$_DFFE_PP__2154  (.L_HI(net2154));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][4]$_DFFE_PP__2155  (.L_HI(net2155));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][5]$_DFFE_PP__2156  (.L_HI(net2156));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][6]$_DFFE_PP__2157  (.L_HI(net2157));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][7]$_DFFE_PP__2158  (.L_HI(net2158));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][8]$_DFFE_PP__2159  (.L_HI(net2159));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][9]$_DFFE_PP__2160  (.L_HI(net2160));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][0]$_DFFE_PP__2161  (.L_HI(net2161));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][10]$_DFFE_PP__2162  (.L_HI(net2162));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][11]$_DFFE_PP__2163  (.L_HI(net2163));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][1]$_DFFE_PP__2164  (.L_HI(net2164));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][2]$_DFFE_PP__2165  (.L_HI(net2165));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][3]$_DFFE_PP__2166  (.L_HI(net2166));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][4]$_DFFE_PP__2167  (.L_HI(net2167));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][5]$_DFFE_PP__2168  (.L_HI(net2168));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][6]$_DFFE_PP__2169  (.L_HI(net2169));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][7]$_DFFE_PP__2170  (.L_HI(net2170));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][8]$_DFFE_PP__2171  (.L_HI(net2171));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][9]$_DFFE_PP__2172  (.L_HI(net2172));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][0]$_DFFE_PP__2173  (.L_HI(net2173));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][10]$_DFFE_PP__2174  (.L_HI(net2174));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][11]$_DFFE_PP__2175  (.L_HI(net2175));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][1]$_DFFE_PP__2176  (.L_HI(net2176));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][2]$_DFFE_PP__2177  (.L_HI(net2177));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][3]$_DFFE_PP__2178  (.L_HI(net2178));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][4]$_DFFE_PP__2179  (.L_HI(net2179));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][5]$_DFFE_PP__2180  (.L_HI(net2180));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][6]$_DFFE_PP__2181  (.L_HI(net2181));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][7]$_DFFE_PP__2182  (.L_HI(net2182));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][8]$_DFFE_PP__2183  (.L_HI(net2183));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][9]$_DFFE_PP__2184  (.L_HI(net2184));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][0]$_DFFE_PP__2185  (.L_HI(net2185));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][10]$_DFFE_PP__2186  (.L_HI(net2186));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][11]$_DFFE_PP__2187  (.L_HI(net2187));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][1]$_DFFE_PP__2188  (.L_HI(net2188));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][2]$_DFFE_PP__2189  (.L_HI(net2189));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][3]$_DFFE_PP__2190  (.L_HI(net2190));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][4]$_DFFE_PP__2191  (.L_HI(net2191));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][5]$_DFFE_PP__2192  (.L_HI(net2192));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][6]$_DFFE_PP__2193  (.L_HI(net2193));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][7]$_DFFE_PP__2194  (.L_HI(net2194));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][8]$_DFFE_PP__2195  (.L_HI(net2195));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][9]$_DFFE_PP__2196  (.L_HI(net2196));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][0]$_DFFE_PP__2197  (.L_HI(net2197));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][10]$_DFFE_PP__2198  (.L_HI(net2198));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][11]$_DFFE_PP__2199  (.L_HI(net2199));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][1]$_DFFE_PP__2200  (.L_HI(net2200));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][2]$_DFFE_PP__2201  (.L_HI(net2201));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][3]$_DFFE_PP__2202  (.L_HI(net2202));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][4]$_DFFE_PP__2203  (.L_HI(net2203));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][5]$_DFFE_PP__2204  (.L_HI(net2204));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][6]$_DFFE_PP__2205  (.L_HI(net2205));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][7]$_DFFE_PP__2206  (.L_HI(net2206));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][8]$_DFFE_PP__2207  (.L_HI(net2207));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][9]$_DFFE_PP__2208  (.L_HI(net2208));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][0]$_DFFE_PP__2209  (.L_HI(net2209));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][10]$_DFFE_PP__2210  (.L_HI(net2210));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][11]$_DFFE_PP__2211  (.L_HI(net2211));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][1]$_DFFE_PP__2212  (.L_HI(net2212));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][2]$_DFFE_PP__2213  (.L_HI(net2213));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][3]$_DFFE_PP__2214  (.L_HI(net2214));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][4]$_DFFE_PP__2215  (.L_HI(net2215));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][5]$_DFFE_PP__2216  (.L_HI(net2216));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][6]$_DFFE_PP__2217  (.L_HI(net2217));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][7]$_DFFE_PP__2218  (.L_HI(net2218));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][8]$_DFFE_PP__2219  (.L_HI(net2219));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][9]$_DFFE_PP__2220  (.L_HI(net2220));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][0]$_DFFE_PP__2221  (.L_HI(net2221));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][10]$_DFFE_PP__2222  (.L_HI(net2222));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][11]$_DFFE_PP__2223  (.L_HI(net2223));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][1]$_DFFE_PP__2224  (.L_HI(net2224));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][2]$_DFFE_PP__2225  (.L_HI(net2225));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][3]$_DFFE_PP__2226  (.L_HI(net2226));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][4]$_DFFE_PP__2227  (.L_HI(net2227));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][5]$_DFFE_PP__2228  (.L_HI(net2228));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][6]$_DFFE_PP__2229  (.L_HI(net2229));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][7]$_DFFE_PP__2230  (.L_HI(net2230));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][8]$_DFFE_PP__2231  (.L_HI(net2231));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][9]$_DFFE_PP__2232  (.L_HI(net2232));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][0]$_DFFE_PP__2233  (.L_HI(net2233));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][10]$_DFFE_PP__2234  (.L_HI(net2234));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][11]$_DFFE_PP__2235  (.L_HI(net2235));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][1]$_DFFE_PP__2236  (.L_HI(net2236));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][2]$_DFFE_PP__2237  (.L_HI(net2237));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][3]$_DFFE_PP__2238  (.L_HI(net2238));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][4]$_DFFE_PP__2239  (.L_HI(net2239));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][5]$_DFFE_PP__2240  (.L_HI(net2240));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][6]$_DFFE_PP__2241  (.L_HI(net2241));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][7]$_DFFE_PP__2242  (.L_HI(net2242));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][8]$_DFFE_PP__2243  (.L_HI(net2243));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][9]$_DFFE_PP__2244  (.L_HI(net2244));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][0]$_DFFE_PP__2245  (.L_HI(net2245));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][10]$_DFFE_PP__2246  (.L_HI(net2246));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][11]$_DFFE_PP__2247  (.L_HI(net2247));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][1]$_DFFE_PP__2248  (.L_HI(net2248));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][2]$_DFFE_PP__2249  (.L_HI(net2249));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][3]$_DFFE_PP__2250  (.L_HI(net2250));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][4]$_DFFE_PP__2251  (.L_HI(net2251));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][5]$_DFFE_PP__2252  (.L_HI(net2252));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][6]$_DFFE_PP__2253  (.L_HI(net2253));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][7]$_DFFE_PP__2254  (.L_HI(net2254));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][8]$_DFFE_PP__2255  (.L_HI(net2255));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][9]$_DFFE_PP__2256  (.L_HI(net2256));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][0]$_DFFE_PP__2257  (.L_HI(net2257));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][10]$_DFFE_PP__2258  (.L_HI(net2258));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][11]$_DFFE_PP__2259  (.L_HI(net2259));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][1]$_DFFE_PP__2260  (.L_HI(net2260));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][2]$_DFFE_PP__2261  (.L_HI(net2261));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][3]$_DFFE_PP__2262  (.L_HI(net2262));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][4]$_DFFE_PP__2263  (.L_HI(net2263));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][5]$_DFFE_PP__2264  (.L_HI(net2264));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][6]$_DFFE_PP__2265  (.L_HI(net2265));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][7]$_DFFE_PP__2266  (.L_HI(net2266));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][8]$_DFFE_PP__2267  (.L_HI(net2267));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][9]$_DFFE_PP__2268  (.L_HI(net2268));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][0]$_DFFE_PP__2269  (.L_HI(net2269));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][10]$_DFFE_PP__2270  (.L_HI(net2270));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][11]$_DFFE_PP__2271  (.L_HI(net2271));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][1]$_DFFE_PP__2272  (.L_HI(net2272));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][2]$_DFFE_PP__2273  (.L_HI(net2273));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][3]$_DFFE_PP__2274  (.L_HI(net2274));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][4]$_DFFE_PP__2275  (.L_HI(net2275));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][5]$_DFFE_PP__2276  (.L_HI(net2276));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][6]$_DFFE_PP__2277  (.L_HI(net2277));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][7]$_DFFE_PP__2278  (.L_HI(net2278));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][8]$_DFFE_PP__2279  (.L_HI(net2279));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][9]$_DFFE_PP__2280  (.L_HI(net2280));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][0]$_DFFE_PP__2281  (.L_HI(net2281));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][10]$_DFFE_PP__2282  (.L_HI(net2282));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][11]$_DFFE_PP__2283  (.L_HI(net2283));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][1]$_DFFE_PP__2284  (.L_HI(net2284));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][2]$_DFFE_PP__2285  (.L_HI(net2285));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][3]$_DFFE_PP__2286  (.L_HI(net2286));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][4]$_DFFE_PP__2287  (.L_HI(net2287));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][5]$_DFFE_PP__2288  (.L_HI(net2288));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][6]$_DFFE_PP__2289  (.L_HI(net2289));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][7]$_DFFE_PP__2290  (.L_HI(net2290));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][8]$_DFFE_PP__2291  (.L_HI(net2291));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][9]$_DFFE_PP__2292  (.L_HI(net2292));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][0]$_DFFE_PP__2293  (.L_HI(net2293));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][10]$_DFFE_PP__2294  (.L_HI(net2294));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][11]$_DFFE_PP__2295  (.L_HI(net2295));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][1]$_DFFE_PP__2296  (.L_HI(net2296));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][2]$_DFFE_PP__2297  (.L_HI(net2297));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][3]$_DFFE_PP__2298  (.L_HI(net2298));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][4]$_DFFE_PP__2299  (.L_HI(net2299));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][5]$_DFFE_PP__2300  (.L_HI(net2300));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][6]$_DFFE_PP__2301  (.L_HI(net2301));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][7]$_DFFE_PP__2302  (.L_HI(net2302));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][8]$_DFFE_PP__2303  (.L_HI(net2303));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][9]$_DFFE_PP__2304  (.L_HI(net2304));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][0]$_DFFE_PP__2305  (.L_HI(net2305));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][10]$_DFFE_PP__2306  (.L_HI(net2306));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][11]$_DFFE_PP__2307  (.L_HI(net2307));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][1]$_DFFE_PP__2308  (.L_HI(net2308));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][2]$_DFFE_PP__2309  (.L_HI(net2309));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][3]$_DFFE_PP__2310  (.L_HI(net2310));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][4]$_DFFE_PP__2311  (.L_HI(net2311));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][5]$_DFFE_PP__2312  (.L_HI(net2312));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][6]$_DFFE_PP__2313  (.L_HI(net2313));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][7]$_DFFE_PP__2314  (.L_HI(net2314));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][8]$_DFFE_PP__2315  (.L_HI(net2315));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][9]$_DFFE_PP__2316  (.L_HI(net2316));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][0]$_DFFE_PP__2317  (.L_HI(net2317));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][10]$_DFFE_PP__2318  (.L_HI(net2318));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][11]$_DFFE_PP__2319  (.L_HI(net2319));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][1]$_DFFE_PP__2320  (.L_HI(net2320));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][2]$_DFFE_PP__2321  (.L_HI(net2321));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][3]$_DFFE_PP__2322  (.L_HI(net2322));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][4]$_DFFE_PP__2323  (.L_HI(net2323));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][5]$_DFFE_PP__2324  (.L_HI(net2324));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][6]$_DFFE_PP__2325  (.L_HI(net2325));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][7]$_DFFE_PP__2326  (.L_HI(net2326));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][8]$_DFFE_PP__2327  (.L_HI(net2327));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][9]$_DFFE_PP__2328  (.L_HI(net2328));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][0]$_DFFE_PP__2329  (.L_HI(net2329));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][10]$_DFFE_PP__2330  (.L_HI(net2330));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][11]$_DFFE_PP__2331  (.L_HI(net2331));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][1]$_DFFE_PP__2332  (.L_HI(net2332));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][2]$_DFFE_PP__2333  (.L_HI(net2333));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][3]$_DFFE_PP__2334  (.L_HI(net2334));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][4]$_DFFE_PP__2335  (.L_HI(net2335));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][5]$_DFFE_PP__2336  (.L_HI(net2336));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][6]$_DFFE_PP__2337  (.L_HI(net2337));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][7]$_DFFE_PP__2338  (.L_HI(net2338));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][8]$_DFFE_PP__2339  (.L_HI(net2339));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][9]$_DFFE_PP__2340  (.L_HI(net2340));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][0]$_DFFE_PP__2341  (.L_HI(net2341));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][10]$_DFFE_PP__2342  (.L_HI(net2342));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][11]$_DFFE_PP__2343  (.L_HI(net2343));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][1]$_DFFE_PP__2344  (.L_HI(net2344));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][2]$_DFFE_PP__2345  (.L_HI(net2345));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][3]$_DFFE_PP__2346  (.L_HI(net2346));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][4]$_DFFE_PP__2347  (.L_HI(net2347));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][5]$_DFFE_PP__2348  (.L_HI(net2348));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][6]$_DFFE_PP__2349  (.L_HI(net2349));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][7]$_DFFE_PP__2350  (.L_HI(net2350));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][8]$_DFFE_PP__2351  (.L_HI(net2351));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][9]$_DFFE_PP__2352  (.L_HI(net2352));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][0]$_DFFE_PP__2353  (.L_HI(net2353));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][10]$_DFFE_PP__2354  (.L_HI(net2354));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][11]$_DFFE_PP__2355  (.L_HI(net2355));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][1]$_DFFE_PP__2356  (.L_HI(net2356));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][2]$_DFFE_PP__2357  (.L_HI(net2357));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][3]$_DFFE_PP__2358  (.L_HI(net2358));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][4]$_DFFE_PP__2359  (.L_HI(net2359));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][5]$_DFFE_PP__2360  (.L_HI(net2360));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][6]$_DFFE_PP__2361  (.L_HI(net2361));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][7]$_DFFE_PP__2362  (.L_HI(net2362));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][8]$_DFFE_PP__2363  (.L_HI(net2363));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][9]$_DFFE_PP__2364  (.L_HI(net2364));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][0]$_DFFE_PP__2365  (.L_HI(net2365));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][10]$_DFFE_PP__2366  (.L_HI(net2366));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][11]$_DFFE_PP__2367  (.L_HI(net2367));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][1]$_DFFE_PP__2368  (.L_HI(net2368));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][2]$_DFFE_PP__2369  (.L_HI(net2369));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][3]$_DFFE_PP__2370  (.L_HI(net2370));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][4]$_DFFE_PP__2371  (.L_HI(net2371));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][5]$_DFFE_PP__2372  (.L_HI(net2372));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][6]$_DFFE_PP__2373  (.L_HI(net2373));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][7]$_DFFE_PP__2374  (.L_HI(net2374));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][8]$_DFFE_PP__2375  (.L_HI(net2375));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][9]$_DFFE_PP__2376  (.L_HI(net2376));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][0]$_DFFE_PP__2377  (.L_HI(net2377));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][10]$_DFFE_PP__2378  (.L_HI(net2378));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][11]$_DFFE_PP__2379  (.L_HI(net2379));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][1]$_DFFE_PP__2380  (.L_HI(net2380));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][2]$_DFFE_PP__2381  (.L_HI(net2381));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][3]$_DFFE_PP__2382  (.L_HI(net2382));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][4]$_DFFE_PP__2383  (.L_HI(net2383));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][5]$_DFFE_PP__2384  (.L_HI(net2384));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][6]$_DFFE_PP__2385  (.L_HI(net2385));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][7]$_DFFE_PP__2386  (.L_HI(net2386));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][8]$_DFFE_PP__2387  (.L_HI(net2387));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][9]$_DFFE_PP__2388  (.L_HI(net2388));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][0]$_DFFE_PP__2389  (.L_HI(net2389));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][10]$_DFFE_PP__2390  (.L_HI(net2390));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][11]$_DFFE_PP__2391  (.L_HI(net2391));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][1]$_DFFE_PP__2392  (.L_HI(net2392));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][2]$_DFFE_PP__2393  (.L_HI(net2393));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][3]$_DFFE_PP__2394  (.L_HI(net2394));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][4]$_DFFE_PP__2395  (.L_HI(net2395));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][5]$_DFFE_PP__2396  (.L_HI(net2396));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][6]$_DFFE_PP__2397  (.L_HI(net2397));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][7]$_DFFE_PP__2398  (.L_HI(net2398));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][8]$_DFFE_PP__2399  (.L_HI(net2399));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][9]$_DFFE_PP__2400  (.L_HI(net2400));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][0]$_DFFE_PP__2401  (.L_HI(net2401));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][10]$_DFFE_PP__2402  (.L_HI(net2402));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][11]$_DFFE_PP__2403  (.L_HI(net2403));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][1]$_DFFE_PP__2404  (.L_HI(net2404));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][2]$_DFFE_PP__2405  (.L_HI(net2405));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][3]$_DFFE_PP__2406  (.L_HI(net2406));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][4]$_DFFE_PP__2407  (.L_HI(net2407));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][5]$_DFFE_PP__2408  (.L_HI(net2408));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][6]$_DFFE_PP__2409  (.L_HI(net2409));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][7]$_DFFE_PP__2410  (.L_HI(net2410));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][8]$_DFFE_PP__2411  (.L_HI(net2411));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][9]$_DFFE_PP__2412  (.L_HI(net2412));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][0]$_DFFE_PP__2413  (.L_HI(net2413));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][10]$_DFFE_PP__2414  (.L_HI(net2414));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][11]$_DFFE_PP__2415  (.L_HI(net2415));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][1]$_DFFE_PP__2416  (.L_HI(net2416));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][2]$_DFFE_PP__2417  (.L_HI(net2417));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][3]$_DFFE_PP__2418  (.L_HI(net2418));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][4]$_DFFE_PP__2419  (.L_HI(net2419));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][5]$_DFFE_PP__2420  (.L_HI(net2420));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][6]$_DFFE_PP__2421  (.L_HI(net2421));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][7]$_DFFE_PP__2422  (.L_HI(net2422));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][8]$_DFFE_PP__2423  (.L_HI(net2423));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][9]$_DFFE_PP__2424  (.L_HI(net2424));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][0]$_DFFE_PP__2425  (.L_HI(net2425));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][10]$_DFFE_PP__2426  (.L_HI(net2426));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][11]$_DFFE_PP__2427  (.L_HI(net2427));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][1]$_DFFE_PP__2428  (.L_HI(net2428));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][2]$_DFFE_PP__2429  (.L_HI(net2429));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][3]$_DFFE_PP__2430  (.L_HI(net2430));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][4]$_DFFE_PP__2431  (.L_HI(net2431));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][5]$_DFFE_PP__2432  (.L_HI(net2432));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][6]$_DFFE_PP__2433  (.L_HI(net2433));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][7]$_DFFE_PP__2434  (.L_HI(net2434));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][8]$_DFFE_PP__2435  (.L_HI(net2435));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][9]$_DFFE_PP__2436  (.L_HI(net2436));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][0]$_DFFE_PP__2437  (.L_HI(net2437));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][10]$_DFFE_PP__2438  (.L_HI(net2438));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][11]$_DFFE_PP__2439  (.L_HI(net2439));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][1]$_DFFE_PP__2440  (.L_HI(net2440));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][2]$_DFFE_PP__2441  (.L_HI(net2441));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][3]$_DFFE_PP__2442  (.L_HI(net2442));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][4]$_DFFE_PP__2443  (.L_HI(net2443));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][5]$_DFFE_PP__2444  (.L_HI(net2444));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][6]$_DFFE_PP__2445  (.L_HI(net2445));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][7]$_DFFE_PP__2446  (.L_HI(net2446));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][8]$_DFFE_PP__2447  (.L_HI(net2447));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][9]$_DFFE_PP__2448  (.L_HI(net2448));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][0]$_DFFE_PP__2449  (.L_HI(net2449));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][10]$_DFFE_PP__2450  (.L_HI(net2450));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][11]$_DFFE_PP__2451  (.L_HI(net2451));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][1]$_DFFE_PP__2452  (.L_HI(net2452));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][2]$_DFFE_PP__2453  (.L_HI(net2453));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][3]$_DFFE_PP__2454  (.L_HI(net2454));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][4]$_DFFE_PP__2455  (.L_HI(net2455));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][5]$_DFFE_PP__2456  (.L_HI(net2456));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][6]$_DFFE_PP__2457  (.L_HI(net2457));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][7]$_DFFE_PP__2458  (.L_HI(net2458));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][8]$_DFFE_PP__2459  (.L_HI(net2459));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][9]$_DFFE_PP__2460  (.L_HI(net2460));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][0]$_DFFE_PP__2461  (.L_HI(net2461));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][10]$_DFFE_PP__2462  (.L_HI(net2462));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][11]$_DFFE_PP__2463  (.L_HI(net2463));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][1]$_DFFE_PP__2464  (.L_HI(net2464));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][2]$_DFFE_PP__2465  (.L_HI(net2465));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][3]$_DFFE_PP__2466  (.L_HI(net2466));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][4]$_DFFE_PP__2467  (.L_HI(net2467));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][5]$_DFFE_PP__2468  (.L_HI(net2468));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][6]$_DFFE_PP__2469  (.L_HI(net2469));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][7]$_DFFE_PP__2470  (.L_HI(net2470));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][8]$_DFFE_PP__2471  (.L_HI(net2471));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][9]$_DFFE_PP__2472  (.L_HI(net2472));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][0]$_DFFE_PP__2473  (.L_HI(net2473));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][10]$_DFFE_PP__2474  (.L_HI(net2474));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][11]$_DFFE_PP__2475  (.L_HI(net2475));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][1]$_DFFE_PP__2476  (.L_HI(net2476));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][2]$_DFFE_PP__2477  (.L_HI(net2477));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][3]$_DFFE_PP__2478  (.L_HI(net2478));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][4]$_DFFE_PP__2479  (.L_HI(net2479));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][5]$_DFFE_PP__2480  (.L_HI(net2480));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][6]$_DFFE_PP__2481  (.L_HI(net2481));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][7]$_DFFE_PP__2482  (.L_HI(net2482));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][8]$_DFFE_PP__2483  (.L_HI(net2483));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][9]$_DFFE_PP__2484  (.L_HI(net2484));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][0]$_DFFE_PP__2485  (.L_HI(net2485));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][10]$_DFFE_PP__2486  (.L_HI(net2486));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][11]$_DFFE_PP__2487  (.L_HI(net2487));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][1]$_DFFE_PP__2488  (.L_HI(net2488));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][2]$_DFFE_PP__2489  (.L_HI(net2489));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][3]$_DFFE_PP__2490  (.L_HI(net2490));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][4]$_DFFE_PP__2491  (.L_HI(net2491));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][5]$_DFFE_PP__2492  (.L_HI(net2492));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][6]$_DFFE_PP__2493  (.L_HI(net2493));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][7]$_DFFE_PP__2494  (.L_HI(net2494));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][8]$_DFFE_PP__2495  (.L_HI(net2495));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][9]$_DFFE_PP__2496  (.L_HI(net2496));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][0]$_DFFE_PP__2497  (.L_HI(net2497));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][10]$_DFFE_PP__2498  (.L_HI(net2498));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][11]$_DFFE_PP__2499  (.L_HI(net2499));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][1]$_DFFE_PP__2500  (.L_HI(net2500));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][2]$_DFFE_PP__2501  (.L_HI(net2501));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][3]$_DFFE_PP__2502  (.L_HI(net2502));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][4]$_DFFE_PP__2503  (.L_HI(net2503));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][5]$_DFFE_PP__2504  (.L_HI(net2504));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][6]$_DFFE_PP__2505  (.L_HI(net2505));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][7]$_DFFE_PP__2506  (.L_HI(net2506));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][8]$_DFFE_PP__2507  (.L_HI(net2507));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][9]$_DFFE_PP__2508  (.L_HI(net2508));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][0]$_DFFE_PP__2509  (.L_HI(net2509));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][10]$_DFFE_PP__2510  (.L_HI(net2510));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][11]$_DFFE_PP__2511  (.L_HI(net2511));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][1]$_DFFE_PP__2512  (.L_HI(net2512));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][2]$_DFFE_PP__2513  (.L_HI(net2513));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][3]$_DFFE_PP__2514  (.L_HI(net2514));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][4]$_DFFE_PP__2515  (.L_HI(net2515));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][5]$_DFFE_PP__2516  (.L_HI(net2516));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][6]$_DFFE_PP__2517  (.L_HI(net2517));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][7]$_DFFE_PP__2518  (.L_HI(net2518));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][8]$_DFFE_PP__2519  (.L_HI(net2519));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][9]$_DFFE_PP__2520  (.L_HI(net2520));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][0]$_DFFE_PP__2521  (.L_HI(net2521));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][10]$_DFFE_PP__2522  (.L_HI(net2522));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][11]$_DFFE_PP__2523  (.L_HI(net2523));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][1]$_DFFE_PP__2524  (.L_HI(net2524));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][2]$_DFFE_PP__2525  (.L_HI(net2525));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][3]$_DFFE_PP__2526  (.L_HI(net2526));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][4]$_DFFE_PP__2527  (.L_HI(net2527));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][5]$_DFFE_PP__2528  (.L_HI(net2528));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][6]$_DFFE_PP__2529  (.L_HI(net2529));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][7]$_DFFE_PP__2530  (.L_HI(net2530));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][8]$_DFFE_PP__2531  (.L_HI(net2531));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][9]$_DFFE_PP__2532  (.L_HI(net2532));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][0]$_DFFE_PP__2533  (.L_HI(net2533));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][10]$_DFFE_PP__2534  (.L_HI(net2534));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][11]$_DFFE_PP__2535  (.L_HI(net2535));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][1]$_DFFE_PP__2536  (.L_HI(net2536));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][2]$_DFFE_PP__2537  (.L_HI(net2537));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][3]$_DFFE_PP__2538  (.L_HI(net2538));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][4]$_DFFE_PP__2539  (.L_HI(net2539));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][5]$_DFFE_PP__2540  (.L_HI(net2540));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][6]$_DFFE_PP__2541  (.L_HI(net2541));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][7]$_DFFE_PP__2542  (.L_HI(net2542));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][8]$_DFFE_PP__2543  (.L_HI(net2543));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][9]$_DFFE_PP__2544  (.L_HI(net2544));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][0]$_DFFE_PP__2545  (.L_HI(net2545));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][10]$_DFFE_PP__2546  (.L_HI(net2546));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][11]$_DFFE_PP__2547  (.L_HI(net2547));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][1]$_DFFE_PP__2548  (.L_HI(net2548));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][2]$_DFFE_PP__2549  (.L_HI(net2549));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][3]$_DFFE_PP__2550  (.L_HI(net2550));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][4]$_DFFE_PP__2551  (.L_HI(net2551));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][5]$_DFFE_PP__2552  (.L_HI(net2552));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][6]$_DFFE_PP__2553  (.L_HI(net2553));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][7]$_DFFE_PP__2554  (.L_HI(net2554));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][8]$_DFFE_PP__2555  (.L_HI(net2555));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][9]$_DFFE_PP__2556  (.L_HI(net2556));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][0]$_DFFE_PP__2557  (.L_HI(net2557));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][10]$_DFFE_PP__2558  (.L_HI(net2558));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][11]$_DFFE_PP__2559  (.L_HI(net2559));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][1]$_DFFE_PP__2560  (.L_HI(net2560));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][2]$_DFFE_PP__2561  (.L_HI(net2561));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][3]$_DFFE_PP__2562  (.L_HI(net2562));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][4]$_DFFE_PP__2563  (.L_HI(net2563));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][5]$_DFFE_PP__2564  (.L_HI(net2564));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][6]$_DFFE_PP__2565  (.L_HI(net2565));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][7]$_DFFE_PP__2566  (.L_HI(net2566));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][8]$_DFFE_PP__2567  (.L_HI(net2567));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][9]$_DFFE_PP__2568  (.L_HI(net2568));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][0]$_DFFE_PP__2569  (.L_HI(net2569));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][10]$_DFFE_PP__2570  (.L_HI(net2570));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][11]$_DFFE_PP__2571  (.L_HI(net2571));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][1]$_DFFE_PP__2572  (.L_HI(net2572));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][2]$_DFFE_PP__2573  (.L_HI(net2573));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][3]$_DFFE_PP__2574  (.L_HI(net2574));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][4]$_DFFE_PP__2575  (.L_HI(net2575));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][5]$_DFFE_PP__2576  (.L_HI(net2576));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][6]$_DFFE_PP__2577  (.L_HI(net2577));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][7]$_DFFE_PP__2578  (.L_HI(net2578));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][8]$_DFFE_PP__2579  (.L_HI(net2579));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][9]$_DFFE_PP__2580  (.L_HI(net2580));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][0]$_DFFE_PP__2581  (.L_HI(net2581));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][10]$_DFFE_PP__2582  (.L_HI(net2582));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][11]$_DFFE_PP__2583  (.L_HI(net2583));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][1]$_DFFE_PP__2584  (.L_HI(net2584));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][2]$_DFFE_PP__2585  (.L_HI(net2585));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][3]$_DFFE_PP__2586  (.L_HI(net2586));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][4]$_DFFE_PP__2587  (.L_HI(net2587));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][5]$_DFFE_PP__2588  (.L_HI(net2588));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][6]$_DFFE_PP__2589  (.L_HI(net2589));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][7]$_DFFE_PP__2590  (.L_HI(net2590));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][8]$_DFFE_PP__2591  (.L_HI(net2591));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][9]$_DFFE_PP__2592  (.L_HI(net2592));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][0]$_DFFE_PP__2593  (.L_HI(net2593));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][10]$_DFFE_PP__2594  (.L_HI(net2594));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][11]$_DFFE_PP__2595  (.L_HI(net2595));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][1]$_DFFE_PP__2596  (.L_HI(net2596));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][2]$_DFFE_PP__2597  (.L_HI(net2597));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][3]$_DFFE_PP__2598  (.L_HI(net2598));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][4]$_DFFE_PP__2599  (.L_HI(net2599));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][5]$_DFFE_PP__2600  (.L_HI(net2600));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][6]$_DFFE_PP__2601  (.L_HI(net2601));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][7]$_DFFE_PP__2602  (.L_HI(net2602));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][8]$_DFFE_PP__2603  (.L_HI(net2603));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][9]$_DFFE_PP__2604  (.L_HI(net2604));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][0]$_DFFE_PP__2605  (.L_HI(net2605));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][10]$_DFFE_PP__2606  (.L_HI(net2606));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][11]$_DFFE_PP__2607  (.L_HI(net2607));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][1]$_DFFE_PP__2608  (.L_HI(net2608));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][2]$_DFFE_PP__2609  (.L_HI(net2609));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][3]$_DFFE_PP__2610  (.L_HI(net2610));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][4]$_DFFE_PP__2611  (.L_HI(net2611));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][5]$_DFFE_PP__2612  (.L_HI(net2612));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][6]$_DFFE_PP__2613  (.L_HI(net2613));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][7]$_DFFE_PP__2614  (.L_HI(net2614));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][8]$_DFFE_PP__2615  (.L_HI(net2615));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][9]$_DFFE_PP__2616  (.L_HI(net2616));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][0]$_DFFE_PP__2617  (.L_HI(net2617));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][10]$_DFFE_PP__2618  (.L_HI(net2618));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][11]$_DFFE_PP__2619  (.L_HI(net2619));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][1]$_DFFE_PP__2620  (.L_HI(net2620));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][2]$_DFFE_PP__2621  (.L_HI(net2621));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][3]$_DFFE_PP__2622  (.L_HI(net2622));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][4]$_DFFE_PP__2623  (.L_HI(net2623));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][5]$_DFFE_PP__2624  (.L_HI(net2624));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][6]$_DFFE_PP__2625  (.L_HI(net2625));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][7]$_DFFE_PP__2626  (.L_HI(net2626));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][8]$_DFFE_PP__2627  (.L_HI(net2627));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][9]$_DFFE_PP__2628  (.L_HI(net2628));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][0]$_DFFE_PP__2629  (.L_HI(net2629));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][10]$_DFFE_PP__2630  (.L_HI(net2630));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][11]$_DFFE_PP__2631  (.L_HI(net2631));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][1]$_DFFE_PP__2632  (.L_HI(net2632));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][2]$_DFFE_PP__2633  (.L_HI(net2633));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][3]$_DFFE_PP__2634  (.L_HI(net2634));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][4]$_DFFE_PP__2635  (.L_HI(net2635));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][5]$_DFFE_PP__2636  (.L_HI(net2636));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][6]$_DFFE_PP__2637  (.L_HI(net2637));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][7]$_DFFE_PP__2638  (.L_HI(net2638));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][8]$_DFFE_PP__2639  (.L_HI(net2639));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][9]$_DFFE_PP__2640  (.L_HI(net2640));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][0]$_DFFE_PP__2641  (.L_HI(net2641));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][10]$_DFFE_PP__2642  (.L_HI(net2642));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][11]$_DFFE_PP__2643  (.L_HI(net2643));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][1]$_DFFE_PP__2644  (.L_HI(net2644));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][2]$_DFFE_PP__2645  (.L_HI(net2645));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][3]$_DFFE_PP__2646  (.L_HI(net2646));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][4]$_DFFE_PP__2647  (.L_HI(net2647));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][5]$_DFFE_PP__2648  (.L_HI(net2648));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][6]$_DFFE_PP__2649  (.L_HI(net2649));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][7]$_DFFE_PP__2650  (.L_HI(net2650));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][8]$_DFFE_PP__2651  (.L_HI(net2651));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][9]$_DFFE_PP__2652  (.L_HI(net2652));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][0]$_DFFE_PP__2653  (.L_HI(net2653));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][10]$_DFFE_PP__2654  (.L_HI(net2654));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][11]$_DFFE_PP__2655  (.L_HI(net2655));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][1]$_DFFE_PP__2656  (.L_HI(net2656));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][2]$_DFFE_PP__2657  (.L_HI(net2657));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][3]$_DFFE_PP__2658  (.L_HI(net2658));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][4]$_DFFE_PP__2659  (.L_HI(net2659));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][5]$_DFFE_PP__2660  (.L_HI(net2660));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][6]$_DFFE_PP__2661  (.L_HI(net2661));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][7]$_DFFE_PP__2662  (.L_HI(net2662));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][8]$_DFFE_PP__2663  (.L_HI(net2663));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][9]$_DFFE_PP__2664  (.L_HI(net2664));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][0]$_DFFE_PP__2665  (.L_HI(net2665));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][10]$_DFFE_PP__2666  (.L_HI(net2666));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][11]$_DFFE_PP__2667  (.L_HI(net2667));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][1]$_DFFE_PP__2668  (.L_HI(net2668));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][2]$_DFFE_PP__2669  (.L_HI(net2669));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][3]$_DFFE_PP__2670  (.L_HI(net2670));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][4]$_DFFE_PP__2671  (.L_HI(net2671));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][5]$_DFFE_PP__2672  (.L_HI(net2672));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][6]$_DFFE_PP__2673  (.L_HI(net2673));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][7]$_DFFE_PP__2674  (.L_HI(net2674));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][8]$_DFFE_PP__2675  (.L_HI(net2675));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][9]$_DFFE_PP__2676  (.L_HI(net2676));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][0]$_DFFE_PP__2677  (.L_HI(net2677));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][10]$_DFFE_PP__2678  (.L_HI(net2678));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][11]$_DFFE_PP__2679  (.L_HI(net2679));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][1]$_DFFE_PP__2680  (.L_HI(net2680));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][2]$_DFFE_PP__2681  (.L_HI(net2681));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][3]$_DFFE_PP__2682  (.L_HI(net2682));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][4]$_DFFE_PP__2683  (.L_HI(net2683));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][5]$_DFFE_PP__2684  (.L_HI(net2684));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][6]$_DFFE_PP__2685  (.L_HI(net2685));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][7]$_DFFE_PP__2686  (.L_HI(net2686));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][8]$_DFFE_PP__2687  (.L_HI(net2687));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][9]$_DFFE_PP__2688  (.L_HI(net2688));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][0]$_DFFE_PP__2689  (.L_HI(net2689));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][10]$_DFFE_PP__2690  (.L_HI(net2690));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][11]$_DFFE_PP__2691  (.L_HI(net2691));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][1]$_DFFE_PP__2692  (.L_HI(net2692));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][2]$_DFFE_PP__2693  (.L_HI(net2693));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][3]$_DFFE_PP__2694  (.L_HI(net2694));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][4]$_DFFE_PP__2695  (.L_HI(net2695));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][5]$_DFFE_PP__2696  (.L_HI(net2696));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][6]$_DFFE_PP__2697  (.L_HI(net2697));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][7]$_DFFE_PP__2698  (.L_HI(net2698));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][8]$_DFFE_PP__2699  (.L_HI(net2699));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][9]$_DFFE_PP__2700  (.L_HI(net2700));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][0]$_DFFE_PP__2701  (.L_HI(net2701));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][10]$_DFFE_PP__2702  (.L_HI(net2702));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][11]$_DFFE_PP__2703  (.L_HI(net2703));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][1]$_DFFE_PP__2704  (.L_HI(net2704));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][2]$_DFFE_PP__2705  (.L_HI(net2705));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][3]$_DFFE_PP__2706  (.L_HI(net2706));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][4]$_DFFE_PP__2707  (.L_HI(net2707));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][5]$_DFFE_PP__2708  (.L_HI(net2708));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][6]$_DFFE_PP__2709  (.L_HI(net2709));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][7]$_DFFE_PP__2710  (.L_HI(net2710));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][8]$_DFFE_PP__2711  (.L_HI(net2711));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][9]$_DFFE_PP__2712  (.L_HI(net2712));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][0]$_DFFE_PP__2713  (.L_HI(net2713));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][10]$_DFFE_PP__2714  (.L_HI(net2714));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][11]$_DFFE_PP__2715  (.L_HI(net2715));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][1]$_DFFE_PP__2716  (.L_HI(net2716));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][2]$_DFFE_PP__2717  (.L_HI(net2717));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][3]$_DFFE_PP__2718  (.L_HI(net2718));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][4]$_DFFE_PP__2719  (.L_HI(net2719));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][5]$_DFFE_PP__2720  (.L_HI(net2720));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][6]$_DFFE_PP__2721  (.L_HI(net2721));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][7]$_DFFE_PP__2722  (.L_HI(net2722));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][8]$_DFFE_PP__2723  (.L_HI(net2723));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][9]$_DFFE_PP__2724  (.L_HI(net2724));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][0]$_DFFE_PP__2725  (.L_HI(net2725));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][10]$_DFFE_PP__2726  (.L_HI(net2726));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][11]$_DFFE_PP__2727  (.L_HI(net2727));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][1]$_DFFE_PP__2728  (.L_HI(net2728));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][2]$_DFFE_PP__2729  (.L_HI(net2729));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][3]$_DFFE_PP__2730  (.L_HI(net2730));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][4]$_DFFE_PP__2731  (.L_HI(net2731));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][5]$_DFFE_PP__2732  (.L_HI(net2732));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][6]$_DFFE_PP__2733  (.L_HI(net2733));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][7]$_DFFE_PP__2734  (.L_HI(net2734));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][8]$_DFFE_PP__2735  (.L_HI(net2735));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][9]$_DFFE_PP__2736  (.L_HI(net2736));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][0]$_DFFE_PP__2737  (.L_HI(net2737));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][10]$_DFFE_PP__2738  (.L_HI(net2738));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][11]$_DFFE_PP__2739  (.L_HI(net2739));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][1]$_DFFE_PP__2740  (.L_HI(net2740));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][2]$_DFFE_PP__2741  (.L_HI(net2741));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][3]$_DFFE_PP__2742  (.L_HI(net2742));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][4]$_DFFE_PP__2743  (.L_HI(net2743));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][5]$_DFFE_PP__2744  (.L_HI(net2744));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][6]$_DFFE_PP__2745  (.L_HI(net2745));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][7]$_DFFE_PP__2746  (.L_HI(net2746));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][8]$_DFFE_PP__2747  (.L_HI(net2747));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][9]$_DFFE_PP__2748  (.L_HI(net2748));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[0]$_DFFE_PP__2749  (.L_HI(net2749));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[10]$_DFFE_PP__2750  (.L_HI(net2750));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[11]$_DFFE_PP__2751  (.L_HI(net2751));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[12]$_DFFE_PP__2752  (.L_HI(net2752));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[13]$_DFFE_PP__2753  (.L_HI(net2753));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[14]$_DFFE_PP__2754  (.L_HI(net2754));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[15]$_DFFE_PP__2755  (.L_HI(net2755));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[16]$_DFFE_PP__2756  (.L_HI(net2756));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[17]$_DFFE_PP__2757  (.L_HI(net2757));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[18]$_DFFE_PP__2758  (.L_HI(net2758));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[19]$_DFFE_PP__2759  (.L_HI(net2759));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[1]$_DFFE_PP__2760  (.L_HI(net2760));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[20]$_DFFE_PP__2761  (.L_HI(net2761));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[21]$_DFFE_PP__2762  (.L_HI(net2762));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[22]$_DFFE_PP__2763  (.L_HI(net2763));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[23]$_DFFE_PP__2764  (.L_HI(net2764));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[24]$_DFFE_PP__2765  (.L_HI(net2765));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[25]$_DFFE_PP__2766  (.L_HI(net2766));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[26]$_DFFE_PP__2767  (.L_HI(net2767));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[27]$_DFFE_PP__2768  (.L_HI(net2768));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[28]$_DFFE_PP__2769  (.L_HI(net2769));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[29]$_DFFE_PP__2770  (.L_HI(net2770));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[2]$_DFFE_PP__2771  (.L_HI(net2771));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[30]$_DFFE_PP__2772  (.L_HI(net2772));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[31]$_DFFE_PP__2773  (.L_HI(net2773));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[3]$_DFFE_PP__2774  (.L_HI(net2774));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[4]$_DFFE_PP__2775  (.L_HI(net2775));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[5]$_DFFE_PP__2776  (.L_HI(net2776));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[6]$_DFFE_PP__2777  (.L_HI(net2777));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[7]$_DFFE_PP__2778  (.L_HI(net2778));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[8]$_DFFE_PP__2779  (.L_HI(net2779));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[9]$_DFFE_PP__2780  (.L_HI(net2780));
 sg13g2_tiehi \cpu.gpio.r_enable_in[0]$_SDFFE_PN0P__2781  (.L_HI(net2781));
 sg13g2_tiehi \cpu.gpio.r_enable_in[1]$_SDFFE_PN0P__2782  (.L_HI(net2782));
 sg13g2_tiehi \cpu.gpio.r_enable_in[2]$_SDFFE_PN0P__2783  (.L_HI(net2783));
 sg13g2_tiehi \cpu.gpio.r_enable_in[3]$_SDFFE_PN0P__2784  (.L_HI(net2784));
 sg13g2_tiehi \cpu.gpio.r_enable_in[4]$_SDFFE_PN0P__2785  (.L_HI(net2785));
 sg13g2_tiehi \cpu.gpio.r_enable_in[5]$_SDFFE_PN0P__2786  (.L_HI(net2786));
 sg13g2_tiehi \cpu.gpio.r_enable_in[6]$_SDFFE_PN0P__2787  (.L_HI(net2787));
 sg13g2_tiehi \cpu.gpio.r_enable_in[7]$_SDFFE_PN0P__2788  (.L_HI(net2788));
 sg13g2_tiehi \cpu.gpio.r_enable_io[0]$_SDFFE_PN0P__2789  (.L_HI(net2789));
 sg13g2_tiehi \cpu.gpio.r_enable_io[1]$_SDFFE_PN0P__2790  (.L_HI(net2790));
 sg13g2_tiehi \cpu.gpio.r_enable_io[2]$_SDFFE_PN0P__2791  (.L_HI(net2791));
 sg13g2_tiehi \cpu.gpio.r_enable_io[3]$_SDFFE_PN0P__2792  (.L_HI(net2792));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[0]$_SDFFE_PN0P__2793  (.L_HI(net2793));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[1]$_SDFFE_PN0P__2794  (.L_HI(net2794));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[2]$_SDFFE_PN0P__2795  (.L_HI(net2795));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[3]$_SDFFE_PN0P__2796  (.L_HI(net2796));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[0]$_DFFE_PP__2797  (.L_HI(net2797));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[1]$_DFFE_PP__2798  (.L_HI(net2798));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[2]$_DFFE_PP__2799  (.L_HI(net2799));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[3]$_DFFE_PP__2800  (.L_HI(net2800));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[0]$_DFFE_PP__2801  (.L_HI(net2801));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[1]$_DFFE_PP__2802  (.L_HI(net2802));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[2]$_DFFE_PP__2803  (.L_HI(net2803));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[3]$_DFFE_PP__2804  (.L_HI(net2804));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[4]$_DFFE_PP__2805  (.L_HI(net2805));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][0]$_DFFE_PP__2806  (.L_HI(net2806));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][1]$_DFFE_PP__2807  (.L_HI(net2807));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][2]$_DFFE_PP__2808  (.L_HI(net2808));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][3]$_DFFE_PP__2809  (.L_HI(net2809));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][0]$_DFFE_PP__2810  (.L_HI(net2810));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][1]$_DFFE_PP__2811  (.L_HI(net2811));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][2]$_DFFE_PP__2812  (.L_HI(net2812));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][3]$_DFFE_PP__2813  (.L_HI(net2813));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][0]$_DFFE_PP__2814  (.L_HI(net2814));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][1]$_DFFE_PP__2815  (.L_HI(net2815));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][2]$_DFFE_PP__2816  (.L_HI(net2816));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][3]$_DFFE_PP__2817  (.L_HI(net2817));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][0]$_DFFE_PP__2818  (.L_HI(net2818));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][1]$_DFFE_PP__2819  (.L_HI(net2819));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][2]$_DFFE_PP__2820  (.L_HI(net2820));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][3]$_DFFE_PP__2821  (.L_HI(net2821));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][0]$_DFFE_PP__2822  (.L_HI(net2822));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][1]$_DFFE_PP__2823  (.L_HI(net2823));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][2]$_DFFE_PP__2824  (.L_HI(net2824));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][3]$_DFFE_PP__2825  (.L_HI(net2825));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][0]$_DFFE_PP__2826  (.L_HI(net2826));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][1]$_DFFE_PP__2827  (.L_HI(net2827));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][2]$_DFFE_PP__2828  (.L_HI(net2828));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][3]$_DFFE_PP__2829  (.L_HI(net2829));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][0]$_DFFE_PP__2830  (.L_HI(net2830));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][1]$_DFFE_PP__2831  (.L_HI(net2831));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][2]$_DFFE_PP__2832  (.L_HI(net2832));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][3]$_DFFE_PP__2833  (.L_HI(net2833));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][0]$_DFFE_PP__2834  (.L_HI(net2834));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][1]$_DFFE_PP__2835  (.L_HI(net2835));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][2]$_DFFE_PP__2836  (.L_HI(net2836));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][3]$_DFFE_PP__2837  (.L_HI(net2837));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][0]$_DFFE_PP__2838  (.L_HI(net2838));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][1]$_DFFE_PP__2839  (.L_HI(net2839));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][2]$_DFFE_PP__2840  (.L_HI(net2840));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][3]$_DFFE_PP__2841  (.L_HI(net2841));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][0]$_SDFFE_PN1P__2842  (.L_HI(net2842));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][1]$_SDFFE_PN0P__2843  (.L_HI(net2843));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][2]$_SDFFE_PN0P__2844  (.L_HI(net2844));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][3]$_SDFFE_PN0P__2845  (.L_HI(net2845));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][0]$_DFFE_PP__2846  (.L_HI(net2846));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][1]$_DFFE_PP__2847  (.L_HI(net2847));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][2]$_DFFE_PP__2848  (.L_HI(net2848));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][3]$_DFFE_PP__2849  (.L_HI(net2849));
 sg13g2_tiehi \cpu.gpio.r_uart_rx_src[0]$_SDFFE_PN0P__2850  (.L_HI(net2850));
 sg13g2_tiehi \cpu.gpio.r_uart_rx_src[1]$_SDFFE_PN0P__2851  (.L_HI(net2851));
 sg13g2_tiehi \cpu.gpio.r_uart_rx_src[2]$_SDFFE_PN0P__2852  (.L_HI(net2852));
 sg13g2_tiehi \cpu.icache.r_data[0][0]$_DFFE_PP__2853  (.L_HI(net2853));
 sg13g2_tiehi \cpu.icache.r_data[0][10]$_DFFE_PP__2854  (.L_HI(net2854));
 sg13g2_tiehi \cpu.icache.r_data[0][11]$_DFFE_PP__2855  (.L_HI(net2855));
 sg13g2_tiehi \cpu.icache.r_data[0][12]$_DFFE_PP__2856  (.L_HI(net2856));
 sg13g2_tiehi \cpu.icache.r_data[0][13]$_DFFE_PP__2857  (.L_HI(net2857));
 sg13g2_tiehi \cpu.icache.r_data[0][14]$_DFFE_PP__2858  (.L_HI(net2858));
 sg13g2_tiehi \cpu.icache.r_data[0][15]$_DFFE_PP__2859  (.L_HI(net2859));
 sg13g2_tiehi \cpu.icache.r_data[0][16]$_DFFE_PP__2860  (.L_HI(net2860));
 sg13g2_tiehi \cpu.icache.r_data[0][17]$_DFFE_PP__2861  (.L_HI(net2861));
 sg13g2_tiehi \cpu.icache.r_data[0][18]$_DFFE_PP__2862  (.L_HI(net2862));
 sg13g2_tiehi \cpu.icache.r_data[0][19]$_DFFE_PP__2863  (.L_HI(net2863));
 sg13g2_tiehi \cpu.icache.r_data[0][1]$_DFFE_PP__2864  (.L_HI(net2864));
 sg13g2_tiehi \cpu.icache.r_data[0][20]$_DFFE_PP__2865  (.L_HI(net2865));
 sg13g2_tiehi \cpu.icache.r_data[0][21]$_DFFE_PP__2866  (.L_HI(net2866));
 sg13g2_tiehi \cpu.icache.r_data[0][22]$_DFFE_PP__2867  (.L_HI(net2867));
 sg13g2_tiehi \cpu.icache.r_data[0][23]$_DFFE_PP__2868  (.L_HI(net2868));
 sg13g2_tiehi \cpu.icache.r_data[0][24]$_DFFE_PP__2869  (.L_HI(net2869));
 sg13g2_tiehi \cpu.icache.r_data[0][25]$_DFFE_PP__2870  (.L_HI(net2870));
 sg13g2_tiehi \cpu.icache.r_data[0][26]$_DFFE_PP__2871  (.L_HI(net2871));
 sg13g2_tiehi \cpu.icache.r_data[0][27]$_DFFE_PP__2872  (.L_HI(net2872));
 sg13g2_tiehi \cpu.icache.r_data[0][28]$_DFFE_PP__2873  (.L_HI(net2873));
 sg13g2_tiehi \cpu.icache.r_data[0][29]$_DFFE_PP__2874  (.L_HI(net2874));
 sg13g2_tiehi \cpu.icache.r_data[0][2]$_DFFE_PP__2875  (.L_HI(net2875));
 sg13g2_tiehi \cpu.icache.r_data[0][30]$_DFFE_PP__2876  (.L_HI(net2876));
 sg13g2_tiehi \cpu.icache.r_data[0][31]$_DFFE_PP__2877  (.L_HI(net2877));
 sg13g2_tiehi \cpu.icache.r_data[0][3]$_DFFE_PP__2878  (.L_HI(net2878));
 sg13g2_tiehi \cpu.icache.r_data[0][4]$_DFFE_PP__2879  (.L_HI(net2879));
 sg13g2_tiehi \cpu.icache.r_data[0][5]$_DFFE_PP__2880  (.L_HI(net2880));
 sg13g2_tiehi \cpu.icache.r_data[0][6]$_DFFE_PP__2881  (.L_HI(net2881));
 sg13g2_tiehi \cpu.icache.r_data[0][7]$_DFFE_PP__2882  (.L_HI(net2882));
 sg13g2_tiehi \cpu.icache.r_data[0][8]$_DFFE_PP__2883  (.L_HI(net2883));
 sg13g2_tiehi \cpu.icache.r_data[0][9]$_DFFE_PP__2884  (.L_HI(net2884));
 sg13g2_tiehi \cpu.icache.r_data[1][0]$_DFFE_PP__2885  (.L_HI(net2885));
 sg13g2_tiehi \cpu.icache.r_data[1][10]$_DFFE_PP__2886  (.L_HI(net2886));
 sg13g2_tiehi \cpu.icache.r_data[1][11]$_DFFE_PP__2887  (.L_HI(net2887));
 sg13g2_tiehi \cpu.icache.r_data[1][12]$_DFFE_PP__2888  (.L_HI(net2888));
 sg13g2_tiehi \cpu.icache.r_data[1][13]$_DFFE_PP__2889  (.L_HI(net2889));
 sg13g2_tiehi \cpu.icache.r_data[1][14]$_DFFE_PP__2890  (.L_HI(net2890));
 sg13g2_tiehi \cpu.icache.r_data[1][15]$_DFFE_PP__2891  (.L_HI(net2891));
 sg13g2_tiehi \cpu.icache.r_data[1][16]$_DFFE_PP__2892  (.L_HI(net2892));
 sg13g2_tiehi \cpu.icache.r_data[1][17]$_DFFE_PP__2893  (.L_HI(net2893));
 sg13g2_tiehi \cpu.icache.r_data[1][18]$_DFFE_PP__2894  (.L_HI(net2894));
 sg13g2_tiehi \cpu.icache.r_data[1][19]$_DFFE_PP__2895  (.L_HI(net2895));
 sg13g2_tiehi \cpu.icache.r_data[1][1]$_DFFE_PP__2896  (.L_HI(net2896));
 sg13g2_tiehi \cpu.icache.r_data[1][20]$_DFFE_PP__2897  (.L_HI(net2897));
 sg13g2_tiehi \cpu.icache.r_data[1][21]$_DFFE_PP__2898  (.L_HI(net2898));
 sg13g2_tiehi \cpu.icache.r_data[1][22]$_DFFE_PP__2899  (.L_HI(net2899));
 sg13g2_tiehi \cpu.icache.r_data[1][23]$_DFFE_PP__2900  (.L_HI(net2900));
 sg13g2_tiehi \cpu.icache.r_data[1][24]$_DFFE_PP__2901  (.L_HI(net2901));
 sg13g2_tiehi \cpu.icache.r_data[1][25]$_DFFE_PP__2902  (.L_HI(net2902));
 sg13g2_tiehi \cpu.icache.r_data[1][26]$_DFFE_PP__2903  (.L_HI(net2903));
 sg13g2_tiehi \cpu.icache.r_data[1][27]$_DFFE_PP__2904  (.L_HI(net2904));
 sg13g2_tiehi \cpu.icache.r_data[1][28]$_DFFE_PP__2905  (.L_HI(net2905));
 sg13g2_tiehi \cpu.icache.r_data[1][29]$_DFFE_PP__2906  (.L_HI(net2906));
 sg13g2_tiehi \cpu.icache.r_data[1][2]$_DFFE_PP__2907  (.L_HI(net2907));
 sg13g2_tiehi \cpu.icache.r_data[1][30]$_DFFE_PP__2908  (.L_HI(net2908));
 sg13g2_tiehi \cpu.icache.r_data[1][31]$_DFFE_PP__2909  (.L_HI(net2909));
 sg13g2_tiehi \cpu.icache.r_data[1][3]$_DFFE_PP__2910  (.L_HI(net2910));
 sg13g2_tiehi \cpu.icache.r_data[1][4]$_DFFE_PP__2911  (.L_HI(net2911));
 sg13g2_tiehi \cpu.icache.r_data[1][5]$_DFFE_PP__2912  (.L_HI(net2912));
 sg13g2_tiehi \cpu.icache.r_data[1][6]$_DFFE_PP__2913  (.L_HI(net2913));
 sg13g2_tiehi \cpu.icache.r_data[1][7]$_DFFE_PP__2914  (.L_HI(net2914));
 sg13g2_tiehi \cpu.icache.r_data[1][8]$_DFFE_PP__2915  (.L_HI(net2915));
 sg13g2_tiehi \cpu.icache.r_data[1][9]$_DFFE_PP__2916  (.L_HI(net2916));
 sg13g2_tiehi \cpu.icache.r_data[2][0]$_DFFE_PP__2917  (.L_HI(net2917));
 sg13g2_tiehi \cpu.icache.r_data[2][10]$_DFFE_PP__2918  (.L_HI(net2918));
 sg13g2_tiehi \cpu.icache.r_data[2][11]$_DFFE_PP__2919  (.L_HI(net2919));
 sg13g2_tiehi \cpu.icache.r_data[2][12]$_DFFE_PP__2920  (.L_HI(net2920));
 sg13g2_tiehi \cpu.icache.r_data[2][13]$_DFFE_PP__2921  (.L_HI(net2921));
 sg13g2_tiehi \cpu.icache.r_data[2][14]$_DFFE_PP__2922  (.L_HI(net2922));
 sg13g2_tiehi \cpu.icache.r_data[2][15]$_DFFE_PP__2923  (.L_HI(net2923));
 sg13g2_tiehi \cpu.icache.r_data[2][16]$_DFFE_PP__2924  (.L_HI(net2924));
 sg13g2_tiehi \cpu.icache.r_data[2][17]$_DFFE_PP__2925  (.L_HI(net2925));
 sg13g2_tiehi \cpu.icache.r_data[2][18]$_DFFE_PP__2926  (.L_HI(net2926));
 sg13g2_tiehi \cpu.icache.r_data[2][19]$_DFFE_PP__2927  (.L_HI(net2927));
 sg13g2_tiehi \cpu.icache.r_data[2][1]$_DFFE_PP__2928  (.L_HI(net2928));
 sg13g2_tiehi \cpu.icache.r_data[2][20]$_DFFE_PP__2929  (.L_HI(net2929));
 sg13g2_tiehi \cpu.icache.r_data[2][21]$_DFFE_PP__2930  (.L_HI(net2930));
 sg13g2_tiehi \cpu.icache.r_data[2][22]$_DFFE_PP__2931  (.L_HI(net2931));
 sg13g2_tiehi \cpu.icache.r_data[2][23]$_DFFE_PP__2932  (.L_HI(net2932));
 sg13g2_tiehi \cpu.icache.r_data[2][24]$_DFFE_PP__2933  (.L_HI(net2933));
 sg13g2_tiehi \cpu.icache.r_data[2][25]$_DFFE_PP__2934  (.L_HI(net2934));
 sg13g2_tiehi \cpu.icache.r_data[2][26]$_DFFE_PP__2935  (.L_HI(net2935));
 sg13g2_tiehi \cpu.icache.r_data[2][27]$_DFFE_PP__2936  (.L_HI(net2936));
 sg13g2_tiehi \cpu.icache.r_data[2][28]$_DFFE_PP__2937  (.L_HI(net2937));
 sg13g2_tiehi \cpu.icache.r_data[2][29]$_DFFE_PP__2938  (.L_HI(net2938));
 sg13g2_tiehi \cpu.icache.r_data[2][2]$_DFFE_PP__2939  (.L_HI(net2939));
 sg13g2_tiehi \cpu.icache.r_data[2][30]$_DFFE_PP__2940  (.L_HI(net2940));
 sg13g2_tiehi \cpu.icache.r_data[2][31]$_DFFE_PP__2941  (.L_HI(net2941));
 sg13g2_tiehi \cpu.icache.r_data[2][3]$_DFFE_PP__2942  (.L_HI(net2942));
 sg13g2_tiehi \cpu.icache.r_data[2][4]$_DFFE_PP__2943  (.L_HI(net2943));
 sg13g2_tiehi \cpu.icache.r_data[2][5]$_DFFE_PP__2944  (.L_HI(net2944));
 sg13g2_tiehi \cpu.icache.r_data[2][6]$_DFFE_PP__2945  (.L_HI(net2945));
 sg13g2_tiehi \cpu.icache.r_data[2][7]$_DFFE_PP__2946  (.L_HI(net2946));
 sg13g2_tiehi \cpu.icache.r_data[2][8]$_DFFE_PP__2947  (.L_HI(net2947));
 sg13g2_tiehi \cpu.icache.r_data[2][9]$_DFFE_PP__2948  (.L_HI(net2948));
 sg13g2_tiehi \cpu.icache.r_data[3][0]$_DFFE_PP__2949  (.L_HI(net2949));
 sg13g2_tiehi \cpu.icache.r_data[3][10]$_DFFE_PP__2950  (.L_HI(net2950));
 sg13g2_tiehi \cpu.icache.r_data[3][11]$_DFFE_PP__2951  (.L_HI(net2951));
 sg13g2_tiehi \cpu.icache.r_data[3][12]$_DFFE_PP__2952  (.L_HI(net2952));
 sg13g2_tiehi \cpu.icache.r_data[3][13]$_DFFE_PP__2953  (.L_HI(net2953));
 sg13g2_tiehi \cpu.icache.r_data[3][14]$_DFFE_PP__2954  (.L_HI(net2954));
 sg13g2_tiehi \cpu.icache.r_data[3][15]$_DFFE_PP__2955  (.L_HI(net2955));
 sg13g2_tiehi \cpu.icache.r_data[3][16]$_DFFE_PP__2956  (.L_HI(net2956));
 sg13g2_tiehi \cpu.icache.r_data[3][17]$_DFFE_PP__2957  (.L_HI(net2957));
 sg13g2_tiehi \cpu.icache.r_data[3][18]$_DFFE_PP__2958  (.L_HI(net2958));
 sg13g2_tiehi \cpu.icache.r_data[3][19]$_DFFE_PP__2959  (.L_HI(net2959));
 sg13g2_tiehi \cpu.icache.r_data[3][1]$_DFFE_PP__2960  (.L_HI(net2960));
 sg13g2_tiehi \cpu.icache.r_data[3][20]$_DFFE_PP__2961  (.L_HI(net2961));
 sg13g2_tiehi \cpu.icache.r_data[3][21]$_DFFE_PP__2962  (.L_HI(net2962));
 sg13g2_tiehi \cpu.icache.r_data[3][22]$_DFFE_PP__2963  (.L_HI(net2963));
 sg13g2_tiehi \cpu.icache.r_data[3][23]$_DFFE_PP__2964  (.L_HI(net2964));
 sg13g2_tiehi \cpu.icache.r_data[3][24]$_DFFE_PP__2965  (.L_HI(net2965));
 sg13g2_tiehi \cpu.icache.r_data[3][25]$_DFFE_PP__2966  (.L_HI(net2966));
 sg13g2_tiehi \cpu.icache.r_data[3][26]$_DFFE_PP__2967  (.L_HI(net2967));
 sg13g2_tiehi \cpu.icache.r_data[3][27]$_DFFE_PP__2968  (.L_HI(net2968));
 sg13g2_tiehi \cpu.icache.r_data[3][28]$_DFFE_PP__2969  (.L_HI(net2969));
 sg13g2_tiehi \cpu.icache.r_data[3][29]$_DFFE_PP__2970  (.L_HI(net2970));
 sg13g2_tiehi \cpu.icache.r_data[3][2]$_DFFE_PP__2971  (.L_HI(net2971));
 sg13g2_tiehi \cpu.icache.r_data[3][30]$_DFFE_PP__2972  (.L_HI(net2972));
 sg13g2_tiehi \cpu.icache.r_data[3][31]$_DFFE_PP__2973  (.L_HI(net2973));
 sg13g2_tiehi \cpu.icache.r_data[3][3]$_DFFE_PP__2974  (.L_HI(net2974));
 sg13g2_tiehi \cpu.icache.r_data[3][4]$_DFFE_PP__2975  (.L_HI(net2975));
 sg13g2_tiehi \cpu.icache.r_data[3][5]$_DFFE_PP__2976  (.L_HI(net2976));
 sg13g2_tiehi \cpu.icache.r_data[3][6]$_DFFE_PP__2977  (.L_HI(net2977));
 sg13g2_tiehi \cpu.icache.r_data[3][7]$_DFFE_PP__2978  (.L_HI(net2978));
 sg13g2_tiehi \cpu.icache.r_data[3][8]$_DFFE_PP__2979  (.L_HI(net2979));
 sg13g2_tiehi \cpu.icache.r_data[3][9]$_DFFE_PP__2980  (.L_HI(net2980));
 sg13g2_tiehi \cpu.icache.r_data[4][0]$_DFFE_PP__2981  (.L_HI(net2981));
 sg13g2_tiehi \cpu.icache.r_data[4][10]$_DFFE_PP__2982  (.L_HI(net2982));
 sg13g2_tiehi \cpu.icache.r_data[4][11]$_DFFE_PP__2983  (.L_HI(net2983));
 sg13g2_tiehi \cpu.icache.r_data[4][12]$_DFFE_PP__2984  (.L_HI(net2984));
 sg13g2_tiehi \cpu.icache.r_data[4][13]$_DFFE_PP__2985  (.L_HI(net2985));
 sg13g2_tiehi \cpu.icache.r_data[4][14]$_DFFE_PP__2986  (.L_HI(net2986));
 sg13g2_tiehi \cpu.icache.r_data[4][15]$_DFFE_PP__2987  (.L_HI(net2987));
 sg13g2_tiehi \cpu.icache.r_data[4][16]$_DFFE_PP__2988  (.L_HI(net2988));
 sg13g2_tiehi \cpu.icache.r_data[4][17]$_DFFE_PP__2989  (.L_HI(net2989));
 sg13g2_tiehi \cpu.icache.r_data[4][18]$_DFFE_PP__2990  (.L_HI(net2990));
 sg13g2_tiehi \cpu.icache.r_data[4][19]$_DFFE_PP__2991  (.L_HI(net2991));
 sg13g2_tiehi \cpu.icache.r_data[4][1]$_DFFE_PP__2992  (.L_HI(net2992));
 sg13g2_tiehi \cpu.icache.r_data[4][20]$_DFFE_PP__2993  (.L_HI(net2993));
 sg13g2_tiehi \cpu.icache.r_data[4][21]$_DFFE_PP__2994  (.L_HI(net2994));
 sg13g2_tiehi \cpu.icache.r_data[4][22]$_DFFE_PP__2995  (.L_HI(net2995));
 sg13g2_tiehi \cpu.icache.r_data[4][23]$_DFFE_PP__2996  (.L_HI(net2996));
 sg13g2_tiehi \cpu.icache.r_data[4][24]$_DFFE_PP__2997  (.L_HI(net2997));
 sg13g2_tiehi \cpu.icache.r_data[4][25]$_DFFE_PP__2998  (.L_HI(net2998));
 sg13g2_tiehi \cpu.icache.r_data[4][26]$_DFFE_PP__2999  (.L_HI(net2999));
 sg13g2_tiehi \cpu.icache.r_data[4][27]$_DFFE_PP__3000  (.L_HI(net3000));
 sg13g2_tiehi \cpu.icache.r_data[4][28]$_DFFE_PP__3001  (.L_HI(net3001));
 sg13g2_tiehi \cpu.icache.r_data[4][29]$_DFFE_PP__3002  (.L_HI(net3002));
 sg13g2_tiehi \cpu.icache.r_data[4][2]$_DFFE_PP__3003  (.L_HI(net3003));
 sg13g2_tiehi \cpu.icache.r_data[4][30]$_DFFE_PP__3004  (.L_HI(net3004));
 sg13g2_tiehi \cpu.icache.r_data[4][31]$_DFFE_PP__3005  (.L_HI(net3005));
 sg13g2_tiehi \cpu.icache.r_data[4][3]$_DFFE_PP__3006  (.L_HI(net3006));
 sg13g2_tiehi \cpu.icache.r_data[4][4]$_DFFE_PP__3007  (.L_HI(net3007));
 sg13g2_tiehi \cpu.icache.r_data[4][5]$_DFFE_PP__3008  (.L_HI(net3008));
 sg13g2_tiehi \cpu.icache.r_data[4][6]$_DFFE_PP__3009  (.L_HI(net3009));
 sg13g2_tiehi \cpu.icache.r_data[4][7]$_DFFE_PP__3010  (.L_HI(net3010));
 sg13g2_tiehi \cpu.icache.r_data[4][8]$_DFFE_PP__3011  (.L_HI(net3011));
 sg13g2_tiehi \cpu.icache.r_data[4][9]$_DFFE_PP__3012  (.L_HI(net3012));
 sg13g2_tiehi \cpu.icache.r_data[5][0]$_DFFE_PP__3013  (.L_HI(net3013));
 sg13g2_tiehi \cpu.icache.r_data[5][10]$_DFFE_PP__3014  (.L_HI(net3014));
 sg13g2_tiehi \cpu.icache.r_data[5][11]$_DFFE_PP__3015  (.L_HI(net3015));
 sg13g2_tiehi \cpu.icache.r_data[5][12]$_DFFE_PP__3016  (.L_HI(net3016));
 sg13g2_tiehi \cpu.icache.r_data[5][13]$_DFFE_PP__3017  (.L_HI(net3017));
 sg13g2_tiehi \cpu.icache.r_data[5][14]$_DFFE_PP__3018  (.L_HI(net3018));
 sg13g2_tiehi \cpu.icache.r_data[5][15]$_DFFE_PP__3019  (.L_HI(net3019));
 sg13g2_tiehi \cpu.icache.r_data[5][16]$_DFFE_PP__3020  (.L_HI(net3020));
 sg13g2_tiehi \cpu.icache.r_data[5][17]$_DFFE_PP__3021  (.L_HI(net3021));
 sg13g2_tiehi \cpu.icache.r_data[5][18]$_DFFE_PP__3022  (.L_HI(net3022));
 sg13g2_tiehi \cpu.icache.r_data[5][19]$_DFFE_PP__3023  (.L_HI(net3023));
 sg13g2_tiehi \cpu.icache.r_data[5][1]$_DFFE_PP__3024  (.L_HI(net3024));
 sg13g2_tiehi \cpu.icache.r_data[5][20]$_DFFE_PP__3025  (.L_HI(net3025));
 sg13g2_tiehi \cpu.icache.r_data[5][21]$_DFFE_PP__3026  (.L_HI(net3026));
 sg13g2_tiehi \cpu.icache.r_data[5][22]$_DFFE_PP__3027  (.L_HI(net3027));
 sg13g2_tiehi \cpu.icache.r_data[5][23]$_DFFE_PP__3028  (.L_HI(net3028));
 sg13g2_tiehi \cpu.icache.r_data[5][24]$_DFFE_PP__3029  (.L_HI(net3029));
 sg13g2_tiehi \cpu.icache.r_data[5][25]$_DFFE_PP__3030  (.L_HI(net3030));
 sg13g2_tiehi \cpu.icache.r_data[5][26]$_DFFE_PP__3031  (.L_HI(net3031));
 sg13g2_tiehi \cpu.icache.r_data[5][27]$_DFFE_PP__3032  (.L_HI(net3032));
 sg13g2_tiehi \cpu.icache.r_data[5][28]$_DFFE_PP__3033  (.L_HI(net3033));
 sg13g2_tiehi \cpu.icache.r_data[5][29]$_DFFE_PP__3034  (.L_HI(net3034));
 sg13g2_tiehi \cpu.icache.r_data[5][2]$_DFFE_PP__3035  (.L_HI(net3035));
 sg13g2_tiehi \cpu.icache.r_data[5][30]$_DFFE_PP__3036  (.L_HI(net3036));
 sg13g2_tiehi \cpu.icache.r_data[5][31]$_DFFE_PP__3037  (.L_HI(net3037));
 sg13g2_tiehi \cpu.icache.r_data[5][3]$_DFFE_PP__3038  (.L_HI(net3038));
 sg13g2_tiehi \cpu.icache.r_data[5][4]$_DFFE_PP__3039  (.L_HI(net3039));
 sg13g2_tiehi \cpu.icache.r_data[5][5]$_DFFE_PP__3040  (.L_HI(net3040));
 sg13g2_tiehi \cpu.icache.r_data[5][6]$_DFFE_PP__3041  (.L_HI(net3041));
 sg13g2_tiehi \cpu.icache.r_data[5][7]$_DFFE_PP__3042  (.L_HI(net3042));
 sg13g2_tiehi \cpu.icache.r_data[5][8]$_DFFE_PP__3043  (.L_HI(net3043));
 sg13g2_tiehi \cpu.icache.r_data[5][9]$_DFFE_PP__3044  (.L_HI(net3044));
 sg13g2_tiehi \cpu.icache.r_data[6][0]$_DFFE_PP__3045  (.L_HI(net3045));
 sg13g2_tiehi \cpu.icache.r_data[6][10]$_DFFE_PP__3046  (.L_HI(net3046));
 sg13g2_tiehi \cpu.icache.r_data[6][11]$_DFFE_PP__3047  (.L_HI(net3047));
 sg13g2_tiehi \cpu.icache.r_data[6][12]$_DFFE_PP__3048  (.L_HI(net3048));
 sg13g2_tiehi \cpu.icache.r_data[6][13]$_DFFE_PP__3049  (.L_HI(net3049));
 sg13g2_tiehi \cpu.icache.r_data[6][14]$_DFFE_PP__3050  (.L_HI(net3050));
 sg13g2_tiehi \cpu.icache.r_data[6][15]$_DFFE_PP__3051  (.L_HI(net3051));
 sg13g2_tiehi \cpu.icache.r_data[6][16]$_DFFE_PP__3052  (.L_HI(net3052));
 sg13g2_tiehi \cpu.icache.r_data[6][17]$_DFFE_PP__3053  (.L_HI(net3053));
 sg13g2_tiehi \cpu.icache.r_data[6][18]$_DFFE_PP__3054  (.L_HI(net3054));
 sg13g2_tiehi \cpu.icache.r_data[6][19]$_DFFE_PP__3055  (.L_HI(net3055));
 sg13g2_tiehi \cpu.icache.r_data[6][1]$_DFFE_PP__3056  (.L_HI(net3056));
 sg13g2_tiehi \cpu.icache.r_data[6][20]$_DFFE_PP__3057  (.L_HI(net3057));
 sg13g2_tiehi \cpu.icache.r_data[6][21]$_DFFE_PP__3058  (.L_HI(net3058));
 sg13g2_tiehi \cpu.icache.r_data[6][22]$_DFFE_PP__3059  (.L_HI(net3059));
 sg13g2_tiehi \cpu.icache.r_data[6][23]$_DFFE_PP__3060  (.L_HI(net3060));
 sg13g2_tiehi \cpu.icache.r_data[6][24]$_DFFE_PP__3061  (.L_HI(net3061));
 sg13g2_tiehi \cpu.icache.r_data[6][25]$_DFFE_PP__3062  (.L_HI(net3062));
 sg13g2_tiehi \cpu.icache.r_data[6][26]$_DFFE_PP__3063  (.L_HI(net3063));
 sg13g2_tiehi \cpu.icache.r_data[6][27]$_DFFE_PP__3064  (.L_HI(net3064));
 sg13g2_tiehi \cpu.icache.r_data[6][28]$_DFFE_PP__3065  (.L_HI(net3065));
 sg13g2_tiehi \cpu.icache.r_data[6][29]$_DFFE_PP__3066  (.L_HI(net3066));
 sg13g2_tiehi \cpu.icache.r_data[6][2]$_DFFE_PP__3067  (.L_HI(net3067));
 sg13g2_tiehi \cpu.icache.r_data[6][30]$_DFFE_PP__3068  (.L_HI(net3068));
 sg13g2_tiehi \cpu.icache.r_data[6][31]$_DFFE_PP__3069  (.L_HI(net3069));
 sg13g2_tiehi \cpu.icache.r_data[6][3]$_DFFE_PP__3070  (.L_HI(net3070));
 sg13g2_tiehi \cpu.icache.r_data[6][4]$_DFFE_PP__3071  (.L_HI(net3071));
 sg13g2_tiehi \cpu.icache.r_data[6][5]$_DFFE_PP__3072  (.L_HI(net3072));
 sg13g2_tiehi \cpu.icache.r_data[6][6]$_DFFE_PP__3073  (.L_HI(net3073));
 sg13g2_tiehi \cpu.icache.r_data[6][7]$_DFFE_PP__3074  (.L_HI(net3074));
 sg13g2_tiehi \cpu.icache.r_data[6][8]$_DFFE_PP__3075  (.L_HI(net3075));
 sg13g2_tiehi \cpu.icache.r_data[6][9]$_DFFE_PP__3076  (.L_HI(net3076));
 sg13g2_tiehi \cpu.icache.r_data[7][0]$_DFFE_PP__3077  (.L_HI(net3077));
 sg13g2_tiehi \cpu.icache.r_data[7][10]$_DFFE_PP__3078  (.L_HI(net3078));
 sg13g2_tiehi \cpu.icache.r_data[7][11]$_DFFE_PP__3079  (.L_HI(net3079));
 sg13g2_tiehi \cpu.icache.r_data[7][12]$_DFFE_PP__3080  (.L_HI(net3080));
 sg13g2_tiehi \cpu.icache.r_data[7][13]$_DFFE_PP__3081  (.L_HI(net3081));
 sg13g2_tiehi \cpu.icache.r_data[7][14]$_DFFE_PP__3082  (.L_HI(net3082));
 sg13g2_tiehi \cpu.icache.r_data[7][15]$_DFFE_PP__3083  (.L_HI(net3083));
 sg13g2_tiehi \cpu.icache.r_data[7][16]$_DFFE_PP__3084  (.L_HI(net3084));
 sg13g2_tiehi \cpu.icache.r_data[7][17]$_DFFE_PP__3085  (.L_HI(net3085));
 sg13g2_tiehi \cpu.icache.r_data[7][18]$_DFFE_PP__3086  (.L_HI(net3086));
 sg13g2_tiehi \cpu.icache.r_data[7][19]$_DFFE_PP__3087  (.L_HI(net3087));
 sg13g2_tiehi \cpu.icache.r_data[7][1]$_DFFE_PP__3088  (.L_HI(net3088));
 sg13g2_tiehi \cpu.icache.r_data[7][20]$_DFFE_PP__3089  (.L_HI(net3089));
 sg13g2_tiehi \cpu.icache.r_data[7][21]$_DFFE_PP__3090  (.L_HI(net3090));
 sg13g2_tiehi \cpu.icache.r_data[7][22]$_DFFE_PP__3091  (.L_HI(net3091));
 sg13g2_tiehi \cpu.icache.r_data[7][23]$_DFFE_PP__3092  (.L_HI(net3092));
 sg13g2_tiehi \cpu.icache.r_data[7][24]$_DFFE_PP__3093  (.L_HI(net3093));
 sg13g2_tiehi \cpu.icache.r_data[7][25]$_DFFE_PP__3094  (.L_HI(net3094));
 sg13g2_tiehi \cpu.icache.r_data[7][26]$_DFFE_PP__3095  (.L_HI(net3095));
 sg13g2_tiehi \cpu.icache.r_data[7][27]$_DFFE_PP__3096  (.L_HI(net3096));
 sg13g2_tiehi \cpu.icache.r_data[7][28]$_DFFE_PP__3097  (.L_HI(net3097));
 sg13g2_tiehi \cpu.icache.r_data[7][29]$_DFFE_PP__3098  (.L_HI(net3098));
 sg13g2_tiehi \cpu.icache.r_data[7][2]$_DFFE_PP__3099  (.L_HI(net3099));
 sg13g2_tiehi \cpu.icache.r_data[7][30]$_DFFE_PP__3100  (.L_HI(net3100));
 sg13g2_tiehi \cpu.icache.r_data[7][31]$_DFFE_PP__3101  (.L_HI(net3101));
 sg13g2_tiehi \cpu.icache.r_data[7][3]$_DFFE_PP__3102  (.L_HI(net3102));
 sg13g2_tiehi \cpu.icache.r_data[7][4]$_DFFE_PP__3103  (.L_HI(net3103));
 sg13g2_tiehi \cpu.icache.r_data[7][5]$_DFFE_PP__3104  (.L_HI(net3104));
 sg13g2_tiehi \cpu.icache.r_data[7][6]$_DFFE_PP__3105  (.L_HI(net3105));
 sg13g2_tiehi \cpu.icache.r_data[7][7]$_DFFE_PP__3106  (.L_HI(net3106));
 sg13g2_tiehi \cpu.icache.r_data[7][8]$_DFFE_PP__3107  (.L_HI(net3107));
 sg13g2_tiehi \cpu.icache.r_data[7][9]$_DFFE_PP__3108  (.L_HI(net3108));
 sg13g2_tiehi \cpu.icache.r_offset[0]$_SDFF_PN0__3109  (.L_HI(net3109));
 sg13g2_tiehi \cpu.icache.r_offset[1]$_SDFF_PN0__3110  (.L_HI(net3110));
 sg13g2_tiehi \cpu.icache.r_offset[2]$_SDFF_PN0__3111  (.L_HI(net3111));
 sg13g2_tiehi \cpu.icache.r_tag[0][0]$_DFFE_PP__3112  (.L_HI(net3112));
 sg13g2_tiehi \cpu.icache.r_tag[0][10]$_DFFE_PP__3113  (.L_HI(net3113));
 sg13g2_tiehi \cpu.icache.r_tag[0][11]$_DFFE_PP__3114  (.L_HI(net3114));
 sg13g2_tiehi \cpu.icache.r_tag[0][12]$_DFFE_PP__3115  (.L_HI(net3115));
 sg13g2_tiehi \cpu.icache.r_tag[0][13]$_DFFE_PP__3116  (.L_HI(net3116));
 sg13g2_tiehi \cpu.icache.r_tag[0][14]$_DFFE_PP__3117  (.L_HI(net3117));
 sg13g2_tiehi \cpu.icache.r_tag[0][15]$_DFFE_PP__3118  (.L_HI(net3118));
 sg13g2_tiehi \cpu.icache.r_tag[0][16]$_DFFE_PP__3119  (.L_HI(net3119));
 sg13g2_tiehi \cpu.icache.r_tag[0][17]$_DFFE_PP__3120  (.L_HI(net3120));
 sg13g2_tiehi \cpu.icache.r_tag[0][18]$_DFFE_PP__3121  (.L_HI(net3121));
 sg13g2_tiehi \cpu.icache.r_tag[0][1]$_DFFE_PP__3122  (.L_HI(net3122));
 sg13g2_tiehi \cpu.icache.r_tag[0][2]$_DFFE_PP__3123  (.L_HI(net3123));
 sg13g2_tiehi \cpu.icache.r_tag[0][3]$_DFFE_PP__3124  (.L_HI(net3124));
 sg13g2_tiehi \cpu.icache.r_tag[0][4]$_DFFE_PP__3125  (.L_HI(net3125));
 sg13g2_tiehi \cpu.icache.r_tag[0][5]$_DFFE_PP__3126  (.L_HI(net3126));
 sg13g2_tiehi \cpu.icache.r_tag[0][6]$_DFFE_PP__3127  (.L_HI(net3127));
 sg13g2_tiehi \cpu.icache.r_tag[0][7]$_DFFE_PP__3128  (.L_HI(net3128));
 sg13g2_tiehi \cpu.icache.r_tag[0][8]$_DFFE_PP__3129  (.L_HI(net3129));
 sg13g2_tiehi \cpu.icache.r_tag[0][9]$_DFFE_PP__3130  (.L_HI(net3130));
 sg13g2_tiehi \cpu.icache.r_tag[1][0]$_DFFE_PP__3131  (.L_HI(net3131));
 sg13g2_tiehi \cpu.icache.r_tag[1][10]$_DFFE_PP__3132  (.L_HI(net3132));
 sg13g2_tiehi \cpu.icache.r_tag[1][11]$_DFFE_PP__3133  (.L_HI(net3133));
 sg13g2_tiehi \cpu.icache.r_tag[1][12]$_DFFE_PP__3134  (.L_HI(net3134));
 sg13g2_tiehi \cpu.icache.r_tag[1][13]$_DFFE_PP__3135  (.L_HI(net3135));
 sg13g2_tiehi \cpu.icache.r_tag[1][14]$_DFFE_PP__3136  (.L_HI(net3136));
 sg13g2_tiehi \cpu.icache.r_tag[1][15]$_DFFE_PP__3137  (.L_HI(net3137));
 sg13g2_tiehi \cpu.icache.r_tag[1][16]$_DFFE_PP__3138  (.L_HI(net3138));
 sg13g2_tiehi \cpu.icache.r_tag[1][17]$_DFFE_PP__3139  (.L_HI(net3139));
 sg13g2_tiehi \cpu.icache.r_tag[1][18]$_DFFE_PP__3140  (.L_HI(net3140));
 sg13g2_tiehi \cpu.icache.r_tag[1][1]$_DFFE_PP__3141  (.L_HI(net3141));
 sg13g2_tiehi \cpu.icache.r_tag[1][2]$_DFFE_PP__3142  (.L_HI(net3142));
 sg13g2_tiehi \cpu.icache.r_tag[1][3]$_DFFE_PP__3143  (.L_HI(net3143));
 sg13g2_tiehi \cpu.icache.r_tag[1][4]$_DFFE_PP__3144  (.L_HI(net3144));
 sg13g2_tiehi \cpu.icache.r_tag[1][5]$_DFFE_PP__3145  (.L_HI(net3145));
 sg13g2_tiehi \cpu.icache.r_tag[1][6]$_DFFE_PP__3146  (.L_HI(net3146));
 sg13g2_tiehi \cpu.icache.r_tag[1][7]$_DFFE_PP__3147  (.L_HI(net3147));
 sg13g2_tiehi \cpu.icache.r_tag[1][8]$_DFFE_PP__3148  (.L_HI(net3148));
 sg13g2_tiehi \cpu.icache.r_tag[1][9]$_DFFE_PP__3149  (.L_HI(net3149));
 sg13g2_tiehi \cpu.icache.r_tag[2][0]$_DFFE_PP__3150  (.L_HI(net3150));
 sg13g2_tiehi \cpu.icache.r_tag[2][10]$_DFFE_PP__3151  (.L_HI(net3151));
 sg13g2_tiehi \cpu.icache.r_tag[2][11]$_DFFE_PP__3152  (.L_HI(net3152));
 sg13g2_tiehi \cpu.icache.r_tag[2][12]$_DFFE_PP__3153  (.L_HI(net3153));
 sg13g2_tiehi \cpu.icache.r_tag[2][13]$_DFFE_PP__3154  (.L_HI(net3154));
 sg13g2_tiehi \cpu.icache.r_tag[2][14]$_DFFE_PP__3155  (.L_HI(net3155));
 sg13g2_tiehi \cpu.icache.r_tag[2][15]$_DFFE_PP__3156  (.L_HI(net3156));
 sg13g2_tiehi \cpu.icache.r_tag[2][16]$_DFFE_PP__3157  (.L_HI(net3157));
 sg13g2_tiehi \cpu.icache.r_tag[2][17]$_DFFE_PP__3158  (.L_HI(net3158));
 sg13g2_tiehi \cpu.icache.r_tag[2][18]$_DFFE_PP__3159  (.L_HI(net3159));
 sg13g2_tiehi \cpu.icache.r_tag[2][1]$_DFFE_PP__3160  (.L_HI(net3160));
 sg13g2_tiehi \cpu.icache.r_tag[2][2]$_DFFE_PP__3161  (.L_HI(net3161));
 sg13g2_tiehi \cpu.icache.r_tag[2][3]$_DFFE_PP__3162  (.L_HI(net3162));
 sg13g2_tiehi \cpu.icache.r_tag[2][4]$_DFFE_PP__3163  (.L_HI(net3163));
 sg13g2_tiehi \cpu.icache.r_tag[2][5]$_DFFE_PP__3164  (.L_HI(net3164));
 sg13g2_tiehi \cpu.icache.r_tag[2][6]$_DFFE_PP__3165  (.L_HI(net3165));
 sg13g2_tiehi \cpu.icache.r_tag[2][7]$_DFFE_PP__3166  (.L_HI(net3166));
 sg13g2_tiehi \cpu.icache.r_tag[2][8]$_DFFE_PP__3167  (.L_HI(net3167));
 sg13g2_tiehi \cpu.icache.r_tag[2][9]$_DFFE_PP__3168  (.L_HI(net3168));
 sg13g2_tiehi \cpu.icache.r_tag[3][0]$_DFFE_PP__3169  (.L_HI(net3169));
 sg13g2_tiehi \cpu.icache.r_tag[3][10]$_DFFE_PP__3170  (.L_HI(net3170));
 sg13g2_tiehi \cpu.icache.r_tag[3][11]$_DFFE_PP__3171  (.L_HI(net3171));
 sg13g2_tiehi \cpu.icache.r_tag[3][12]$_DFFE_PP__3172  (.L_HI(net3172));
 sg13g2_tiehi \cpu.icache.r_tag[3][13]$_DFFE_PP__3173  (.L_HI(net3173));
 sg13g2_tiehi \cpu.icache.r_tag[3][14]$_DFFE_PP__3174  (.L_HI(net3174));
 sg13g2_tiehi \cpu.icache.r_tag[3][15]$_DFFE_PP__3175  (.L_HI(net3175));
 sg13g2_tiehi \cpu.icache.r_tag[3][16]$_DFFE_PP__3176  (.L_HI(net3176));
 sg13g2_tiehi \cpu.icache.r_tag[3][17]$_DFFE_PP__3177  (.L_HI(net3177));
 sg13g2_tiehi \cpu.icache.r_tag[3][18]$_DFFE_PP__3178  (.L_HI(net3178));
 sg13g2_tiehi \cpu.icache.r_tag[3][1]$_DFFE_PP__3179  (.L_HI(net3179));
 sg13g2_tiehi \cpu.icache.r_tag[3][2]$_DFFE_PP__3180  (.L_HI(net3180));
 sg13g2_tiehi \cpu.icache.r_tag[3][3]$_DFFE_PP__3181  (.L_HI(net3181));
 sg13g2_tiehi \cpu.icache.r_tag[3][4]$_DFFE_PP__3182  (.L_HI(net3182));
 sg13g2_tiehi \cpu.icache.r_tag[3][5]$_DFFE_PP__3183  (.L_HI(net3183));
 sg13g2_tiehi \cpu.icache.r_tag[3][6]$_DFFE_PP__3184  (.L_HI(net3184));
 sg13g2_tiehi \cpu.icache.r_tag[3][7]$_DFFE_PP__3185  (.L_HI(net3185));
 sg13g2_tiehi \cpu.icache.r_tag[3][8]$_DFFE_PP__3186  (.L_HI(net3186));
 sg13g2_tiehi \cpu.icache.r_tag[3][9]$_DFFE_PP__3187  (.L_HI(net3187));
 sg13g2_tiehi \cpu.icache.r_tag[4][0]$_DFFE_PP__3188  (.L_HI(net3188));
 sg13g2_tiehi \cpu.icache.r_tag[4][10]$_DFFE_PP__3189  (.L_HI(net3189));
 sg13g2_tiehi \cpu.icache.r_tag[4][11]$_DFFE_PP__3190  (.L_HI(net3190));
 sg13g2_tiehi \cpu.icache.r_tag[4][12]$_DFFE_PP__3191  (.L_HI(net3191));
 sg13g2_tiehi \cpu.icache.r_tag[4][13]$_DFFE_PP__3192  (.L_HI(net3192));
 sg13g2_tiehi \cpu.icache.r_tag[4][14]$_DFFE_PP__3193  (.L_HI(net3193));
 sg13g2_tiehi \cpu.icache.r_tag[4][15]$_DFFE_PP__3194  (.L_HI(net3194));
 sg13g2_tiehi \cpu.icache.r_tag[4][16]$_DFFE_PP__3195  (.L_HI(net3195));
 sg13g2_tiehi \cpu.icache.r_tag[4][17]$_DFFE_PP__3196  (.L_HI(net3196));
 sg13g2_tiehi \cpu.icache.r_tag[4][18]$_DFFE_PP__3197  (.L_HI(net3197));
 sg13g2_tiehi \cpu.icache.r_tag[4][1]$_DFFE_PP__3198  (.L_HI(net3198));
 sg13g2_tiehi \cpu.icache.r_tag[4][2]$_DFFE_PP__3199  (.L_HI(net3199));
 sg13g2_tiehi \cpu.icache.r_tag[4][3]$_DFFE_PP__3200  (.L_HI(net3200));
 sg13g2_tiehi \cpu.icache.r_tag[4][4]$_DFFE_PP__3201  (.L_HI(net3201));
 sg13g2_tiehi \cpu.icache.r_tag[4][5]$_DFFE_PP__3202  (.L_HI(net3202));
 sg13g2_tiehi \cpu.icache.r_tag[4][6]$_DFFE_PP__3203  (.L_HI(net3203));
 sg13g2_tiehi \cpu.icache.r_tag[4][7]$_DFFE_PP__3204  (.L_HI(net3204));
 sg13g2_tiehi \cpu.icache.r_tag[4][8]$_DFFE_PP__3205  (.L_HI(net3205));
 sg13g2_tiehi \cpu.icache.r_tag[4][9]$_DFFE_PP__3206  (.L_HI(net3206));
 sg13g2_tiehi \cpu.icache.r_tag[5][0]$_DFFE_PP__3207  (.L_HI(net3207));
 sg13g2_tiehi \cpu.icache.r_tag[5][10]$_DFFE_PP__3208  (.L_HI(net3208));
 sg13g2_tiehi \cpu.icache.r_tag[5][11]$_DFFE_PP__3209  (.L_HI(net3209));
 sg13g2_tiehi \cpu.icache.r_tag[5][12]$_DFFE_PP__3210  (.L_HI(net3210));
 sg13g2_tiehi \cpu.icache.r_tag[5][13]$_DFFE_PP__3211  (.L_HI(net3211));
 sg13g2_tiehi \cpu.icache.r_tag[5][14]$_DFFE_PP__3212  (.L_HI(net3212));
 sg13g2_tiehi \cpu.icache.r_tag[5][15]$_DFFE_PP__3213  (.L_HI(net3213));
 sg13g2_tiehi \cpu.icache.r_tag[5][16]$_DFFE_PP__3214  (.L_HI(net3214));
 sg13g2_tiehi \cpu.icache.r_tag[5][17]$_DFFE_PP__3215  (.L_HI(net3215));
 sg13g2_tiehi \cpu.icache.r_tag[5][18]$_DFFE_PP__3216  (.L_HI(net3216));
 sg13g2_tiehi \cpu.icache.r_tag[5][1]$_DFFE_PP__3217  (.L_HI(net3217));
 sg13g2_tiehi \cpu.icache.r_tag[5][2]$_DFFE_PP__3218  (.L_HI(net3218));
 sg13g2_tiehi \cpu.icache.r_tag[5][3]$_DFFE_PP__3219  (.L_HI(net3219));
 sg13g2_tiehi \cpu.icache.r_tag[5][4]$_DFFE_PP__3220  (.L_HI(net3220));
 sg13g2_tiehi \cpu.icache.r_tag[5][5]$_DFFE_PP__3221  (.L_HI(net3221));
 sg13g2_tiehi \cpu.icache.r_tag[5][6]$_DFFE_PP__3222  (.L_HI(net3222));
 sg13g2_tiehi \cpu.icache.r_tag[5][7]$_DFFE_PP__3223  (.L_HI(net3223));
 sg13g2_tiehi \cpu.icache.r_tag[5][8]$_DFFE_PP__3224  (.L_HI(net3224));
 sg13g2_tiehi \cpu.icache.r_tag[5][9]$_DFFE_PP__3225  (.L_HI(net3225));
 sg13g2_tiehi \cpu.icache.r_tag[6][0]$_DFFE_PP__3226  (.L_HI(net3226));
 sg13g2_tiehi \cpu.icache.r_tag[6][10]$_DFFE_PP__3227  (.L_HI(net3227));
 sg13g2_tiehi \cpu.icache.r_tag[6][11]$_DFFE_PP__3228  (.L_HI(net3228));
 sg13g2_tiehi \cpu.icache.r_tag[6][12]$_DFFE_PP__3229  (.L_HI(net3229));
 sg13g2_tiehi \cpu.icache.r_tag[6][13]$_DFFE_PP__3230  (.L_HI(net3230));
 sg13g2_tiehi \cpu.icache.r_tag[6][14]$_DFFE_PP__3231  (.L_HI(net3231));
 sg13g2_tiehi \cpu.icache.r_tag[6][15]$_DFFE_PP__3232  (.L_HI(net3232));
 sg13g2_tiehi \cpu.icache.r_tag[6][16]$_DFFE_PP__3233  (.L_HI(net3233));
 sg13g2_tiehi \cpu.icache.r_tag[6][17]$_DFFE_PP__3234  (.L_HI(net3234));
 sg13g2_tiehi \cpu.icache.r_tag[6][18]$_DFFE_PP__3235  (.L_HI(net3235));
 sg13g2_tiehi \cpu.icache.r_tag[6][1]$_DFFE_PP__3236  (.L_HI(net3236));
 sg13g2_tiehi \cpu.icache.r_tag[6][2]$_DFFE_PP__3237  (.L_HI(net3237));
 sg13g2_tiehi \cpu.icache.r_tag[6][3]$_DFFE_PP__3238  (.L_HI(net3238));
 sg13g2_tiehi \cpu.icache.r_tag[6][4]$_DFFE_PP__3239  (.L_HI(net3239));
 sg13g2_tiehi \cpu.icache.r_tag[6][5]$_DFFE_PP__3240  (.L_HI(net3240));
 sg13g2_tiehi \cpu.icache.r_tag[6][6]$_DFFE_PP__3241  (.L_HI(net3241));
 sg13g2_tiehi \cpu.icache.r_tag[6][7]$_DFFE_PP__3242  (.L_HI(net3242));
 sg13g2_tiehi \cpu.icache.r_tag[6][8]$_DFFE_PP__3243  (.L_HI(net3243));
 sg13g2_tiehi \cpu.icache.r_tag[6][9]$_DFFE_PP__3244  (.L_HI(net3244));
 sg13g2_tiehi \cpu.icache.r_tag[7][0]$_DFFE_PP__3245  (.L_HI(net3245));
 sg13g2_tiehi \cpu.icache.r_tag[7][10]$_DFFE_PP__3246  (.L_HI(net3246));
 sg13g2_tiehi \cpu.icache.r_tag[7][11]$_DFFE_PP__3247  (.L_HI(net3247));
 sg13g2_tiehi \cpu.icache.r_tag[7][12]$_DFFE_PP__3248  (.L_HI(net3248));
 sg13g2_tiehi \cpu.icache.r_tag[7][13]$_DFFE_PP__3249  (.L_HI(net3249));
 sg13g2_tiehi \cpu.icache.r_tag[7][14]$_DFFE_PP__3250  (.L_HI(net3250));
 sg13g2_tiehi \cpu.icache.r_tag[7][15]$_DFFE_PP__3251  (.L_HI(net3251));
 sg13g2_tiehi \cpu.icache.r_tag[7][16]$_DFFE_PP__3252  (.L_HI(net3252));
 sg13g2_tiehi \cpu.icache.r_tag[7][17]$_DFFE_PP__3253  (.L_HI(net3253));
 sg13g2_tiehi \cpu.icache.r_tag[7][18]$_DFFE_PP__3254  (.L_HI(net3254));
 sg13g2_tiehi \cpu.icache.r_tag[7][1]$_DFFE_PP__3255  (.L_HI(net3255));
 sg13g2_tiehi \cpu.icache.r_tag[7][2]$_DFFE_PP__3256  (.L_HI(net3256));
 sg13g2_tiehi \cpu.icache.r_tag[7][3]$_DFFE_PP__3257  (.L_HI(net3257));
 sg13g2_tiehi \cpu.icache.r_tag[7][4]$_DFFE_PP__3258  (.L_HI(net3258));
 sg13g2_tiehi \cpu.icache.r_tag[7][5]$_DFFE_PP__3259  (.L_HI(net3259));
 sg13g2_tiehi \cpu.icache.r_tag[7][6]$_DFFE_PP__3260  (.L_HI(net3260));
 sg13g2_tiehi \cpu.icache.r_tag[7][7]$_DFFE_PP__3261  (.L_HI(net3261));
 sg13g2_tiehi \cpu.icache.r_tag[7][8]$_DFFE_PP__3262  (.L_HI(net3262));
 sg13g2_tiehi \cpu.icache.r_tag[7][9]$_DFFE_PP__3263  (.L_HI(net3263));
 sg13g2_tiehi \cpu.icache.r_valid[0]$_SDFFE_PP0P__3264  (.L_HI(net3264));
 sg13g2_tiehi \cpu.icache.r_valid[1]$_SDFFE_PP0P__3265  (.L_HI(net3265));
 sg13g2_tiehi \cpu.icache.r_valid[2]$_SDFFE_PP0P__3266  (.L_HI(net3266));
 sg13g2_tiehi \cpu.icache.r_valid[3]$_SDFFE_PP0P__3267  (.L_HI(net3267));
 sg13g2_tiehi \cpu.icache.r_valid[4]$_SDFFE_PP0P__3268  (.L_HI(net3268));
 sg13g2_tiehi \cpu.icache.r_valid[5]$_SDFFE_PP0P__3269  (.L_HI(net3269));
 sg13g2_tiehi \cpu.icache.r_valid[6]$_SDFFE_PP0P__3270  (.L_HI(net3270));
 sg13g2_tiehi \cpu.icache.r_valid[7]$_SDFFE_PP0P__3271  (.L_HI(net3271));
 sg13g2_tiehi \cpu.intr.r_clock$_SDFFE_PN0P__3272  (.L_HI(net3272));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[0]$_DFFE_PP__3273  (.L_HI(net3273));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[10]$_DFFE_PP__3274  (.L_HI(net3274));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[11]$_DFFE_PP__3275  (.L_HI(net3275));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[12]$_DFFE_PP__3276  (.L_HI(net3276));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[13]$_DFFE_PP__3277  (.L_HI(net3277));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[14]$_DFFE_PP__3278  (.L_HI(net3278));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[15]$_DFFE_PP__3279  (.L_HI(net3279));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[16]$_DFFE_PP__3280  (.L_HI(net3280));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[17]$_DFFE_PP__3281  (.L_HI(net3281));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[18]$_DFFE_PP__3282  (.L_HI(net3282));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[19]$_DFFE_PP__3283  (.L_HI(net3283));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[1]$_DFFE_PP__3284  (.L_HI(net3284));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[20]$_DFFE_PP__3285  (.L_HI(net3285));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[21]$_DFFE_PP__3286  (.L_HI(net3286));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[22]$_DFFE_PP__3287  (.L_HI(net3287));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[23]$_DFFE_PP__3288  (.L_HI(net3288));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[24]$_DFFE_PP__3289  (.L_HI(net3289));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[25]$_DFFE_PP__3290  (.L_HI(net3290));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[26]$_DFFE_PP__3291  (.L_HI(net3291));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[27]$_DFFE_PP__3292  (.L_HI(net3292));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[28]$_DFFE_PP__3293  (.L_HI(net3293));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[29]$_DFFE_PP__3294  (.L_HI(net3294));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[2]$_DFFE_PP__3295  (.L_HI(net3295));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[30]$_DFFE_PP__3296  (.L_HI(net3296));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[31]$_DFFE_PP__3297  (.L_HI(net3297));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[3]$_DFFE_PP__3298  (.L_HI(net3298));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[4]$_DFFE_PP__3299  (.L_HI(net3299));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[5]$_DFFE_PP__3300  (.L_HI(net3300));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[6]$_DFFE_PP__3301  (.L_HI(net3301));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[7]$_DFFE_PP__3302  (.L_HI(net3302));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[8]$_DFFE_PP__3303  (.L_HI(net3303));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[9]$_DFFE_PP__3304  (.L_HI(net3304));
 sg13g2_tiehi \cpu.intr.r_clock_count[0]$_DFF_P__3305  (.L_HI(net3305));
 sg13g2_tiehi \cpu.intr.r_clock_count[10]$_DFF_P__3306  (.L_HI(net3306));
 sg13g2_tiehi \cpu.intr.r_clock_count[11]$_DFF_P__3307  (.L_HI(net3307));
 sg13g2_tiehi \cpu.intr.r_clock_count[12]$_DFF_P__3308  (.L_HI(net3308));
 sg13g2_tiehi \cpu.intr.r_clock_count[13]$_DFF_P__3309  (.L_HI(net3309));
 sg13g2_tiehi \cpu.intr.r_clock_count[14]$_DFF_P__3310  (.L_HI(net3310));
 sg13g2_tiehi \cpu.intr.r_clock_count[15]$_DFF_P__3311  (.L_HI(net3311));
 sg13g2_tiehi \cpu.intr.r_clock_count[16]$_DFFE_PN__3312  (.L_HI(net3312));
 sg13g2_tiehi \cpu.intr.r_clock_count[17]$_DFFE_PN__3313  (.L_HI(net3313));
 sg13g2_tiehi \cpu.intr.r_clock_count[18]$_DFFE_PN__3314  (.L_HI(net3314));
 sg13g2_tiehi \cpu.intr.r_clock_count[19]$_DFFE_PN__3315  (.L_HI(net3315));
 sg13g2_tiehi \cpu.intr.r_clock_count[1]$_DFF_P__3316  (.L_HI(net3316));
 sg13g2_tiehi \cpu.intr.r_clock_count[20]$_DFFE_PN__3317  (.L_HI(net3317));
 sg13g2_tiehi \cpu.intr.r_clock_count[21]$_DFFE_PN__3318  (.L_HI(net3318));
 sg13g2_tiehi \cpu.intr.r_clock_count[22]$_DFFE_PN__3319  (.L_HI(net3319));
 sg13g2_tiehi \cpu.intr.r_clock_count[23]$_DFFE_PN__3320  (.L_HI(net3320));
 sg13g2_tiehi \cpu.intr.r_clock_count[24]$_DFFE_PN__3321  (.L_HI(net3321));
 sg13g2_tiehi \cpu.intr.r_clock_count[25]$_DFFE_PN__3322  (.L_HI(net3322));
 sg13g2_tiehi \cpu.intr.r_clock_count[26]$_DFFE_PN__3323  (.L_HI(net3323));
 sg13g2_tiehi \cpu.intr.r_clock_count[27]$_DFFE_PN__3324  (.L_HI(net3324));
 sg13g2_tiehi \cpu.intr.r_clock_count[28]$_DFFE_PN__3325  (.L_HI(net3325));
 sg13g2_tiehi \cpu.intr.r_clock_count[29]$_DFFE_PN__3326  (.L_HI(net3326));
 sg13g2_tiehi \cpu.intr.r_clock_count[2]$_DFF_P__3327  (.L_HI(net3327));
 sg13g2_tiehi \cpu.intr.r_clock_count[30]$_DFFE_PN__3328  (.L_HI(net3328));
 sg13g2_tiehi \cpu.intr.r_clock_count[31]$_DFFE_PN__3329  (.L_HI(net3329));
 sg13g2_tiehi \cpu.intr.r_clock_count[3]$_DFF_P__3330  (.L_HI(net3330));
 sg13g2_tiehi \cpu.intr.r_clock_count[4]$_DFF_P__3331  (.L_HI(net3331));
 sg13g2_tiehi \cpu.intr.r_clock_count[5]$_DFF_P__3332  (.L_HI(net3332));
 sg13g2_tiehi \cpu.intr.r_clock_count[6]$_DFF_P__3333  (.L_HI(net3333));
 sg13g2_tiehi \cpu.intr.r_clock_count[7]$_DFF_P__3334  (.L_HI(net3334));
 sg13g2_tiehi \cpu.intr.r_clock_count[8]$_DFF_P__3335  (.L_HI(net3335));
 sg13g2_tiehi \cpu.intr.r_clock_count[9]$_DFF_P__3336  (.L_HI(net3336));
 sg13g2_tiehi \cpu.intr.r_enable[0]$_SDFFE_PN0P__3337  (.L_HI(net3337));
 sg13g2_tiehi \cpu.intr.r_enable[1]$_SDFFE_PN0P__3338  (.L_HI(net3338));
 sg13g2_tiehi \cpu.intr.r_enable[2]$_SDFFE_PN0P__3339  (.L_HI(net3339));
 sg13g2_tiehi \cpu.intr.r_enable[3]$_SDFFE_PN0P__3340  (.L_HI(net3340));
 sg13g2_tiehi \cpu.intr.r_enable[4]$_SDFFE_PN0P__3341  (.L_HI(net3341));
 sg13g2_tiehi \cpu.intr.r_enable[5]$_SDFFE_PN0P__3342  (.L_HI(net3342));
 sg13g2_tiehi \cpu.intr.r_timer$_SDFFE_PN0P__3343  (.L_HI(net3343));
 sg13g2_tiehi \cpu.intr.r_timer_count[0]$_DFF_P__3344  (.L_HI(net3344));
 sg13g2_tiehi \cpu.intr.r_timer_count[10]$_DFF_P__3345  (.L_HI(net3345));
 sg13g2_tiehi \cpu.intr.r_timer_count[11]$_DFF_P__3346  (.L_HI(net3346));
 sg13g2_tiehi \cpu.intr.r_timer_count[12]$_DFF_P__3347  (.L_HI(net3347));
 sg13g2_tiehi \cpu.intr.r_timer_count[13]$_DFF_P__3348  (.L_HI(net3348));
 sg13g2_tiehi \cpu.intr.r_timer_count[14]$_DFF_P__3349  (.L_HI(net3349));
 sg13g2_tiehi \cpu.intr.r_timer_count[15]$_DFF_P__3350  (.L_HI(net3350));
 sg13g2_tiehi \cpu.intr.r_timer_count[16]$_DFF_P__3351  (.L_HI(net3351));
 sg13g2_tiehi \cpu.intr.r_timer_count[17]$_DFF_P__3352  (.L_HI(net3352));
 sg13g2_tiehi \cpu.intr.r_timer_count[18]$_DFF_P__3353  (.L_HI(net3353));
 sg13g2_tiehi \cpu.intr.r_timer_count[19]$_DFF_P__3354  (.L_HI(net3354));
 sg13g2_tiehi \cpu.intr.r_timer_count[1]$_DFF_P__3355  (.L_HI(net3355));
 sg13g2_tiehi \cpu.intr.r_timer_count[20]$_DFF_P__3356  (.L_HI(net3356));
 sg13g2_tiehi \cpu.intr.r_timer_count[21]$_DFF_P__3357  (.L_HI(net3357));
 sg13g2_tiehi \cpu.intr.r_timer_count[22]$_DFF_P__3358  (.L_HI(net3358));
 sg13g2_tiehi \cpu.intr.r_timer_count[23]$_DFF_P__3359  (.L_HI(net3359));
 sg13g2_tiehi \cpu.intr.r_timer_count[2]$_DFF_P__3360  (.L_HI(net3360));
 sg13g2_tiehi \cpu.intr.r_timer_count[3]$_DFF_P__3361  (.L_HI(net3361));
 sg13g2_tiehi \cpu.intr.r_timer_count[4]$_DFF_P__3362  (.L_HI(net3362));
 sg13g2_tiehi \cpu.intr.r_timer_count[5]$_DFF_P__3363  (.L_HI(net3363));
 sg13g2_tiehi \cpu.intr.r_timer_count[6]$_DFF_P__3364  (.L_HI(net3364));
 sg13g2_tiehi \cpu.intr.r_timer_count[7]$_DFF_P__3365  (.L_HI(net3365));
 sg13g2_tiehi \cpu.intr.r_timer_count[8]$_DFF_P__3366  (.L_HI(net3366));
 sg13g2_tiehi \cpu.intr.r_timer_count[9]$_DFF_P__3367  (.L_HI(net3367));
 sg13g2_tiehi \cpu.intr.r_timer_reload[0]$_DFFE_PP__3368  (.L_HI(net3368));
 sg13g2_tiehi \cpu.intr.r_timer_reload[10]$_DFFE_PP__3369  (.L_HI(net3369));
 sg13g2_tiehi \cpu.intr.r_timer_reload[11]$_DFFE_PP__3370  (.L_HI(net3370));
 sg13g2_tiehi \cpu.intr.r_timer_reload[12]$_DFFE_PP__3371  (.L_HI(net3371));
 sg13g2_tiehi \cpu.intr.r_timer_reload[13]$_DFFE_PP__3372  (.L_HI(net3372));
 sg13g2_tiehi \cpu.intr.r_timer_reload[14]$_DFFE_PP__3373  (.L_HI(net3373));
 sg13g2_tiehi \cpu.intr.r_timer_reload[15]$_DFFE_PP__3374  (.L_HI(net3374));
 sg13g2_tiehi \cpu.intr.r_timer_reload[16]$_DFFE_PP__3375  (.L_HI(net3375));
 sg13g2_tiehi \cpu.intr.r_timer_reload[17]$_DFFE_PP__3376  (.L_HI(net3376));
 sg13g2_tiehi \cpu.intr.r_timer_reload[18]$_DFFE_PP__3377  (.L_HI(net3377));
 sg13g2_tiehi \cpu.intr.r_timer_reload[19]$_DFFE_PP__3378  (.L_HI(net3378));
 sg13g2_tiehi \cpu.intr.r_timer_reload[1]$_DFFE_PP__3379  (.L_HI(net3379));
 sg13g2_tiehi \cpu.intr.r_timer_reload[20]$_DFFE_PP__3380  (.L_HI(net3380));
 sg13g2_tiehi \cpu.intr.r_timer_reload[21]$_DFFE_PP__3381  (.L_HI(net3381));
 sg13g2_tiehi \cpu.intr.r_timer_reload[22]$_DFFE_PP__3382  (.L_HI(net3382));
 sg13g2_tiehi \cpu.intr.r_timer_reload[23]$_DFFE_PP__3383  (.L_HI(net3383));
 sg13g2_tiehi \cpu.intr.r_timer_reload[2]$_DFFE_PP__3384  (.L_HI(net3384));
 sg13g2_tiehi \cpu.intr.r_timer_reload[3]$_DFFE_PP__3385  (.L_HI(net3385));
 sg13g2_tiehi \cpu.intr.r_timer_reload[4]$_DFFE_PP__3386  (.L_HI(net3386));
 sg13g2_tiehi \cpu.intr.r_timer_reload[5]$_DFFE_PP__3387  (.L_HI(net3387));
 sg13g2_tiehi \cpu.intr.r_timer_reload[6]$_DFFE_PP__3388  (.L_HI(net3388));
 sg13g2_tiehi \cpu.intr.r_timer_reload[7]$_DFFE_PP__3389  (.L_HI(net3389));
 sg13g2_tiehi \cpu.intr.r_timer_reload[8]$_DFFE_PP__3390  (.L_HI(net3390));
 sg13g2_tiehi \cpu.intr.r_timer_reload[9]$_DFFE_PP__3391  (.L_HI(net3391));
 sg13g2_tiehi \cpu.qspi.r_count[0]$_DFFE_PP__3392  (.L_HI(net3392));
 sg13g2_tiehi \cpu.qspi.r_count[1]$_DFFE_PP__3393  (.L_HI(net3393));
 sg13g2_tiehi \cpu.qspi.r_count[2]$_DFFE_PP__3394  (.L_HI(net3394));
 sg13g2_tiehi \cpu.qspi.r_count[3]$_DFFE_PP__3395  (.L_HI(net3395));
 sg13g2_tiehi \cpu.qspi.r_count[4]$_DFFE_PP__3396  (.L_HI(net3396));
 sg13g2_tiehi \cpu.qspi.r_cs[0]$_SDFFE_PN1P__3397  (.L_HI(net3397));
 sg13g2_tiehi \cpu.qspi.r_cs[1]$_SDFFE_PN1P__3398  (.L_HI(net3398));
 sg13g2_tiehi \cpu.qspi.r_cs[2]$_SDFFE_PN1P__3399  (.L_HI(net3399));
 sg13g2_tiehi \cpu.qspi.r_ind$_SDFFE_PN0N__3400  (.L_HI(net3400));
 sg13g2_tiehi \cpu.qspi.r_mask[0]$_SDFFE_PN0P__3401  (.L_HI(net3401));
 sg13g2_tiehi \cpu.qspi.r_mask[1]$_SDFFE_PN1P__3402  (.L_HI(net3402));
 sg13g2_tiehi \cpu.qspi.r_mask[2]$_SDFFE_PN0P__3403  (.L_HI(net3403));
 sg13g2_tiehi \cpu.qspi.r_quad[0]$_SDFFE_PN1P__3404  (.L_HI(net3404));
 sg13g2_tiehi \cpu.qspi.r_quad[1]$_SDFFE_PN0P__3405  (.L_HI(net3405));
 sg13g2_tiehi \cpu.qspi.r_quad[2]$_SDFFE_PN1P__3406  (.L_HI(net3406));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][0]$_SDFFCE_PN0P__3407  (.L_HI(net3407));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][1]$_SDFFCE_PN0P__3408  (.L_HI(net3408));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][2]$_SDFFCE_PN1P__3409  (.L_HI(net3409));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][3]$_SDFFCE_PN0P__3410  (.L_HI(net3410));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][0]$_SDFFCE_PN0P__3411  (.L_HI(net3411));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][1]$_SDFFCE_PN0P__3412  (.L_HI(net3412));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][2]$_SDFFCE_PN1P__3413  (.L_HI(net3413));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][3]$_SDFFCE_PN0P__3414  (.L_HI(net3414));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][0]$_SDFFCE_PN0P__3415  (.L_HI(net3415));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][1]$_SDFFCE_PN0P__3416  (.L_HI(net3416));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][2]$_SDFFCE_PN1P__3417  (.L_HI(net3417));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][3]$_SDFFCE_PN0P__3418  (.L_HI(net3418));
 sg13g2_tiehi \cpu.qspi.r_rom_mode[0]$_SDFFE_PN1P__3419  (.L_HI(net3419));
 sg13g2_tiehi \cpu.qspi.r_rom_mode[1]$_SDFFE_PN1P__3420  (.L_HI(net3420));
 sg13g2_tiehi \cpu.qspi.r_rstrobe_d$_DFF_P__3421  (.L_HI(net3421));
 sg13g2_tiehi \cpu.qspi.r_state[0]$_DFF_P__3422  (.L_HI(net3422));
 sg13g2_tiehi \cpu.qspi.r_state[10]$_DFF_P__3423  (.L_HI(net3423));
 sg13g2_tiehi \cpu.qspi.r_state[11]$_DFF_P__3424  (.L_HI(net3424));
 sg13g2_tiehi \cpu.qspi.r_state[12]$_DFF_P__3425  (.L_HI(net3425));
 sg13g2_tiehi \cpu.qspi.r_state[13]$_DFF_P__3426  (.L_HI(net3426));
 sg13g2_tiehi \cpu.qspi.r_state[14]$_DFF_P__3427  (.L_HI(net3427));
 sg13g2_tiehi \cpu.qspi.r_state[15]$_DFF_P__3428  (.L_HI(net3428));
 sg13g2_tiehi \cpu.qspi.r_state[16]$_DFF_P__3429  (.L_HI(net3429));
 sg13g2_tiehi \cpu.qspi.r_state[17]$_DFF_P__3430  (.L_HI(net3430));
 sg13g2_tiehi \cpu.qspi.r_state[1]$_DFF_P__3431  (.L_HI(net3431));
 sg13g2_tiehi \cpu.qspi.r_state[2]$_DFF_P__3432  (.L_HI(net3432));
 sg13g2_tiehi \cpu.qspi.r_state[3]$_DFF_P__3433  (.L_HI(net3433));
 sg13g2_tiehi \cpu.qspi.r_state[4]$_DFF_P__3434  (.L_HI(net3434));
 sg13g2_tiehi \cpu.qspi.r_state[5]$_DFF_P__3435  (.L_HI(net3435));
 sg13g2_tiehi \cpu.qspi.r_state[6]$_DFF_P__3436  (.L_HI(net3436));
 sg13g2_tiehi \cpu.qspi.r_state[7]$_DFF_P__3437  (.L_HI(net3437));
 sg13g2_tiehi \cpu.qspi.r_state[8]$_DFF_P__3438  (.L_HI(net3438));
 sg13g2_tiehi \cpu.qspi.r_state[9]$_DFF_P__3439  (.L_HI(net3439));
 sg13g2_tiehi \cpu.qspi.r_uio_oe[0]$_SDFFE_PN0P__3440  (.L_HI(net3440));
 sg13g2_tiehi \cpu.qspi.r_uio_oe[1]$_SDFFE_PN0P__3441  (.L_HI(net3441));
 sg13g2_tiehi \cpu.qspi.r_uio_out[0]$_DFFE_PP__3442  (.L_HI(net3442));
 sg13g2_tiehi \cpu.qspi.r_uio_out[1]$_DFFE_PP__3443  (.L_HI(net3443));
 sg13g2_tiehi \cpu.qspi.r_uio_out[2]$_DFFE_PP__3444  (.L_HI(net3444));
 sg13g2_tiehi \cpu.qspi.r_uio_out[3]$_DFFE_PP__3445  (.L_HI(net3445));
 sg13g2_tiehi \cpu.qspi.r_wstrobe_d$_DFF_P__3446  (.L_HI(net3446));
 sg13g2_tiehi \cpu.qspi.r_wstrobe_i$_DFF_P__3447  (.L_HI(net3447));
 sg13g2_tiehi \cpu.r_clk_invert$_DFFE_PN__3448  (.L_HI(net3448));
 sg13g2_tiehi \cpu.spi.r_bits[0]$_SDFFE_PN1P__3449  (.L_HI(net3449));
 sg13g2_tiehi \cpu.spi.r_bits[1]$_SDFFE_PN1P__3450  (.L_HI(net3450));
 sg13g2_tiehi \cpu.spi.r_bits[2]$_SDFFE_PN1P__3451  (.L_HI(net3451));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][0]$_DFFE_PP__3452  (.L_HI(net3452));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][1]$_DFFE_PP__3453  (.L_HI(net3453));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][2]$_DFFE_PP__3454  (.L_HI(net3454));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][3]$_DFFE_PP__3455  (.L_HI(net3455));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][4]$_DFFE_PP__3456  (.L_HI(net3456));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][5]$_DFFE_PP__3457  (.L_HI(net3457));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][6]$_DFFE_PP__3458  (.L_HI(net3458));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][7]$_DFFE_PP__3459  (.L_HI(net3459));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][0]$_DFFE_PP__3460  (.L_HI(net3460));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][1]$_DFFE_PP__3461  (.L_HI(net3461));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][2]$_DFFE_PP__3462  (.L_HI(net3462));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][3]$_DFFE_PP__3463  (.L_HI(net3463));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][4]$_DFFE_PP__3464  (.L_HI(net3464));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][5]$_DFFE_PP__3465  (.L_HI(net3465));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][6]$_DFFE_PP__3466  (.L_HI(net3466));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][7]$_DFFE_PP__3467  (.L_HI(net3467));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][0]$_DFFE_PP__3468  (.L_HI(net3468));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][1]$_DFFE_PP__3469  (.L_HI(net3469));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][2]$_DFFE_PP__3470  (.L_HI(net3470));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][3]$_DFFE_PP__3471  (.L_HI(net3471));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][4]$_DFFE_PP__3472  (.L_HI(net3472));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][5]$_DFFE_PP__3473  (.L_HI(net3473));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][6]$_DFFE_PP__3474  (.L_HI(net3474));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][7]$_DFFE_PP__3475  (.L_HI(net3475));
 sg13g2_tiehi \cpu.spi.r_count[0]$_DFFE_PP__3476  (.L_HI(net3476));
 sg13g2_tiehi \cpu.spi.r_count[1]$_DFFE_PP__3477  (.L_HI(net3477));
 sg13g2_tiehi \cpu.spi.r_count[2]$_DFFE_PP__3478  (.L_HI(net3478));
 sg13g2_tiehi \cpu.spi.r_count[3]$_DFFE_PP__3479  (.L_HI(net3479));
 sg13g2_tiehi \cpu.spi.r_count[4]$_DFFE_PP__3480  (.L_HI(net3480));
 sg13g2_tiehi \cpu.spi.r_count[5]$_DFFE_PP__3481  (.L_HI(net3481));
 sg13g2_tiehi \cpu.spi.r_count[6]$_DFFE_PP__3482  (.L_HI(net3482));
 sg13g2_tiehi \cpu.spi.r_count[7]$_DFFE_PP__3483  (.L_HI(net3483));
 sg13g2_tiehi \cpu.spi.r_cs[0]$_SDFFE_PN1P__3484  (.L_HI(net3484));
 sg13g2_tiehi \cpu.spi.r_cs[1]$_SDFFE_PN1P__3485  (.L_HI(net3485));
 sg13g2_tiehi \cpu.spi.r_cs[2]$_SDFFE_PN1P__3486  (.L_HI(net3486));
 sg13g2_tiehi \cpu.spi.r_in[0]$_DFFE_PP__3487  (.L_HI(net3487));
 sg13g2_tiehi \cpu.spi.r_in[1]$_DFFE_PP__3488  (.L_HI(net3488));
 sg13g2_tiehi \cpu.spi.r_in[2]$_DFFE_PP__3489  (.L_HI(net3489));
 sg13g2_tiehi \cpu.spi.r_in[3]$_DFFE_PP__3490  (.L_HI(net3490));
 sg13g2_tiehi \cpu.spi.r_in[4]$_DFFE_PP__3491  (.L_HI(net3491));
 sg13g2_tiehi \cpu.spi.r_in[5]$_DFFE_PP__3492  (.L_HI(net3492));
 sg13g2_tiehi \cpu.spi.r_in[6]$_DFFE_PP__3493  (.L_HI(net3493));
 sg13g2_tiehi \cpu.spi.r_in[7]$_DFFE_PP__3494  (.L_HI(net3494));
 sg13g2_tiehi \cpu.spi.r_interrupt$_SDFFE_PN0P__3495  (.L_HI(net3495));
 sg13g2_tiehi \cpu.spi.r_mode[0][0]$_DFFE_PP__3496  (.L_HI(net3496));
 sg13g2_tiehi \cpu.spi.r_mode[0][1]$_DFFE_PP__3497  (.L_HI(net3497));
 sg13g2_tiehi \cpu.spi.r_mode[1][0]$_DFFE_PP__3498  (.L_HI(net3498));
 sg13g2_tiehi \cpu.spi.r_mode[1][1]$_DFFE_PP__3499  (.L_HI(net3499));
 sg13g2_tiehi \cpu.spi.r_mode[2][0]$_DFFE_PP__3500  (.L_HI(net3500));
 sg13g2_tiehi \cpu.spi.r_mode[2][1]$_DFFE_PP__3501  (.L_HI(net3501));
 sg13g2_tiehi \cpu.spi.r_out[0]$_DFFE_PP__3502  (.L_HI(net3502));
 sg13g2_tiehi \cpu.spi.r_out[1]$_DFFE_PP__3503  (.L_HI(net3503));
 sg13g2_tiehi \cpu.spi.r_out[2]$_DFFE_PP__3504  (.L_HI(net3504));
 sg13g2_tiehi \cpu.spi.r_out[3]$_DFFE_PP__3505  (.L_HI(net3505));
 sg13g2_tiehi \cpu.spi.r_out[4]$_DFFE_PP__3506  (.L_HI(net3506));
 sg13g2_tiehi \cpu.spi.r_out[5]$_DFFE_PP__3507  (.L_HI(net3507));
 sg13g2_tiehi \cpu.spi.r_out[6]$_DFFE_PP__3508  (.L_HI(net3508));
 sg13g2_tiehi \cpu.spi.r_out[7]$_DFFE_PP__3509  (.L_HI(net3509));
 sg13g2_tiehi \cpu.spi.r_ready$_SDFFE_PN1P__3510  (.L_HI(net3510));
 sg13g2_tiehi \cpu.spi.r_searching$_SDFFE_PN0P__3511  (.L_HI(net3511));
 sg13g2_tiehi \cpu.spi.r_sel[0]$_DFFE_PP__3512  (.L_HI(net3512));
 sg13g2_tiehi \cpu.spi.r_sel[1]$_DFFE_PP__3513  (.L_HI(net3513));
 sg13g2_tiehi \cpu.spi.r_src[0]$_DFFE_PP__3514  (.L_HI(net3514));
 sg13g2_tiehi \cpu.spi.r_src[1]$_DFFE_PP__3515  (.L_HI(net3515));
 sg13g2_tiehi \cpu.spi.r_src[2]$_DFFE_PP__3516  (.L_HI(net3516));
 sg13g2_tiehi \cpu.spi.r_state[0]$_DFF_P__3517  (.L_HI(net3517));
 sg13g2_tiehi \cpu.spi.r_state[1]$_DFF_P__3518  (.L_HI(net3518));
 sg13g2_tiehi \cpu.spi.r_state[2]$_DFF_P__3519  (.L_HI(net3519));
 sg13g2_tiehi \cpu.spi.r_state[3]$_DFF_P__3520  (.L_HI(net3520));
 sg13g2_tiehi \cpu.spi.r_state[4]$_DFF_P__3521  (.L_HI(net3521));
 sg13g2_tiehi \cpu.spi.r_state[5]$_DFF_P__3522  (.L_HI(net3522));
 sg13g2_tiehi \cpu.spi.r_state[6]$_DFF_P__3523  (.L_HI(net3523));
 sg13g2_tiehi \cpu.spi.r_timeout[0]$_DFFE_PP__3524  (.L_HI(net3524));
 sg13g2_tiehi \cpu.spi.r_timeout[1]$_DFFE_PP__3525  (.L_HI(net3525));
 sg13g2_tiehi \cpu.spi.r_timeout[2]$_DFFE_PP__3526  (.L_HI(net3526));
 sg13g2_tiehi \cpu.spi.r_timeout[3]$_DFFE_PP__3527  (.L_HI(net3527));
 sg13g2_tiehi \cpu.spi.r_timeout[4]$_DFFE_PP__3528  (.L_HI(net3528));
 sg13g2_tiehi \cpu.spi.r_timeout[5]$_DFFE_PP__3529  (.L_HI(net3529));
 sg13g2_tiehi \cpu.spi.r_timeout[6]$_DFFE_PP__3530  (.L_HI(net3530));
 sg13g2_tiehi \cpu.spi.r_timeout[7]$_DFFE_PP__3531  (.L_HI(net3531));
 sg13g2_tiehi \cpu.spi.r_timeout_count[0]$_DFFE_PP__3532  (.L_HI(net3532));
 sg13g2_tiehi \cpu.spi.r_timeout_count[1]$_DFFE_PP__3533  (.L_HI(net3533));
 sg13g2_tiehi \cpu.spi.r_timeout_count[2]$_DFFE_PP__3534  (.L_HI(net3534));
 sg13g2_tiehi \cpu.spi.r_timeout_count[3]$_DFFE_PP__3535  (.L_HI(net3535));
 sg13g2_tiehi \cpu.spi.r_timeout_count[4]$_DFFE_PP__3536  (.L_HI(net3536));
 sg13g2_tiehi \cpu.spi.r_timeout_count[5]$_DFFE_PP__3537  (.L_HI(net3537));
 sg13g2_tiehi \cpu.spi.r_timeout_count[6]$_DFFE_PP__3538  (.L_HI(net3538));
 sg13g2_tiehi \cpu.spi.r_timeout_count[7]$_DFFE_PP__3539  (.L_HI(net3539));
 sg13g2_tiehi \cpu.uart.r_div[0]$_DFF_P__3540  (.L_HI(net3540));
 sg13g2_tiehi \cpu.uart.r_div[10]$_DFF_P__3541  (.L_HI(net3541));
 sg13g2_tiehi \cpu.uart.r_div[11]$_DFF_P__3542  (.L_HI(net3542));
 sg13g2_tiehi \cpu.uart.r_div[1]$_DFF_P__3543  (.L_HI(net3543));
 sg13g2_tiehi \cpu.uart.r_div[2]$_DFF_P__3544  (.L_HI(net3544));
 sg13g2_tiehi \cpu.uart.r_div[3]$_DFF_P__3545  (.L_HI(net3545));
 sg13g2_tiehi \cpu.uart.r_div[4]$_DFF_P__3546  (.L_HI(net3546));
 sg13g2_tiehi \cpu.uart.r_div[5]$_DFF_P__3547  (.L_HI(net3547));
 sg13g2_tiehi \cpu.uart.r_div[6]$_DFF_P__3548  (.L_HI(net3548));
 sg13g2_tiehi \cpu.uart.r_div[7]$_DFF_P__3549  (.L_HI(net3549));
 sg13g2_tiehi \cpu.uart.r_div[8]$_DFF_P__3550  (.L_HI(net3550));
 sg13g2_tiehi \cpu.uart.r_div[9]$_DFF_P__3551  (.L_HI(net3551));
 sg13g2_tiehi \cpu.uart.r_div_value[0]$_SDFFE_PN1P__3552  (.L_HI(net3552));
 sg13g2_tiehi \cpu.uart.r_div_value[10]$_SDFFE_PN0P__3553  (.L_HI(net3553));
 sg13g2_tiehi \cpu.uart.r_div_value[11]$_SDFFE_PN0P__3554  (.L_HI(net3554));
 sg13g2_tiehi \cpu.uart.r_div_value[1]$_SDFFE_PN0P__3555  (.L_HI(net3555));
 sg13g2_tiehi \cpu.uart.r_div_value[2]$_SDFFE_PN0P__3556  (.L_HI(net3556));
 sg13g2_tiehi \cpu.uart.r_div_value[3]$_SDFFE_PN0P__3557  (.L_HI(net3557));
 sg13g2_tiehi \cpu.uart.r_div_value[4]$_SDFFE_PN0P__3558  (.L_HI(net3558));
 sg13g2_tiehi \cpu.uart.r_div_value[5]$_SDFFE_PN0P__3559  (.L_HI(net3559));
 sg13g2_tiehi \cpu.uart.r_div_value[6]$_SDFFE_PN0P__3560  (.L_HI(net3560));
 sg13g2_tiehi \cpu.uart.r_div_value[7]$_SDFFE_PN0P__3561  (.L_HI(net3561));
 sg13g2_tiehi \cpu.uart.r_div_value[8]$_SDFFE_PN0P__3562  (.L_HI(net3562));
 sg13g2_tiehi \cpu.uart.r_div_value[9]$_SDFFE_PN0P__3563  (.L_HI(net3563));
 sg13g2_tiehi \cpu.uart.r_ib[0]$_DFFE_PP__3564  (.L_HI(net3564));
 sg13g2_tiehi \cpu.uart.r_ib[1]$_DFFE_PP__3565  (.L_HI(net3565));
 sg13g2_tiehi \cpu.uart.r_ib[2]$_DFFE_PP__3566  (.L_HI(net3566));
 sg13g2_tiehi \cpu.uart.r_ib[3]$_DFFE_PP__3567  (.L_HI(net3567));
 sg13g2_tiehi \cpu.uart.r_ib[4]$_DFFE_PP__3568  (.L_HI(net3568));
 sg13g2_tiehi \cpu.uart.r_ib[5]$_DFFE_PP__3569  (.L_HI(net3569));
 sg13g2_tiehi \cpu.uart.r_ib[6]$_DFFE_PP__3570  (.L_HI(net3570));
 sg13g2_tiehi \cpu.uart.r_in[0]$_DFFE_PP__3571  (.L_HI(net3571));
 sg13g2_tiehi \cpu.uart.r_in[1]$_DFFE_PP__3572  (.L_HI(net3572));
 sg13g2_tiehi \cpu.uart.r_in[2]$_DFFE_PP__3573  (.L_HI(net3573));
 sg13g2_tiehi \cpu.uart.r_in[3]$_DFFE_PP__3574  (.L_HI(net3574));
 sg13g2_tiehi \cpu.uart.r_in[4]$_DFFE_PP__3575  (.L_HI(net3575));
 sg13g2_tiehi \cpu.uart.r_in[5]$_DFFE_PP__3576  (.L_HI(net3576));
 sg13g2_tiehi \cpu.uart.r_in[6]$_DFFE_PP__3577  (.L_HI(net3577));
 sg13g2_tiehi \cpu.uart.r_in[7]$_DFFE_PP__3578  (.L_HI(net3578));
 sg13g2_tiehi \cpu.uart.r_out[0]$_DFFE_PP__3579  (.L_HI(net3579));
 sg13g2_tiehi \cpu.uart.r_out[1]$_DFFE_PP__3580  (.L_HI(net3580));
 sg13g2_tiehi \cpu.uart.r_out[2]$_DFFE_PP__3581  (.L_HI(net3581));
 sg13g2_tiehi \cpu.uart.r_out[3]$_DFFE_PP__3582  (.L_HI(net3582));
 sg13g2_tiehi \cpu.uart.r_out[4]$_DFFE_PP__3583  (.L_HI(net3583));
 sg13g2_tiehi \cpu.uart.r_out[5]$_DFFE_PP__3584  (.L_HI(net3584));
 sg13g2_tiehi \cpu.uart.r_out[6]$_DFFE_PP__3585  (.L_HI(net3585));
 sg13g2_tiehi \cpu.uart.r_out[7]$_DFFE_PP__3586  (.L_HI(net3586));
 sg13g2_tiehi \cpu.uart.r_r$_DFF_P__3587  (.L_HI(net3587));
 sg13g2_tiehi \cpu.uart.r_r_int$_SDFFE_PN0P__3588  (.L_HI(net3588));
 sg13g2_tiehi \cpu.uart.r_r_invert$_SDFFE_PN0P__3589  (.L_HI(net3589));
 sg13g2_tiehi \cpu.uart.r_rcnt[0]$_DFFE_PP__3590  (.L_HI(net3590));
 sg13g2_tiehi \cpu.uart.r_rcnt[1]$_DFFE_PP__3591  (.L_HI(net3591));
 sg13g2_tiehi \cpu.uart.r_rstate[0]$_SDFFE_PN0P__3592  (.L_HI(net3592));
 sg13g2_tiehi \cpu.uart.r_rstate[1]$_SDFFE_PN0P__3593  (.L_HI(net3593));
 sg13g2_tiehi \cpu.uart.r_rstate[2]$_SDFFE_PN0P__3594  (.L_HI(net3594));
 sg13g2_tiehi \cpu.uart.r_rstate[3]$_SDFFE_PN0P__3595  (.L_HI(net3595));
 sg13g2_tiehi \cpu.uart.r_x$_DFFE_PP__3596  (.L_HI(net3596));
 sg13g2_tiehi \cpu.uart.r_x_int$_SDFFE_PN0P__3597  (.L_HI(net3597));
 sg13g2_tiehi \cpu.uart.r_x_invert$_SDFFE_PN0P__3598  (.L_HI(net3598));
 sg13g2_tiehi \cpu.uart.r_xcnt[0]$_DFFE_PP__3599  (.L_HI(net3599));
 sg13g2_tiehi \cpu.uart.r_xcnt[1]$_DFFE_PP__3600  (.L_HI(net3600));
 sg13g2_tiehi \cpu.uart.r_xstate[0]$_SDFFE_PN0P__3601  (.L_HI(net3601));
 sg13g2_tiehi \cpu.uart.r_xstate[1]$_SDFFE_PN0P__3602  (.L_HI(net3602));
 sg13g2_tiehi \cpu.uart.r_xstate[2]$_SDFFE_PN0P__3603  (.L_HI(net3603));
 sg13g2_tiehi \cpu.uart.r_xstate[3]$_SDFFE_PN0P__3604  (.L_HI(net3604));
 sg13g2_tiehi \r_reset$_DFF_P__3605  (.L_HI(net3605));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_8 clkbuf_leaf_78_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_8 clkbuf_leaf_79_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_8 clkbuf_leaf_80_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_8 clkbuf_leaf_81_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_8 clkbuf_leaf_82_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_8 clkbuf_leaf_83_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_8 clkbuf_leaf_84_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_8 clkbuf_leaf_85_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_8 clkbuf_leaf_86_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_8 clkbuf_leaf_87_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_8 clkbuf_leaf_88_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_8 clkbuf_leaf_89_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_8 clkbuf_leaf_90_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_8 clkbuf_leaf_91_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_8 clkbuf_leaf_92_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_8 clkbuf_leaf_93_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_8 clkbuf_leaf_94_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_8 clkbuf_leaf_95_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_8 clkbuf_leaf_96_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_8 clkbuf_leaf_97_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_8 clkbuf_leaf_98_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_8 clkbuf_leaf_99_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_8 clkbuf_leaf_100_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_8 clkbuf_leaf_101_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_8 clkbuf_leaf_102_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_8 clkbuf_leaf_103_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_8 clkbuf_leaf_104_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_8 clkbuf_leaf_105_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_8 clkbuf_leaf_106_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_8 clkbuf_leaf_107_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_8 clkbuf_leaf_108_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_8 clkbuf_leaf_109_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_8 clkbuf_leaf_110_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_8 clkbuf_leaf_111_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_8 clkbuf_leaf_112_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_8 clkbuf_leaf_113_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_8 clkbuf_leaf_114_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_8 clkbuf_leaf_115_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_8 clkbuf_leaf_116_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_8 clkbuf_leaf_117_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_8 clkbuf_leaf_118_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_8 clkbuf_leaf_119_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_8 clkbuf_leaf_120_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_8 clkbuf_leaf_121_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_8 clkbuf_leaf_122_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_8 clkbuf_leaf_123_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_8 clkbuf_leaf_124_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_8 clkbuf_leaf_125_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_8 clkbuf_leaf_126_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_8 clkbuf_leaf_127_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_8 clkbuf_leaf_128_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_8 clkbuf_leaf_129_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_8 clkbuf_leaf_130_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_8 clkbuf_leaf_131_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_8 clkbuf_leaf_132_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_8 clkbuf_leaf_133_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_8 clkbuf_leaf_134_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_8 clkbuf_leaf_135_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_8 clkbuf_leaf_136_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_8 clkbuf_leaf_137_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_8 clkbuf_leaf_138_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_8 clkbuf_leaf_139_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_8 clkbuf_leaf_140_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_8 clkbuf_leaf_141_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_8 clkbuf_leaf_142_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_8 clkbuf_leaf_143_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_8 clkbuf_leaf_144_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_144_clk));
 sg13g2_buf_8 clkbuf_leaf_145_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_8 clkbuf_leaf_146_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_146_clk));
 sg13g2_buf_8 clkbuf_leaf_147_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_147_clk));
 sg13g2_buf_8 clkbuf_leaf_148_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_148_clk));
 sg13g2_buf_8 clkbuf_leaf_149_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_149_clk));
 sg13g2_buf_8 clkbuf_leaf_150_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_150_clk));
 sg13g2_buf_8 clkbuf_leaf_151_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_151_clk));
 sg13g2_buf_8 clkbuf_leaf_152_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_152_clk));
 sg13g2_buf_8 clkbuf_leaf_153_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_153_clk));
 sg13g2_buf_8 clkbuf_leaf_154_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_154_clk));
 sg13g2_buf_8 clkbuf_leaf_155_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_155_clk));
 sg13g2_buf_8 clkbuf_leaf_156_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_156_clk));
 sg13g2_buf_8 clkbuf_leaf_157_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_157_clk));
 sg13g2_buf_8 clkbuf_leaf_158_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_158_clk));
 sg13g2_buf_8 clkbuf_leaf_159_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_159_clk));
 sg13g2_buf_8 clkbuf_leaf_160_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_160_clk));
 sg13g2_buf_8 clkbuf_leaf_161_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_161_clk));
 sg13g2_buf_8 clkbuf_leaf_162_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_162_clk));
 sg13g2_buf_8 clkbuf_leaf_163_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_163_clk));
 sg13g2_buf_8 clkbuf_leaf_164_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_164_clk));
 sg13g2_buf_8 clkbuf_leaf_165_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_165_clk));
 sg13g2_buf_8 clkbuf_leaf_166_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_166_clk));
 sg13g2_buf_8 clkbuf_leaf_167_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_167_clk));
 sg13g2_buf_8 clkbuf_leaf_168_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_168_clk));
 sg13g2_buf_8 clkbuf_leaf_169_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_169_clk));
 sg13g2_buf_8 clkbuf_leaf_170_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_170_clk));
 sg13g2_buf_8 clkbuf_leaf_171_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_171_clk));
 sg13g2_buf_8 clkbuf_leaf_172_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_172_clk));
 sg13g2_buf_8 clkbuf_leaf_173_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_173_clk));
 sg13g2_buf_8 clkbuf_leaf_174_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_174_clk));
 sg13g2_buf_8 clkbuf_leaf_175_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_175_clk));
 sg13g2_buf_8 clkbuf_leaf_176_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_176_clk));
 sg13g2_buf_8 clkbuf_leaf_177_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_177_clk));
 sg13g2_buf_8 clkbuf_leaf_178_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_178_clk));
 sg13g2_buf_8 clkbuf_leaf_179_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_179_clk));
 sg13g2_buf_8 clkbuf_leaf_180_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_180_clk));
 sg13g2_buf_8 clkbuf_leaf_181_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_181_clk));
 sg13g2_buf_8 clkbuf_leaf_182_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_182_clk));
 sg13g2_buf_8 clkbuf_leaf_183_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_183_clk));
 sg13g2_buf_8 clkbuf_leaf_184_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_184_clk));
 sg13g2_buf_8 clkbuf_leaf_185_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_185_clk));
 sg13g2_buf_8 clkbuf_leaf_186_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_186_clk));
 sg13g2_buf_8 clkbuf_leaf_187_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_187_clk));
 sg13g2_buf_8 clkbuf_leaf_188_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_188_clk));
 sg13g2_buf_8 clkbuf_leaf_189_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_189_clk));
 sg13g2_buf_8 clkbuf_leaf_190_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_190_clk));
 sg13g2_buf_8 clkbuf_leaf_191_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_191_clk));
 sg13g2_buf_8 clkbuf_leaf_192_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_192_clk));
 sg13g2_buf_8 clkbuf_leaf_193_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_193_clk));
 sg13g2_buf_8 clkbuf_leaf_194_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_194_clk));
 sg13g2_buf_8 clkbuf_leaf_195_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_195_clk));
 sg13g2_buf_8 clkbuf_leaf_196_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_196_clk));
 sg13g2_buf_8 clkbuf_leaf_197_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_197_clk));
 sg13g2_buf_8 clkbuf_leaf_198_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_198_clk));
 sg13g2_buf_8 clkbuf_leaf_199_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_199_clk));
 sg13g2_buf_8 clkbuf_leaf_200_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_200_clk));
 sg13g2_buf_8 clkbuf_leaf_201_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_201_clk));
 sg13g2_buf_8 clkbuf_leaf_202_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_202_clk));
 sg13g2_buf_8 clkbuf_leaf_203_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_203_clk));
 sg13g2_buf_8 clkbuf_leaf_204_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_204_clk));
 sg13g2_buf_8 clkbuf_leaf_205_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_205_clk));
 sg13g2_buf_8 clkbuf_leaf_206_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_206_clk));
 sg13g2_buf_8 clkbuf_leaf_207_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_207_clk));
 sg13g2_buf_8 clkbuf_leaf_208_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_208_clk));
 sg13g2_buf_8 clkbuf_leaf_209_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_209_clk));
 sg13g2_buf_8 clkbuf_leaf_210_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_210_clk));
 sg13g2_buf_8 clkbuf_leaf_211_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_211_clk));
 sg13g2_buf_8 clkbuf_leaf_212_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_212_clk));
 sg13g2_buf_8 clkbuf_leaf_213_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_213_clk));
 sg13g2_buf_8 clkbuf_leaf_214_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_214_clk));
 sg13g2_buf_8 clkbuf_leaf_215_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_215_clk));
 sg13g2_buf_8 clkbuf_leaf_216_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_216_clk));
 sg13g2_buf_8 clkbuf_leaf_217_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_217_clk));
 sg13g2_buf_8 clkbuf_leaf_218_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_218_clk));
 sg13g2_buf_8 clkbuf_leaf_219_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_219_clk));
 sg13g2_buf_8 clkbuf_leaf_220_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_220_clk));
 sg13g2_buf_8 clkbuf_leaf_221_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_221_clk));
 sg13g2_buf_8 clkbuf_leaf_222_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_222_clk));
 sg13g2_buf_8 clkbuf_leaf_223_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_223_clk));
 sg13g2_buf_8 clkbuf_leaf_224_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_224_clk));
 sg13g2_buf_8 clkbuf_leaf_225_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_225_clk));
 sg13g2_buf_8 clkbuf_leaf_226_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_226_clk));
 sg13g2_buf_8 clkbuf_leaf_227_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_227_clk));
 sg13g2_buf_8 clkbuf_leaf_228_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_228_clk));
 sg13g2_buf_8 clkbuf_leaf_229_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_229_clk));
 sg13g2_buf_8 clkbuf_leaf_230_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_230_clk));
 sg13g2_buf_8 clkbuf_leaf_231_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_231_clk));
 sg13g2_buf_8 clkbuf_leaf_232_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_232_clk));
 sg13g2_buf_8 clkbuf_leaf_233_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_233_clk));
 sg13g2_buf_8 clkbuf_leaf_234_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_234_clk));
 sg13g2_buf_8 clkbuf_leaf_235_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_235_clk));
 sg13g2_buf_8 clkbuf_leaf_236_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_236_clk));
 sg13g2_buf_8 clkbuf_leaf_237_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_237_clk));
 sg13g2_buf_8 clkbuf_leaf_238_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_238_clk));
 sg13g2_buf_8 clkbuf_leaf_239_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_239_clk));
 sg13g2_buf_8 clkbuf_leaf_240_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_240_clk));
 sg13g2_buf_8 clkbuf_leaf_241_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_241_clk));
 sg13g2_buf_8 clkbuf_leaf_242_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_242_clk));
 sg13g2_buf_8 clkbuf_leaf_243_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_243_clk));
 sg13g2_buf_8 clkbuf_leaf_244_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_244_clk));
 sg13g2_buf_8 clkbuf_leaf_245_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_245_clk));
 sg13g2_buf_8 clkbuf_leaf_246_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_246_clk));
 sg13g2_buf_8 clkbuf_leaf_247_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_247_clk));
 sg13g2_buf_8 clkbuf_leaf_248_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_248_clk));
 sg13g2_buf_8 clkbuf_leaf_249_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_249_clk));
 sg13g2_buf_8 clkbuf_leaf_250_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_250_clk));
 sg13g2_buf_8 clkbuf_leaf_251_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_251_clk));
 sg13g2_buf_8 clkbuf_leaf_252_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_252_clk));
 sg13g2_buf_8 clkbuf_leaf_253_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_253_clk));
 sg13g2_buf_8 clkbuf_leaf_254_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_254_clk));
 sg13g2_buf_8 clkbuf_leaf_255_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_255_clk));
 sg13g2_buf_8 clkbuf_leaf_256_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_256_clk));
 sg13g2_buf_8 clkbuf_leaf_257_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_257_clk));
 sg13g2_buf_8 clkbuf_leaf_258_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_258_clk));
 sg13g2_buf_8 clkbuf_leaf_259_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_259_clk));
 sg13g2_buf_8 clkbuf_leaf_260_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_260_clk));
 sg13g2_buf_8 clkbuf_leaf_261_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_261_clk));
 sg13g2_buf_8 clkbuf_leaf_262_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_262_clk));
 sg13g2_buf_8 clkbuf_leaf_263_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_263_clk));
 sg13g2_buf_8 clkbuf_leaf_264_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_264_clk));
 sg13g2_buf_8 clkbuf_leaf_265_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_265_clk));
 sg13g2_buf_8 clkbuf_leaf_266_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_266_clk));
 sg13g2_buf_8 clkbuf_leaf_267_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_267_clk));
 sg13g2_buf_8 clkbuf_leaf_268_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_268_clk));
 sg13g2_buf_8 clkbuf_leaf_269_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_269_clk));
 sg13g2_buf_8 clkbuf_leaf_270_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_270_clk));
 sg13g2_buf_8 clkbuf_leaf_271_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_271_clk));
 sg13g2_buf_8 clkbuf_leaf_272_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_272_clk));
 sg13g2_buf_8 clkbuf_leaf_273_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_273_clk));
 sg13g2_buf_8 clkbuf_leaf_274_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_274_clk));
 sg13g2_buf_8 clkbuf_leaf_275_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_275_clk));
 sg13g2_buf_8 clkbuf_leaf_276_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_276_clk));
 sg13g2_buf_8 clkbuf_leaf_277_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_277_clk));
 sg13g2_buf_8 clkbuf_leaf_278_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_278_clk));
 sg13g2_buf_8 clkbuf_leaf_279_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_279_clk));
 sg13g2_buf_8 clkbuf_leaf_280_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_280_clk));
 sg13g2_buf_8 clkbuf_leaf_281_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_281_clk));
 sg13g2_buf_8 clkbuf_leaf_282_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_282_clk));
 sg13g2_buf_8 clkbuf_leaf_283_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_283_clk));
 sg13g2_buf_8 clkbuf_leaf_284_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_284_clk));
 sg13g2_buf_8 clkbuf_leaf_285_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_285_clk));
 sg13g2_buf_8 clkbuf_leaf_286_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_286_clk));
 sg13g2_buf_8 clkbuf_leaf_287_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_287_clk));
 sg13g2_buf_8 clkbuf_leaf_288_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_288_clk));
 sg13g2_buf_8 clkbuf_leaf_289_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_289_clk));
 sg13g2_buf_8 clkbuf_leaf_290_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_290_clk));
 sg13g2_buf_8 clkbuf_leaf_291_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_291_clk));
 sg13g2_buf_8 clkbuf_leaf_292_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_292_clk));
 sg13g2_buf_8 clkbuf_leaf_293_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_293_clk));
 sg13g2_buf_8 clkbuf_leaf_294_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_294_clk));
 sg13g2_buf_8 clkbuf_leaf_295_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_295_clk));
 sg13g2_buf_8 clkbuf_leaf_296_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_296_clk));
 sg13g2_buf_8 clkbuf_leaf_297_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_297_clk));
 sg13g2_buf_8 clkbuf_leaf_298_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_298_clk));
 sg13g2_buf_8 clkbuf_leaf_299_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_299_clk));
 sg13g2_buf_8 clkbuf_leaf_300_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_300_clk));
 sg13g2_buf_8 clkbuf_leaf_301_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_301_clk));
 sg13g2_buf_8 clkbuf_leaf_302_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_302_clk));
 sg13g2_buf_8 clkbuf_leaf_303_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_303_clk));
 sg13g2_buf_8 clkbuf_leaf_304_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_304_clk));
 sg13g2_buf_8 clkbuf_leaf_305_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_305_clk));
 sg13g2_buf_8 clkbuf_leaf_306_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_306_clk));
 sg13g2_buf_8 clkbuf_leaf_307_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_307_clk));
 sg13g2_buf_8 clkbuf_leaf_308_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_308_clk));
 sg13g2_buf_8 clkbuf_leaf_309_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_309_clk));
 sg13g2_buf_8 clkbuf_leaf_310_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_310_clk));
 sg13g2_buf_8 clkbuf_leaf_311_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_311_clk));
 sg13g2_buf_8 clkbuf_leaf_312_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_312_clk));
 sg13g2_buf_8 clkbuf_leaf_313_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_313_clk));
 sg13g2_buf_4 clkbuf_0_clk (.X(clknet_0_clk),
    .A(clk));
 sg13g2_buf_8 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sg13g2_buf_8 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sg13g2_buf_8 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sg13g2_buf_8 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sg13g2_buf_8 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sg13g2_buf_8 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sg13g2_buf_8 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sg13g2_buf_8 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_0__f_clk (.X(clknet_6_0__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_1__f_clk (.X(clknet_6_1__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_2__f_clk (.X(clknet_6_2__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_3__f_clk (.X(clknet_6_3__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_4__f_clk (.X(clknet_6_4__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_5__f_clk (.X(clknet_6_5__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_6__f_clk (.X(clknet_6_6__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_7__f_clk (.X(clknet_6_7__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_8__f_clk (.X(clknet_6_8__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_9__f_clk (.X(clknet_6_9__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_10__f_clk (.X(clknet_6_10__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_11__f_clk (.X(clknet_6_11__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_12__f_clk (.X(clknet_6_12__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_13__f_clk (.X(clknet_6_13__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_14__f_clk (.X(clknet_6_14__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_15__f_clk (.X(clknet_6_15__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_16__f_clk (.X(clknet_6_16__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_17__f_clk (.X(clknet_6_17__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_18__f_clk (.X(clknet_6_18__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_19__f_clk (.X(clknet_6_19__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_20__f_clk (.X(clknet_6_20__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_21__f_clk (.X(clknet_6_21__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_22__f_clk (.X(clknet_6_22__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_23__f_clk (.X(clknet_6_23__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_24__f_clk (.X(clknet_6_24__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_25__f_clk (.X(clknet_6_25__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_26__f_clk (.X(clknet_6_26__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_27__f_clk (.X(clknet_6_27__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_28__f_clk (.X(clknet_6_28__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_29__f_clk (.X(clknet_6_29__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_30__f_clk (.X(clknet_6_30__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_31__f_clk (.X(clknet_6_31__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_32__f_clk (.X(clknet_6_32__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_33__f_clk (.X(clknet_6_33__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_34__f_clk (.X(clknet_6_34__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_35__f_clk (.X(clknet_6_35__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_36__f_clk (.X(clknet_6_36__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_37__f_clk (.X(clknet_6_37__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_38__f_clk (.X(clknet_6_38__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_39__f_clk (.X(clknet_6_39__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_40__f_clk (.X(clknet_6_40__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_41__f_clk (.X(clknet_6_41__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_42__f_clk (.X(clknet_6_42__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_43__f_clk (.X(clknet_6_43__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_44__f_clk (.X(clknet_6_44__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_45__f_clk (.X(clknet_6_45__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_46__f_clk (.X(clknet_6_46__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_47__f_clk (.X(clknet_6_47__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_48__f_clk (.X(clknet_6_48__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_49__f_clk (.X(clknet_6_49__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_50__f_clk (.X(clknet_6_50__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_51__f_clk (.X(clknet_6_51__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_52__f_clk (.X(clknet_6_52__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_53__f_clk (.X(clknet_6_53__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_54__f_clk (.X(clknet_6_54__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_55__f_clk (.X(clknet_6_55__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_56__f_clk (.X(clknet_6_56__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_57__f_clk (.X(clknet_6_57__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_58__f_clk (.X(clknet_6_58__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_59__f_clk (.X(clknet_6_59__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_60__f_clk (.X(clknet_6_60__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_61__f_clk (.X(clknet_6_61__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_62__f_clk (.X(clknet_6_62__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_63__f_clk (.X(clknet_6_63__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_6_15__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_6_23__leaf_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_6_31__leaf_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_6_47__leaf_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_6_55__leaf_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_6_63__leaf_clk));
 sg13g2_buf_8 clkload6 (.A(clknet_leaf_313_clk));
 sg13g2_buf_8 clkload7 (.A(clknet_leaf_106_clk));
 sg13g2_inv_4 clkload8 (.A(clknet_leaf_97_clk));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_253_clk));
 sg13g2_buf_16 clkload10 (.A(clknet_leaf_260_clk));
 sg13g2_inv_2 clkload11 (.A(clknet_leaf_175_clk));
 sg13g2_buf_16 clkload12 (.A(clknet_leaf_114_clk));
 sg13g2_inv_2 clkload13 (.A(clknet_leaf_112_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_00054_));
 sg13g2_antennanp ANTENNA_2 (.A(_00054_));
 sg13g2_antennanp ANTENNA_3 (.A(_00201_));
 sg13g2_antennanp ANTENNA_4 (.A(_00207_));
 sg13g2_antennanp ANTENNA_5 (.A(_00235_));
 sg13g2_antennanp ANTENNA_6 (.A(_00769_));
 sg13g2_antennanp ANTENNA_7 (.A(_00905_));
 sg13g2_antennanp ANTENNA_8 (.A(_00923_));
 sg13g2_antennanp ANTENNA_9 (.A(_00923_));
 sg13g2_antennanp ANTENNA_10 (.A(_00964_));
 sg13g2_antennanp ANTENNA_11 (.A(_00964_));
 sg13g2_antennanp ANTENNA_12 (.A(_01012_));
 sg13g2_antennanp ANTENNA_13 (.A(_01012_));
 sg13g2_antennanp ANTENNA_14 (.A(_01048_));
 sg13g2_antennanp ANTENNA_15 (.A(_02918_));
 sg13g2_antennanp ANTENNA_16 (.A(_02918_));
 sg13g2_antennanp ANTENNA_17 (.A(_02918_));
 sg13g2_antennanp ANTENNA_18 (.A(_02918_));
 sg13g2_antennanp ANTENNA_19 (.A(_02918_));
 sg13g2_antennanp ANTENNA_20 (.A(_02918_));
 sg13g2_antennanp ANTENNA_21 (.A(_02918_));
 sg13g2_antennanp ANTENNA_22 (.A(_02918_));
 sg13g2_antennanp ANTENNA_23 (.A(_02918_));
 sg13g2_antennanp ANTENNA_24 (.A(_02963_));
 sg13g2_antennanp ANTENNA_25 (.A(_02963_));
 sg13g2_antennanp ANTENNA_26 (.A(_02963_));
 sg13g2_antennanp ANTENNA_27 (.A(_02963_));
 sg13g2_antennanp ANTENNA_28 (.A(_02963_));
 sg13g2_antennanp ANTENNA_29 (.A(_02963_));
 sg13g2_antennanp ANTENNA_30 (.A(_03057_));
 sg13g2_antennanp ANTENNA_31 (.A(_03057_));
 sg13g2_antennanp ANTENNA_32 (.A(_03057_));
 sg13g2_antennanp ANTENNA_33 (.A(_03093_));
 sg13g2_antennanp ANTENNA_34 (.A(_03093_));
 sg13g2_antennanp ANTENNA_35 (.A(_03093_));
 sg13g2_antennanp ANTENNA_36 (.A(_03093_));
 sg13g2_antennanp ANTENNA_37 (.A(_03093_));
 sg13g2_antennanp ANTENNA_38 (.A(_03093_));
 sg13g2_antennanp ANTENNA_39 (.A(_03093_));
 sg13g2_antennanp ANTENNA_40 (.A(_03093_));
 sg13g2_antennanp ANTENNA_41 (.A(_03093_));
 sg13g2_antennanp ANTENNA_42 (.A(_03093_));
 sg13g2_antennanp ANTENNA_43 (.A(_03096_));
 sg13g2_antennanp ANTENNA_44 (.A(_03096_));
 sg13g2_antennanp ANTENNA_45 (.A(_03096_));
 sg13g2_antennanp ANTENNA_46 (.A(_03096_));
 sg13g2_antennanp ANTENNA_47 (.A(_03096_));
 sg13g2_antennanp ANTENNA_48 (.A(_03096_));
 sg13g2_antennanp ANTENNA_49 (.A(_03096_));
 sg13g2_antennanp ANTENNA_50 (.A(_03096_));
 sg13g2_antennanp ANTENNA_51 (.A(_03096_));
 sg13g2_antennanp ANTENNA_52 (.A(_03096_));
 sg13g2_antennanp ANTENNA_53 (.A(_03107_));
 sg13g2_antennanp ANTENNA_54 (.A(_03107_));
 sg13g2_antennanp ANTENNA_55 (.A(_03107_));
 sg13g2_antennanp ANTENNA_56 (.A(_03107_));
 sg13g2_antennanp ANTENNA_57 (.A(_03107_));
 sg13g2_antennanp ANTENNA_58 (.A(_03108_));
 sg13g2_antennanp ANTENNA_59 (.A(_03108_));
 sg13g2_antennanp ANTENNA_60 (.A(_03108_));
 sg13g2_antennanp ANTENNA_61 (.A(_03108_));
 sg13g2_antennanp ANTENNA_62 (.A(_03108_));
 sg13g2_antennanp ANTENNA_63 (.A(_03108_));
 sg13g2_antennanp ANTENNA_64 (.A(_03108_));
 sg13g2_antennanp ANTENNA_65 (.A(_03108_));
 sg13g2_antennanp ANTENNA_66 (.A(_03108_));
 sg13g2_antennanp ANTENNA_67 (.A(_03109_));
 sg13g2_antennanp ANTENNA_68 (.A(_03109_));
 sg13g2_antennanp ANTENNA_69 (.A(_03109_));
 sg13g2_antennanp ANTENNA_70 (.A(_03133_));
 sg13g2_antennanp ANTENNA_71 (.A(_03133_));
 sg13g2_antennanp ANTENNA_72 (.A(_03133_));
 sg13g2_antennanp ANTENNA_73 (.A(_03133_));
 sg13g2_antennanp ANTENNA_74 (.A(_03137_));
 sg13g2_antennanp ANTENNA_75 (.A(_03137_));
 sg13g2_antennanp ANTENNA_76 (.A(_03137_));
 sg13g2_antennanp ANTENNA_77 (.A(_03137_));
 sg13g2_antennanp ANTENNA_78 (.A(_03137_));
 sg13g2_antennanp ANTENNA_79 (.A(_03212_));
 sg13g2_antennanp ANTENNA_80 (.A(_03229_));
 sg13g2_antennanp ANTENNA_81 (.A(_03642_));
 sg13g2_antennanp ANTENNA_82 (.A(_03642_));
 sg13g2_antennanp ANTENNA_83 (.A(_03642_));
 sg13g2_antennanp ANTENNA_84 (.A(_03647_));
 sg13g2_antennanp ANTENNA_85 (.A(_03647_));
 sg13g2_antennanp ANTENNA_86 (.A(_03647_));
 sg13g2_antennanp ANTENNA_87 (.A(_03647_));
 sg13g2_antennanp ANTENNA_88 (.A(_03653_));
 sg13g2_antennanp ANTENNA_89 (.A(_03653_));
 sg13g2_antennanp ANTENNA_90 (.A(_03653_));
 sg13g2_antennanp ANTENNA_91 (.A(_03653_));
 sg13g2_antennanp ANTENNA_92 (.A(_03653_));
 sg13g2_antennanp ANTENNA_93 (.A(_03653_));
 sg13g2_antennanp ANTENNA_94 (.A(_03653_));
 sg13g2_antennanp ANTENNA_95 (.A(_03653_));
 sg13g2_antennanp ANTENNA_96 (.A(_03653_));
 sg13g2_antennanp ANTENNA_97 (.A(_03656_));
 sg13g2_antennanp ANTENNA_98 (.A(_03656_));
 sg13g2_antennanp ANTENNA_99 (.A(_03656_));
 sg13g2_antennanp ANTENNA_100 (.A(_03657_));
 sg13g2_antennanp ANTENNA_101 (.A(_03657_));
 sg13g2_antennanp ANTENNA_102 (.A(_03657_));
 sg13g2_antennanp ANTENNA_103 (.A(_03657_));
 sg13g2_antennanp ANTENNA_104 (.A(_03657_));
 sg13g2_antennanp ANTENNA_105 (.A(_03657_));
 sg13g2_antennanp ANTENNA_106 (.A(_03657_));
 sg13g2_antennanp ANTENNA_107 (.A(_03657_));
 sg13g2_antennanp ANTENNA_108 (.A(_03657_));
 sg13g2_antennanp ANTENNA_109 (.A(_04770_));
 sg13g2_antennanp ANTENNA_110 (.A(_04770_));
 sg13g2_antennanp ANTENNA_111 (.A(_04770_));
 sg13g2_antennanp ANTENNA_112 (.A(_04770_));
 sg13g2_antennanp ANTENNA_113 (.A(_04771_));
 sg13g2_antennanp ANTENNA_114 (.A(_04771_));
 sg13g2_antennanp ANTENNA_115 (.A(_04771_));
 sg13g2_antennanp ANTENNA_116 (.A(_04771_));
 sg13g2_antennanp ANTENNA_117 (.A(_04848_));
 sg13g2_antennanp ANTENNA_118 (.A(_04848_));
 sg13g2_antennanp ANTENNA_119 (.A(_05001_));
 sg13g2_antennanp ANTENNA_120 (.A(_05431_));
 sg13g2_antennanp ANTENNA_121 (.A(_05642_));
 sg13g2_antennanp ANTENNA_122 (.A(_05735_));
 sg13g2_antennanp ANTENNA_123 (.A(_05753_));
 sg13g2_antennanp ANTENNA_124 (.A(_05753_));
 sg13g2_antennanp ANTENNA_125 (.A(_05753_));
 sg13g2_antennanp ANTENNA_126 (.A(_05753_));
 sg13g2_antennanp ANTENNA_127 (.A(_05754_));
 sg13g2_antennanp ANTENNA_128 (.A(_05754_));
 sg13g2_antennanp ANTENNA_129 (.A(_05754_));
 sg13g2_antennanp ANTENNA_130 (.A(_05754_));
 sg13g2_antennanp ANTENNA_131 (.A(_05766_));
 sg13g2_antennanp ANTENNA_132 (.A(_05771_));
 sg13g2_antennanp ANTENNA_133 (.A(_05773_));
 sg13g2_antennanp ANTENNA_134 (.A(_05778_));
 sg13g2_antennanp ANTENNA_135 (.A(_05782_));
 sg13g2_antennanp ANTENNA_136 (.A(_05782_));
 sg13g2_antennanp ANTENNA_137 (.A(_05782_));
 sg13g2_antennanp ANTENNA_138 (.A(_05782_));
 sg13g2_antennanp ANTENNA_139 (.A(_05786_));
 sg13g2_antennanp ANTENNA_140 (.A(_05791_));
 sg13g2_antennanp ANTENNA_141 (.A(_06092_));
 sg13g2_antennanp ANTENNA_142 (.A(_06092_));
 sg13g2_antennanp ANTENNA_143 (.A(_06092_));
 sg13g2_antennanp ANTENNA_144 (.A(_06092_));
 sg13g2_antennanp ANTENNA_145 (.A(_06092_));
 sg13g2_antennanp ANTENNA_146 (.A(_06137_));
 sg13g2_antennanp ANTENNA_147 (.A(_06137_));
 sg13g2_antennanp ANTENNA_148 (.A(_06137_));
 sg13g2_antennanp ANTENNA_149 (.A(_06137_));
 sg13g2_antennanp ANTENNA_150 (.A(_06137_));
 sg13g2_antennanp ANTENNA_151 (.A(_06137_));
 sg13g2_antennanp ANTENNA_152 (.A(_06304_));
 sg13g2_antennanp ANTENNA_153 (.A(_06304_));
 sg13g2_antennanp ANTENNA_154 (.A(_06304_));
 sg13g2_antennanp ANTENNA_155 (.A(_06304_));
 sg13g2_antennanp ANTENNA_156 (.A(_06386_));
 sg13g2_antennanp ANTENNA_157 (.A(_06386_));
 sg13g2_antennanp ANTENNA_158 (.A(_06386_));
 sg13g2_antennanp ANTENNA_159 (.A(_06386_));
 sg13g2_antennanp ANTENNA_160 (.A(_06386_));
 sg13g2_antennanp ANTENNA_161 (.A(_06386_));
 sg13g2_antennanp ANTENNA_162 (.A(_06386_));
 sg13g2_antennanp ANTENNA_163 (.A(_06386_));
 sg13g2_antennanp ANTENNA_164 (.A(_06386_));
 sg13g2_antennanp ANTENNA_165 (.A(_07450_));
 sg13g2_antennanp ANTENNA_166 (.A(_07450_));
 sg13g2_antennanp ANTENNA_167 (.A(_07450_));
 sg13g2_antennanp ANTENNA_168 (.A(_07729_));
 sg13g2_antennanp ANTENNA_169 (.A(_07729_));
 sg13g2_antennanp ANTENNA_170 (.A(_07729_));
 sg13g2_antennanp ANTENNA_171 (.A(_07729_));
 sg13g2_antennanp ANTENNA_172 (.A(_07729_));
 sg13g2_antennanp ANTENNA_173 (.A(_07729_));
 sg13g2_antennanp ANTENNA_174 (.A(_07729_));
 sg13g2_antennanp ANTENNA_175 (.A(_07729_));
 sg13g2_antennanp ANTENNA_176 (.A(_07729_));
 sg13g2_antennanp ANTENNA_177 (.A(_08126_));
 sg13g2_antennanp ANTENNA_178 (.A(_08126_));
 sg13g2_antennanp ANTENNA_179 (.A(_08126_));
 sg13g2_antennanp ANTENNA_180 (.A(_08126_));
 sg13g2_antennanp ANTENNA_181 (.A(_08133_));
 sg13g2_antennanp ANTENNA_182 (.A(_08133_));
 sg13g2_antennanp ANTENNA_183 (.A(_08133_));
 sg13g2_antennanp ANTENNA_184 (.A(_08133_));
 sg13g2_antennanp ANTENNA_185 (.A(_08133_));
 sg13g2_antennanp ANTENNA_186 (.A(_08133_));
 sg13g2_antennanp ANTENNA_187 (.A(_08181_));
 sg13g2_antennanp ANTENNA_188 (.A(_08181_));
 sg13g2_antennanp ANTENNA_189 (.A(_08181_));
 sg13g2_antennanp ANTENNA_190 (.A(_08181_));
 sg13g2_antennanp ANTENNA_191 (.A(_08181_));
 sg13g2_antennanp ANTENNA_192 (.A(_08181_));
 sg13g2_antennanp ANTENNA_193 (.A(_08181_));
 sg13g2_antennanp ANTENNA_194 (.A(_08190_));
 sg13g2_antennanp ANTENNA_195 (.A(_08190_));
 sg13g2_antennanp ANTENNA_196 (.A(_08190_));
 sg13g2_antennanp ANTENNA_197 (.A(_08190_));
 sg13g2_antennanp ANTENNA_198 (.A(_08190_));
 sg13g2_antennanp ANTENNA_199 (.A(_08190_));
 sg13g2_antennanp ANTENNA_200 (.A(_08190_));
 sg13g2_antennanp ANTENNA_201 (.A(_08190_));
 sg13g2_antennanp ANTENNA_202 (.A(_08192_));
 sg13g2_antennanp ANTENNA_203 (.A(_08273_));
 sg13g2_antennanp ANTENNA_204 (.A(_08273_));
 sg13g2_antennanp ANTENNA_205 (.A(_08273_));
 sg13g2_antennanp ANTENNA_206 (.A(_08273_));
 sg13g2_antennanp ANTENNA_207 (.A(_08285_));
 sg13g2_antennanp ANTENNA_208 (.A(_08285_));
 sg13g2_antennanp ANTENNA_209 (.A(_08285_));
 sg13g2_antennanp ANTENNA_210 (.A(_08285_));
 sg13g2_antennanp ANTENNA_211 (.A(_08285_));
 sg13g2_antennanp ANTENNA_212 (.A(_08285_));
 sg13g2_antennanp ANTENNA_213 (.A(_08302_));
 sg13g2_antennanp ANTENNA_214 (.A(_08302_));
 sg13g2_antennanp ANTENNA_215 (.A(_08302_));
 sg13g2_antennanp ANTENNA_216 (.A(_08302_));
 sg13g2_antennanp ANTENNA_217 (.A(_08302_));
 sg13g2_antennanp ANTENNA_218 (.A(_08302_));
 sg13g2_antennanp ANTENNA_219 (.A(_08356_));
 sg13g2_antennanp ANTENNA_220 (.A(_08356_));
 sg13g2_antennanp ANTENNA_221 (.A(_08356_));
 sg13g2_antennanp ANTENNA_222 (.A(_08356_));
 sg13g2_antennanp ANTENNA_223 (.A(_08356_));
 sg13g2_antennanp ANTENNA_224 (.A(_08356_));
 sg13g2_antennanp ANTENNA_225 (.A(_08356_));
 sg13g2_antennanp ANTENNA_226 (.A(_08356_));
 sg13g2_antennanp ANTENNA_227 (.A(_08356_));
 sg13g2_antennanp ANTENNA_228 (.A(_08447_));
 sg13g2_antennanp ANTENNA_229 (.A(_08447_));
 sg13g2_antennanp ANTENNA_230 (.A(_08447_));
 sg13g2_antennanp ANTENNA_231 (.A(_08473_));
 sg13g2_antennanp ANTENNA_232 (.A(_08473_));
 sg13g2_antennanp ANTENNA_233 (.A(_08473_));
 sg13g2_antennanp ANTENNA_234 (.A(_08494_));
 sg13g2_antennanp ANTENNA_235 (.A(_08494_));
 sg13g2_antennanp ANTENNA_236 (.A(_08494_));
 sg13g2_antennanp ANTENNA_237 (.A(_08557_));
 sg13g2_antennanp ANTENNA_238 (.A(_08557_));
 sg13g2_antennanp ANTENNA_239 (.A(_08557_));
 sg13g2_antennanp ANTENNA_240 (.A(_08705_));
 sg13g2_antennanp ANTENNA_241 (.A(_08705_));
 sg13g2_antennanp ANTENNA_242 (.A(_08705_));
 sg13g2_antennanp ANTENNA_243 (.A(_08708_));
 sg13g2_antennanp ANTENNA_244 (.A(_08708_));
 sg13g2_antennanp ANTENNA_245 (.A(_08708_));
 sg13g2_antennanp ANTENNA_246 (.A(_08709_));
 sg13g2_antennanp ANTENNA_247 (.A(_08709_));
 sg13g2_antennanp ANTENNA_248 (.A(_08709_));
 sg13g2_antennanp ANTENNA_249 (.A(_08709_));
 sg13g2_antennanp ANTENNA_250 (.A(_08801_));
 sg13g2_antennanp ANTENNA_251 (.A(_08801_));
 sg13g2_antennanp ANTENNA_252 (.A(_08964_));
 sg13g2_antennanp ANTENNA_253 (.A(_08964_));
 sg13g2_antennanp ANTENNA_254 (.A(_08964_));
 sg13g2_antennanp ANTENNA_255 (.A(_08964_));
 sg13g2_antennanp ANTENNA_256 (.A(_08979_));
 sg13g2_antennanp ANTENNA_257 (.A(_08979_));
 sg13g2_antennanp ANTENNA_258 (.A(_08979_));
 sg13g2_antennanp ANTENNA_259 (.A(_08979_));
 sg13g2_antennanp ANTENNA_260 (.A(_08979_));
 sg13g2_antennanp ANTENNA_261 (.A(_09008_));
 sg13g2_antennanp ANTENNA_262 (.A(_09008_));
 sg13g2_antennanp ANTENNA_263 (.A(_09008_));
 sg13g2_antennanp ANTENNA_264 (.A(_09008_));
 sg13g2_antennanp ANTENNA_265 (.A(_09008_));
 sg13g2_antennanp ANTENNA_266 (.A(_09008_));
 sg13g2_antennanp ANTENNA_267 (.A(_09022_));
 sg13g2_antennanp ANTENNA_268 (.A(_09022_));
 sg13g2_antennanp ANTENNA_269 (.A(_09022_));
 sg13g2_antennanp ANTENNA_270 (.A(_09025_));
 sg13g2_antennanp ANTENNA_271 (.A(_09025_));
 sg13g2_antennanp ANTENNA_272 (.A(_09025_));
 sg13g2_antennanp ANTENNA_273 (.A(_09025_));
 sg13g2_antennanp ANTENNA_274 (.A(_09025_));
 sg13g2_antennanp ANTENNA_275 (.A(_09025_));
 sg13g2_antennanp ANTENNA_276 (.A(_09025_));
 sg13g2_antennanp ANTENNA_277 (.A(_09025_));
 sg13g2_antennanp ANTENNA_278 (.A(_09025_));
 sg13g2_antennanp ANTENNA_279 (.A(_09026_));
 sg13g2_antennanp ANTENNA_280 (.A(_09026_));
 sg13g2_antennanp ANTENNA_281 (.A(_09026_));
 sg13g2_antennanp ANTENNA_282 (.A(_09026_));
 sg13g2_antennanp ANTENNA_283 (.A(_09026_));
 sg13g2_antennanp ANTENNA_284 (.A(_09026_));
 sg13g2_antennanp ANTENNA_285 (.A(_09026_));
 sg13g2_antennanp ANTENNA_286 (.A(_09026_));
 sg13g2_antennanp ANTENNA_287 (.A(_09026_));
 sg13g2_antennanp ANTENNA_288 (.A(_09045_));
 sg13g2_antennanp ANTENNA_289 (.A(_09050_));
 sg13g2_antennanp ANTENNA_290 (.A(_09050_));
 sg13g2_antennanp ANTENNA_291 (.A(_09050_));
 sg13g2_antennanp ANTENNA_292 (.A(_09052_));
 sg13g2_antennanp ANTENNA_293 (.A(_09052_));
 sg13g2_antennanp ANTENNA_294 (.A(_09052_));
 sg13g2_antennanp ANTENNA_295 (.A(_09052_));
 sg13g2_antennanp ANTENNA_296 (.A(_09118_));
 sg13g2_antennanp ANTENNA_297 (.A(_09118_));
 sg13g2_antennanp ANTENNA_298 (.A(_09118_));
 sg13g2_antennanp ANTENNA_299 (.A(_09118_));
 sg13g2_antennanp ANTENNA_300 (.A(_09122_));
 sg13g2_antennanp ANTENNA_301 (.A(_09122_));
 sg13g2_antennanp ANTENNA_302 (.A(_09122_));
 sg13g2_antennanp ANTENNA_303 (.A(_09124_));
 sg13g2_antennanp ANTENNA_304 (.A(_09124_));
 sg13g2_antennanp ANTENNA_305 (.A(_09124_));
 sg13g2_antennanp ANTENNA_306 (.A(_09124_));
 sg13g2_antennanp ANTENNA_307 (.A(_09124_));
 sg13g2_antennanp ANTENNA_308 (.A(_09124_));
 sg13g2_antennanp ANTENNA_309 (.A(_09124_));
 sg13g2_antennanp ANTENNA_310 (.A(_09124_));
 sg13g2_antennanp ANTENNA_311 (.A(_09124_));
 sg13g2_antennanp ANTENNA_312 (.A(_09124_));
 sg13g2_antennanp ANTENNA_313 (.A(_09166_));
 sg13g2_antennanp ANTENNA_314 (.A(_09166_));
 sg13g2_antennanp ANTENNA_315 (.A(_09166_));
 sg13g2_antennanp ANTENNA_316 (.A(_09166_));
 sg13g2_antennanp ANTENNA_317 (.A(_09207_));
 sg13g2_antennanp ANTENNA_318 (.A(_09251_));
 sg13g2_antennanp ANTENNA_319 (.A(_09273_));
 sg13g2_antennanp ANTENNA_320 (.A(_09273_));
 sg13g2_antennanp ANTENNA_321 (.A(_09273_));
 sg13g2_antennanp ANTENNA_322 (.A(_09273_));
 sg13g2_antennanp ANTENNA_323 (.A(_09273_));
 sg13g2_antennanp ANTENNA_324 (.A(_09273_));
 sg13g2_antennanp ANTENNA_325 (.A(_09273_));
 sg13g2_antennanp ANTENNA_326 (.A(_09273_));
 sg13g2_antennanp ANTENNA_327 (.A(_09293_));
 sg13g2_antennanp ANTENNA_328 (.A(_09328_));
 sg13g2_antennanp ANTENNA_329 (.A(_09340_));
 sg13g2_antennanp ANTENNA_330 (.A(_09340_));
 sg13g2_antennanp ANTENNA_331 (.A(_09340_));
 sg13g2_antennanp ANTENNA_332 (.A(_09361_));
 sg13g2_antennanp ANTENNA_333 (.A(_09361_));
 sg13g2_antennanp ANTENNA_334 (.A(_09398_));
 sg13g2_antennanp ANTENNA_335 (.A(_09417_));
 sg13g2_antennanp ANTENNA_336 (.A(_09417_));
 sg13g2_antennanp ANTENNA_337 (.A(_09417_));
 sg13g2_antennanp ANTENNA_338 (.A(_09417_));
 sg13g2_antennanp ANTENNA_339 (.A(_09445_));
 sg13g2_antennanp ANTENNA_340 (.A(_09445_));
 sg13g2_antennanp ANTENNA_341 (.A(_09485_));
 sg13g2_antennanp ANTENNA_342 (.A(_09499_));
 sg13g2_antennanp ANTENNA_343 (.A(_09501_));
 sg13g2_antennanp ANTENNA_344 (.A(_09606_));
 sg13g2_antennanp ANTENNA_345 (.A(_09606_));
 sg13g2_antennanp ANTENNA_346 (.A(_09637_));
 sg13g2_antennanp ANTENNA_347 (.A(_09875_));
 sg13g2_antennanp ANTENNA_348 (.A(_09875_));
 sg13g2_antennanp ANTENNA_349 (.A(_09875_));
 sg13g2_antennanp ANTENNA_350 (.A(_09875_));
 sg13g2_antennanp ANTENNA_351 (.A(_09875_));
 sg13g2_antennanp ANTENNA_352 (.A(_09875_));
 sg13g2_antennanp ANTENNA_353 (.A(_09875_));
 sg13g2_antennanp ANTENNA_354 (.A(_09875_));
 sg13g2_antennanp ANTENNA_355 (.A(_09875_));
 sg13g2_antennanp ANTENNA_356 (.A(_09927_));
 sg13g2_antennanp ANTENNA_357 (.A(_09927_));
 sg13g2_antennanp ANTENNA_358 (.A(_09927_));
 sg13g2_antennanp ANTENNA_359 (.A(_09991_));
 sg13g2_antennanp ANTENNA_360 (.A(_09991_));
 sg13g2_antennanp ANTENNA_361 (.A(_09991_));
 sg13g2_antennanp ANTENNA_362 (.A(_09991_));
 sg13g2_antennanp ANTENNA_363 (.A(_09991_));
 sg13g2_antennanp ANTENNA_364 (.A(_09991_));
 sg13g2_antennanp ANTENNA_365 (.A(_09991_));
 sg13g2_antennanp ANTENNA_366 (.A(_09991_));
 sg13g2_antennanp ANTENNA_367 (.A(_09991_));
 sg13g2_antennanp ANTENNA_368 (.A(_09991_));
 sg13g2_antennanp ANTENNA_369 (.A(_09991_));
 sg13g2_antennanp ANTENNA_370 (.A(_09991_));
 sg13g2_antennanp ANTENNA_371 (.A(_09991_));
 sg13g2_antennanp ANTENNA_372 (.A(_10110_));
 sg13g2_antennanp ANTENNA_373 (.A(_10423_));
 sg13g2_antennanp ANTENNA_374 (.A(_10423_));
 sg13g2_antennanp ANTENNA_375 (.A(_10423_));
 sg13g2_antennanp ANTENNA_376 (.A(_10423_));
 sg13g2_antennanp ANTENNA_377 (.A(_10831_));
 sg13g2_antennanp ANTENNA_378 (.A(_10831_));
 sg13g2_antennanp ANTENNA_379 (.A(_10831_));
 sg13g2_antennanp ANTENNA_380 (.A(_10831_));
 sg13g2_antennanp ANTENNA_381 (.A(_10831_));
 sg13g2_antennanp ANTENNA_382 (.A(_10831_));
 sg13g2_antennanp ANTENNA_383 (.A(_10831_));
 sg13g2_antennanp ANTENNA_384 (.A(_10831_));
 sg13g2_antennanp ANTENNA_385 (.A(_10831_));
 sg13g2_antennanp ANTENNA_386 (.A(_10831_));
 sg13g2_antennanp ANTENNA_387 (.A(_10831_));
 sg13g2_antennanp ANTENNA_388 (.A(_10831_));
 sg13g2_antennanp ANTENNA_389 (.A(_10831_));
 sg13g2_antennanp ANTENNA_390 (.A(_10831_));
 sg13g2_antennanp ANTENNA_391 (.A(_10831_));
 sg13g2_antennanp ANTENNA_392 (.A(_10831_));
 sg13g2_antennanp ANTENNA_393 (.A(_10831_));
 sg13g2_antennanp ANTENNA_394 (.A(_10831_));
 sg13g2_antennanp ANTENNA_395 (.A(_10831_));
 sg13g2_antennanp ANTENNA_396 (.A(_10831_));
 sg13g2_antennanp ANTENNA_397 (.A(_10831_));
 sg13g2_antennanp ANTENNA_398 (.A(_10831_));
 sg13g2_antennanp ANTENNA_399 (.A(_10831_));
 sg13g2_antennanp ANTENNA_400 (.A(_10963_));
 sg13g2_antennanp ANTENNA_401 (.A(_10963_));
 sg13g2_antennanp ANTENNA_402 (.A(_10963_));
 sg13g2_antennanp ANTENNA_403 (.A(_10963_));
 sg13g2_antennanp ANTENNA_404 (.A(_10963_));
 sg13g2_antennanp ANTENNA_405 (.A(_10963_));
 sg13g2_antennanp ANTENNA_406 (.A(_11495_));
 sg13g2_antennanp ANTENNA_407 (.A(_11495_));
 sg13g2_antennanp ANTENNA_408 (.A(_11495_));
 sg13g2_antennanp ANTENNA_409 (.A(_11495_));
 sg13g2_antennanp ANTENNA_410 (.A(_11495_));
 sg13g2_antennanp ANTENNA_411 (.A(_11900_));
 sg13g2_antennanp ANTENNA_412 (.A(_11900_));
 sg13g2_antennanp ANTENNA_413 (.A(_11900_));
 sg13g2_antennanp ANTENNA_414 (.A(_11900_));
 sg13g2_antennanp ANTENNA_415 (.A(_11988_));
 sg13g2_antennanp ANTENNA_416 (.A(_11988_));
 sg13g2_antennanp ANTENNA_417 (.A(_11988_));
 sg13g2_antennanp ANTENNA_418 (.A(_11988_));
 sg13g2_antennanp ANTENNA_419 (.A(_11988_));
 sg13g2_antennanp ANTENNA_420 (.A(_11988_));
 sg13g2_antennanp ANTENNA_421 (.A(_11988_));
 sg13g2_antennanp ANTENNA_422 (.A(_11988_));
 sg13g2_antennanp ANTENNA_423 (.A(_11988_));
 sg13g2_antennanp ANTENNA_424 (.A(_11988_));
 sg13g2_antennanp ANTENNA_425 (.A(_12007_));
 sg13g2_antennanp ANTENNA_426 (.A(_12007_));
 sg13g2_antennanp ANTENNA_427 (.A(_12007_));
 sg13g2_antennanp ANTENNA_428 (.A(_12007_));
 sg13g2_antennanp ANTENNA_429 (.A(_12007_));
 sg13g2_antennanp ANTENNA_430 (.A(_12007_));
 sg13g2_antennanp ANTENNA_431 (.A(_12007_));
 sg13g2_antennanp ANTENNA_432 (.A(_12007_));
 sg13g2_antennanp ANTENNA_433 (.A(_12007_));
 sg13g2_antennanp ANTENNA_434 (.A(_12031_));
 sg13g2_antennanp ANTENNA_435 (.A(_12031_));
 sg13g2_antennanp ANTENNA_436 (.A(_12031_));
 sg13g2_antennanp ANTENNA_437 (.A(_12031_));
 sg13g2_antennanp ANTENNA_438 (.A(_12031_));
 sg13g2_antennanp ANTENNA_439 (.A(_12031_));
 sg13g2_antennanp ANTENNA_440 (.A(_12031_));
 sg13g2_antennanp ANTENNA_441 (.A(_12031_));
 sg13g2_antennanp ANTENNA_442 (.A(_12031_));
 sg13g2_antennanp ANTENNA_443 (.A(_12047_));
 sg13g2_antennanp ANTENNA_444 (.A(_12047_));
 sg13g2_antennanp ANTENNA_445 (.A(_12047_));
 sg13g2_antennanp ANTENNA_446 (.A(_12047_));
 sg13g2_antennanp ANTENNA_447 (.A(_12067_));
 sg13g2_antennanp ANTENNA_448 (.A(_12067_));
 sg13g2_antennanp ANTENNA_449 (.A(_12067_));
 sg13g2_antennanp ANTENNA_450 (.A(_12067_));
 sg13g2_antennanp ANTENNA_451 (.A(_12067_));
 sg13g2_antennanp ANTENNA_452 (.A(_12067_));
 sg13g2_antennanp ANTENNA_453 (.A(_12067_));
 sg13g2_antennanp ANTENNA_454 (.A(_12067_));
 sg13g2_antennanp ANTENNA_455 (.A(_12067_));
 sg13g2_antennanp ANTENNA_456 (.A(_12107_));
 sg13g2_antennanp ANTENNA_457 (.A(_12107_));
 sg13g2_antennanp ANTENNA_458 (.A(_12107_));
 sg13g2_antennanp ANTENNA_459 (.A(_12107_));
 sg13g2_antennanp ANTENNA_460 (.A(_12107_));
 sg13g2_antennanp ANTENNA_461 (.A(_12107_));
 sg13g2_antennanp ANTENNA_462 (.A(_12107_));
 sg13g2_antennanp ANTENNA_463 (.A(_12107_));
 sg13g2_antennanp ANTENNA_464 (.A(_12107_));
 sg13g2_antennanp ANTENNA_465 (.A(_12136_));
 sg13g2_antennanp ANTENNA_466 (.A(_12136_));
 sg13g2_antennanp ANTENNA_467 (.A(_12136_));
 sg13g2_antennanp ANTENNA_468 (.A(\cpu.dec.r_trap ));
 sg13g2_antennanp ANTENNA_469 (.A(\cpu.ex.pc[2] ));
 sg13g2_antennanp ANTENNA_470 (.A(\cpu.gpio.uart_rx ));
 sg13g2_antennanp ANTENNA_471 (.A(\cpu.gpio.uart_rx ));
 sg13g2_antennanp ANTENNA_472 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_473 (.A(net3));
 sg13g2_antennanp ANTENNA_474 (.A(net3));
 sg13g2_antennanp ANTENNA_475 (.A(net3));
 sg13g2_antennanp ANTENNA_476 (.A(net11));
 sg13g2_antennanp ANTENNA_477 (.A(net11));
 sg13g2_antennanp ANTENNA_478 (.A(net11));
 sg13g2_antennanp ANTENNA_479 (.A(net12));
 sg13g2_antennanp ANTENNA_480 (.A(net12));
 sg13g2_antennanp ANTENNA_481 (.A(net12));
 sg13g2_antennanp ANTENNA_482 (.A(net13));
 sg13g2_antennanp ANTENNA_483 (.A(net13));
 sg13g2_antennanp ANTENNA_484 (.A(net13));
 sg13g2_antennanp ANTENNA_485 (.A(net410));
 sg13g2_antennanp ANTENNA_486 (.A(net410));
 sg13g2_antennanp ANTENNA_487 (.A(net410));
 sg13g2_antennanp ANTENNA_488 (.A(net410));
 sg13g2_antennanp ANTENNA_489 (.A(net410));
 sg13g2_antennanp ANTENNA_490 (.A(net410));
 sg13g2_antennanp ANTENNA_491 (.A(net410));
 sg13g2_antennanp ANTENNA_492 (.A(net410));
 sg13g2_antennanp ANTENNA_493 (.A(net410));
 sg13g2_antennanp ANTENNA_494 (.A(net410));
 sg13g2_antennanp ANTENNA_495 (.A(net410));
 sg13g2_antennanp ANTENNA_496 (.A(net410));
 sg13g2_antennanp ANTENNA_497 (.A(net410));
 sg13g2_antennanp ANTENNA_498 (.A(net410));
 sg13g2_antennanp ANTENNA_499 (.A(net410));
 sg13g2_antennanp ANTENNA_500 (.A(net410));
 sg13g2_antennanp ANTENNA_501 (.A(net410));
 sg13g2_antennanp ANTENNA_502 (.A(net410));
 sg13g2_antennanp ANTENNA_503 (.A(net410));
 sg13g2_antennanp ANTENNA_504 (.A(net410));
 sg13g2_antennanp ANTENNA_505 (.A(net410));
 sg13g2_antennanp ANTENNA_506 (.A(net566));
 sg13g2_antennanp ANTENNA_507 (.A(net566));
 sg13g2_antennanp ANTENNA_508 (.A(net566));
 sg13g2_antennanp ANTENNA_509 (.A(net566));
 sg13g2_antennanp ANTENNA_510 (.A(net566));
 sg13g2_antennanp ANTENNA_511 (.A(net566));
 sg13g2_antennanp ANTENNA_512 (.A(net566));
 sg13g2_antennanp ANTENNA_513 (.A(net566));
 sg13g2_antennanp ANTENNA_514 (.A(net566));
 sg13g2_antennanp ANTENNA_515 (.A(net577));
 sg13g2_antennanp ANTENNA_516 (.A(net577));
 sg13g2_antennanp ANTENNA_517 (.A(net577));
 sg13g2_antennanp ANTENNA_518 (.A(net577));
 sg13g2_antennanp ANTENNA_519 (.A(net577));
 sg13g2_antennanp ANTENNA_520 (.A(net577));
 sg13g2_antennanp ANTENNA_521 (.A(net577));
 sg13g2_antennanp ANTENNA_522 (.A(net577));
 sg13g2_antennanp ANTENNA_523 (.A(net577));
 sg13g2_antennanp ANTENNA_524 (.A(net607));
 sg13g2_antennanp ANTENNA_525 (.A(net607));
 sg13g2_antennanp ANTENNA_526 (.A(net607));
 sg13g2_antennanp ANTENNA_527 (.A(net607));
 sg13g2_antennanp ANTENNA_528 (.A(net607));
 sg13g2_antennanp ANTENNA_529 (.A(net607));
 sg13g2_antennanp ANTENNA_530 (.A(net607));
 sg13g2_antennanp ANTENNA_531 (.A(net607));
 sg13g2_antennanp ANTENNA_532 (.A(net639));
 sg13g2_antennanp ANTENNA_533 (.A(net639));
 sg13g2_antennanp ANTENNA_534 (.A(net639));
 sg13g2_antennanp ANTENNA_535 (.A(net639));
 sg13g2_antennanp ANTENNA_536 (.A(net639));
 sg13g2_antennanp ANTENNA_537 (.A(net639));
 sg13g2_antennanp ANTENNA_538 (.A(net639));
 sg13g2_antennanp ANTENNA_539 (.A(net639));
 sg13g2_antennanp ANTENNA_540 (.A(net639));
 sg13g2_antennanp ANTENNA_541 (.A(net639));
 sg13g2_antennanp ANTENNA_542 (.A(net639));
 sg13g2_antennanp ANTENNA_543 (.A(net639));
 sg13g2_antennanp ANTENNA_544 (.A(net639));
 sg13g2_antennanp ANTENNA_545 (.A(net678));
 sg13g2_antennanp ANTENNA_546 (.A(net678));
 sg13g2_antennanp ANTENNA_547 (.A(net678));
 sg13g2_antennanp ANTENNA_548 (.A(net678));
 sg13g2_antennanp ANTENNA_549 (.A(net678));
 sg13g2_antennanp ANTENNA_550 (.A(net678));
 sg13g2_antennanp ANTENNA_551 (.A(net678));
 sg13g2_antennanp ANTENNA_552 (.A(net678));
 sg13g2_antennanp ANTENNA_553 (.A(net678));
 sg13g2_antennanp ANTENNA_554 (.A(net679));
 sg13g2_antennanp ANTENNA_555 (.A(net679));
 sg13g2_antennanp ANTENNA_556 (.A(net679));
 sg13g2_antennanp ANTENNA_557 (.A(net679));
 sg13g2_antennanp ANTENNA_558 (.A(net679));
 sg13g2_antennanp ANTENNA_559 (.A(net679));
 sg13g2_antennanp ANTENNA_560 (.A(net679));
 sg13g2_antennanp ANTENNA_561 (.A(net679));
 sg13g2_antennanp ANTENNA_562 (.A(net679));
 sg13g2_antennanp ANTENNA_563 (.A(net679));
 sg13g2_antennanp ANTENNA_564 (.A(net679));
 sg13g2_antennanp ANTENNA_565 (.A(net679));
 sg13g2_antennanp ANTENNA_566 (.A(net679));
 sg13g2_antennanp ANTENNA_567 (.A(net679));
 sg13g2_antennanp ANTENNA_568 (.A(net679));
 sg13g2_antennanp ANTENNA_569 (.A(net684));
 sg13g2_antennanp ANTENNA_570 (.A(net684));
 sg13g2_antennanp ANTENNA_571 (.A(net684));
 sg13g2_antennanp ANTENNA_572 (.A(net684));
 sg13g2_antennanp ANTENNA_573 (.A(net684));
 sg13g2_antennanp ANTENNA_574 (.A(net684));
 sg13g2_antennanp ANTENNA_575 (.A(net684));
 sg13g2_antennanp ANTENNA_576 (.A(net684));
 sg13g2_antennanp ANTENNA_577 (.A(net684));
 sg13g2_antennanp ANTENNA_578 (.A(net732));
 sg13g2_antennanp ANTENNA_579 (.A(net732));
 sg13g2_antennanp ANTENNA_580 (.A(net732));
 sg13g2_antennanp ANTENNA_581 (.A(net732));
 sg13g2_antennanp ANTENNA_582 (.A(net732));
 sg13g2_antennanp ANTENNA_583 (.A(net732));
 sg13g2_antennanp ANTENNA_584 (.A(net732));
 sg13g2_antennanp ANTENNA_585 (.A(net732));
 sg13g2_antennanp ANTENNA_586 (.A(net779));
 sg13g2_antennanp ANTENNA_587 (.A(net779));
 sg13g2_antennanp ANTENNA_588 (.A(net779));
 sg13g2_antennanp ANTENNA_589 (.A(net779));
 sg13g2_antennanp ANTENNA_590 (.A(net779));
 sg13g2_antennanp ANTENNA_591 (.A(net779));
 sg13g2_antennanp ANTENNA_592 (.A(net779));
 sg13g2_antennanp ANTENNA_593 (.A(net779));
 sg13g2_antennanp ANTENNA_594 (.A(net783));
 sg13g2_antennanp ANTENNA_595 (.A(net783));
 sg13g2_antennanp ANTENNA_596 (.A(net783));
 sg13g2_antennanp ANTENNA_597 (.A(net783));
 sg13g2_antennanp ANTENNA_598 (.A(net783));
 sg13g2_antennanp ANTENNA_599 (.A(net783));
 sg13g2_antennanp ANTENNA_600 (.A(net783));
 sg13g2_antennanp ANTENNA_601 (.A(net783));
 sg13g2_antennanp ANTENNA_602 (.A(net783));
 sg13g2_antennanp ANTENNA_603 (.A(net783));
 sg13g2_antennanp ANTENNA_604 (.A(net783));
 sg13g2_antennanp ANTENNA_605 (.A(net783));
 sg13g2_antennanp ANTENNA_606 (.A(net783));
 sg13g2_antennanp ANTENNA_607 (.A(net788));
 sg13g2_antennanp ANTENNA_608 (.A(net788));
 sg13g2_antennanp ANTENNA_609 (.A(net788));
 sg13g2_antennanp ANTENNA_610 (.A(net788));
 sg13g2_antennanp ANTENNA_611 (.A(net788));
 sg13g2_antennanp ANTENNA_612 (.A(net788));
 sg13g2_antennanp ANTENNA_613 (.A(net788));
 sg13g2_antennanp ANTENNA_614 (.A(net788));
 sg13g2_antennanp ANTENNA_615 (.A(net789));
 sg13g2_antennanp ANTENNA_616 (.A(net789));
 sg13g2_antennanp ANTENNA_617 (.A(net789));
 sg13g2_antennanp ANTENNA_618 (.A(net789));
 sg13g2_antennanp ANTENNA_619 (.A(net789));
 sg13g2_antennanp ANTENNA_620 (.A(net789));
 sg13g2_antennanp ANTENNA_621 (.A(net789));
 sg13g2_antennanp ANTENNA_622 (.A(net789));
 sg13g2_antennanp ANTENNA_623 (.A(net789));
 sg13g2_antennanp ANTENNA_624 (.A(net890));
 sg13g2_antennanp ANTENNA_625 (.A(net890));
 sg13g2_antennanp ANTENNA_626 (.A(net890));
 sg13g2_antennanp ANTENNA_627 (.A(net890));
 sg13g2_antennanp ANTENNA_628 (.A(net890));
 sg13g2_antennanp ANTENNA_629 (.A(net890));
 sg13g2_antennanp ANTENNA_630 (.A(net890));
 sg13g2_antennanp ANTENNA_631 (.A(net890));
 sg13g2_antennanp ANTENNA_632 (.A(net890));
 sg13g2_antennanp ANTENNA_633 (.A(net890));
 sg13g2_antennanp ANTENNA_634 (.A(net890));
 sg13g2_antennanp ANTENNA_635 (.A(net890));
 sg13g2_antennanp ANTENNA_636 (.A(net890));
 sg13g2_antennanp ANTENNA_637 (.A(net890));
 sg13g2_antennanp ANTENNA_638 (.A(net897));
 sg13g2_antennanp ANTENNA_639 (.A(net897));
 sg13g2_antennanp ANTENNA_640 (.A(net897));
 sg13g2_antennanp ANTENNA_641 (.A(net897));
 sg13g2_antennanp ANTENNA_642 (.A(net897));
 sg13g2_antennanp ANTENNA_643 (.A(net897));
 sg13g2_antennanp ANTENNA_644 (.A(net897));
 sg13g2_antennanp ANTENNA_645 (.A(net897));
 sg13g2_antennanp ANTENNA_646 (.A(net897));
 sg13g2_antennanp ANTENNA_647 (.A(net961));
 sg13g2_antennanp ANTENNA_648 (.A(net961));
 sg13g2_antennanp ANTENNA_649 (.A(net961));
 sg13g2_antennanp ANTENNA_650 (.A(net961));
 sg13g2_antennanp ANTENNA_651 (.A(net961));
 sg13g2_antennanp ANTENNA_652 (.A(net961));
 sg13g2_antennanp ANTENNA_653 (.A(net961));
 sg13g2_antennanp ANTENNA_654 (.A(net961));
 sg13g2_antennanp ANTENNA_655 (.A(net961));
 sg13g2_antennanp ANTENNA_656 (.A(net961));
 sg13g2_antennanp ANTENNA_657 (.A(net961));
 sg13g2_antennanp ANTENNA_658 (.A(net961));
 sg13g2_antennanp ANTENNA_659 (.A(net961));
 sg13g2_antennanp ANTENNA_660 (.A(net961));
 sg13g2_antennanp ANTENNA_661 (.A(net961));
 sg13g2_antennanp ANTENNA_662 (.A(net966));
 sg13g2_antennanp ANTENNA_663 (.A(net966));
 sg13g2_antennanp ANTENNA_664 (.A(net966));
 sg13g2_antennanp ANTENNA_665 (.A(net966));
 sg13g2_antennanp ANTENNA_666 (.A(net966));
 sg13g2_antennanp ANTENNA_667 (.A(net966));
 sg13g2_antennanp ANTENNA_668 (.A(net966));
 sg13g2_antennanp ANTENNA_669 (.A(net966));
 sg13g2_antennanp ANTENNA_670 (.A(net988));
 sg13g2_antennanp ANTENNA_671 (.A(net988));
 sg13g2_antennanp ANTENNA_672 (.A(net988));
 sg13g2_antennanp ANTENNA_673 (.A(net988));
 sg13g2_antennanp ANTENNA_674 (.A(net988));
 sg13g2_antennanp ANTENNA_675 (.A(net988));
 sg13g2_antennanp ANTENNA_676 (.A(net988));
 sg13g2_antennanp ANTENNA_677 (.A(net988));
 sg13g2_antennanp ANTENNA_678 (.A(net988));
 sg13g2_antennanp ANTENNA_679 (.A(net988));
 sg13g2_antennanp ANTENNA_680 (.A(net988));
 sg13g2_antennanp ANTENNA_681 (.A(net988));
 sg13g2_antennanp ANTENNA_682 (.A(net988));
 sg13g2_antennanp ANTENNA_683 (.A(net988));
 sg13g2_antennanp ANTENNA_684 (.A(net988));
 sg13g2_antennanp ANTENNA_685 (.A(net988));
 sg13g2_antennanp ANTENNA_686 (.A(net988));
 sg13g2_antennanp ANTENNA_687 (.A(net988));
 sg13g2_antennanp ANTENNA_688 (.A(net988));
 sg13g2_antennanp ANTENNA_689 (.A(net988));
 sg13g2_antennanp ANTENNA_690 (.A(net988));
 sg13g2_antennanp ANTENNA_691 (.A(net988));
 sg13g2_antennanp ANTENNA_692 (.A(net988));
 sg13g2_antennanp ANTENNA_693 (.A(net988));
 sg13g2_antennanp ANTENNA_694 (.A(net992));
 sg13g2_antennanp ANTENNA_695 (.A(net992));
 sg13g2_antennanp ANTENNA_696 (.A(net992));
 sg13g2_antennanp ANTENNA_697 (.A(net992));
 sg13g2_antennanp ANTENNA_698 (.A(net992));
 sg13g2_antennanp ANTENNA_699 (.A(net992));
 sg13g2_antennanp ANTENNA_700 (.A(net992));
 sg13g2_antennanp ANTENNA_701 (.A(net992));
 sg13g2_antennanp ANTENNA_702 (.A(net992));
 sg13g2_antennanp ANTENNA_703 (.A(net992));
 sg13g2_antennanp ANTENNA_704 (.A(net992));
 sg13g2_antennanp ANTENNA_705 (.A(net992));
 sg13g2_antennanp ANTENNA_706 (.A(net992));
 sg13g2_antennanp ANTENNA_707 (.A(net992));
 sg13g2_antennanp ANTENNA_708 (.A(net992));
 sg13g2_antennanp ANTENNA_709 (.A(net1056));
 sg13g2_antennanp ANTENNA_710 (.A(net1056));
 sg13g2_antennanp ANTENNA_711 (.A(net1056));
 sg13g2_antennanp ANTENNA_712 (.A(net1056));
 sg13g2_antennanp ANTENNA_713 (.A(net1056));
 sg13g2_antennanp ANTENNA_714 (.A(net1056));
 sg13g2_antennanp ANTENNA_715 (.A(net1056));
 sg13g2_antennanp ANTENNA_716 (.A(net1056));
 sg13g2_antennanp ANTENNA_717 (.A(net1056));
 sg13g2_antennanp ANTENNA_718 (.A(net1056));
 sg13g2_antennanp ANTENNA_719 (.A(net1056));
 sg13g2_antennanp ANTENNA_720 (.A(net1056));
 sg13g2_antennanp ANTENNA_721 (.A(net1056));
 sg13g2_antennanp ANTENNA_722 (.A(net1056));
 sg13g2_antennanp ANTENNA_723 (.A(net1057));
 sg13g2_antennanp ANTENNA_724 (.A(net1057));
 sg13g2_antennanp ANTENNA_725 (.A(net1057));
 sg13g2_antennanp ANTENNA_726 (.A(net1057));
 sg13g2_antennanp ANTENNA_727 (.A(net1057));
 sg13g2_antennanp ANTENNA_728 (.A(net1057));
 sg13g2_antennanp ANTENNA_729 (.A(net1057));
 sg13g2_antennanp ANTENNA_730 (.A(net1057));
 sg13g2_antennanp ANTENNA_731 (.A(net1057));
 sg13g2_antennanp ANTENNA_732 (.A(net1095));
 sg13g2_antennanp ANTENNA_733 (.A(net1095));
 sg13g2_antennanp ANTENNA_734 (.A(net1095));
 sg13g2_antennanp ANTENNA_735 (.A(net1095));
 sg13g2_antennanp ANTENNA_736 (.A(net1095));
 sg13g2_antennanp ANTENNA_737 (.A(net1095));
 sg13g2_antennanp ANTENNA_738 (.A(net1095));
 sg13g2_antennanp ANTENNA_739 (.A(net1095));
 sg13g2_antennanp ANTENNA_740 (.A(net1095));
 sg13g2_antennanp ANTENNA_741 (.A(net1095));
 sg13g2_antennanp ANTENNA_742 (.A(net1095));
 sg13g2_antennanp ANTENNA_743 (.A(net1095));
 sg13g2_antennanp ANTENNA_744 (.A(net1095));
 sg13g2_antennanp ANTENNA_745 (.A(net1095));
 sg13g2_antennanp ANTENNA_746 (.A(net1095));
 sg13g2_antennanp ANTENNA_747 (.A(net1095));
 sg13g2_antennanp ANTENNA_748 (.A(net1095));
 sg13g2_antennanp ANTENNA_749 (.A(net1095));
 sg13g2_antennanp ANTENNA_750 (.A(net1095));
 sg13g2_antennanp ANTENNA_751 (.A(net1095));
 sg13g2_antennanp ANTENNA_752 (.A(net1095));
 sg13g2_antennanp ANTENNA_753 (.A(net1095));
 sg13g2_antennanp ANTENNA_754 (.A(net1095));
 sg13g2_antennanp ANTENNA_755 (.A(net1095));
 sg13g2_antennanp ANTENNA_756 (.A(net1095));
 sg13g2_antennanp ANTENNA_757 (.A(net1095));
 sg13g2_antennanp ANTENNA_758 (.A(net1095));
 sg13g2_antennanp ANTENNA_759 (.A(net1095));
 sg13g2_antennanp ANTENNA_760 (.A(net1095));
 sg13g2_antennanp ANTENNA_761 (.A(net1095));
 sg13g2_antennanp ANTENNA_762 (.A(net1095));
 sg13g2_antennanp ANTENNA_763 (.A(net1095));
 sg13g2_antennanp ANTENNA_764 (.A(_00054_));
 sg13g2_antennanp ANTENNA_765 (.A(_00201_));
 sg13g2_antennanp ANTENNA_766 (.A(_00207_));
 sg13g2_antennanp ANTENNA_767 (.A(_00235_));
 sg13g2_antennanp ANTENNA_768 (.A(_00905_));
 sg13g2_antennanp ANTENNA_769 (.A(_00964_));
 sg13g2_antennanp ANTENNA_770 (.A(_00964_));
 sg13g2_antennanp ANTENNA_771 (.A(_01048_));
 sg13g2_antennanp ANTENNA_772 (.A(_02918_));
 sg13g2_antennanp ANTENNA_773 (.A(_02918_));
 sg13g2_antennanp ANTENNA_774 (.A(_02918_));
 sg13g2_antennanp ANTENNA_775 (.A(_02918_));
 sg13g2_antennanp ANTENNA_776 (.A(_02918_));
 sg13g2_antennanp ANTENNA_777 (.A(_02918_));
 sg13g2_antennanp ANTENNA_778 (.A(_02918_));
 sg13g2_antennanp ANTENNA_779 (.A(_02918_));
 sg13g2_antennanp ANTENNA_780 (.A(_02918_));
 sg13g2_antennanp ANTENNA_781 (.A(_02963_));
 sg13g2_antennanp ANTENNA_782 (.A(_02963_));
 sg13g2_antennanp ANTENNA_783 (.A(_02963_));
 sg13g2_antennanp ANTENNA_784 (.A(_02963_));
 sg13g2_antennanp ANTENNA_785 (.A(_02963_));
 sg13g2_antennanp ANTENNA_786 (.A(_02963_));
 sg13g2_antennanp ANTENNA_787 (.A(_03057_));
 sg13g2_antennanp ANTENNA_788 (.A(_03057_));
 sg13g2_antennanp ANTENNA_789 (.A(_03057_));
 sg13g2_antennanp ANTENNA_790 (.A(_03093_));
 sg13g2_antennanp ANTENNA_791 (.A(_03093_));
 sg13g2_antennanp ANTENNA_792 (.A(_03093_));
 sg13g2_antennanp ANTENNA_793 (.A(_03093_));
 sg13g2_antennanp ANTENNA_794 (.A(_03093_));
 sg13g2_antennanp ANTENNA_795 (.A(_03093_));
 sg13g2_antennanp ANTENNA_796 (.A(_03093_));
 sg13g2_antennanp ANTENNA_797 (.A(_03093_));
 sg13g2_antennanp ANTENNA_798 (.A(_03093_));
 sg13g2_antennanp ANTENNA_799 (.A(_03093_));
 sg13g2_antennanp ANTENNA_800 (.A(_03096_));
 sg13g2_antennanp ANTENNA_801 (.A(_03096_));
 sg13g2_antennanp ANTENNA_802 (.A(_03096_));
 sg13g2_antennanp ANTENNA_803 (.A(_03096_));
 sg13g2_antennanp ANTENNA_804 (.A(_03096_));
 sg13g2_antennanp ANTENNA_805 (.A(_03096_));
 sg13g2_antennanp ANTENNA_806 (.A(_03096_));
 sg13g2_antennanp ANTENNA_807 (.A(_03096_));
 sg13g2_antennanp ANTENNA_808 (.A(_03096_));
 sg13g2_antennanp ANTENNA_809 (.A(_03096_));
 sg13g2_antennanp ANTENNA_810 (.A(_03107_));
 sg13g2_antennanp ANTENNA_811 (.A(_03107_));
 sg13g2_antennanp ANTENNA_812 (.A(_03107_));
 sg13g2_antennanp ANTENNA_813 (.A(_03107_));
 sg13g2_antennanp ANTENNA_814 (.A(_03107_));
 sg13g2_antennanp ANTENNA_815 (.A(_03107_));
 sg13g2_antennanp ANTENNA_816 (.A(_03107_));
 sg13g2_antennanp ANTENNA_817 (.A(_03107_));
 sg13g2_antennanp ANTENNA_818 (.A(_03107_));
 sg13g2_antennanp ANTENNA_819 (.A(_03108_));
 sg13g2_antennanp ANTENNA_820 (.A(_03108_));
 sg13g2_antennanp ANTENNA_821 (.A(_03108_));
 sg13g2_antennanp ANTENNA_822 (.A(_03108_));
 sg13g2_antennanp ANTENNA_823 (.A(_03108_));
 sg13g2_antennanp ANTENNA_824 (.A(_03108_));
 sg13g2_antennanp ANTENNA_825 (.A(_03108_));
 sg13g2_antennanp ANTENNA_826 (.A(_03108_));
 sg13g2_antennanp ANTENNA_827 (.A(_03108_));
 sg13g2_antennanp ANTENNA_828 (.A(_03133_));
 sg13g2_antennanp ANTENNA_829 (.A(_03133_));
 sg13g2_antennanp ANTENNA_830 (.A(_03133_));
 sg13g2_antennanp ANTENNA_831 (.A(_03133_));
 sg13g2_antennanp ANTENNA_832 (.A(_03133_));
 sg13g2_antennanp ANTENNA_833 (.A(_03133_));
 sg13g2_antennanp ANTENNA_834 (.A(_03212_));
 sg13g2_antennanp ANTENNA_835 (.A(_03229_));
 sg13g2_antennanp ANTENNA_836 (.A(_03229_));
 sg13g2_antennanp ANTENNA_837 (.A(_03642_));
 sg13g2_antennanp ANTENNA_838 (.A(_03642_));
 sg13g2_antennanp ANTENNA_839 (.A(_03642_));
 sg13g2_antennanp ANTENNA_840 (.A(_03647_));
 sg13g2_antennanp ANTENNA_841 (.A(_03647_));
 sg13g2_antennanp ANTENNA_842 (.A(_03647_));
 sg13g2_antennanp ANTENNA_843 (.A(_03647_));
 sg13g2_antennanp ANTENNA_844 (.A(_03653_));
 sg13g2_antennanp ANTENNA_845 (.A(_03653_));
 sg13g2_antennanp ANTENNA_846 (.A(_03653_));
 sg13g2_antennanp ANTENNA_847 (.A(_03653_));
 sg13g2_antennanp ANTENNA_848 (.A(_03653_));
 sg13g2_antennanp ANTENNA_849 (.A(_03653_));
 sg13g2_antennanp ANTENNA_850 (.A(_03653_));
 sg13g2_antennanp ANTENNA_851 (.A(_03653_));
 sg13g2_antennanp ANTENNA_852 (.A(_03653_));
 sg13g2_antennanp ANTENNA_853 (.A(_03656_));
 sg13g2_antennanp ANTENNA_854 (.A(_03656_));
 sg13g2_antennanp ANTENNA_855 (.A(_03656_));
 sg13g2_antennanp ANTENNA_856 (.A(_03657_));
 sg13g2_antennanp ANTENNA_857 (.A(_03657_));
 sg13g2_antennanp ANTENNA_858 (.A(_03657_));
 sg13g2_antennanp ANTENNA_859 (.A(_03657_));
 sg13g2_antennanp ANTENNA_860 (.A(_03657_));
 sg13g2_antennanp ANTENNA_861 (.A(_03657_));
 sg13g2_antennanp ANTENNA_862 (.A(_03657_));
 sg13g2_antennanp ANTENNA_863 (.A(_03657_));
 sg13g2_antennanp ANTENNA_864 (.A(_03657_));
 sg13g2_antennanp ANTENNA_865 (.A(_03657_));
 sg13g2_antennanp ANTENNA_866 (.A(_03657_));
 sg13g2_antennanp ANTENNA_867 (.A(_03657_));
 sg13g2_antennanp ANTENNA_868 (.A(_03657_));
 sg13g2_antennanp ANTENNA_869 (.A(_03657_));
 sg13g2_antennanp ANTENNA_870 (.A(_04770_));
 sg13g2_antennanp ANTENNA_871 (.A(_04770_));
 sg13g2_antennanp ANTENNA_872 (.A(_04770_));
 sg13g2_antennanp ANTENNA_873 (.A(_04770_));
 sg13g2_antennanp ANTENNA_874 (.A(_04771_));
 sg13g2_antennanp ANTENNA_875 (.A(_04771_));
 sg13g2_antennanp ANTENNA_876 (.A(_04771_));
 sg13g2_antennanp ANTENNA_877 (.A(_04771_));
 sg13g2_antennanp ANTENNA_878 (.A(_04848_));
 sg13g2_antennanp ANTENNA_879 (.A(_04848_));
 sg13g2_antennanp ANTENNA_880 (.A(_05001_));
 sg13g2_antennanp ANTENNA_881 (.A(_05431_));
 sg13g2_antennanp ANTENNA_882 (.A(_05642_));
 sg13g2_antennanp ANTENNA_883 (.A(_05753_));
 sg13g2_antennanp ANTENNA_884 (.A(_05753_));
 sg13g2_antennanp ANTENNA_885 (.A(_05753_));
 sg13g2_antennanp ANTENNA_886 (.A(_05753_));
 sg13g2_antennanp ANTENNA_887 (.A(_05766_));
 sg13g2_antennanp ANTENNA_888 (.A(_05771_));
 sg13g2_antennanp ANTENNA_889 (.A(_05773_));
 sg13g2_antennanp ANTENNA_890 (.A(_05778_));
 sg13g2_antennanp ANTENNA_891 (.A(_05782_));
 sg13g2_antennanp ANTENNA_892 (.A(_05782_));
 sg13g2_antennanp ANTENNA_893 (.A(_05782_));
 sg13g2_antennanp ANTENNA_894 (.A(_05782_));
 sg13g2_antennanp ANTENNA_895 (.A(_05786_));
 sg13g2_antennanp ANTENNA_896 (.A(_05791_));
 sg13g2_antennanp ANTENNA_897 (.A(_06137_));
 sg13g2_antennanp ANTENNA_898 (.A(_06137_));
 sg13g2_antennanp ANTENNA_899 (.A(_06137_));
 sg13g2_antennanp ANTENNA_900 (.A(_06137_));
 sg13g2_antennanp ANTENNA_901 (.A(_06137_));
 sg13g2_antennanp ANTENNA_902 (.A(_06137_));
 sg13g2_antennanp ANTENNA_903 (.A(_06304_));
 sg13g2_antennanp ANTENNA_904 (.A(_06304_));
 sg13g2_antennanp ANTENNA_905 (.A(_06304_));
 sg13g2_antennanp ANTENNA_906 (.A(_06304_));
 sg13g2_antennanp ANTENNA_907 (.A(_06386_));
 sg13g2_antennanp ANTENNA_908 (.A(_06386_));
 sg13g2_antennanp ANTENNA_909 (.A(_06386_));
 sg13g2_antennanp ANTENNA_910 (.A(_06386_));
 sg13g2_antennanp ANTENNA_911 (.A(_06386_));
 sg13g2_antennanp ANTENNA_912 (.A(_06386_));
 sg13g2_antennanp ANTENNA_913 (.A(_06386_));
 sg13g2_antennanp ANTENNA_914 (.A(_06386_));
 sg13g2_antennanp ANTENNA_915 (.A(_06386_));
 sg13g2_antennanp ANTENNA_916 (.A(_07450_));
 sg13g2_antennanp ANTENNA_917 (.A(_07450_));
 sg13g2_antennanp ANTENNA_918 (.A(_07450_));
 sg13g2_antennanp ANTENNA_919 (.A(_07729_));
 sg13g2_antennanp ANTENNA_920 (.A(_07729_));
 sg13g2_antennanp ANTENNA_921 (.A(_07729_));
 sg13g2_antennanp ANTENNA_922 (.A(_07729_));
 sg13g2_antennanp ANTENNA_923 (.A(_07729_));
 sg13g2_antennanp ANTENNA_924 (.A(_07729_));
 sg13g2_antennanp ANTENNA_925 (.A(_07729_));
 sg13g2_antennanp ANTENNA_926 (.A(_07729_));
 sg13g2_antennanp ANTENNA_927 (.A(_07729_));
 sg13g2_antennanp ANTENNA_928 (.A(_08126_));
 sg13g2_antennanp ANTENNA_929 (.A(_08126_));
 sg13g2_antennanp ANTENNA_930 (.A(_08126_));
 sg13g2_antennanp ANTENNA_931 (.A(_08126_));
 sg13g2_antennanp ANTENNA_932 (.A(_08181_));
 sg13g2_antennanp ANTENNA_933 (.A(_08181_));
 sg13g2_antennanp ANTENNA_934 (.A(_08181_));
 sg13g2_antennanp ANTENNA_935 (.A(_08181_));
 sg13g2_antennanp ANTENNA_936 (.A(_08181_));
 sg13g2_antennanp ANTENNA_937 (.A(_08181_));
 sg13g2_antennanp ANTENNA_938 (.A(_08181_));
 sg13g2_antennanp ANTENNA_939 (.A(_08184_));
 sg13g2_antennanp ANTENNA_940 (.A(_08184_));
 sg13g2_antennanp ANTENNA_941 (.A(_08184_));
 sg13g2_antennanp ANTENNA_942 (.A(_08184_));
 sg13g2_antennanp ANTENNA_943 (.A(_08192_));
 sg13g2_antennanp ANTENNA_944 (.A(_08285_));
 sg13g2_antennanp ANTENNA_945 (.A(_08285_));
 sg13g2_antennanp ANTENNA_946 (.A(_08285_));
 sg13g2_antennanp ANTENNA_947 (.A(_08285_));
 sg13g2_antennanp ANTENNA_948 (.A(_08356_));
 sg13g2_antennanp ANTENNA_949 (.A(_08356_));
 sg13g2_antennanp ANTENNA_950 (.A(_08356_));
 sg13g2_antennanp ANTENNA_951 (.A(_08447_));
 sg13g2_antennanp ANTENNA_952 (.A(_08447_));
 sg13g2_antennanp ANTENNA_953 (.A(_08447_));
 sg13g2_antennanp ANTENNA_954 (.A(_08494_));
 sg13g2_antennanp ANTENNA_955 (.A(_08494_));
 sg13g2_antennanp ANTENNA_956 (.A(_08494_));
 sg13g2_antennanp ANTENNA_957 (.A(_08557_));
 sg13g2_antennanp ANTENNA_958 (.A(_08557_));
 sg13g2_antennanp ANTENNA_959 (.A(_08557_));
 sg13g2_antennanp ANTENNA_960 (.A(_08708_));
 sg13g2_antennanp ANTENNA_961 (.A(_08708_));
 sg13g2_antennanp ANTENNA_962 (.A(_08708_));
 sg13g2_antennanp ANTENNA_963 (.A(_08709_));
 sg13g2_antennanp ANTENNA_964 (.A(_08709_));
 sg13g2_antennanp ANTENNA_965 (.A(_08709_));
 sg13g2_antennanp ANTENNA_966 (.A(_08709_));
 sg13g2_antennanp ANTENNA_967 (.A(_08801_));
 sg13g2_antennanp ANTENNA_968 (.A(_08801_));
 sg13g2_antennanp ANTENNA_969 (.A(_08877_));
 sg13g2_antennanp ANTENNA_970 (.A(_08877_));
 sg13g2_antennanp ANTENNA_971 (.A(_08877_));
 sg13g2_antennanp ANTENNA_972 (.A(_08901_));
 sg13g2_antennanp ANTENNA_973 (.A(_08901_));
 sg13g2_antennanp ANTENNA_974 (.A(_08901_));
 sg13g2_antennanp ANTENNA_975 (.A(_08901_));
 sg13g2_antennanp ANTENNA_976 (.A(_08964_));
 sg13g2_antennanp ANTENNA_977 (.A(_08964_));
 sg13g2_antennanp ANTENNA_978 (.A(_08964_));
 sg13g2_antennanp ANTENNA_979 (.A(_08964_));
 sg13g2_antennanp ANTENNA_980 (.A(_08979_));
 sg13g2_antennanp ANTENNA_981 (.A(_08979_));
 sg13g2_antennanp ANTENNA_982 (.A(_08979_));
 sg13g2_antennanp ANTENNA_983 (.A(_08979_));
 sg13g2_antennanp ANTENNA_984 (.A(_08979_));
 sg13g2_antennanp ANTENNA_985 (.A(_09008_));
 sg13g2_antennanp ANTENNA_986 (.A(_09008_));
 sg13g2_antennanp ANTENNA_987 (.A(_09008_));
 sg13g2_antennanp ANTENNA_988 (.A(_09008_));
 sg13g2_antennanp ANTENNA_989 (.A(_09008_));
 sg13g2_antennanp ANTENNA_990 (.A(_09008_));
 sg13g2_antennanp ANTENNA_991 (.A(_09022_));
 sg13g2_antennanp ANTENNA_992 (.A(_09022_));
 sg13g2_antennanp ANTENNA_993 (.A(_09022_));
 sg13g2_antennanp ANTENNA_994 (.A(_09022_));
 sg13g2_antennanp ANTENNA_995 (.A(_09022_));
 sg13g2_antennanp ANTENNA_996 (.A(_09022_));
 sg13g2_antennanp ANTENNA_997 (.A(_09025_));
 sg13g2_antennanp ANTENNA_998 (.A(_09025_));
 sg13g2_antennanp ANTENNA_999 (.A(_09025_));
 sg13g2_antennanp ANTENNA_1000 (.A(_09025_));
 sg13g2_antennanp ANTENNA_1001 (.A(_09025_));
 sg13g2_antennanp ANTENNA_1002 (.A(_09025_));
 sg13g2_antennanp ANTENNA_1003 (.A(_09026_));
 sg13g2_antennanp ANTENNA_1004 (.A(_09026_));
 sg13g2_antennanp ANTENNA_1005 (.A(_09026_));
 sg13g2_antennanp ANTENNA_1006 (.A(_09026_));
 sg13g2_antennanp ANTENNA_1007 (.A(_09026_));
 sg13g2_antennanp ANTENNA_1008 (.A(_09026_));
 sg13g2_antennanp ANTENNA_1009 (.A(_09026_));
 sg13g2_antennanp ANTENNA_1010 (.A(_09026_));
 sg13g2_antennanp ANTENNA_1011 (.A(_09026_));
 sg13g2_antennanp ANTENNA_1012 (.A(_09036_));
 sg13g2_antennanp ANTENNA_1013 (.A(_09036_));
 sg13g2_antennanp ANTENNA_1014 (.A(_09036_));
 sg13g2_antennanp ANTENNA_1015 (.A(_09036_));
 sg13g2_antennanp ANTENNA_1016 (.A(_09045_));
 sg13g2_antennanp ANTENNA_1017 (.A(_09045_));
 sg13g2_antennanp ANTENNA_1018 (.A(_09106_));
 sg13g2_antennanp ANTENNA_1019 (.A(_09106_));
 sg13g2_antennanp ANTENNA_1020 (.A(_09106_));
 sg13g2_antennanp ANTENNA_1021 (.A(_09118_));
 sg13g2_antennanp ANTENNA_1022 (.A(_09118_));
 sg13g2_antennanp ANTENNA_1023 (.A(_09118_));
 sg13g2_antennanp ANTENNA_1024 (.A(_09118_));
 sg13g2_antennanp ANTENNA_1025 (.A(_09118_));
 sg13g2_antennanp ANTENNA_1026 (.A(_09122_));
 sg13g2_antennanp ANTENNA_1027 (.A(_09122_));
 sg13g2_antennanp ANTENNA_1028 (.A(_09122_));
 sg13g2_antennanp ANTENNA_1029 (.A(_09124_));
 sg13g2_antennanp ANTENNA_1030 (.A(_09124_));
 sg13g2_antennanp ANTENNA_1031 (.A(_09124_));
 sg13g2_antennanp ANTENNA_1032 (.A(_09124_));
 sg13g2_antennanp ANTENNA_1033 (.A(_09124_));
 sg13g2_antennanp ANTENNA_1034 (.A(_09124_));
 sg13g2_antennanp ANTENNA_1035 (.A(_09124_));
 sg13g2_antennanp ANTENNA_1036 (.A(_09124_));
 sg13g2_antennanp ANTENNA_1037 (.A(_09124_));
 sg13g2_antennanp ANTENNA_1038 (.A(_09124_));
 sg13g2_antennanp ANTENNA_1039 (.A(_09166_));
 sg13g2_antennanp ANTENNA_1040 (.A(_09166_));
 sg13g2_antennanp ANTENNA_1041 (.A(_09166_));
 sg13g2_antennanp ANTENNA_1042 (.A(_09166_));
 sg13g2_antennanp ANTENNA_1043 (.A(_09207_));
 sg13g2_antennanp ANTENNA_1044 (.A(_09251_));
 sg13g2_antennanp ANTENNA_1045 (.A(_09251_));
 sg13g2_antennanp ANTENNA_1046 (.A(_09273_));
 sg13g2_antennanp ANTENNA_1047 (.A(_09273_));
 sg13g2_antennanp ANTENNA_1048 (.A(_09273_));
 sg13g2_antennanp ANTENNA_1049 (.A(_09273_));
 sg13g2_antennanp ANTENNA_1050 (.A(_09273_));
 sg13g2_antennanp ANTENNA_1051 (.A(_09273_));
 sg13g2_antennanp ANTENNA_1052 (.A(_09273_));
 sg13g2_antennanp ANTENNA_1053 (.A(_09273_));
 sg13g2_antennanp ANTENNA_1054 (.A(_09293_));
 sg13g2_antennanp ANTENNA_1055 (.A(_09328_));
 sg13g2_antennanp ANTENNA_1056 (.A(_09340_));
 sg13g2_antennanp ANTENNA_1057 (.A(_09340_));
 sg13g2_antennanp ANTENNA_1058 (.A(_09340_));
 sg13g2_antennanp ANTENNA_1059 (.A(_09361_));
 sg13g2_antennanp ANTENNA_1060 (.A(_09398_));
 sg13g2_antennanp ANTENNA_1061 (.A(_09445_));
 sg13g2_antennanp ANTENNA_1062 (.A(_09485_));
 sg13g2_antennanp ANTENNA_1063 (.A(_09499_));
 sg13g2_antennanp ANTENNA_1064 (.A(_09606_));
 sg13g2_antennanp ANTENNA_1065 (.A(_09637_));
 sg13g2_antennanp ANTENNA_1066 (.A(_09872_));
 sg13g2_antennanp ANTENNA_1067 (.A(_09872_));
 sg13g2_antennanp ANTENNA_1068 (.A(_09872_));
 sg13g2_antennanp ANTENNA_1069 (.A(_09872_));
 sg13g2_antennanp ANTENNA_1070 (.A(_09872_));
 sg13g2_antennanp ANTENNA_1071 (.A(_09872_));
 sg13g2_antennanp ANTENNA_1072 (.A(_09872_));
 sg13g2_antennanp ANTENNA_1073 (.A(_09872_));
 sg13g2_antennanp ANTENNA_1074 (.A(_09872_));
 sg13g2_antennanp ANTENNA_1075 (.A(_09872_));
 sg13g2_antennanp ANTENNA_1076 (.A(_09872_));
 sg13g2_antennanp ANTENNA_1077 (.A(_09872_));
 sg13g2_antennanp ANTENNA_1078 (.A(_09872_));
 sg13g2_antennanp ANTENNA_1079 (.A(_09872_));
 sg13g2_antennanp ANTENNA_1080 (.A(_09875_));
 sg13g2_antennanp ANTENNA_1081 (.A(_09875_));
 sg13g2_antennanp ANTENNA_1082 (.A(_09875_));
 sg13g2_antennanp ANTENNA_1083 (.A(_09875_));
 sg13g2_antennanp ANTENNA_1084 (.A(_09875_));
 sg13g2_antennanp ANTENNA_1085 (.A(_09875_));
 sg13g2_antennanp ANTENNA_1086 (.A(_09875_));
 sg13g2_antennanp ANTENNA_1087 (.A(_09875_));
 sg13g2_antennanp ANTENNA_1088 (.A(_09875_));
 sg13g2_antennanp ANTENNA_1089 (.A(_09991_));
 sg13g2_antennanp ANTENNA_1090 (.A(_09991_));
 sg13g2_antennanp ANTENNA_1091 (.A(_09991_));
 sg13g2_antennanp ANTENNA_1092 (.A(_09991_));
 sg13g2_antennanp ANTENNA_1093 (.A(_09991_));
 sg13g2_antennanp ANTENNA_1094 (.A(_09991_));
 sg13g2_antennanp ANTENNA_1095 (.A(_09991_));
 sg13g2_antennanp ANTENNA_1096 (.A(_09991_));
 sg13g2_antennanp ANTENNA_1097 (.A(_10110_));
 sg13g2_antennanp ANTENNA_1098 (.A(_10423_));
 sg13g2_antennanp ANTENNA_1099 (.A(_10423_));
 sg13g2_antennanp ANTENNA_1100 (.A(_10423_));
 sg13g2_antennanp ANTENNA_1101 (.A(_10963_));
 sg13g2_antennanp ANTENNA_1102 (.A(_10963_));
 sg13g2_antennanp ANTENNA_1103 (.A(_10963_));
 sg13g2_antennanp ANTENNA_1104 (.A(_10963_));
 sg13g2_antennanp ANTENNA_1105 (.A(_11495_));
 sg13g2_antennanp ANTENNA_1106 (.A(_11495_));
 sg13g2_antennanp ANTENNA_1107 (.A(_11495_));
 sg13g2_antennanp ANTENNA_1108 (.A(_11495_));
 sg13g2_antennanp ANTENNA_1109 (.A(_11495_));
 sg13g2_antennanp ANTENNA_1110 (.A(_11900_));
 sg13g2_antennanp ANTENNA_1111 (.A(_11900_));
 sg13g2_antennanp ANTENNA_1112 (.A(_11900_));
 sg13g2_antennanp ANTENNA_1113 (.A(_11988_));
 sg13g2_antennanp ANTENNA_1114 (.A(_11988_));
 sg13g2_antennanp ANTENNA_1115 (.A(_11988_));
 sg13g2_antennanp ANTENNA_1116 (.A(_12007_));
 sg13g2_antennanp ANTENNA_1117 (.A(_12007_));
 sg13g2_antennanp ANTENNA_1118 (.A(_12007_));
 sg13g2_antennanp ANTENNA_1119 (.A(_12007_));
 sg13g2_antennanp ANTENNA_1120 (.A(_12007_));
 sg13g2_antennanp ANTENNA_1121 (.A(_12007_));
 sg13g2_antennanp ANTENNA_1122 (.A(_12007_));
 sg13g2_antennanp ANTENNA_1123 (.A(_12007_));
 sg13g2_antennanp ANTENNA_1124 (.A(_12007_));
 sg13g2_antennanp ANTENNA_1125 (.A(_12007_));
 sg13g2_antennanp ANTENNA_1126 (.A(_12007_));
 sg13g2_antennanp ANTENNA_1127 (.A(_12007_));
 sg13g2_antennanp ANTENNA_1128 (.A(_12007_));
 sg13g2_antennanp ANTENNA_1129 (.A(_12007_));
 sg13g2_antennanp ANTENNA_1130 (.A(_12007_));
 sg13g2_antennanp ANTENNA_1131 (.A(_12007_));
 sg13g2_antennanp ANTENNA_1132 (.A(_12007_));
 sg13g2_antennanp ANTENNA_1133 (.A(_12007_));
 sg13g2_antennanp ANTENNA_1134 (.A(_12031_));
 sg13g2_antennanp ANTENNA_1135 (.A(_12031_));
 sg13g2_antennanp ANTENNA_1136 (.A(_12031_));
 sg13g2_antennanp ANTENNA_1137 (.A(_12031_));
 sg13g2_antennanp ANTENNA_1138 (.A(_12031_));
 sg13g2_antennanp ANTENNA_1139 (.A(_12031_));
 sg13g2_antennanp ANTENNA_1140 (.A(_12031_));
 sg13g2_antennanp ANTENNA_1141 (.A(_12031_));
 sg13g2_antennanp ANTENNA_1142 (.A(_12031_));
 sg13g2_antennanp ANTENNA_1143 (.A(_12047_));
 sg13g2_antennanp ANTENNA_1144 (.A(_12047_));
 sg13g2_antennanp ANTENNA_1145 (.A(_12047_));
 sg13g2_antennanp ANTENNA_1146 (.A(_12047_));
 sg13g2_antennanp ANTENNA_1147 (.A(_12047_));
 sg13g2_antennanp ANTENNA_1148 (.A(_12047_));
 sg13g2_antennanp ANTENNA_1149 (.A(_12047_));
 sg13g2_antennanp ANTENNA_1150 (.A(_12047_));
 sg13g2_antennanp ANTENNA_1151 (.A(_12047_));
 sg13g2_antennanp ANTENNA_1152 (.A(_12067_));
 sg13g2_antennanp ANTENNA_1153 (.A(_12067_));
 sg13g2_antennanp ANTENNA_1154 (.A(_12067_));
 sg13g2_antennanp ANTENNA_1155 (.A(_12067_));
 sg13g2_antennanp ANTENNA_1156 (.A(_12067_));
 sg13g2_antennanp ANTENNA_1157 (.A(_12067_));
 sg13g2_antennanp ANTENNA_1158 (.A(_12067_));
 sg13g2_antennanp ANTENNA_1159 (.A(_12067_));
 sg13g2_antennanp ANTENNA_1160 (.A(_12067_));
 sg13g2_antennanp ANTENNA_1161 (.A(_12107_));
 sg13g2_antennanp ANTENNA_1162 (.A(_12107_));
 sg13g2_antennanp ANTENNA_1163 (.A(_12107_));
 sg13g2_antennanp ANTENNA_1164 (.A(_12107_));
 sg13g2_antennanp ANTENNA_1165 (.A(_12107_));
 sg13g2_antennanp ANTENNA_1166 (.A(_12107_));
 sg13g2_antennanp ANTENNA_1167 (.A(_12107_));
 sg13g2_antennanp ANTENNA_1168 (.A(_12107_));
 sg13g2_antennanp ANTENNA_1169 (.A(_12107_));
 sg13g2_antennanp ANTENNA_1170 (.A(_12136_));
 sg13g2_antennanp ANTENNA_1171 (.A(_12136_));
 sg13g2_antennanp ANTENNA_1172 (.A(_12136_));
 sg13g2_antennanp ANTENNA_1173 (.A(\cpu.dec.r_trap ));
 sg13g2_antennanp ANTENNA_1174 (.A(\cpu.ex.pc[2] ));
 sg13g2_antennanp ANTENNA_1175 (.A(\cpu.gpio.uart_rx ));
 sg13g2_antennanp ANTENNA_1176 (.A(\cpu.gpio.uart_rx ));
 sg13g2_antennanp ANTENNA_1177 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_1178 (.A(net3));
 sg13g2_antennanp ANTENNA_1179 (.A(net3));
 sg13g2_antennanp ANTENNA_1180 (.A(net3));
 sg13g2_antennanp ANTENNA_1181 (.A(net11));
 sg13g2_antennanp ANTENNA_1182 (.A(net11));
 sg13g2_antennanp ANTENNA_1183 (.A(net11));
 sg13g2_antennanp ANTENNA_1184 (.A(net12));
 sg13g2_antennanp ANTENNA_1185 (.A(net12));
 sg13g2_antennanp ANTENNA_1186 (.A(net12));
 sg13g2_antennanp ANTENNA_1187 (.A(net13));
 sg13g2_antennanp ANTENNA_1188 (.A(net13));
 sg13g2_antennanp ANTENNA_1189 (.A(net13));
 sg13g2_antennanp ANTENNA_1190 (.A(net566));
 sg13g2_antennanp ANTENNA_1191 (.A(net566));
 sg13g2_antennanp ANTENNA_1192 (.A(net566));
 sg13g2_antennanp ANTENNA_1193 (.A(net566));
 sg13g2_antennanp ANTENNA_1194 (.A(net566));
 sg13g2_antennanp ANTENNA_1195 (.A(net566));
 sg13g2_antennanp ANTENNA_1196 (.A(net566));
 sg13g2_antennanp ANTENNA_1197 (.A(net566));
 sg13g2_antennanp ANTENNA_1198 (.A(net566));
 sg13g2_antennanp ANTENNA_1199 (.A(net577));
 sg13g2_antennanp ANTENNA_1200 (.A(net577));
 sg13g2_antennanp ANTENNA_1201 (.A(net577));
 sg13g2_antennanp ANTENNA_1202 (.A(net577));
 sg13g2_antennanp ANTENNA_1203 (.A(net577));
 sg13g2_antennanp ANTENNA_1204 (.A(net577));
 sg13g2_antennanp ANTENNA_1205 (.A(net577));
 sg13g2_antennanp ANTENNA_1206 (.A(net577));
 sg13g2_antennanp ANTENNA_1207 (.A(net577));
 sg13g2_antennanp ANTENNA_1208 (.A(net589));
 sg13g2_antennanp ANTENNA_1209 (.A(net589));
 sg13g2_antennanp ANTENNA_1210 (.A(net589));
 sg13g2_antennanp ANTENNA_1211 (.A(net589));
 sg13g2_antennanp ANTENNA_1212 (.A(net589));
 sg13g2_antennanp ANTENNA_1213 (.A(net589));
 sg13g2_antennanp ANTENNA_1214 (.A(net589));
 sg13g2_antennanp ANTENNA_1215 (.A(net589));
 sg13g2_antennanp ANTENNA_1216 (.A(net589));
 sg13g2_antennanp ANTENNA_1217 (.A(net589));
 sg13g2_antennanp ANTENNA_1218 (.A(net589));
 sg13g2_antennanp ANTENNA_1219 (.A(net589));
 sg13g2_antennanp ANTENNA_1220 (.A(net589));
 sg13g2_antennanp ANTENNA_1221 (.A(net589));
 sg13g2_antennanp ANTENNA_1222 (.A(net589));
 sg13g2_antennanp ANTENNA_1223 (.A(net589));
 sg13g2_antennanp ANTENNA_1224 (.A(net639));
 sg13g2_antennanp ANTENNA_1225 (.A(net639));
 sg13g2_antennanp ANTENNA_1226 (.A(net639));
 sg13g2_antennanp ANTENNA_1227 (.A(net639));
 sg13g2_antennanp ANTENNA_1228 (.A(net639));
 sg13g2_antennanp ANTENNA_1229 (.A(net639));
 sg13g2_antennanp ANTENNA_1230 (.A(net639));
 sg13g2_antennanp ANTENNA_1231 (.A(net639));
 sg13g2_antennanp ANTENNA_1232 (.A(net639));
 sg13g2_antennanp ANTENNA_1233 (.A(net639));
 sg13g2_antennanp ANTENNA_1234 (.A(net639));
 sg13g2_antennanp ANTENNA_1235 (.A(net639));
 sg13g2_antennanp ANTENNA_1236 (.A(net639));
 sg13g2_antennanp ANTENNA_1237 (.A(net639));
 sg13g2_antennanp ANTENNA_1238 (.A(net639));
 sg13g2_antennanp ANTENNA_1239 (.A(net639));
 sg13g2_antennanp ANTENNA_1240 (.A(net639));
 sg13g2_antennanp ANTENNA_1241 (.A(net639));
 sg13g2_antennanp ANTENNA_1242 (.A(net639));
 sg13g2_antennanp ANTENNA_1243 (.A(net639));
 sg13g2_antennanp ANTENNA_1244 (.A(net639));
 sg13g2_antennanp ANTENNA_1245 (.A(net639));
 sg13g2_antennanp ANTENNA_1246 (.A(net639));
 sg13g2_antennanp ANTENNA_1247 (.A(net639));
 sg13g2_antennanp ANTENNA_1248 (.A(net640));
 sg13g2_antennanp ANTENNA_1249 (.A(net640));
 sg13g2_antennanp ANTENNA_1250 (.A(net640));
 sg13g2_antennanp ANTENNA_1251 (.A(net640));
 sg13g2_antennanp ANTENNA_1252 (.A(net640));
 sg13g2_antennanp ANTENNA_1253 (.A(net640));
 sg13g2_antennanp ANTENNA_1254 (.A(net640));
 sg13g2_antennanp ANTENNA_1255 (.A(net640));
 sg13g2_antennanp ANTENNA_1256 (.A(net640));
 sg13g2_antennanp ANTENNA_1257 (.A(net640));
 sg13g2_antennanp ANTENNA_1258 (.A(net640));
 sg13g2_antennanp ANTENNA_1259 (.A(net640));
 sg13g2_antennanp ANTENNA_1260 (.A(net640));
 sg13g2_antennanp ANTENNA_1261 (.A(net640));
 sg13g2_antennanp ANTENNA_1262 (.A(net640));
 sg13g2_antennanp ANTENNA_1263 (.A(net640));
 sg13g2_antennanp ANTENNA_1264 (.A(net640));
 sg13g2_antennanp ANTENNA_1265 (.A(net640));
 sg13g2_antennanp ANTENNA_1266 (.A(net640));
 sg13g2_antennanp ANTENNA_1267 (.A(net640));
 sg13g2_antennanp ANTENNA_1268 (.A(net640));
 sg13g2_antennanp ANTENNA_1269 (.A(net640));
 sg13g2_antennanp ANTENNA_1270 (.A(net640));
 sg13g2_antennanp ANTENNA_1271 (.A(net640));
 sg13g2_antennanp ANTENNA_1272 (.A(net640));
 sg13g2_antennanp ANTENNA_1273 (.A(net640));
 sg13g2_antennanp ANTENNA_1274 (.A(net640));
 sg13g2_antennanp ANTENNA_1275 (.A(net640));
 sg13g2_antennanp ANTENNA_1276 (.A(net640));
 sg13g2_antennanp ANTENNA_1277 (.A(net640));
 sg13g2_antennanp ANTENNA_1278 (.A(net640));
 sg13g2_antennanp ANTENNA_1279 (.A(net640));
 sg13g2_antennanp ANTENNA_1280 (.A(net640));
 sg13g2_antennanp ANTENNA_1281 (.A(net673));
 sg13g2_antennanp ANTENNA_1282 (.A(net673));
 sg13g2_antennanp ANTENNA_1283 (.A(net673));
 sg13g2_antennanp ANTENNA_1284 (.A(net673));
 sg13g2_antennanp ANTENNA_1285 (.A(net673));
 sg13g2_antennanp ANTENNA_1286 (.A(net673));
 sg13g2_antennanp ANTENNA_1287 (.A(net673));
 sg13g2_antennanp ANTENNA_1288 (.A(net673));
 sg13g2_antennanp ANTENNA_1289 (.A(net673));
 sg13g2_antennanp ANTENNA_1290 (.A(net673));
 sg13g2_antennanp ANTENNA_1291 (.A(net673));
 sg13g2_antennanp ANTENNA_1292 (.A(net673));
 sg13g2_antennanp ANTENNA_1293 (.A(net673));
 sg13g2_antennanp ANTENNA_1294 (.A(net673));
 sg13g2_antennanp ANTENNA_1295 (.A(net673));
 sg13g2_antennanp ANTENNA_1296 (.A(net673));
 sg13g2_antennanp ANTENNA_1297 (.A(net673));
 sg13g2_antennanp ANTENNA_1298 (.A(net673));
 sg13g2_antennanp ANTENNA_1299 (.A(net673));
 sg13g2_antennanp ANTENNA_1300 (.A(net673));
 sg13g2_antennanp ANTENNA_1301 (.A(net679));
 sg13g2_antennanp ANTENNA_1302 (.A(net679));
 sg13g2_antennanp ANTENNA_1303 (.A(net679));
 sg13g2_antennanp ANTENNA_1304 (.A(net679));
 sg13g2_antennanp ANTENNA_1305 (.A(net679));
 sg13g2_antennanp ANTENNA_1306 (.A(net679));
 sg13g2_antennanp ANTENNA_1307 (.A(net679));
 sg13g2_antennanp ANTENNA_1308 (.A(net679));
 sg13g2_antennanp ANTENNA_1309 (.A(net679));
 sg13g2_antennanp ANTENNA_1310 (.A(net679));
 sg13g2_antennanp ANTENNA_1311 (.A(net679));
 sg13g2_antennanp ANTENNA_1312 (.A(net679));
 sg13g2_antennanp ANTENNA_1313 (.A(net679));
 sg13g2_antennanp ANTENNA_1314 (.A(net679));
 sg13g2_antennanp ANTENNA_1315 (.A(net679));
 sg13g2_antennanp ANTENNA_1316 (.A(net684));
 sg13g2_antennanp ANTENNA_1317 (.A(net684));
 sg13g2_antennanp ANTENNA_1318 (.A(net684));
 sg13g2_antennanp ANTENNA_1319 (.A(net684));
 sg13g2_antennanp ANTENNA_1320 (.A(net684));
 sg13g2_antennanp ANTENNA_1321 (.A(net684));
 sg13g2_antennanp ANTENNA_1322 (.A(net684));
 sg13g2_antennanp ANTENNA_1323 (.A(net684));
 sg13g2_antennanp ANTENNA_1324 (.A(net684));
 sg13g2_antennanp ANTENNA_1325 (.A(net789));
 sg13g2_antennanp ANTENNA_1326 (.A(net789));
 sg13g2_antennanp ANTENNA_1327 (.A(net789));
 sg13g2_antennanp ANTENNA_1328 (.A(net789));
 sg13g2_antennanp ANTENNA_1329 (.A(net789));
 sg13g2_antennanp ANTENNA_1330 (.A(net789));
 sg13g2_antennanp ANTENNA_1331 (.A(net789));
 sg13g2_antennanp ANTENNA_1332 (.A(net789));
 sg13g2_antennanp ANTENNA_1333 (.A(net789));
 sg13g2_antennanp ANTENNA_1334 (.A(net855));
 sg13g2_antennanp ANTENNA_1335 (.A(net855));
 sg13g2_antennanp ANTENNA_1336 (.A(net855));
 sg13g2_antennanp ANTENNA_1337 (.A(net855));
 sg13g2_antennanp ANTENNA_1338 (.A(net855));
 sg13g2_antennanp ANTENNA_1339 (.A(net855));
 sg13g2_antennanp ANTENNA_1340 (.A(net855));
 sg13g2_antennanp ANTENNA_1341 (.A(net855));
 sg13g2_antennanp ANTENNA_1342 (.A(net855));
 sg13g2_antennanp ANTENNA_1343 (.A(net961));
 sg13g2_antennanp ANTENNA_1344 (.A(net961));
 sg13g2_antennanp ANTENNA_1345 (.A(net961));
 sg13g2_antennanp ANTENNA_1346 (.A(net961));
 sg13g2_antennanp ANTENNA_1347 (.A(net961));
 sg13g2_antennanp ANTENNA_1348 (.A(net961));
 sg13g2_antennanp ANTENNA_1349 (.A(net961));
 sg13g2_antennanp ANTENNA_1350 (.A(net961));
 sg13g2_antennanp ANTENNA_1351 (.A(net992));
 sg13g2_antennanp ANTENNA_1352 (.A(net992));
 sg13g2_antennanp ANTENNA_1353 (.A(net992));
 sg13g2_antennanp ANTENNA_1354 (.A(net992));
 sg13g2_antennanp ANTENNA_1355 (.A(net992));
 sg13g2_antennanp ANTENNA_1356 (.A(net992));
 sg13g2_antennanp ANTENNA_1357 (.A(net992));
 sg13g2_antennanp ANTENNA_1358 (.A(net992));
 sg13g2_antennanp ANTENNA_1359 (.A(net992));
 sg13g2_antennanp ANTENNA_1360 (.A(net992));
 sg13g2_antennanp ANTENNA_1361 (.A(net992));
 sg13g2_antennanp ANTENNA_1362 (.A(net992));
 sg13g2_antennanp ANTENNA_1363 (.A(net992));
 sg13g2_antennanp ANTENNA_1364 (.A(net992));
 sg13g2_antennanp ANTENNA_1365 (.A(net992));
 sg13g2_antennanp ANTENNA_1366 (.A(net1046));
 sg13g2_antennanp ANTENNA_1367 (.A(net1046));
 sg13g2_antennanp ANTENNA_1368 (.A(net1046));
 sg13g2_antennanp ANTENNA_1369 (.A(net1046));
 sg13g2_antennanp ANTENNA_1370 (.A(net1046));
 sg13g2_antennanp ANTENNA_1371 (.A(net1046));
 sg13g2_antennanp ANTENNA_1372 (.A(net1046));
 sg13g2_antennanp ANTENNA_1373 (.A(net1046));
 sg13g2_antennanp ANTENNA_1374 (.A(net1056));
 sg13g2_antennanp ANTENNA_1375 (.A(net1056));
 sg13g2_antennanp ANTENNA_1376 (.A(net1056));
 sg13g2_antennanp ANTENNA_1377 (.A(net1056));
 sg13g2_antennanp ANTENNA_1378 (.A(net1056));
 sg13g2_antennanp ANTENNA_1379 (.A(net1056));
 sg13g2_antennanp ANTENNA_1380 (.A(net1056));
 sg13g2_antennanp ANTENNA_1381 (.A(net1056));
 sg13g2_antennanp ANTENNA_1382 (.A(net1056));
 sg13g2_antennanp ANTENNA_1383 (.A(net1056));
 sg13g2_antennanp ANTENNA_1384 (.A(net1056));
 sg13g2_antennanp ANTENNA_1385 (.A(net1056));
 sg13g2_antennanp ANTENNA_1386 (.A(net1056));
 sg13g2_antennanp ANTENNA_1387 (.A(net1057));
 sg13g2_antennanp ANTENNA_1388 (.A(net1057));
 sg13g2_antennanp ANTENNA_1389 (.A(net1057));
 sg13g2_antennanp ANTENNA_1390 (.A(net1057));
 sg13g2_antennanp ANTENNA_1391 (.A(net1057));
 sg13g2_antennanp ANTENNA_1392 (.A(net1057));
 sg13g2_antennanp ANTENNA_1393 (.A(net1057));
 sg13g2_antennanp ANTENNA_1394 (.A(net1057));
 sg13g2_antennanp ANTENNA_1395 (.A(net1057));
 sg13g2_antennanp ANTENNA_1396 (.A(net1095));
 sg13g2_antennanp ANTENNA_1397 (.A(net1095));
 sg13g2_antennanp ANTENNA_1398 (.A(net1095));
 sg13g2_antennanp ANTENNA_1399 (.A(net1095));
 sg13g2_antennanp ANTENNA_1400 (.A(net1095));
 sg13g2_antennanp ANTENNA_1401 (.A(net1095));
 sg13g2_antennanp ANTENNA_1402 (.A(net1095));
 sg13g2_antennanp ANTENNA_1403 (.A(net1095));
 sg13g2_antennanp ANTENNA_1404 (.A(net1095));
 sg13g2_antennanp ANTENNA_1405 (.A(_00054_));
 sg13g2_antennanp ANTENNA_1406 (.A(_00201_));
 sg13g2_antennanp ANTENNA_1407 (.A(_00207_));
 sg13g2_antennanp ANTENNA_1408 (.A(_00235_));
 sg13g2_antennanp ANTENNA_1409 (.A(_00727_));
 sg13g2_antennanp ANTENNA_1410 (.A(_00769_));
 sg13g2_antennanp ANTENNA_1411 (.A(_00905_));
 sg13g2_antennanp ANTENNA_1412 (.A(_00964_));
 sg13g2_antennanp ANTENNA_1413 (.A(_00964_));
 sg13g2_antennanp ANTENNA_1414 (.A(_01048_));
 sg13g2_antennanp ANTENNA_1415 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1416 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1417 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1418 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1419 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1420 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1421 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1422 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1423 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1424 (.A(_02963_));
 sg13g2_antennanp ANTENNA_1425 (.A(_02963_));
 sg13g2_antennanp ANTENNA_1426 (.A(_02963_));
 sg13g2_antennanp ANTENNA_1427 (.A(_03093_));
 sg13g2_antennanp ANTENNA_1428 (.A(_03093_));
 sg13g2_antennanp ANTENNA_1429 (.A(_03093_));
 sg13g2_antennanp ANTENNA_1430 (.A(_03093_));
 sg13g2_antennanp ANTENNA_1431 (.A(_03093_));
 sg13g2_antennanp ANTENNA_1432 (.A(_03093_));
 sg13g2_antennanp ANTENNA_1433 (.A(_03093_));
 sg13g2_antennanp ANTENNA_1434 (.A(_03093_));
 sg13g2_antennanp ANTENNA_1435 (.A(_03093_));
 sg13g2_antennanp ANTENNA_1436 (.A(_03093_));
 sg13g2_antennanp ANTENNA_1437 (.A(_03096_));
 sg13g2_antennanp ANTENNA_1438 (.A(_03096_));
 sg13g2_antennanp ANTENNA_1439 (.A(_03096_));
 sg13g2_antennanp ANTENNA_1440 (.A(_03096_));
 sg13g2_antennanp ANTENNA_1441 (.A(_03096_));
 sg13g2_antennanp ANTENNA_1442 (.A(_03096_));
 sg13g2_antennanp ANTENNA_1443 (.A(_03096_));
 sg13g2_antennanp ANTENNA_1444 (.A(_03096_));
 sg13g2_antennanp ANTENNA_1445 (.A(_03096_));
 sg13g2_antennanp ANTENNA_1446 (.A(_03096_));
 sg13g2_antennanp ANTENNA_1447 (.A(_03107_));
 sg13g2_antennanp ANTENNA_1448 (.A(_03107_));
 sg13g2_antennanp ANTENNA_1449 (.A(_03107_));
 sg13g2_antennanp ANTENNA_1450 (.A(_03107_));
 sg13g2_antennanp ANTENNA_1451 (.A(_03107_));
 sg13g2_antennanp ANTENNA_1452 (.A(_03107_));
 sg13g2_antennanp ANTENNA_1453 (.A(_03107_));
 sg13g2_antennanp ANTENNA_1454 (.A(_03107_));
 sg13g2_antennanp ANTENNA_1455 (.A(_03107_));
 sg13g2_antennanp ANTENNA_1456 (.A(_03108_));
 sg13g2_antennanp ANTENNA_1457 (.A(_03108_));
 sg13g2_antennanp ANTENNA_1458 (.A(_03108_));
 sg13g2_antennanp ANTENNA_1459 (.A(_03108_));
 sg13g2_antennanp ANTENNA_1460 (.A(_03108_));
 sg13g2_antennanp ANTENNA_1461 (.A(_03108_));
 sg13g2_antennanp ANTENNA_1462 (.A(_03108_));
 sg13g2_antennanp ANTENNA_1463 (.A(_03108_));
 sg13g2_antennanp ANTENNA_1464 (.A(_03108_));
 sg13g2_antennanp ANTENNA_1465 (.A(_03133_));
 sg13g2_antennanp ANTENNA_1466 (.A(_03133_));
 sg13g2_antennanp ANTENNA_1467 (.A(_03133_));
 sg13g2_antennanp ANTENNA_1468 (.A(_03133_));
 sg13g2_antennanp ANTENNA_1469 (.A(_03133_));
 sg13g2_antennanp ANTENNA_1470 (.A(_03133_));
 sg13g2_antennanp ANTENNA_1471 (.A(_03133_));
 sg13g2_antennanp ANTENNA_1472 (.A(_03133_));
 sg13g2_antennanp ANTENNA_1473 (.A(_03133_));
 sg13g2_antennanp ANTENNA_1474 (.A(_03212_));
 sg13g2_antennanp ANTENNA_1475 (.A(_03229_));
 sg13g2_antennanp ANTENNA_1476 (.A(_03229_));
 sg13g2_antennanp ANTENNA_1477 (.A(_03642_));
 sg13g2_antennanp ANTENNA_1478 (.A(_03642_));
 sg13g2_antennanp ANTENNA_1479 (.A(_03642_));
 sg13g2_antennanp ANTENNA_1480 (.A(_03647_));
 sg13g2_antennanp ANTENNA_1481 (.A(_03647_));
 sg13g2_antennanp ANTENNA_1482 (.A(_03647_));
 sg13g2_antennanp ANTENNA_1483 (.A(_03647_));
 sg13g2_antennanp ANTENNA_1484 (.A(_03653_));
 sg13g2_antennanp ANTENNA_1485 (.A(_03653_));
 sg13g2_antennanp ANTENNA_1486 (.A(_03653_));
 sg13g2_antennanp ANTENNA_1487 (.A(_03653_));
 sg13g2_antennanp ANTENNA_1488 (.A(_03653_));
 sg13g2_antennanp ANTENNA_1489 (.A(_03653_));
 sg13g2_antennanp ANTENNA_1490 (.A(_03653_));
 sg13g2_antennanp ANTENNA_1491 (.A(_03653_));
 sg13g2_antennanp ANTENNA_1492 (.A(_03653_));
 sg13g2_antennanp ANTENNA_1493 (.A(_03656_));
 sg13g2_antennanp ANTENNA_1494 (.A(_03656_));
 sg13g2_antennanp ANTENNA_1495 (.A(_03656_));
 sg13g2_antennanp ANTENNA_1496 (.A(_03657_));
 sg13g2_antennanp ANTENNA_1497 (.A(_03657_));
 sg13g2_antennanp ANTENNA_1498 (.A(_03657_));
 sg13g2_antennanp ANTENNA_1499 (.A(_03657_));
 sg13g2_antennanp ANTENNA_1500 (.A(_03657_));
 sg13g2_antennanp ANTENNA_1501 (.A(_03657_));
 sg13g2_antennanp ANTENNA_1502 (.A(_03657_));
 sg13g2_antennanp ANTENNA_1503 (.A(_03657_));
 sg13g2_antennanp ANTENNA_1504 (.A(_03657_));
 sg13g2_antennanp ANTENNA_1505 (.A(_04770_));
 sg13g2_antennanp ANTENNA_1506 (.A(_04770_));
 sg13g2_antennanp ANTENNA_1507 (.A(_04770_));
 sg13g2_antennanp ANTENNA_1508 (.A(_04770_));
 sg13g2_antennanp ANTENNA_1509 (.A(_04848_));
 sg13g2_antennanp ANTENNA_1510 (.A(_04848_));
 sg13g2_antennanp ANTENNA_1511 (.A(_05001_));
 sg13g2_antennanp ANTENNA_1512 (.A(_05642_));
 sg13g2_antennanp ANTENNA_1513 (.A(_05753_));
 sg13g2_antennanp ANTENNA_1514 (.A(_05753_));
 sg13g2_antennanp ANTENNA_1515 (.A(_05753_));
 sg13g2_antennanp ANTENNA_1516 (.A(_05753_));
 sg13g2_antennanp ANTENNA_1517 (.A(_05766_));
 sg13g2_antennanp ANTENNA_1518 (.A(_05771_));
 sg13g2_antennanp ANTENNA_1519 (.A(_05771_));
 sg13g2_antennanp ANTENNA_1520 (.A(_05773_));
 sg13g2_antennanp ANTENNA_1521 (.A(_05778_));
 sg13g2_antennanp ANTENNA_1522 (.A(_05782_));
 sg13g2_antennanp ANTENNA_1523 (.A(_05782_));
 sg13g2_antennanp ANTENNA_1524 (.A(_05782_));
 sg13g2_antennanp ANTENNA_1525 (.A(_05782_));
 sg13g2_antennanp ANTENNA_1526 (.A(_05786_));
 sg13g2_antennanp ANTENNA_1527 (.A(_05791_));
 sg13g2_antennanp ANTENNA_1528 (.A(_06137_));
 sg13g2_antennanp ANTENNA_1529 (.A(_06137_));
 sg13g2_antennanp ANTENNA_1530 (.A(_06137_));
 sg13g2_antennanp ANTENNA_1531 (.A(_06137_));
 sg13g2_antennanp ANTENNA_1532 (.A(_06137_));
 sg13g2_antennanp ANTENNA_1533 (.A(_06137_));
 sg13g2_antennanp ANTENNA_1534 (.A(_06386_));
 sg13g2_antennanp ANTENNA_1535 (.A(_06386_));
 sg13g2_antennanp ANTENNA_1536 (.A(_06386_));
 sg13g2_antennanp ANTENNA_1537 (.A(_06386_));
 sg13g2_antennanp ANTENNA_1538 (.A(_06386_));
 sg13g2_antennanp ANTENNA_1539 (.A(_06386_));
 sg13g2_antennanp ANTENNA_1540 (.A(_06386_));
 sg13g2_antennanp ANTENNA_1541 (.A(_06386_));
 sg13g2_antennanp ANTENNA_1542 (.A(_06386_));
 sg13g2_antennanp ANTENNA_1543 (.A(_07450_));
 sg13g2_antennanp ANTENNA_1544 (.A(_07450_));
 sg13g2_antennanp ANTENNA_1545 (.A(_07450_));
 sg13g2_antennanp ANTENNA_1546 (.A(_07450_));
 sg13g2_antennanp ANTENNA_1547 (.A(_07729_));
 sg13g2_antennanp ANTENNA_1548 (.A(_07729_));
 sg13g2_antennanp ANTENNA_1549 (.A(_07729_));
 sg13g2_antennanp ANTENNA_1550 (.A(_07729_));
 sg13g2_antennanp ANTENNA_1551 (.A(_07729_));
 sg13g2_antennanp ANTENNA_1552 (.A(_07729_));
 sg13g2_antennanp ANTENNA_1553 (.A(_07729_));
 sg13g2_antennanp ANTENNA_1554 (.A(_07729_));
 sg13g2_antennanp ANTENNA_1555 (.A(_07729_));
 sg13g2_antennanp ANTENNA_1556 (.A(_08184_));
 sg13g2_antennanp ANTENNA_1557 (.A(_08184_));
 sg13g2_antennanp ANTENNA_1558 (.A(_08184_));
 sg13g2_antennanp ANTENNA_1559 (.A(_08184_));
 sg13g2_antennanp ANTENNA_1560 (.A(_08192_));
 sg13g2_antennanp ANTENNA_1561 (.A(_08285_));
 sg13g2_antennanp ANTENNA_1562 (.A(_08285_));
 sg13g2_antennanp ANTENNA_1563 (.A(_08285_));
 sg13g2_antennanp ANTENNA_1564 (.A(_08285_));
 sg13g2_antennanp ANTENNA_1565 (.A(_08447_));
 sg13g2_antennanp ANTENNA_1566 (.A(_08447_));
 sg13g2_antennanp ANTENNA_1567 (.A(_08447_));
 sg13g2_antennanp ANTENNA_1568 (.A(_08494_));
 sg13g2_antennanp ANTENNA_1569 (.A(_08494_));
 sg13g2_antennanp ANTENNA_1570 (.A(_08494_));
 sg13g2_antennanp ANTENNA_1571 (.A(_08708_));
 sg13g2_antennanp ANTENNA_1572 (.A(_08708_));
 sg13g2_antennanp ANTENNA_1573 (.A(_08708_));
 sg13g2_antennanp ANTENNA_1574 (.A(_08709_));
 sg13g2_antennanp ANTENNA_1575 (.A(_08709_));
 sg13g2_antennanp ANTENNA_1576 (.A(_08709_));
 sg13g2_antennanp ANTENNA_1577 (.A(_08709_));
 sg13g2_antennanp ANTENNA_1578 (.A(_08801_));
 sg13g2_antennanp ANTENNA_1579 (.A(_08801_));
 sg13g2_antennanp ANTENNA_1580 (.A(_08901_));
 sg13g2_antennanp ANTENNA_1581 (.A(_08901_));
 sg13g2_antennanp ANTENNA_1582 (.A(_08901_));
 sg13g2_antennanp ANTENNA_1583 (.A(_08901_));
 sg13g2_antennanp ANTENNA_1584 (.A(_08964_));
 sg13g2_antennanp ANTENNA_1585 (.A(_08964_));
 sg13g2_antennanp ANTENNA_1586 (.A(_08964_));
 sg13g2_antennanp ANTENNA_1587 (.A(_08964_));
 sg13g2_antennanp ANTENNA_1588 (.A(_08979_));
 sg13g2_antennanp ANTENNA_1589 (.A(_08979_));
 sg13g2_antennanp ANTENNA_1590 (.A(_08979_));
 sg13g2_antennanp ANTENNA_1591 (.A(_08979_));
 sg13g2_antennanp ANTENNA_1592 (.A(_08979_));
 sg13g2_antennanp ANTENNA_1593 (.A(_09008_));
 sg13g2_antennanp ANTENNA_1594 (.A(_09008_));
 sg13g2_antennanp ANTENNA_1595 (.A(_09008_));
 sg13g2_antennanp ANTENNA_1596 (.A(_09008_));
 sg13g2_antennanp ANTENNA_1597 (.A(_09008_));
 sg13g2_antennanp ANTENNA_1598 (.A(_09008_));
 sg13g2_antennanp ANTENNA_1599 (.A(_09022_));
 sg13g2_antennanp ANTENNA_1600 (.A(_09022_));
 sg13g2_antennanp ANTENNA_1601 (.A(_09022_));
 sg13g2_antennanp ANTENNA_1602 (.A(_09025_));
 sg13g2_antennanp ANTENNA_1603 (.A(_09025_));
 sg13g2_antennanp ANTENNA_1604 (.A(_09025_));
 sg13g2_antennanp ANTENNA_1605 (.A(_09025_));
 sg13g2_antennanp ANTENNA_1606 (.A(_09025_));
 sg13g2_antennanp ANTENNA_1607 (.A(_09025_));
 sg13g2_antennanp ANTENNA_1608 (.A(_09025_));
 sg13g2_antennanp ANTENNA_1609 (.A(_09025_));
 sg13g2_antennanp ANTENNA_1610 (.A(_09025_));
 sg13g2_antennanp ANTENNA_1611 (.A(_09036_));
 sg13g2_antennanp ANTENNA_1612 (.A(_09036_));
 sg13g2_antennanp ANTENNA_1613 (.A(_09036_));
 sg13g2_antennanp ANTENNA_1614 (.A(_09036_));
 sg13g2_antennanp ANTENNA_1615 (.A(_09045_));
 sg13g2_antennanp ANTENNA_1616 (.A(_09045_));
 sg13g2_antennanp ANTENNA_1617 (.A(_09052_));
 sg13g2_antennanp ANTENNA_1618 (.A(_09052_));
 sg13g2_antennanp ANTENNA_1619 (.A(_09052_));
 sg13g2_antennanp ANTENNA_1620 (.A(_09052_));
 sg13g2_antennanp ANTENNA_1621 (.A(_09052_));
 sg13g2_antennanp ANTENNA_1622 (.A(_09052_));
 sg13g2_antennanp ANTENNA_1623 (.A(_09052_));
 sg13g2_antennanp ANTENNA_1624 (.A(_09052_));
 sg13g2_antennanp ANTENNA_1625 (.A(_09052_));
 sg13g2_antennanp ANTENNA_1626 (.A(_09052_));
 sg13g2_antennanp ANTENNA_1627 (.A(_09118_));
 sg13g2_antennanp ANTENNA_1628 (.A(_09118_));
 sg13g2_antennanp ANTENNA_1629 (.A(_09118_));
 sg13g2_antennanp ANTENNA_1630 (.A(_09122_));
 sg13g2_antennanp ANTENNA_1631 (.A(_09122_));
 sg13g2_antennanp ANTENNA_1632 (.A(_09122_));
 sg13g2_antennanp ANTENNA_1633 (.A(_09124_));
 sg13g2_antennanp ANTENNA_1634 (.A(_09124_));
 sg13g2_antennanp ANTENNA_1635 (.A(_09124_));
 sg13g2_antennanp ANTENNA_1636 (.A(_09124_));
 sg13g2_antennanp ANTENNA_1637 (.A(_09124_));
 sg13g2_antennanp ANTENNA_1638 (.A(_09124_));
 sg13g2_antennanp ANTENNA_1639 (.A(_09124_));
 sg13g2_antennanp ANTENNA_1640 (.A(_09124_));
 sg13g2_antennanp ANTENNA_1641 (.A(_09124_));
 sg13g2_antennanp ANTENNA_1642 (.A(_09166_));
 sg13g2_antennanp ANTENNA_1643 (.A(_09166_));
 sg13g2_antennanp ANTENNA_1644 (.A(_09166_));
 sg13g2_antennanp ANTENNA_1645 (.A(_09166_));
 sg13g2_antennanp ANTENNA_1646 (.A(_09207_));
 sg13g2_antennanp ANTENNA_1647 (.A(_09251_));
 sg13g2_antennanp ANTENNA_1648 (.A(_09273_));
 sg13g2_antennanp ANTENNA_1649 (.A(_09273_));
 sg13g2_antennanp ANTENNA_1650 (.A(_09273_));
 sg13g2_antennanp ANTENNA_1651 (.A(_09273_));
 sg13g2_antennanp ANTENNA_1652 (.A(_09273_));
 sg13g2_antennanp ANTENNA_1653 (.A(_09273_));
 sg13g2_antennanp ANTENNA_1654 (.A(_09273_));
 sg13g2_antennanp ANTENNA_1655 (.A(_09273_));
 sg13g2_antennanp ANTENNA_1656 (.A(_09328_));
 sg13g2_antennanp ANTENNA_1657 (.A(_09361_));
 sg13g2_antennanp ANTENNA_1658 (.A(_09398_));
 sg13g2_antennanp ANTENNA_1659 (.A(_09445_));
 sg13g2_antennanp ANTENNA_1660 (.A(_09485_));
 sg13g2_antennanp ANTENNA_1661 (.A(_09499_));
 sg13g2_antennanp ANTENNA_1662 (.A(_09606_));
 sg13g2_antennanp ANTENNA_1663 (.A(_09637_));
 sg13g2_antennanp ANTENNA_1664 (.A(_09875_));
 sg13g2_antennanp ANTENNA_1665 (.A(_09875_));
 sg13g2_antennanp ANTENNA_1666 (.A(_09875_));
 sg13g2_antennanp ANTENNA_1667 (.A(_09875_));
 sg13g2_antennanp ANTENNA_1668 (.A(_09875_));
 sg13g2_antennanp ANTENNA_1669 (.A(_09875_));
 sg13g2_antennanp ANTENNA_1670 (.A(_09875_));
 sg13g2_antennanp ANTENNA_1671 (.A(_09875_));
 sg13g2_antennanp ANTENNA_1672 (.A(_09875_));
 sg13g2_antennanp ANTENNA_1673 (.A(_09907_));
 sg13g2_antennanp ANTENNA_1674 (.A(_09907_));
 sg13g2_antennanp ANTENNA_1675 (.A(_09907_));
 sg13g2_antennanp ANTENNA_1676 (.A(_09907_));
 sg13g2_antennanp ANTENNA_1677 (.A(_09907_));
 sg13g2_antennanp ANTENNA_1678 (.A(_09907_));
 sg13g2_antennanp ANTENNA_1679 (.A(_09907_));
 sg13g2_antennanp ANTENNA_1680 (.A(_10110_));
 sg13g2_antennanp ANTENNA_1681 (.A(_10831_));
 sg13g2_antennanp ANTENNA_1682 (.A(_10831_));
 sg13g2_antennanp ANTENNA_1683 (.A(_10831_));
 sg13g2_antennanp ANTENNA_1684 (.A(_10831_));
 sg13g2_antennanp ANTENNA_1685 (.A(_10831_));
 sg13g2_antennanp ANTENNA_1686 (.A(_10831_));
 sg13g2_antennanp ANTENNA_1687 (.A(_10831_));
 sg13g2_antennanp ANTENNA_1688 (.A(_10831_));
 sg13g2_antennanp ANTENNA_1689 (.A(_10831_));
 sg13g2_antennanp ANTENNA_1690 (.A(_10963_));
 sg13g2_antennanp ANTENNA_1691 (.A(_10963_));
 sg13g2_antennanp ANTENNA_1692 (.A(_10963_));
 sg13g2_antennanp ANTENNA_1693 (.A(_10963_));
 sg13g2_antennanp ANTENNA_1694 (.A(_11495_));
 sg13g2_antennanp ANTENNA_1695 (.A(_11495_));
 sg13g2_antennanp ANTENNA_1696 (.A(_11495_));
 sg13g2_antennanp ANTENNA_1697 (.A(_11495_));
 sg13g2_antennanp ANTENNA_1698 (.A(_11495_));
 sg13g2_antennanp ANTENNA_1699 (.A(_12007_));
 sg13g2_antennanp ANTENNA_1700 (.A(_12007_));
 sg13g2_antennanp ANTENNA_1701 (.A(_12007_));
 sg13g2_antennanp ANTENNA_1702 (.A(_12007_));
 sg13g2_antennanp ANTENNA_1703 (.A(_12007_));
 sg13g2_antennanp ANTENNA_1704 (.A(_12007_));
 sg13g2_antennanp ANTENNA_1705 (.A(_12007_));
 sg13g2_antennanp ANTENNA_1706 (.A(_12007_));
 sg13g2_antennanp ANTENNA_1707 (.A(_12007_));
 sg13g2_antennanp ANTENNA_1708 (.A(_12031_));
 sg13g2_antennanp ANTENNA_1709 (.A(_12031_));
 sg13g2_antennanp ANTENNA_1710 (.A(_12031_));
 sg13g2_antennanp ANTENNA_1711 (.A(_12031_));
 sg13g2_antennanp ANTENNA_1712 (.A(_12031_));
 sg13g2_antennanp ANTENNA_1713 (.A(_12031_));
 sg13g2_antennanp ANTENNA_1714 (.A(_12031_));
 sg13g2_antennanp ANTENNA_1715 (.A(_12031_));
 sg13g2_antennanp ANTENNA_1716 (.A(_12031_));
 sg13g2_antennanp ANTENNA_1717 (.A(_12047_));
 sg13g2_antennanp ANTENNA_1718 (.A(_12047_));
 sg13g2_antennanp ANTENNA_1719 (.A(_12047_));
 sg13g2_antennanp ANTENNA_1720 (.A(_12047_));
 sg13g2_antennanp ANTENNA_1721 (.A(_12047_));
 sg13g2_antennanp ANTENNA_1722 (.A(_12047_));
 sg13g2_antennanp ANTENNA_1723 (.A(_12047_));
 sg13g2_antennanp ANTENNA_1724 (.A(_12047_));
 sg13g2_antennanp ANTENNA_1725 (.A(_12047_));
 sg13g2_antennanp ANTENNA_1726 (.A(_12067_));
 sg13g2_antennanp ANTENNA_1727 (.A(_12067_));
 sg13g2_antennanp ANTENNA_1728 (.A(_12067_));
 sg13g2_antennanp ANTENNA_1729 (.A(_12067_));
 sg13g2_antennanp ANTENNA_1730 (.A(_12067_));
 sg13g2_antennanp ANTENNA_1731 (.A(_12067_));
 sg13g2_antennanp ANTENNA_1732 (.A(_12067_));
 sg13g2_antennanp ANTENNA_1733 (.A(_12067_));
 sg13g2_antennanp ANTENNA_1734 (.A(_12067_));
 sg13g2_antennanp ANTENNA_1735 (.A(_12107_));
 sg13g2_antennanp ANTENNA_1736 (.A(_12107_));
 sg13g2_antennanp ANTENNA_1737 (.A(_12107_));
 sg13g2_antennanp ANTENNA_1738 (.A(_12107_));
 sg13g2_antennanp ANTENNA_1739 (.A(_12107_));
 sg13g2_antennanp ANTENNA_1740 (.A(_12107_));
 sg13g2_antennanp ANTENNA_1741 (.A(_12107_));
 sg13g2_antennanp ANTENNA_1742 (.A(_12107_));
 sg13g2_antennanp ANTENNA_1743 (.A(_12107_));
 sg13g2_antennanp ANTENNA_1744 (.A(_12136_));
 sg13g2_antennanp ANTENNA_1745 (.A(_12136_));
 sg13g2_antennanp ANTENNA_1746 (.A(_12136_));
 sg13g2_antennanp ANTENNA_1747 (.A(\cpu.dec.r_trap ));
 sg13g2_antennanp ANTENNA_1748 (.A(\cpu.ex.pc[2] ));
 sg13g2_antennanp ANTENNA_1749 (.A(\cpu.gpio.uart_rx ));
 sg13g2_antennanp ANTENNA_1750 (.A(\cpu.gpio.uart_rx ));
 sg13g2_antennanp ANTENNA_1751 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_1752 (.A(net11));
 sg13g2_antennanp ANTENNA_1753 (.A(net11));
 sg13g2_antennanp ANTENNA_1754 (.A(net11));
 sg13g2_antennanp ANTENNA_1755 (.A(net12));
 sg13g2_antennanp ANTENNA_1756 (.A(net12));
 sg13g2_antennanp ANTENNA_1757 (.A(net12));
 sg13g2_antennanp ANTENNA_1758 (.A(net13));
 sg13g2_antennanp ANTENNA_1759 (.A(net13));
 sg13g2_antennanp ANTENNA_1760 (.A(net410));
 sg13g2_antennanp ANTENNA_1761 (.A(net410));
 sg13g2_antennanp ANTENNA_1762 (.A(net410));
 sg13g2_antennanp ANTENNA_1763 (.A(net410));
 sg13g2_antennanp ANTENNA_1764 (.A(net410));
 sg13g2_antennanp ANTENNA_1765 (.A(net410));
 sg13g2_antennanp ANTENNA_1766 (.A(net410));
 sg13g2_antennanp ANTENNA_1767 (.A(net410));
 sg13g2_antennanp ANTENNA_1768 (.A(net566));
 sg13g2_antennanp ANTENNA_1769 (.A(net566));
 sg13g2_antennanp ANTENNA_1770 (.A(net566));
 sg13g2_antennanp ANTENNA_1771 (.A(net566));
 sg13g2_antennanp ANTENNA_1772 (.A(net566));
 sg13g2_antennanp ANTENNA_1773 (.A(net566));
 sg13g2_antennanp ANTENNA_1774 (.A(net566));
 sg13g2_antennanp ANTENNA_1775 (.A(net566));
 sg13g2_antennanp ANTENNA_1776 (.A(net566));
 sg13g2_antennanp ANTENNA_1777 (.A(net577));
 sg13g2_antennanp ANTENNA_1778 (.A(net577));
 sg13g2_antennanp ANTENNA_1779 (.A(net577));
 sg13g2_antennanp ANTENNA_1780 (.A(net577));
 sg13g2_antennanp ANTENNA_1781 (.A(net577));
 sg13g2_antennanp ANTENNA_1782 (.A(net577));
 sg13g2_antennanp ANTENNA_1783 (.A(net577));
 sg13g2_antennanp ANTENNA_1784 (.A(net577));
 sg13g2_antennanp ANTENNA_1785 (.A(net577));
 sg13g2_antennanp ANTENNA_1786 (.A(net589));
 sg13g2_antennanp ANTENNA_1787 (.A(net589));
 sg13g2_antennanp ANTENNA_1788 (.A(net589));
 sg13g2_antennanp ANTENNA_1789 (.A(net589));
 sg13g2_antennanp ANTENNA_1790 (.A(net589));
 sg13g2_antennanp ANTENNA_1791 (.A(net589));
 sg13g2_antennanp ANTENNA_1792 (.A(net589));
 sg13g2_antennanp ANTENNA_1793 (.A(net589));
 sg13g2_antennanp ANTENNA_1794 (.A(net589));
 sg13g2_antennanp ANTENNA_1795 (.A(net589));
 sg13g2_antennanp ANTENNA_1796 (.A(net589));
 sg13g2_antennanp ANTENNA_1797 (.A(net589));
 sg13g2_antennanp ANTENNA_1798 (.A(net589));
 sg13g2_antennanp ANTENNA_1799 (.A(net589));
 sg13g2_antennanp ANTENNA_1800 (.A(net589));
 sg13g2_antennanp ANTENNA_1801 (.A(net589));
 sg13g2_antennanp ANTENNA_1802 (.A(net639));
 sg13g2_antennanp ANTENNA_1803 (.A(net639));
 sg13g2_antennanp ANTENNA_1804 (.A(net639));
 sg13g2_antennanp ANTENNA_1805 (.A(net639));
 sg13g2_antennanp ANTENNA_1806 (.A(net639));
 sg13g2_antennanp ANTENNA_1807 (.A(net639));
 sg13g2_antennanp ANTENNA_1808 (.A(net639));
 sg13g2_antennanp ANTENNA_1809 (.A(net639));
 sg13g2_antennanp ANTENNA_1810 (.A(net673));
 sg13g2_antennanp ANTENNA_1811 (.A(net673));
 sg13g2_antennanp ANTENNA_1812 (.A(net673));
 sg13g2_antennanp ANTENNA_1813 (.A(net673));
 sg13g2_antennanp ANTENNA_1814 (.A(net673));
 sg13g2_antennanp ANTENNA_1815 (.A(net673));
 sg13g2_antennanp ANTENNA_1816 (.A(net673));
 sg13g2_antennanp ANTENNA_1817 (.A(net673));
 sg13g2_antennanp ANTENNA_1818 (.A(net679));
 sg13g2_antennanp ANTENNA_1819 (.A(net679));
 sg13g2_antennanp ANTENNA_1820 (.A(net679));
 sg13g2_antennanp ANTENNA_1821 (.A(net679));
 sg13g2_antennanp ANTENNA_1822 (.A(net679));
 sg13g2_antennanp ANTENNA_1823 (.A(net679));
 sg13g2_antennanp ANTENNA_1824 (.A(net679));
 sg13g2_antennanp ANTENNA_1825 (.A(net679));
 sg13g2_antennanp ANTENNA_1826 (.A(net679));
 sg13g2_antennanp ANTENNA_1827 (.A(net679));
 sg13g2_antennanp ANTENNA_1828 (.A(net679));
 sg13g2_antennanp ANTENNA_1829 (.A(net679));
 sg13g2_antennanp ANTENNA_1830 (.A(net679));
 sg13g2_antennanp ANTENNA_1831 (.A(net679));
 sg13g2_antennanp ANTENNA_1832 (.A(net679));
 sg13g2_antennanp ANTENNA_1833 (.A(net684));
 sg13g2_antennanp ANTENNA_1834 (.A(net684));
 sg13g2_antennanp ANTENNA_1835 (.A(net684));
 sg13g2_antennanp ANTENNA_1836 (.A(net684));
 sg13g2_antennanp ANTENNA_1837 (.A(net684));
 sg13g2_antennanp ANTENNA_1838 (.A(net684));
 sg13g2_antennanp ANTENNA_1839 (.A(net684));
 sg13g2_antennanp ANTENNA_1840 (.A(net684));
 sg13g2_antennanp ANTENNA_1841 (.A(net684));
 sg13g2_antennanp ANTENNA_1842 (.A(net783));
 sg13g2_antennanp ANTENNA_1843 (.A(net783));
 sg13g2_antennanp ANTENNA_1844 (.A(net783));
 sg13g2_antennanp ANTENNA_1845 (.A(net783));
 sg13g2_antennanp ANTENNA_1846 (.A(net783));
 sg13g2_antennanp ANTENNA_1847 (.A(net783));
 sg13g2_antennanp ANTENNA_1848 (.A(net783));
 sg13g2_antennanp ANTENNA_1849 (.A(net783));
 sg13g2_antennanp ANTENNA_1850 (.A(net783));
 sg13g2_antennanp ANTENNA_1851 (.A(net783));
 sg13g2_antennanp ANTENNA_1852 (.A(net783));
 sg13g2_antennanp ANTENNA_1853 (.A(net783));
 sg13g2_antennanp ANTENNA_1854 (.A(net783));
 sg13g2_antennanp ANTENNA_1855 (.A(net783));
 sg13g2_antennanp ANTENNA_1856 (.A(net783));
 sg13g2_antennanp ANTENNA_1857 (.A(net789));
 sg13g2_antennanp ANTENNA_1858 (.A(net789));
 sg13g2_antennanp ANTENNA_1859 (.A(net789));
 sg13g2_antennanp ANTENNA_1860 (.A(net789));
 sg13g2_antennanp ANTENNA_1861 (.A(net789));
 sg13g2_antennanp ANTENNA_1862 (.A(net789));
 sg13g2_antennanp ANTENNA_1863 (.A(net789));
 sg13g2_antennanp ANTENNA_1864 (.A(net789));
 sg13g2_antennanp ANTENNA_1865 (.A(net789));
 sg13g2_antennanp ANTENNA_1866 (.A(net961));
 sg13g2_antennanp ANTENNA_1867 (.A(net961));
 sg13g2_antennanp ANTENNA_1868 (.A(net961));
 sg13g2_antennanp ANTENNA_1869 (.A(net961));
 sg13g2_antennanp ANTENNA_1870 (.A(net961));
 sg13g2_antennanp ANTENNA_1871 (.A(net961));
 sg13g2_antennanp ANTENNA_1872 (.A(net961));
 sg13g2_antennanp ANTENNA_1873 (.A(net961));
 sg13g2_antennanp ANTENNA_1874 (.A(net1037));
 sg13g2_antennanp ANTENNA_1875 (.A(net1037));
 sg13g2_antennanp ANTENNA_1876 (.A(net1037));
 sg13g2_antennanp ANTENNA_1877 (.A(net1037));
 sg13g2_antennanp ANTENNA_1878 (.A(net1037));
 sg13g2_antennanp ANTENNA_1879 (.A(net1037));
 sg13g2_antennanp ANTENNA_1880 (.A(net1037));
 sg13g2_antennanp ANTENNA_1881 (.A(net1037));
 sg13g2_antennanp ANTENNA_1882 (.A(net1046));
 sg13g2_antennanp ANTENNA_1883 (.A(net1046));
 sg13g2_antennanp ANTENNA_1884 (.A(net1046));
 sg13g2_antennanp ANTENNA_1885 (.A(net1046));
 sg13g2_antennanp ANTENNA_1886 (.A(net1046));
 sg13g2_antennanp ANTENNA_1887 (.A(net1046));
 sg13g2_antennanp ANTENNA_1888 (.A(net1046));
 sg13g2_antennanp ANTENNA_1889 (.A(net1046));
 sg13g2_antennanp ANTENNA_1890 (.A(net1056));
 sg13g2_antennanp ANTENNA_1891 (.A(net1056));
 sg13g2_antennanp ANTENNA_1892 (.A(net1056));
 sg13g2_antennanp ANTENNA_1893 (.A(net1056));
 sg13g2_antennanp ANTENNA_1894 (.A(net1056));
 sg13g2_antennanp ANTENNA_1895 (.A(net1056));
 sg13g2_antennanp ANTENNA_1896 (.A(net1056));
 sg13g2_antennanp ANTENNA_1897 (.A(net1056));
 sg13g2_antennanp ANTENNA_1898 (.A(net1056));
 sg13g2_antennanp ANTENNA_1899 (.A(net1056));
 sg13g2_antennanp ANTENNA_1900 (.A(net1056));
 sg13g2_antennanp ANTENNA_1901 (.A(net1056));
 sg13g2_antennanp ANTENNA_1902 (.A(_00054_));
 sg13g2_antennanp ANTENNA_1903 (.A(_00201_));
 sg13g2_antennanp ANTENNA_1904 (.A(_00207_));
 sg13g2_antennanp ANTENNA_1905 (.A(_00235_));
 sg13g2_antennanp ANTENNA_1906 (.A(_00727_));
 sg13g2_antennanp ANTENNA_1907 (.A(_00769_));
 sg13g2_antennanp ANTENNA_1908 (.A(_00905_));
 sg13g2_antennanp ANTENNA_1909 (.A(_00964_));
 sg13g2_antennanp ANTENNA_1910 (.A(_00964_));
 sg13g2_antennanp ANTENNA_1911 (.A(_01048_));
 sg13g2_antennanp ANTENNA_1912 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1913 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1914 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1915 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1916 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1917 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1918 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1919 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1920 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1921 (.A(_02963_));
 sg13g2_antennanp ANTENNA_1922 (.A(_02963_));
 sg13g2_antennanp ANTENNA_1923 (.A(_02963_));
 sg13g2_antennanp ANTENNA_1924 (.A(_02963_));
 sg13g2_antennanp ANTENNA_1925 (.A(_03093_));
 sg13g2_antennanp ANTENNA_1926 (.A(_03093_));
 sg13g2_antennanp ANTENNA_1927 (.A(_03093_));
 sg13g2_antennanp ANTENNA_1928 (.A(_03093_));
 sg13g2_antennanp ANTENNA_1929 (.A(_03093_));
 sg13g2_antennanp ANTENNA_1930 (.A(_03093_));
 sg13g2_antennanp ANTENNA_1931 (.A(_03093_));
 sg13g2_antennanp ANTENNA_1932 (.A(_03093_));
 sg13g2_antennanp ANTENNA_1933 (.A(_03093_));
 sg13g2_antennanp ANTENNA_1934 (.A(_03096_));
 sg13g2_antennanp ANTENNA_1935 (.A(_03096_));
 sg13g2_antennanp ANTENNA_1936 (.A(_03096_));
 sg13g2_antennanp ANTENNA_1937 (.A(_03096_));
 sg13g2_antennanp ANTENNA_1938 (.A(_03096_));
 sg13g2_antennanp ANTENNA_1939 (.A(_03096_));
 sg13g2_antennanp ANTENNA_1940 (.A(_03096_));
 sg13g2_antennanp ANTENNA_1941 (.A(_03096_));
 sg13g2_antennanp ANTENNA_1942 (.A(_03096_));
 sg13g2_antennanp ANTENNA_1943 (.A(_03107_));
 sg13g2_antennanp ANTENNA_1944 (.A(_03107_));
 sg13g2_antennanp ANTENNA_1945 (.A(_03107_));
 sg13g2_antennanp ANTENNA_1946 (.A(_03107_));
 sg13g2_antennanp ANTENNA_1947 (.A(_03107_));
 sg13g2_antennanp ANTENNA_1948 (.A(_03108_));
 sg13g2_antennanp ANTENNA_1949 (.A(_03108_));
 sg13g2_antennanp ANTENNA_1950 (.A(_03108_));
 sg13g2_antennanp ANTENNA_1951 (.A(_03108_));
 sg13g2_antennanp ANTENNA_1952 (.A(_03108_));
 sg13g2_antennanp ANTENNA_1953 (.A(_03108_));
 sg13g2_antennanp ANTENNA_1954 (.A(_03108_));
 sg13g2_antennanp ANTENNA_1955 (.A(_03108_));
 sg13g2_antennanp ANTENNA_1956 (.A(_03108_));
 sg13g2_antennanp ANTENNA_1957 (.A(_03133_));
 sg13g2_antennanp ANTENNA_1958 (.A(_03133_));
 sg13g2_antennanp ANTENNA_1959 (.A(_03133_));
 sg13g2_antennanp ANTENNA_1960 (.A(_03133_));
 sg13g2_antennanp ANTENNA_1961 (.A(_03212_));
 sg13g2_antennanp ANTENNA_1962 (.A(_03229_));
 sg13g2_antennanp ANTENNA_1963 (.A(_03229_));
 sg13g2_antennanp ANTENNA_1964 (.A(_03642_));
 sg13g2_antennanp ANTENNA_1965 (.A(_03642_));
 sg13g2_antennanp ANTENNA_1966 (.A(_03642_));
 sg13g2_antennanp ANTENNA_1967 (.A(_03647_));
 sg13g2_antennanp ANTENNA_1968 (.A(_03647_));
 sg13g2_antennanp ANTENNA_1969 (.A(_03647_));
 sg13g2_antennanp ANTENNA_1970 (.A(_03647_));
 sg13g2_antennanp ANTENNA_1971 (.A(_03653_));
 sg13g2_antennanp ANTENNA_1972 (.A(_03653_));
 sg13g2_antennanp ANTENNA_1973 (.A(_03653_));
 sg13g2_antennanp ANTENNA_1974 (.A(_03653_));
 sg13g2_antennanp ANTENNA_1975 (.A(_03653_));
 sg13g2_antennanp ANTENNA_1976 (.A(_03653_));
 sg13g2_antennanp ANTENNA_1977 (.A(_03653_));
 sg13g2_antennanp ANTENNA_1978 (.A(_03653_));
 sg13g2_antennanp ANTENNA_1979 (.A(_03653_));
 sg13g2_antennanp ANTENNA_1980 (.A(_03657_));
 sg13g2_antennanp ANTENNA_1981 (.A(_03657_));
 sg13g2_antennanp ANTENNA_1982 (.A(_03657_));
 sg13g2_antennanp ANTENNA_1983 (.A(_03657_));
 sg13g2_antennanp ANTENNA_1984 (.A(_03657_));
 sg13g2_antennanp ANTENNA_1985 (.A(_03657_));
 sg13g2_antennanp ANTENNA_1986 (.A(_03657_));
 sg13g2_antennanp ANTENNA_1987 (.A(_03657_));
 sg13g2_antennanp ANTENNA_1988 (.A(_03657_));
 sg13g2_antennanp ANTENNA_1989 (.A(_04770_));
 sg13g2_antennanp ANTENNA_1990 (.A(_04770_));
 sg13g2_antennanp ANTENNA_1991 (.A(_04770_));
 sg13g2_antennanp ANTENNA_1992 (.A(_04770_));
 sg13g2_antennanp ANTENNA_1993 (.A(_04848_));
 sg13g2_antennanp ANTENNA_1994 (.A(_04848_));
 sg13g2_antennanp ANTENNA_1995 (.A(_05001_));
 sg13g2_antennanp ANTENNA_1996 (.A(_05431_));
 sg13g2_antennanp ANTENNA_1997 (.A(_05642_));
 sg13g2_antennanp ANTENNA_1998 (.A(_05753_));
 sg13g2_antennanp ANTENNA_1999 (.A(_05753_));
 sg13g2_antennanp ANTENNA_2000 (.A(_05753_));
 sg13g2_antennanp ANTENNA_2001 (.A(_05753_));
 sg13g2_antennanp ANTENNA_2002 (.A(_05754_));
 sg13g2_antennanp ANTENNA_2003 (.A(_05754_));
 sg13g2_antennanp ANTENNA_2004 (.A(_05754_));
 sg13g2_antennanp ANTENNA_2005 (.A(_05754_));
 sg13g2_antennanp ANTENNA_2006 (.A(_05766_));
 sg13g2_antennanp ANTENNA_2007 (.A(_05771_));
 sg13g2_antennanp ANTENNA_2008 (.A(_05773_));
 sg13g2_antennanp ANTENNA_2009 (.A(_05778_));
 sg13g2_antennanp ANTENNA_2010 (.A(_05782_));
 sg13g2_antennanp ANTENNA_2011 (.A(_05782_));
 sg13g2_antennanp ANTENNA_2012 (.A(_05782_));
 sg13g2_antennanp ANTENNA_2013 (.A(_05782_));
 sg13g2_antennanp ANTENNA_2014 (.A(_05786_));
 sg13g2_antennanp ANTENNA_2015 (.A(_05791_));
 sg13g2_antennanp ANTENNA_2016 (.A(_06137_));
 sg13g2_antennanp ANTENNA_2017 (.A(_06137_));
 sg13g2_antennanp ANTENNA_2018 (.A(_06137_));
 sg13g2_antennanp ANTENNA_2019 (.A(_06137_));
 sg13g2_antennanp ANTENNA_2020 (.A(_06137_));
 sg13g2_antennanp ANTENNA_2021 (.A(_06137_));
 sg13g2_antennanp ANTENNA_2022 (.A(_06386_));
 sg13g2_antennanp ANTENNA_2023 (.A(_06386_));
 sg13g2_antennanp ANTENNA_2024 (.A(_06386_));
 sg13g2_antennanp ANTENNA_2025 (.A(_06386_));
 sg13g2_antennanp ANTENNA_2026 (.A(_06386_));
 sg13g2_antennanp ANTENNA_2027 (.A(_06386_));
 sg13g2_antennanp ANTENNA_2028 (.A(_06386_));
 sg13g2_antennanp ANTENNA_2029 (.A(_06386_));
 sg13g2_antennanp ANTENNA_2030 (.A(_06386_));
 sg13g2_antennanp ANTENNA_2031 (.A(_07450_));
 sg13g2_antennanp ANTENNA_2032 (.A(_07450_));
 sg13g2_antennanp ANTENNA_2033 (.A(_07450_));
 sg13g2_antennanp ANTENNA_2034 (.A(_08133_));
 sg13g2_antennanp ANTENNA_2035 (.A(_08133_));
 sg13g2_antennanp ANTENNA_2036 (.A(_08133_));
 sg13g2_antennanp ANTENNA_2037 (.A(_08133_));
 sg13g2_antennanp ANTENNA_2038 (.A(_08133_));
 sg13g2_antennanp ANTENNA_2039 (.A(_08133_));
 sg13g2_antennanp ANTENNA_2040 (.A(_08133_));
 sg13g2_antennanp ANTENNA_2041 (.A(_08181_));
 sg13g2_antennanp ANTENNA_2042 (.A(_08181_));
 sg13g2_antennanp ANTENNA_2043 (.A(_08181_));
 sg13g2_antennanp ANTENNA_2044 (.A(_08181_));
 sg13g2_antennanp ANTENNA_2045 (.A(_08181_));
 sg13g2_antennanp ANTENNA_2046 (.A(_08181_));
 sg13g2_antennanp ANTENNA_2047 (.A(_08181_));
 sg13g2_antennanp ANTENNA_2048 (.A(_08192_));
 sg13g2_antennanp ANTENNA_2049 (.A(_08285_));
 sg13g2_antennanp ANTENNA_2050 (.A(_08285_));
 sg13g2_antennanp ANTENNA_2051 (.A(_08285_));
 sg13g2_antennanp ANTENNA_2052 (.A(_08285_));
 sg13g2_antennanp ANTENNA_2053 (.A(_08494_));
 sg13g2_antennanp ANTENNA_2054 (.A(_08494_));
 sg13g2_antennanp ANTENNA_2055 (.A(_08494_));
 sg13g2_antennanp ANTENNA_2056 (.A(_08708_));
 sg13g2_antennanp ANTENNA_2057 (.A(_08708_));
 sg13g2_antennanp ANTENNA_2058 (.A(_08708_));
 sg13g2_antennanp ANTENNA_2059 (.A(_08709_));
 sg13g2_antennanp ANTENNA_2060 (.A(_08709_));
 sg13g2_antennanp ANTENNA_2061 (.A(_08709_));
 sg13g2_antennanp ANTENNA_2062 (.A(_08709_));
 sg13g2_antennanp ANTENNA_2063 (.A(_08801_));
 sg13g2_antennanp ANTENNA_2064 (.A(_08801_));
 sg13g2_antennanp ANTENNA_2065 (.A(_08877_));
 sg13g2_antennanp ANTENNA_2066 (.A(_08877_));
 sg13g2_antennanp ANTENNA_2067 (.A(_08877_));
 sg13g2_antennanp ANTENNA_2068 (.A(_08901_));
 sg13g2_antennanp ANTENNA_2069 (.A(_08901_));
 sg13g2_antennanp ANTENNA_2070 (.A(_08901_));
 sg13g2_antennanp ANTENNA_2071 (.A(_08901_));
 sg13g2_antennanp ANTENNA_2072 (.A(_08964_));
 sg13g2_antennanp ANTENNA_2073 (.A(_08964_));
 sg13g2_antennanp ANTENNA_2074 (.A(_08964_));
 sg13g2_antennanp ANTENNA_2075 (.A(_08964_));
 sg13g2_antennanp ANTENNA_2076 (.A(_08979_));
 sg13g2_antennanp ANTENNA_2077 (.A(_08979_));
 sg13g2_antennanp ANTENNA_2078 (.A(_08979_));
 sg13g2_antennanp ANTENNA_2079 (.A(_08979_));
 sg13g2_antennanp ANTENNA_2080 (.A(_08979_));
 sg13g2_antennanp ANTENNA_2081 (.A(_09008_));
 sg13g2_antennanp ANTENNA_2082 (.A(_09008_));
 sg13g2_antennanp ANTENNA_2083 (.A(_09008_));
 sg13g2_antennanp ANTENNA_2084 (.A(_09008_));
 sg13g2_antennanp ANTENNA_2085 (.A(_09008_));
 sg13g2_antennanp ANTENNA_2086 (.A(_09008_));
 sg13g2_antennanp ANTENNA_2087 (.A(_09025_));
 sg13g2_antennanp ANTENNA_2088 (.A(_09025_));
 sg13g2_antennanp ANTENNA_2089 (.A(_09025_));
 sg13g2_antennanp ANTENNA_2090 (.A(_09025_));
 sg13g2_antennanp ANTENNA_2091 (.A(_09025_));
 sg13g2_antennanp ANTENNA_2092 (.A(_09025_));
 sg13g2_antennanp ANTENNA_2093 (.A(_09025_));
 sg13g2_antennanp ANTENNA_2094 (.A(_09025_));
 sg13g2_antennanp ANTENNA_2095 (.A(_09025_));
 sg13g2_antennanp ANTENNA_2096 (.A(_09036_));
 sg13g2_antennanp ANTENNA_2097 (.A(_09036_));
 sg13g2_antennanp ANTENNA_2098 (.A(_09036_));
 sg13g2_antennanp ANTENNA_2099 (.A(_09036_));
 sg13g2_antennanp ANTENNA_2100 (.A(_09045_));
 sg13g2_antennanp ANTENNA_2101 (.A(_09045_));
 sg13g2_antennanp ANTENNA_2102 (.A(_09118_));
 sg13g2_antennanp ANTENNA_2103 (.A(_09118_));
 sg13g2_antennanp ANTENNA_2104 (.A(_09118_));
 sg13g2_antennanp ANTENNA_2105 (.A(_09118_));
 sg13g2_antennanp ANTENNA_2106 (.A(_09118_));
 sg13g2_antennanp ANTENNA_2107 (.A(_09118_));
 sg13g2_antennanp ANTENNA_2108 (.A(_09122_));
 sg13g2_antennanp ANTENNA_2109 (.A(_09122_));
 sg13g2_antennanp ANTENNA_2110 (.A(_09122_));
 sg13g2_antennanp ANTENNA_2111 (.A(_09124_));
 sg13g2_antennanp ANTENNA_2112 (.A(_09124_));
 sg13g2_antennanp ANTENNA_2113 (.A(_09124_));
 sg13g2_antennanp ANTENNA_2114 (.A(_09124_));
 sg13g2_antennanp ANTENNA_2115 (.A(_09124_));
 sg13g2_antennanp ANTENNA_2116 (.A(_09124_));
 sg13g2_antennanp ANTENNA_2117 (.A(_09124_));
 sg13g2_antennanp ANTENNA_2118 (.A(_09124_));
 sg13g2_antennanp ANTENNA_2119 (.A(_09124_));
 sg13g2_antennanp ANTENNA_2120 (.A(_09166_));
 sg13g2_antennanp ANTENNA_2121 (.A(_09166_));
 sg13g2_antennanp ANTENNA_2122 (.A(_09166_));
 sg13g2_antennanp ANTENNA_2123 (.A(_09166_));
 sg13g2_antennanp ANTENNA_2124 (.A(_09207_));
 sg13g2_antennanp ANTENNA_2125 (.A(_09251_));
 sg13g2_antennanp ANTENNA_2126 (.A(_09251_));
 sg13g2_antennanp ANTENNA_2127 (.A(_09328_));
 sg13g2_antennanp ANTENNA_2128 (.A(_09361_));
 sg13g2_antennanp ANTENNA_2129 (.A(_09361_));
 sg13g2_antennanp ANTENNA_2130 (.A(_09398_));
 sg13g2_antennanp ANTENNA_2131 (.A(_09445_));
 sg13g2_antennanp ANTENNA_2132 (.A(_09485_));
 sg13g2_antennanp ANTENNA_2133 (.A(_09499_));
 sg13g2_antennanp ANTENNA_2134 (.A(_09606_));
 sg13g2_antennanp ANTENNA_2135 (.A(_09637_));
 sg13g2_antennanp ANTENNA_2136 (.A(_09637_));
 sg13g2_antennanp ANTENNA_2137 (.A(_09875_));
 sg13g2_antennanp ANTENNA_2138 (.A(_09875_));
 sg13g2_antennanp ANTENNA_2139 (.A(_09875_));
 sg13g2_antennanp ANTENNA_2140 (.A(_09875_));
 sg13g2_antennanp ANTENNA_2141 (.A(_09875_));
 sg13g2_antennanp ANTENNA_2142 (.A(_09875_));
 sg13g2_antennanp ANTENNA_2143 (.A(_09875_));
 sg13g2_antennanp ANTENNA_2144 (.A(_09875_));
 sg13g2_antennanp ANTENNA_2145 (.A(_09875_));
 sg13g2_antennanp ANTENNA_2146 (.A(_09991_));
 sg13g2_antennanp ANTENNA_2147 (.A(_09991_));
 sg13g2_antennanp ANTENNA_2148 (.A(_09991_));
 sg13g2_antennanp ANTENNA_2149 (.A(_09991_));
 sg13g2_antennanp ANTENNA_2150 (.A(_09991_));
 sg13g2_antennanp ANTENNA_2151 (.A(_09991_));
 sg13g2_antennanp ANTENNA_2152 (.A(_09991_));
 sg13g2_antennanp ANTENNA_2153 (.A(_09991_));
 sg13g2_antennanp ANTENNA_2154 (.A(_10110_));
 sg13g2_antennanp ANTENNA_2155 (.A(_10423_));
 sg13g2_antennanp ANTENNA_2156 (.A(_10423_));
 sg13g2_antennanp ANTENNA_2157 (.A(_10423_));
 sg13g2_antennanp ANTENNA_2158 (.A(_10423_));
 sg13g2_antennanp ANTENNA_2159 (.A(_10831_));
 sg13g2_antennanp ANTENNA_2160 (.A(_10831_));
 sg13g2_antennanp ANTENNA_2161 (.A(_10831_));
 sg13g2_antennanp ANTENNA_2162 (.A(_10831_));
 sg13g2_antennanp ANTENNA_2163 (.A(_10831_));
 sg13g2_antennanp ANTENNA_2164 (.A(_10831_));
 sg13g2_antennanp ANTENNA_2165 (.A(_10831_));
 sg13g2_antennanp ANTENNA_2166 (.A(_10831_));
 sg13g2_antennanp ANTENNA_2167 (.A(_10831_));
 sg13g2_antennanp ANTENNA_2168 (.A(_10963_));
 sg13g2_antennanp ANTENNA_2169 (.A(_10963_));
 sg13g2_antennanp ANTENNA_2170 (.A(_10963_));
 sg13g2_antennanp ANTENNA_2171 (.A(_10963_));
 sg13g2_antennanp ANTENNA_2172 (.A(_11495_));
 sg13g2_antennanp ANTENNA_2173 (.A(_11495_));
 sg13g2_antennanp ANTENNA_2174 (.A(_11495_));
 sg13g2_antennanp ANTENNA_2175 (.A(_11495_));
 sg13g2_antennanp ANTENNA_2176 (.A(_11495_));
 sg13g2_antennanp ANTENNA_2177 (.A(_12007_));
 sg13g2_antennanp ANTENNA_2178 (.A(_12007_));
 sg13g2_antennanp ANTENNA_2179 (.A(_12007_));
 sg13g2_antennanp ANTENNA_2180 (.A(_12007_));
 sg13g2_antennanp ANTENNA_2181 (.A(_12007_));
 sg13g2_antennanp ANTENNA_2182 (.A(_12007_));
 sg13g2_antennanp ANTENNA_2183 (.A(_12007_));
 sg13g2_antennanp ANTENNA_2184 (.A(_12007_));
 sg13g2_antennanp ANTENNA_2185 (.A(_12007_));
 sg13g2_antennanp ANTENNA_2186 (.A(_12031_));
 sg13g2_antennanp ANTENNA_2187 (.A(_12031_));
 sg13g2_antennanp ANTENNA_2188 (.A(_12031_));
 sg13g2_antennanp ANTENNA_2189 (.A(_12031_));
 sg13g2_antennanp ANTENNA_2190 (.A(_12031_));
 sg13g2_antennanp ANTENNA_2191 (.A(_12031_));
 sg13g2_antennanp ANTENNA_2192 (.A(_12031_));
 sg13g2_antennanp ANTENNA_2193 (.A(_12031_));
 sg13g2_antennanp ANTENNA_2194 (.A(_12031_));
 sg13g2_antennanp ANTENNA_2195 (.A(_12047_));
 sg13g2_antennanp ANTENNA_2196 (.A(_12047_));
 sg13g2_antennanp ANTENNA_2197 (.A(_12047_));
 sg13g2_antennanp ANTENNA_2198 (.A(_12047_));
 sg13g2_antennanp ANTENNA_2199 (.A(_12047_));
 sg13g2_antennanp ANTENNA_2200 (.A(_12067_));
 sg13g2_antennanp ANTENNA_2201 (.A(_12067_));
 sg13g2_antennanp ANTENNA_2202 (.A(_12067_));
 sg13g2_antennanp ANTENNA_2203 (.A(_12067_));
 sg13g2_antennanp ANTENNA_2204 (.A(_12067_));
 sg13g2_antennanp ANTENNA_2205 (.A(_12067_));
 sg13g2_antennanp ANTENNA_2206 (.A(_12067_));
 sg13g2_antennanp ANTENNA_2207 (.A(_12067_));
 sg13g2_antennanp ANTENNA_2208 (.A(_12067_));
 sg13g2_antennanp ANTENNA_2209 (.A(_12107_));
 sg13g2_antennanp ANTENNA_2210 (.A(_12107_));
 sg13g2_antennanp ANTENNA_2211 (.A(_12107_));
 sg13g2_antennanp ANTENNA_2212 (.A(_12107_));
 sg13g2_antennanp ANTENNA_2213 (.A(_12136_));
 sg13g2_antennanp ANTENNA_2214 (.A(_12136_));
 sg13g2_antennanp ANTENNA_2215 (.A(_12136_));
 sg13g2_antennanp ANTENNA_2216 (.A(\cpu.dec.r_trap ));
 sg13g2_antennanp ANTENNA_2217 (.A(\cpu.dec.r_trap ));
 sg13g2_antennanp ANTENNA_2218 (.A(\cpu.ex.pc[2] ));
 sg13g2_antennanp ANTENNA_2219 (.A(\cpu.gpio.uart_rx ));
 sg13g2_antennanp ANTENNA_2220 (.A(\cpu.gpio.uart_rx ));
 sg13g2_antennanp ANTENNA_2221 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_2222 (.A(net11));
 sg13g2_antennanp ANTENNA_2223 (.A(net11));
 sg13g2_antennanp ANTENNA_2224 (.A(net11));
 sg13g2_antennanp ANTENNA_2225 (.A(net12));
 sg13g2_antennanp ANTENNA_2226 (.A(net12));
 sg13g2_antennanp ANTENNA_2227 (.A(net12));
 sg13g2_antennanp ANTENNA_2228 (.A(net577));
 sg13g2_antennanp ANTENNA_2229 (.A(net577));
 sg13g2_antennanp ANTENNA_2230 (.A(net577));
 sg13g2_antennanp ANTENNA_2231 (.A(net577));
 sg13g2_antennanp ANTENNA_2232 (.A(net577));
 sg13g2_antennanp ANTENNA_2233 (.A(net577));
 sg13g2_antennanp ANTENNA_2234 (.A(net577));
 sg13g2_antennanp ANTENNA_2235 (.A(net577));
 sg13g2_antennanp ANTENNA_2236 (.A(net577));
 sg13g2_antennanp ANTENNA_2237 (.A(net639));
 sg13g2_antennanp ANTENNA_2238 (.A(net639));
 sg13g2_antennanp ANTENNA_2239 (.A(net639));
 sg13g2_antennanp ANTENNA_2240 (.A(net639));
 sg13g2_antennanp ANTENNA_2241 (.A(net639));
 sg13g2_antennanp ANTENNA_2242 (.A(net639));
 sg13g2_antennanp ANTENNA_2243 (.A(net639));
 sg13g2_antennanp ANTENNA_2244 (.A(net639));
 sg13g2_antennanp ANTENNA_2245 (.A(net639));
 sg13g2_antennanp ANTENNA_2246 (.A(net679));
 sg13g2_antennanp ANTENNA_2247 (.A(net679));
 sg13g2_antennanp ANTENNA_2248 (.A(net679));
 sg13g2_antennanp ANTENNA_2249 (.A(net679));
 sg13g2_antennanp ANTENNA_2250 (.A(net679));
 sg13g2_antennanp ANTENNA_2251 (.A(net679));
 sg13g2_antennanp ANTENNA_2252 (.A(net679));
 sg13g2_antennanp ANTENNA_2253 (.A(net679));
 sg13g2_antennanp ANTENNA_2254 (.A(net679));
 sg13g2_antennanp ANTENNA_2255 (.A(net732));
 sg13g2_antennanp ANTENNA_2256 (.A(net732));
 sg13g2_antennanp ANTENNA_2257 (.A(net732));
 sg13g2_antennanp ANTENNA_2258 (.A(net732));
 sg13g2_antennanp ANTENNA_2259 (.A(net732));
 sg13g2_antennanp ANTENNA_2260 (.A(net732));
 sg13g2_antennanp ANTENNA_2261 (.A(net732));
 sg13g2_antennanp ANTENNA_2262 (.A(net732));
 sg13g2_antennanp ANTENNA_2263 (.A(net732));
 sg13g2_antennanp ANTENNA_2264 (.A(net789));
 sg13g2_antennanp ANTENNA_2265 (.A(net789));
 sg13g2_antennanp ANTENNA_2266 (.A(net789));
 sg13g2_antennanp ANTENNA_2267 (.A(net789));
 sg13g2_antennanp ANTENNA_2268 (.A(net789));
 sg13g2_antennanp ANTENNA_2269 (.A(net789));
 sg13g2_antennanp ANTENNA_2270 (.A(net789));
 sg13g2_antennanp ANTENNA_2271 (.A(net789));
 sg13g2_antennanp ANTENNA_2272 (.A(net789));
 sg13g2_antennanp ANTENNA_2273 (.A(net966));
 sg13g2_antennanp ANTENNA_2274 (.A(net966));
 sg13g2_antennanp ANTENNA_2275 (.A(net966));
 sg13g2_antennanp ANTENNA_2276 (.A(net966));
 sg13g2_antennanp ANTENNA_2277 (.A(net966));
 sg13g2_antennanp ANTENNA_2278 (.A(net966));
 sg13g2_antennanp ANTENNA_2279 (.A(net966));
 sg13g2_antennanp ANTENNA_2280 (.A(net966));
 sg13g2_antennanp ANTENNA_2281 (.A(net966));
 sg13g2_antennanp ANTENNA_2282 (.A(net966));
 sg13g2_antennanp ANTENNA_2283 (.A(net966));
 sg13g2_antennanp ANTENNA_2284 (.A(net966));
 sg13g2_antennanp ANTENNA_2285 (.A(net966));
 sg13g2_antennanp ANTENNA_2286 (.A(net966));
 sg13g2_antennanp ANTENNA_2287 (.A(net966));
 sg13g2_antennanp ANTENNA_2288 (.A(net966));
 sg13g2_antennanp ANTENNA_2289 (.A(net966));
 sg13g2_antennanp ANTENNA_2290 (.A(net966));
 sg13g2_antennanp ANTENNA_2291 (.A(net966));
 sg13g2_antennanp ANTENNA_2292 (.A(net966));
 sg13g2_antennanp ANTENNA_2293 (.A(net966));
 sg13g2_antennanp ANTENNA_2294 (.A(net966));
 sg13g2_antennanp ANTENNA_2295 (.A(net966));
 sg13g2_antennanp ANTENNA_2296 (.A(net966));
 sg13g2_antennanp ANTENNA_2297 (.A(net966));
 sg13g2_antennanp ANTENNA_2298 (.A(net966));
 sg13g2_antennanp ANTENNA_2299 (.A(net966));
 sg13g2_antennanp ANTENNA_2300 (.A(net966));
 sg13g2_antennanp ANTENNA_2301 (.A(net966));
 sg13g2_antennanp ANTENNA_2302 (.A(net966));
 sg13g2_antennanp ANTENNA_2303 (.A(net966));
 sg13g2_antennanp ANTENNA_2304 (.A(net966));
 sg13g2_antennanp ANTENNA_2305 (.A(net966));
 sg13g2_antennanp ANTENNA_2306 (.A(net1046));
 sg13g2_antennanp ANTENNA_2307 (.A(net1046));
 sg13g2_antennanp ANTENNA_2308 (.A(net1046));
 sg13g2_antennanp ANTENNA_2309 (.A(net1046));
 sg13g2_antennanp ANTENNA_2310 (.A(net1046));
 sg13g2_antennanp ANTENNA_2311 (.A(net1046));
 sg13g2_antennanp ANTENNA_2312 (.A(net1046));
 sg13g2_antennanp ANTENNA_2313 (.A(net1046));
 sg13g2_antennanp ANTENNA_2314 (.A(net1056));
 sg13g2_antennanp ANTENNA_2315 (.A(net1056));
 sg13g2_antennanp ANTENNA_2316 (.A(net1056));
 sg13g2_antennanp ANTENNA_2317 (.A(net1056));
 sg13g2_antennanp ANTENNA_2318 (.A(net1056));
 sg13g2_antennanp ANTENNA_2319 (.A(net1056));
 sg13g2_antennanp ANTENNA_2320 (.A(net1056));
 sg13g2_antennanp ANTENNA_2321 (.A(net1056));
 sg13g2_antennanp ANTENNA_2322 (.A(net1056));
 sg13g2_antennanp ANTENNA_2323 (.A(net1056));
 sg13g2_antennanp ANTENNA_2324 (.A(net1056));
 sg13g2_antennanp ANTENNA_2325 (.A(net1056));
 sg13g2_antennanp ANTENNA_2326 (.A(_00054_));
 sg13g2_antennanp ANTENNA_2327 (.A(_00201_));
 sg13g2_antennanp ANTENNA_2328 (.A(_00207_));
 sg13g2_antennanp ANTENNA_2329 (.A(_00235_));
 sg13g2_antennanp ANTENNA_2330 (.A(_00769_));
 sg13g2_antennanp ANTENNA_2331 (.A(_00905_));
 sg13g2_antennanp ANTENNA_2332 (.A(_00964_));
 sg13g2_antennanp ANTENNA_2333 (.A(_00964_));
 sg13g2_antennanp ANTENNA_2334 (.A(_01048_));
 sg13g2_antennanp ANTENNA_2335 (.A(_02918_));
 sg13g2_antennanp ANTENNA_2336 (.A(_02918_));
 sg13g2_antennanp ANTENNA_2337 (.A(_02918_));
 sg13g2_antennanp ANTENNA_2338 (.A(_02918_));
 sg13g2_antennanp ANTENNA_2339 (.A(_02963_));
 sg13g2_antennanp ANTENNA_2340 (.A(_02963_));
 sg13g2_antennanp ANTENNA_2341 (.A(_02963_));
 sg13g2_antennanp ANTENNA_2342 (.A(_02963_));
 sg13g2_antennanp ANTENNA_2343 (.A(_03093_));
 sg13g2_antennanp ANTENNA_2344 (.A(_03093_));
 sg13g2_antennanp ANTENNA_2345 (.A(_03093_));
 sg13g2_antennanp ANTENNA_2346 (.A(_03093_));
 sg13g2_antennanp ANTENNA_2347 (.A(_03093_));
 sg13g2_antennanp ANTENNA_2348 (.A(_03093_));
 sg13g2_antennanp ANTENNA_2349 (.A(_03093_));
 sg13g2_antennanp ANTENNA_2350 (.A(_03093_));
 sg13g2_antennanp ANTENNA_2351 (.A(_03093_));
 sg13g2_antennanp ANTENNA_2352 (.A(_03093_));
 sg13g2_antennanp ANTENNA_2353 (.A(_03096_));
 sg13g2_antennanp ANTENNA_2354 (.A(_03096_));
 sg13g2_antennanp ANTENNA_2355 (.A(_03096_));
 sg13g2_antennanp ANTENNA_2356 (.A(_03096_));
 sg13g2_antennanp ANTENNA_2357 (.A(_03096_));
 sg13g2_antennanp ANTENNA_2358 (.A(_03096_));
 sg13g2_antennanp ANTENNA_2359 (.A(_03096_));
 sg13g2_antennanp ANTENNA_2360 (.A(_03096_));
 sg13g2_antennanp ANTENNA_2361 (.A(_03096_));
 sg13g2_antennanp ANTENNA_2362 (.A(_03107_));
 sg13g2_antennanp ANTENNA_2363 (.A(_03107_));
 sg13g2_antennanp ANTENNA_2364 (.A(_03107_));
 sg13g2_antennanp ANTENNA_2365 (.A(_03107_));
 sg13g2_antennanp ANTENNA_2366 (.A(_03107_));
 sg13g2_antennanp ANTENNA_2367 (.A(_03108_));
 sg13g2_antennanp ANTENNA_2368 (.A(_03108_));
 sg13g2_antennanp ANTENNA_2369 (.A(_03108_));
 sg13g2_antennanp ANTENNA_2370 (.A(_03108_));
 sg13g2_antennanp ANTENNA_2371 (.A(_03108_));
 sg13g2_antennanp ANTENNA_2372 (.A(_03108_));
 sg13g2_antennanp ANTENNA_2373 (.A(_03108_));
 sg13g2_antennanp ANTENNA_2374 (.A(_03108_));
 sg13g2_antennanp ANTENNA_2375 (.A(_03108_));
 sg13g2_antennanp ANTENNA_2376 (.A(_03133_));
 sg13g2_antennanp ANTENNA_2377 (.A(_03133_));
 sg13g2_antennanp ANTENNA_2378 (.A(_03133_));
 sg13g2_antennanp ANTENNA_2379 (.A(_03133_));
 sg13g2_antennanp ANTENNA_2380 (.A(_03133_));
 sg13g2_antennanp ANTENNA_2381 (.A(_03133_));
 sg13g2_antennanp ANTENNA_2382 (.A(_03133_));
 sg13g2_antennanp ANTENNA_2383 (.A(_03133_));
 sg13g2_antennanp ANTENNA_2384 (.A(_03133_));
 sg13g2_antennanp ANTENNA_2385 (.A(_03212_));
 sg13g2_antennanp ANTENNA_2386 (.A(_03229_));
 sg13g2_antennanp ANTENNA_2387 (.A(_03229_));
 sg13g2_antennanp ANTENNA_2388 (.A(_03642_));
 sg13g2_antennanp ANTENNA_2389 (.A(_03642_));
 sg13g2_antennanp ANTENNA_2390 (.A(_03642_));
 sg13g2_antennanp ANTENNA_2391 (.A(_03647_));
 sg13g2_antennanp ANTENNA_2392 (.A(_03647_));
 sg13g2_antennanp ANTENNA_2393 (.A(_03647_));
 sg13g2_antennanp ANTENNA_2394 (.A(_03647_));
 sg13g2_antennanp ANTENNA_2395 (.A(_03653_));
 sg13g2_antennanp ANTENNA_2396 (.A(_03653_));
 sg13g2_antennanp ANTENNA_2397 (.A(_03653_));
 sg13g2_antennanp ANTENNA_2398 (.A(_03653_));
 sg13g2_antennanp ANTENNA_2399 (.A(_03653_));
 sg13g2_antennanp ANTENNA_2400 (.A(_03653_));
 sg13g2_antennanp ANTENNA_2401 (.A(_03653_));
 sg13g2_antennanp ANTENNA_2402 (.A(_03653_));
 sg13g2_antennanp ANTENNA_2403 (.A(_03653_));
 sg13g2_antennanp ANTENNA_2404 (.A(_03657_));
 sg13g2_antennanp ANTENNA_2405 (.A(_03657_));
 sg13g2_antennanp ANTENNA_2406 (.A(_03657_));
 sg13g2_antennanp ANTENNA_2407 (.A(_03657_));
 sg13g2_antennanp ANTENNA_2408 (.A(_03657_));
 sg13g2_antennanp ANTENNA_2409 (.A(_03657_));
 sg13g2_antennanp ANTENNA_2410 (.A(_03657_));
 sg13g2_antennanp ANTENNA_2411 (.A(_03657_));
 sg13g2_antennanp ANTENNA_2412 (.A(_03657_));
 sg13g2_antennanp ANTENNA_2413 (.A(_04770_));
 sg13g2_antennanp ANTENNA_2414 (.A(_04770_));
 sg13g2_antennanp ANTENNA_2415 (.A(_04770_));
 sg13g2_antennanp ANTENNA_2416 (.A(_04770_));
 sg13g2_antennanp ANTENNA_2417 (.A(_04848_));
 sg13g2_antennanp ANTENNA_2418 (.A(_04848_));
 sg13g2_antennanp ANTENNA_2419 (.A(_05001_));
 sg13g2_antennanp ANTENNA_2420 (.A(_05753_));
 sg13g2_antennanp ANTENNA_2421 (.A(_05753_));
 sg13g2_antennanp ANTENNA_2422 (.A(_05753_));
 sg13g2_antennanp ANTENNA_2423 (.A(_05753_));
 sg13g2_antennanp ANTENNA_2424 (.A(_05766_));
 sg13g2_antennanp ANTENNA_2425 (.A(_05771_));
 sg13g2_antennanp ANTENNA_2426 (.A(_05773_));
 sg13g2_antennanp ANTENNA_2427 (.A(_05778_));
 sg13g2_antennanp ANTENNA_2428 (.A(_05782_));
 sg13g2_antennanp ANTENNA_2429 (.A(_05782_));
 sg13g2_antennanp ANTENNA_2430 (.A(_05782_));
 sg13g2_antennanp ANTENNA_2431 (.A(_05782_));
 sg13g2_antennanp ANTENNA_2432 (.A(_05786_));
 sg13g2_antennanp ANTENNA_2433 (.A(_05791_));
 sg13g2_antennanp ANTENNA_2434 (.A(_06137_));
 sg13g2_antennanp ANTENNA_2435 (.A(_06137_));
 sg13g2_antennanp ANTENNA_2436 (.A(_06137_));
 sg13g2_antennanp ANTENNA_2437 (.A(_06137_));
 sg13g2_antennanp ANTENNA_2438 (.A(_06137_));
 sg13g2_antennanp ANTENNA_2439 (.A(_06137_));
 sg13g2_antennanp ANTENNA_2440 (.A(_06304_));
 sg13g2_antennanp ANTENNA_2441 (.A(_06304_));
 sg13g2_antennanp ANTENNA_2442 (.A(_06304_));
 sg13g2_antennanp ANTENNA_2443 (.A(_06304_));
 sg13g2_antennanp ANTENNA_2444 (.A(_06386_));
 sg13g2_antennanp ANTENNA_2445 (.A(_06386_));
 sg13g2_antennanp ANTENNA_2446 (.A(_06386_));
 sg13g2_antennanp ANTENNA_2447 (.A(_06386_));
 sg13g2_antennanp ANTENNA_2448 (.A(_06386_));
 sg13g2_antennanp ANTENNA_2449 (.A(_06386_));
 sg13g2_antennanp ANTENNA_2450 (.A(_06386_));
 sg13g2_antennanp ANTENNA_2451 (.A(_06386_));
 sg13g2_antennanp ANTENNA_2452 (.A(_06386_));
 sg13g2_antennanp ANTENNA_2453 (.A(_07450_));
 sg13g2_antennanp ANTENNA_2454 (.A(_07450_));
 sg13g2_antennanp ANTENNA_2455 (.A(_07450_));
 sg13g2_antennanp ANTENNA_2456 (.A(_08133_));
 sg13g2_antennanp ANTENNA_2457 (.A(_08133_));
 sg13g2_antennanp ANTENNA_2458 (.A(_08133_));
 sg13g2_antennanp ANTENNA_2459 (.A(_08133_));
 sg13g2_antennanp ANTENNA_2460 (.A(_08133_));
 sg13g2_antennanp ANTENNA_2461 (.A(_08133_));
 sg13g2_antennanp ANTENNA_2462 (.A(_08133_));
 sg13g2_antennanp ANTENNA_2463 (.A(_08181_));
 sg13g2_antennanp ANTENNA_2464 (.A(_08181_));
 sg13g2_antennanp ANTENNA_2465 (.A(_08181_));
 sg13g2_antennanp ANTENNA_2466 (.A(_08181_));
 sg13g2_antennanp ANTENNA_2467 (.A(_08181_));
 sg13g2_antennanp ANTENNA_2468 (.A(_08181_));
 sg13g2_antennanp ANTENNA_2469 (.A(_08181_));
 sg13g2_antennanp ANTENNA_2470 (.A(_08192_));
 sg13g2_antennanp ANTENNA_2471 (.A(_08285_));
 sg13g2_antennanp ANTENNA_2472 (.A(_08285_));
 sg13g2_antennanp ANTENNA_2473 (.A(_08285_));
 sg13g2_antennanp ANTENNA_2474 (.A(_08285_));
 sg13g2_antennanp ANTENNA_2475 (.A(_08447_));
 sg13g2_antennanp ANTENNA_2476 (.A(_08447_));
 sg13g2_antennanp ANTENNA_2477 (.A(_08447_));
 sg13g2_antennanp ANTENNA_2478 (.A(_08494_));
 sg13g2_antennanp ANTENNA_2479 (.A(_08494_));
 sg13g2_antennanp ANTENNA_2480 (.A(_08494_));
 sg13g2_antennanp ANTENNA_2481 (.A(_08705_));
 sg13g2_antennanp ANTENNA_2482 (.A(_08705_));
 sg13g2_antennanp ANTENNA_2483 (.A(_08705_));
 sg13g2_antennanp ANTENNA_2484 (.A(_08708_));
 sg13g2_antennanp ANTENNA_2485 (.A(_08708_));
 sg13g2_antennanp ANTENNA_2486 (.A(_08708_));
 sg13g2_antennanp ANTENNA_2487 (.A(_08709_));
 sg13g2_antennanp ANTENNA_2488 (.A(_08709_));
 sg13g2_antennanp ANTENNA_2489 (.A(_08709_));
 sg13g2_antennanp ANTENNA_2490 (.A(_08709_));
 sg13g2_antennanp ANTENNA_2491 (.A(_08801_));
 sg13g2_antennanp ANTENNA_2492 (.A(_08801_));
 sg13g2_antennanp ANTENNA_2493 (.A(_08901_));
 sg13g2_antennanp ANTENNA_2494 (.A(_08901_));
 sg13g2_antennanp ANTENNA_2495 (.A(_08901_));
 sg13g2_antennanp ANTENNA_2496 (.A(_08901_));
 sg13g2_antennanp ANTENNA_2497 (.A(_08964_));
 sg13g2_antennanp ANTENNA_2498 (.A(_08964_));
 sg13g2_antennanp ANTENNA_2499 (.A(_08964_));
 sg13g2_antennanp ANTENNA_2500 (.A(_08964_));
 sg13g2_antennanp ANTENNA_2501 (.A(_08979_));
 sg13g2_antennanp ANTENNA_2502 (.A(_08979_));
 sg13g2_antennanp ANTENNA_2503 (.A(_08979_));
 sg13g2_antennanp ANTENNA_2504 (.A(_08979_));
 sg13g2_antennanp ANTENNA_2505 (.A(_08979_));
 sg13g2_antennanp ANTENNA_2506 (.A(_09008_));
 sg13g2_antennanp ANTENNA_2507 (.A(_09008_));
 sg13g2_antennanp ANTENNA_2508 (.A(_09008_));
 sg13g2_antennanp ANTENNA_2509 (.A(_09008_));
 sg13g2_antennanp ANTENNA_2510 (.A(_09008_));
 sg13g2_antennanp ANTENNA_2511 (.A(_09008_));
 sg13g2_antennanp ANTENNA_2512 (.A(_09025_));
 sg13g2_antennanp ANTENNA_2513 (.A(_09025_));
 sg13g2_antennanp ANTENNA_2514 (.A(_09025_));
 sg13g2_antennanp ANTENNA_2515 (.A(_09025_));
 sg13g2_antennanp ANTENNA_2516 (.A(_09025_));
 sg13g2_antennanp ANTENNA_2517 (.A(_09025_));
 sg13g2_antennanp ANTENNA_2518 (.A(_09025_));
 sg13g2_antennanp ANTENNA_2519 (.A(_09025_));
 sg13g2_antennanp ANTENNA_2520 (.A(_09025_));
 sg13g2_antennanp ANTENNA_2521 (.A(_09045_));
 sg13g2_antennanp ANTENNA_2522 (.A(_09045_));
 sg13g2_antennanp ANTENNA_2523 (.A(_09118_));
 sg13g2_antennanp ANTENNA_2524 (.A(_09118_));
 sg13g2_antennanp ANTENNA_2525 (.A(_09118_));
 sg13g2_antennanp ANTENNA_2526 (.A(_09118_));
 sg13g2_antennanp ANTENNA_2527 (.A(_09118_));
 sg13g2_antennanp ANTENNA_2528 (.A(_09118_));
 sg13g2_antennanp ANTENNA_2529 (.A(_09118_));
 sg13g2_antennanp ANTENNA_2530 (.A(_09118_));
 sg13g2_antennanp ANTENNA_2531 (.A(_09118_));
 sg13g2_antennanp ANTENNA_2532 (.A(_09118_));
 sg13g2_antennanp ANTENNA_2533 (.A(_09118_));
 sg13g2_antennanp ANTENNA_2534 (.A(_09166_));
 sg13g2_antennanp ANTENNA_2535 (.A(_09166_));
 sg13g2_antennanp ANTENNA_2536 (.A(_09166_));
 sg13g2_antennanp ANTENNA_2537 (.A(_09166_));
 sg13g2_antennanp ANTENNA_2538 (.A(_09251_));
 sg13g2_antennanp ANTENNA_2539 (.A(_09251_));
 sg13g2_antennanp ANTENNA_2540 (.A(_09328_));
 sg13g2_antennanp ANTENNA_2541 (.A(_09361_));
 sg13g2_antennanp ANTENNA_2542 (.A(_09398_));
 sg13g2_antennanp ANTENNA_2543 (.A(_09417_));
 sg13g2_antennanp ANTENNA_2544 (.A(_09417_));
 sg13g2_antennanp ANTENNA_2545 (.A(_09417_));
 sg13g2_antennanp ANTENNA_2546 (.A(_09417_));
 sg13g2_antennanp ANTENNA_2547 (.A(_09445_));
 sg13g2_antennanp ANTENNA_2548 (.A(_09445_));
 sg13g2_antennanp ANTENNA_2549 (.A(_09485_));
 sg13g2_antennanp ANTENNA_2550 (.A(_09606_));
 sg13g2_antennanp ANTENNA_2551 (.A(_09637_));
 sg13g2_antennanp ANTENNA_2552 (.A(_09875_));
 sg13g2_antennanp ANTENNA_2553 (.A(_09875_));
 sg13g2_antennanp ANTENNA_2554 (.A(_09875_));
 sg13g2_antennanp ANTENNA_2555 (.A(_09875_));
 sg13g2_antennanp ANTENNA_2556 (.A(_09875_));
 sg13g2_antennanp ANTENNA_2557 (.A(_09875_));
 sg13g2_antennanp ANTENNA_2558 (.A(_09875_));
 sg13g2_antennanp ANTENNA_2559 (.A(_09875_));
 sg13g2_antennanp ANTENNA_2560 (.A(_09875_));
 sg13g2_antennanp ANTENNA_2561 (.A(_09991_));
 sg13g2_antennanp ANTENNA_2562 (.A(_09991_));
 sg13g2_antennanp ANTENNA_2563 (.A(_09991_));
 sg13g2_antennanp ANTENNA_2564 (.A(_09991_));
 sg13g2_antennanp ANTENNA_2565 (.A(_09991_));
 sg13g2_antennanp ANTENNA_2566 (.A(_09991_));
 sg13g2_antennanp ANTENNA_2567 (.A(_09991_));
 sg13g2_antennanp ANTENNA_2568 (.A(_09991_));
 sg13g2_antennanp ANTENNA_2569 (.A(_10110_));
 sg13g2_antennanp ANTENNA_2570 (.A(_10423_));
 sg13g2_antennanp ANTENNA_2571 (.A(_10423_));
 sg13g2_antennanp ANTENNA_2572 (.A(_10423_));
 sg13g2_antennanp ANTENNA_2573 (.A(_10423_));
 sg13g2_antennanp ANTENNA_2574 (.A(_10831_));
 sg13g2_antennanp ANTENNA_2575 (.A(_10831_));
 sg13g2_antennanp ANTENNA_2576 (.A(_10831_));
 sg13g2_antennanp ANTENNA_2577 (.A(_10831_));
 sg13g2_antennanp ANTENNA_2578 (.A(_10831_));
 sg13g2_antennanp ANTENNA_2579 (.A(_10831_));
 sg13g2_antennanp ANTENNA_2580 (.A(_10831_));
 sg13g2_antennanp ANTENNA_2581 (.A(_10831_));
 sg13g2_antennanp ANTENNA_2582 (.A(_10831_));
 sg13g2_antennanp ANTENNA_2583 (.A(_10831_));
 sg13g2_antennanp ANTENNA_2584 (.A(_10831_));
 sg13g2_antennanp ANTENNA_2585 (.A(_10831_));
 sg13g2_antennanp ANTENNA_2586 (.A(_10831_));
 sg13g2_antennanp ANTENNA_2587 (.A(_10831_));
 sg13g2_antennanp ANTENNA_2588 (.A(_10831_));
 sg13g2_antennanp ANTENNA_2589 (.A(_10831_));
 sg13g2_antennanp ANTENNA_2590 (.A(_10831_));
 sg13g2_antennanp ANTENNA_2591 (.A(_10963_));
 sg13g2_antennanp ANTENNA_2592 (.A(_10963_));
 sg13g2_antennanp ANTENNA_2593 (.A(_10963_));
 sg13g2_antennanp ANTENNA_2594 (.A(_10963_));
 sg13g2_antennanp ANTENNA_2595 (.A(_11495_));
 sg13g2_antennanp ANTENNA_2596 (.A(_11495_));
 sg13g2_antennanp ANTENNA_2597 (.A(_11495_));
 sg13g2_antennanp ANTENNA_2598 (.A(_11495_));
 sg13g2_antennanp ANTENNA_2599 (.A(_11495_));
 sg13g2_antennanp ANTENNA_2600 (.A(_12007_));
 sg13g2_antennanp ANTENNA_2601 (.A(_12007_));
 sg13g2_antennanp ANTENNA_2602 (.A(_12007_));
 sg13g2_antennanp ANTENNA_2603 (.A(_12007_));
 sg13g2_antennanp ANTENNA_2604 (.A(_12007_));
 sg13g2_antennanp ANTENNA_2605 (.A(_12007_));
 sg13g2_antennanp ANTENNA_2606 (.A(_12007_));
 sg13g2_antennanp ANTENNA_2607 (.A(_12007_));
 sg13g2_antennanp ANTENNA_2608 (.A(_12007_));
 sg13g2_antennanp ANTENNA_2609 (.A(_12031_));
 sg13g2_antennanp ANTENNA_2610 (.A(_12031_));
 sg13g2_antennanp ANTENNA_2611 (.A(_12031_));
 sg13g2_antennanp ANTENNA_2612 (.A(_12031_));
 sg13g2_antennanp ANTENNA_2613 (.A(_12031_));
 sg13g2_antennanp ANTENNA_2614 (.A(_12031_));
 sg13g2_antennanp ANTENNA_2615 (.A(_12031_));
 sg13g2_antennanp ANTENNA_2616 (.A(_12031_));
 sg13g2_antennanp ANTENNA_2617 (.A(_12031_));
 sg13g2_antennanp ANTENNA_2618 (.A(_12047_));
 sg13g2_antennanp ANTENNA_2619 (.A(_12047_));
 sg13g2_antennanp ANTENNA_2620 (.A(_12047_));
 sg13g2_antennanp ANTENNA_2621 (.A(_12047_));
 sg13g2_antennanp ANTENNA_2622 (.A(_12047_));
 sg13g2_antennanp ANTENNA_2623 (.A(_12047_));
 sg13g2_antennanp ANTENNA_2624 (.A(_12047_));
 sg13g2_antennanp ANTENNA_2625 (.A(_12047_));
 sg13g2_antennanp ANTENNA_2626 (.A(_12047_));
 sg13g2_antennanp ANTENNA_2627 (.A(_12067_));
 sg13g2_antennanp ANTENNA_2628 (.A(_12067_));
 sg13g2_antennanp ANTENNA_2629 (.A(_12067_));
 sg13g2_antennanp ANTENNA_2630 (.A(_12067_));
 sg13g2_antennanp ANTENNA_2631 (.A(_12067_));
 sg13g2_antennanp ANTENNA_2632 (.A(_12067_));
 sg13g2_antennanp ANTENNA_2633 (.A(_12067_));
 sg13g2_antennanp ANTENNA_2634 (.A(_12067_));
 sg13g2_antennanp ANTENNA_2635 (.A(_12067_));
 sg13g2_antennanp ANTENNA_2636 (.A(_12107_));
 sg13g2_antennanp ANTENNA_2637 (.A(_12107_));
 sg13g2_antennanp ANTENNA_2638 (.A(_12107_));
 sg13g2_antennanp ANTENNA_2639 (.A(_12107_));
 sg13g2_antennanp ANTENNA_2640 (.A(_12107_));
 sg13g2_antennanp ANTENNA_2641 (.A(_12107_));
 sg13g2_antennanp ANTENNA_2642 (.A(_12107_));
 sg13g2_antennanp ANTENNA_2643 (.A(_12107_));
 sg13g2_antennanp ANTENNA_2644 (.A(_12107_));
 sg13g2_antennanp ANTENNA_2645 (.A(_12136_));
 sg13g2_antennanp ANTENNA_2646 (.A(_12136_));
 sg13g2_antennanp ANTENNA_2647 (.A(_12136_));
 sg13g2_antennanp ANTENNA_2648 (.A(\cpu.dec.r_trap ));
 sg13g2_antennanp ANTENNA_2649 (.A(\cpu.ex.pc[2] ));
 sg13g2_antennanp ANTENNA_2650 (.A(\cpu.gpio.uart_rx ));
 sg13g2_antennanp ANTENNA_2651 (.A(\cpu.gpio.uart_rx ));
 sg13g2_antennanp ANTENNA_2652 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_2653 (.A(net11));
 sg13g2_antennanp ANTENNA_2654 (.A(net11));
 sg13g2_antennanp ANTENNA_2655 (.A(net11));
 sg13g2_antennanp ANTENNA_2656 (.A(net12));
 sg13g2_antennanp ANTENNA_2657 (.A(net12));
 sg13g2_antennanp ANTENNA_2658 (.A(net12));
 sg13g2_antennanp ANTENNA_2659 (.A(net13));
 sg13g2_antennanp ANTENNA_2660 (.A(net13));
 sg13g2_antennanp ANTENNA_2661 (.A(net410));
 sg13g2_antennanp ANTENNA_2662 (.A(net410));
 sg13g2_antennanp ANTENNA_2663 (.A(net410));
 sg13g2_antennanp ANTENNA_2664 (.A(net410));
 sg13g2_antennanp ANTENNA_2665 (.A(net410));
 sg13g2_antennanp ANTENNA_2666 (.A(net410));
 sg13g2_antennanp ANTENNA_2667 (.A(net410));
 sg13g2_antennanp ANTENNA_2668 (.A(net410));
 sg13g2_antennanp ANTENNA_2669 (.A(net410));
 sg13g2_antennanp ANTENNA_2670 (.A(net410));
 sg13g2_antennanp ANTENNA_2671 (.A(net410));
 sg13g2_antennanp ANTENNA_2672 (.A(net410));
 sg13g2_antennanp ANTENNA_2673 (.A(net410));
 sg13g2_antennanp ANTENNA_2674 (.A(net410));
 sg13g2_antennanp ANTENNA_2675 (.A(net410));
 sg13g2_antennanp ANTENNA_2676 (.A(net607));
 sg13g2_antennanp ANTENNA_2677 (.A(net607));
 sg13g2_antennanp ANTENNA_2678 (.A(net607));
 sg13g2_antennanp ANTENNA_2679 (.A(net607));
 sg13g2_antennanp ANTENNA_2680 (.A(net607));
 sg13g2_antennanp ANTENNA_2681 (.A(net607));
 sg13g2_antennanp ANTENNA_2682 (.A(net607));
 sg13g2_antennanp ANTENNA_2683 (.A(net607));
 sg13g2_antennanp ANTENNA_2684 (.A(net639));
 sg13g2_antennanp ANTENNA_2685 (.A(net639));
 sg13g2_antennanp ANTENNA_2686 (.A(net639));
 sg13g2_antennanp ANTENNA_2687 (.A(net639));
 sg13g2_antennanp ANTENNA_2688 (.A(net639));
 sg13g2_antennanp ANTENNA_2689 (.A(net639));
 sg13g2_antennanp ANTENNA_2690 (.A(net639));
 sg13g2_antennanp ANTENNA_2691 (.A(net639));
 sg13g2_antennanp ANTENNA_2692 (.A(net639));
 sg13g2_antennanp ANTENNA_2693 (.A(net639));
 sg13g2_antennanp ANTENNA_2694 (.A(net639));
 sg13g2_antennanp ANTENNA_2695 (.A(net639));
 sg13g2_antennanp ANTENNA_2696 (.A(net639));
 sg13g2_antennanp ANTENNA_2697 (.A(net673));
 sg13g2_antennanp ANTENNA_2698 (.A(net673));
 sg13g2_antennanp ANTENNA_2699 (.A(net673));
 sg13g2_antennanp ANTENNA_2700 (.A(net673));
 sg13g2_antennanp ANTENNA_2701 (.A(net673));
 sg13g2_antennanp ANTENNA_2702 (.A(net673));
 sg13g2_antennanp ANTENNA_2703 (.A(net673));
 sg13g2_antennanp ANTENNA_2704 (.A(net673));
 sg13g2_antennanp ANTENNA_2705 (.A(net673));
 sg13g2_antennanp ANTENNA_2706 (.A(net673));
 sg13g2_antennanp ANTENNA_2707 (.A(net673));
 sg13g2_antennanp ANTENNA_2708 (.A(net673));
 sg13g2_antennanp ANTENNA_2709 (.A(net673));
 sg13g2_antennanp ANTENNA_2710 (.A(net673));
 sg13g2_antennanp ANTENNA_2711 (.A(net673));
 sg13g2_antennanp ANTENNA_2712 (.A(net679));
 sg13g2_antennanp ANTENNA_2713 (.A(net679));
 sg13g2_antennanp ANTENNA_2714 (.A(net679));
 sg13g2_antennanp ANTENNA_2715 (.A(net679));
 sg13g2_antennanp ANTENNA_2716 (.A(net679));
 sg13g2_antennanp ANTENNA_2717 (.A(net679));
 sg13g2_antennanp ANTENNA_2718 (.A(net679));
 sg13g2_antennanp ANTENNA_2719 (.A(net679));
 sg13g2_antennanp ANTENNA_2720 (.A(net679));
 sg13g2_antennanp ANTENNA_2721 (.A(net684));
 sg13g2_antennanp ANTENNA_2722 (.A(net684));
 sg13g2_antennanp ANTENNA_2723 (.A(net684));
 sg13g2_antennanp ANTENNA_2724 (.A(net684));
 sg13g2_antennanp ANTENNA_2725 (.A(net684));
 sg13g2_antennanp ANTENNA_2726 (.A(net684));
 sg13g2_antennanp ANTENNA_2727 (.A(net684));
 sg13g2_antennanp ANTENNA_2728 (.A(net684));
 sg13g2_antennanp ANTENNA_2729 (.A(net684));
 sg13g2_antennanp ANTENNA_2730 (.A(net789));
 sg13g2_antennanp ANTENNA_2731 (.A(net789));
 sg13g2_antennanp ANTENNA_2732 (.A(net789));
 sg13g2_antennanp ANTENNA_2733 (.A(net789));
 sg13g2_antennanp ANTENNA_2734 (.A(net789));
 sg13g2_antennanp ANTENNA_2735 (.A(net789));
 sg13g2_antennanp ANTENNA_2736 (.A(net789));
 sg13g2_antennanp ANTENNA_2737 (.A(net789));
 sg13g2_antennanp ANTENNA_2738 (.A(net789));
 sg13g2_antennanp ANTENNA_2739 (.A(net845));
 sg13g2_antennanp ANTENNA_2740 (.A(net845));
 sg13g2_antennanp ANTENNA_2741 (.A(net845));
 sg13g2_antennanp ANTENNA_2742 (.A(net845));
 sg13g2_antennanp ANTENNA_2743 (.A(net845));
 sg13g2_antennanp ANTENNA_2744 (.A(net845));
 sg13g2_antennanp ANTENNA_2745 (.A(net845));
 sg13g2_antennanp ANTENNA_2746 (.A(net845));
 sg13g2_antennanp ANTENNA_2747 (.A(net961));
 sg13g2_antennanp ANTENNA_2748 (.A(net961));
 sg13g2_antennanp ANTENNA_2749 (.A(net961));
 sg13g2_antennanp ANTENNA_2750 (.A(net961));
 sg13g2_antennanp ANTENNA_2751 (.A(net961));
 sg13g2_antennanp ANTENNA_2752 (.A(net961));
 sg13g2_antennanp ANTENNA_2753 (.A(net961));
 sg13g2_antennanp ANTENNA_2754 (.A(net961));
 sg13g2_antennanp ANTENNA_2755 (.A(net966));
 sg13g2_antennanp ANTENNA_2756 (.A(net966));
 sg13g2_antennanp ANTENNA_2757 (.A(net966));
 sg13g2_antennanp ANTENNA_2758 (.A(net966));
 sg13g2_antennanp ANTENNA_2759 (.A(net966));
 sg13g2_antennanp ANTENNA_2760 (.A(net966));
 sg13g2_antennanp ANTENNA_2761 (.A(net966));
 sg13g2_antennanp ANTENNA_2762 (.A(net966));
 sg13g2_antennanp ANTENNA_2763 (.A(net1037));
 sg13g2_antennanp ANTENNA_2764 (.A(net1037));
 sg13g2_antennanp ANTENNA_2765 (.A(net1037));
 sg13g2_antennanp ANTENNA_2766 (.A(net1037));
 sg13g2_antennanp ANTENNA_2767 (.A(net1037));
 sg13g2_antennanp ANTENNA_2768 (.A(net1037));
 sg13g2_antennanp ANTENNA_2769 (.A(net1037));
 sg13g2_antennanp ANTENNA_2770 (.A(net1037));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_fill_2 FILLER_0_77 ();
 sg13g2_fill_1 FILLER_0_79 ();
 sg13g2_decap_8 FILLER_0_106 ();
 sg13g2_decap_8 FILLER_0_113 ();
 sg13g2_decap_8 FILLER_0_120 ();
 sg13g2_decap_8 FILLER_0_127 ();
 sg13g2_decap_8 FILLER_0_134 ();
 sg13g2_decap_8 FILLER_0_141 ();
 sg13g2_decap_4 FILLER_0_148 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_200 ();
 sg13g2_decap_4 FILLER_0_207 ();
 sg13g2_decap_8 FILLER_0_215 ();
 sg13g2_fill_2 FILLER_0_222 ();
 sg13g2_fill_2 FILLER_0_234 ();
 sg13g2_fill_1 FILLER_0_236 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_fill_1 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_286 ();
 sg13g2_decap_4 FILLER_0_293 ();
 sg13g2_fill_1 FILLER_0_297 ();
 sg13g2_decap_8 FILLER_0_324 ();
 sg13g2_decap_8 FILLER_0_331 ();
 sg13g2_decap_8 FILLER_0_338 ();
 sg13g2_decap_8 FILLER_0_345 ();
 sg13g2_decap_8 FILLER_0_352 ();
 sg13g2_decap_8 FILLER_0_359 ();
 sg13g2_decap_8 FILLER_0_366 ();
 sg13g2_decap_4 FILLER_0_373 ();
 sg13g2_fill_1 FILLER_0_377 ();
 sg13g2_decap_8 FILLER_0_404 ();
 sg13g2_decap_8 FILLER_0_411 ();
 sg13g2_decap_8 FILLER_0_418 ();
 sg13g2_decap_8 FILLER_0_425 ();
 sg13g2_decap_8 FILLER_0_432 ();
 sg13g2_decap_8 FILLER_0_439 ();
 sg13g2_decap_8 FILLER_0_446 ();
 sg13g2_decap_8 FILLER_0_479 ();
 sg13g2_decap_8 FILLER_0_486 ();
 sg13g2_decap_4 FILLER_0_493 ();
 sg13g2_fill_1 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_528 ();
 sg13g2_decap_8 FILLER_0_535 ();
 sg13g2_fill_2 FILLER_0_542 ();
 sg13g2_fill_1 FILLER_0_544 ();
 sg13g2_decap_8 FILLER_0_575 ();
 sg13g2_decap_4 FILLER_0_582 ();
 sg13g2_decap_4 FILLER_0_590 ();
 sg13g2_fill_1 FILLER_0_594 ();
 sg13g2_decap_8 FILLER_0_600 ();
 sg13g2_fill_2 FILLER_0_607 ();
 sg13g2_decap_8 FILLER_0_622 ();
 sg13g2_decap_8 FILLER_0_629 ();
 sg13g2_decap_8 FILLER_0_636 ();
 sg13g2_decap_8 FILLER_0_643 ();
 sg13g2_decap_8 FILLER_0_650 ();
 sg13g2_decap_8 FILLER_0_657 ();
 sg13g2_decap_4 FILLER_0_664 ();
 sg13g2_decap_8 FILLER_0_698 ();
 sg13g2_decap_8 FILLER_0_705 ();
 sg13g2_decap_8 FILLER_0_712 ();
 sg13g2_decap_8 FILLER_0_719 ();
 sg13g2_fill_2 FILLER_0_743 ();
 sg13g2_fill_1 FILLER_0_745 ();
 sg13g2_decap_8 FILLER_0_766 ();
 sg13g2_decap_4 FILLER_0_773 ();
 sg13g2_fill_1 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_788 ();
 sg13g2_fill_2 FILLER_0_795 ();
 sg13g2_decap_8 FILLER_0_823 ();
 sg13g2_decap_4 FILLER_0_830 ();
 sg13g2_decap_8 FILLER_0_842 ();
 sg13g2_decap_8 FILLER_0_849 ();
 sg13g2_decap_8 FILLER_0_856 ();
 sg13g2_fill_2 FILLER_0_863 ();
 sg13g2_decap_8 FILLER_0_875 ();
 sg13g2_fill_2 FILLER_0_882 ();
 sg13g2_fill_1 FILLER_0_884 ();
 sg13g2_decap_8 FILLER_0_919 ();
 sg13g2_decap_8 FILLER_0_926 ();
 sg13g2_fill_2 FILLER_0_933 ();
 sg13g2_fill_2 FILLER_0_945 ();
 sg13g2_decap_8 FILLER_0_983 ();
 sg13g2_decap_8 FILLER_0_990 ();
 sg13g2_fill_2 FILLER_0_997 ();
 sg13g2_decap_8 FILLER_0_1019 ();
 sg13g2_decap_8 FILLER_0_1026 ();
 sg13g2_decap_8 FILLER_0_1033 ();
 sg13g2_fill_2 FILLER_0_1040 ();
 sg13g2_fill_1 FILLER_0_1042 ();
 sg13g2_decap_8 FILLER_0_1069 ();
 sg13g2_fill_2 FILLER_0_1076 ();
 sg13g2_decap_4 FILLER_0_1104 ();
 sg13g2_decap_8 FILLER_0_1112 ();
 sg13g2_decap_4 FILLER_0_1119 ();
 sg13g2_fill_2 FILLER_0_1150 ();
 sg13g2_fill_2 FILLER_0_1178 ();
 sg13g2_decap_8 FILLER_0_1184 ();
 sg13g2_decap_8 FILLER_0_1191 ();
 sg13g2_fill_2 FILLER_0_1198 ();
 sg13g2_decap_8 FILLER_0_1226 ();
 sg13g2_decap_8 FILLER_0_1233 ();
 sg13g2_decap_8 FILLER_0_1240 ();
 sg13g2_fill_2 FILLER_0_1247 ();
 sg13g2_decap_8 FILLER_0_1253 ();
 sg13g2_decap_8 FILLER_0_1260 ();
 sg13g2_decap_8 FILLER_0_1267 ();
 sg13g2_decap_8 FILLER_0_1274 ();
 sg13g2_decap_4 FILLER_0_1281 ();
 sg13g2_fill_2 FILLER_0_1289 ();
 sg13g2_decap_8 FILLER_0_1314 ();
 sg13g2_fill_2 FILLER_0_1321 ();
 sg13g2_decap_4 FILLER_0_1331 ();
 sg13g2_fill_2 FILLER_0_1335 ();
 sg13g2_fill_2 FILLER_0_1347 ();
 sg13g2_fill_1 FILLER_0_1349 ();
 sg13g2_decap_8 FILLER_0_1358 ();
 sg13g2_decap_8 FILLER_0_1365 ();
 sg13g2_decap_8 FILLER_0_1372 ();
 sg13g2_decap_8 FILLER_0_1379 ();
 sg13g2_decap_8 FILLER_0_1386 ();
 sg13g2_decap_8 FILLER_0_1393 ();
 sg13g2_decap_8 FILLER_0_1426 ();
 sg13g2_fill_2 FILLER_0_1433 ();
 sg13g2_decap_8 FILLER_0_1461 ();
 sg13g2_decap_8 FILLER_0_1468 ();
 sg13g2_decap_8 FILLER_0_1475 ();
 sg13g2_decap_8 FILLER_0_1508 ();
 sg13g2_decap_8 FILLER_0_1515 ();
 sg13g2_decap_8 FILLER_0_1522 ();
 sg13g2_decap_4 FILLER_0_1529 ();
 sg13g2_decap_8 FILLER_0_1537 ();
 sg13g2_decap_8 FILLER_0_1544 ();
 sg13g2_decap_4 FILLER_0_1551 ();
 sg13g2_fill_1 FILLER_0_1555 ();
 sg13g2_decap_8 FILLER_0_1582 ();
 sg13g2_fill_2 FILLER_0_1589 ();
 sg13g2_fill_1 FILLER_0_1591 ();
 sg13g2_fill_1 FILLER_0_1612 ();
 sg13g2_decap_8 FILLER_0_1652 ();
 sg13g2_decap_8 FILLER_0_1659 ();
 sg13g2_decap_4 FILLER_0_1666 ();
 sg13g2_fill_1 FILLER_0_1700 ();
 sg13g2_fill_2 FILLER_0_1711 ();
 sg13g2_fill_2 FILLER_0_1738 ();
 sg13g2_fill_1 FILLER_0_1740 ();
 sg13g2_decap_8 FILLER_0_1771 ();
 sg13g2_decap_8 FILLER_0_1778 ();
 sg13g2_decap_8 FILLER_0_1785 ();
 sg13g2_decap_8 FILLER_0_1792 ();
 sg13g2_decap_8 FILLER_0_1803 ();
 sg13g2_fill_2 FILLER_0_1810 ();
 sg13g2_fill_1 FILLER_0_1812 ();
 sg13g2_decap_8 FILLER_0_1839 ();
 sg13g2_decap_8 FILLER_0_1846 ();
 sg13g2_decap_8 FILLER_0_1853 ();
 sg13g2_decap_8 FILLER_0_1860 ();
 sg13g2_decap_4 FILLER_0_1867 ();
 sg13g2_fill_2 FILLER_0_1875 ();
 sg13g2_fill_1 FILLER_0_1877 ();
 sg13g2_fill_1 FILLER_0_1882 ();
 sg13g2_decap_8 FILLER_0_1893 ();
 sg13g2_decap_8 FILLER_0_1900 ();
 sg13g2_decap_4 FILLER_0_1907 ();
 sg13g2_decap_8 FILLER_0_1924 ();
 sg13g2_decap_4 FILLER_0_1931 ();
 sg13g2_fill_2 FILLER_0_1935 ();
 sg13g2_decap_8 FILLER_0_1941 ();
 sg13g2_decap_8 FILLER_0_1948 ();
 sg13g2_decap_8 FILLER_0_1955 ();
 sg13g2_decap_4 FILLER_0_1962 ();
 sg13g2_fill_1 FILLER_0_1966 ();
 sg13g2_decap_8 FILLER_0_1997 ();
 sg13g2_decap_8 FILLER_0_2004 ();
 sg13g2_decap_8 FILLER_0_2011 ();
 sg13g2_decap_8 FILLER_0_2018 ();
 sg13g2_decap_8 FILLER_0_2025 ();
 sg13g2_fill_2 FILLER_0_2032 ();
 sg13g2_fill_1 FILLER_0_2038 ();
 sg13g2_decap_8 FILLER_0_2069 ();
 sg13g2_decap_8 FILLER_0_2076 ();
 sg13g2_fill_1 FILLER_0_2083 ();
 sg13g2_decap_4 FILLER_0_2110 ();
 sg13g2_fill_1 FILLER_0_2114 ();
 sg13g2_decap_8 FILLER_0_2119 ();
 sg13g2_decap_8 FILLER_0_2126 ();
 sg13g2_decap_8 FILLER_0_2133 ();
 sg13g2_decap_4 FILLER_0_2140 ();
 sg13g2_fill_2 FILLER_0_2144 ();
 sg13g2_decap_8 FILLER_0_2154 ();
 sg13g2_decap_8 FILLER_0_2165 ();
 sg13g2_decap_8 FILLER_0_2172 ();
 sg13g2_decap_8 FILLER_0_2179 ();
 sg13g2_fill_1 FILLER_0_2186 ();
 sg13g2_decap_8 FILLER_0_2191 ();
 sg13g2_fill_1 FILLER_0_2198 ();
 sg13g2_decap_8 FILLER_0_2207 ();
 sg13g2_decap_8 FILLER_0_2214 ();
 sg13g2_fill_2 FILLER_0_2221 ();
 sg13g2_fill_2 FILLER_0_2233 ();
 sg13g2_fill_1 FILLER_0_2235 ();
 sg13g2_decap_8 FILLER_0_2240 ();
 sg13g2_decap_8 FILLER_0_2247 ();
 sg13g2_decap_8 FILLER_0_2254 ();
 sg13g2_decap_8 FILLER_0_2261 ();
 sg13g2_decap_4 FILLER_0_2268 ();
 sg13g2_fill_1 FILLER_0_2272 ();
 sg13g2_decap_8 FILLER_0_2277 ();
 sg13g2_decap_8 FILLER_0_2284 ();
 sg13g2_decap_8 FILLER_0_2291 ();
 sg13g2_decap_8 FILLER_0_2298 ();
 sg13g2_fill_2 FILLER_0_2305 ();
 sg13g2_decap_8 FILLER_0_2337 ();
 sg13g2_decap_8 FILLER_0_2344 ();
 sg13g2_decap_8 FILLER_0_2351 ();
 sg13g2_decap_8 FILLER_0_2358 ();
 sg13g2_decap_8 FILLER_0_2365 ();
 sg13g2_decap_8 FILLER_0_2372 ();
 sg13g2_decap_4 FILLER_0_2379 ();
 sg13g2_decap_8 FILLER_0_2409 ();
 sg13g2_decap_8 FILLER_0_2416 ();
 sg13g2_decap_8 FILLER_0_2423 ();
 sg13g2_decap_4 FILLER_0_2430 ();
 sg13g2_fill_2 FILLER_0_2434 ();
 sg13g2_decap_8 FILLER_0_2462 ();
 sg13g2_decap_8 FILLER_0_2469 ();
 sg13g2_decap_8 FILLER_0_2476 ();
 sg13g2_decap_4 FILLER_0_2483 ();
 sg13g2_fill_1 FILLER_0_2487 ();
 sg13g2_decap_8 FILLER_0_2501 ();
 sg13g2_fill_1 FILLER_0_2508 ();
 sg13g2_decap_8 FILLER_0_2519 ();
 sg13g2_decap_8 FILLER_0_2526 ();
 sg13g2_decap_8 FILLER_0_2533 ();
 sg13g2_decap_4 FILLER_0_2540 ();
 sg13g2_fill_1 FILLER_0_2544 ();
 sg13g2_decap_8 FILLER_0_2549 ();
 sg13g2_decap_8 FILLER_0_2556 ();
 sg13g2_fill_2 FILLER_0_2563 ();
 sg13g2_decap_8 FILLER_0_2586 ();
 sg13g2_decap_8 FILLER_0_2593 ();
 sg13g2_decap_8 FILLER_0_2600 ();
 sg13g2_decap_8 FILLER_0_2607 ();
 sg13g2_decap_8 FILLER_0_2614 ();
 sg13g2_decap_8 FILLER_0_2621 ();
 sg13g2_decap_8 FILLER_0_2628 ();
 sg13g2_decap_8 FILLER_0_2635 ();
 sg13g2_decap_8 FILLER_0_2642 ();
 sg13g2_decap_8 FILLER_0_2649 ();
 sg13g2_decap_8 FILLER_0_2656 ();
 sg13g2_decap_8 FILLER_0_2663 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_fill_1 FILLER_1_42 ();
 sg13g2_fill_2 FILLER_1_73 ();
 sg13g2_fill_1 FILLER_1_75 ();
 sg13g2_fill_1 FILLER_1_88 ();
 sg13g2_decap_8 FILLER_1_93 ();
 sg13g2_decap_8 FILLER_1_100 ();
 sg13g2_fill_2 FILLER_1_107 ();
 sg13g2_fill_1 FILLER_1_109 ();
 sg13g2_decap_8 FILLER_1_114 ();
 sg13g2_decap_4 FILLER_1_121 ();
 sg13g2_fill_2 FILLER_1_211 ();
 sg13g2_decap_4 FILLER_1_217 ();
 sg13g2_fill_1 FILLER_1_221 ();
 sg13g2_fill_2 FILLER_1_260 ();
 sg13g2_decap_8 FILLER_1_278 ();
 sg13g2_decap_8 FILLER_1_285 ();
 sg13g2_decap_4 FILLER_1_292 ();
 sg13g2_fill_1 FILLER_1_296 ();
 sg13g2_decap_8 FILLER_1_411 ();
 sg13g2_decap_4 FILLER_1_418 ();
 sg13g2_fill_2 FILLER_1_426 ();
 sg13g2_fill_1 FILLER_1_428 ();
 sg13g2_decap_4 FILLER_1_455 ();
 sg13g2_fill_2 FILLER_1_459 ();
 sg13g2_fill_2 FILLER_1_465 ();
 sg13g2_fill_2 FILLER_1_497 ();
 sg13g2_fill_2 FILLER_1_504 ();
 sg13g2_fill_1 FILLER_1_506 ();
 sg13g2_fill_2 FILLER_1_510 ();
 sg13g2_fill_1 FILLER_1_512 ();
 sg13g2_fill_2 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_578 ();
 sg13g2_fill_2 FILLER_1_585 ();
 sg13g2_decap_4 FILLER_1_633 ();
 sg13g2_fill_1 FILLER_1_637 ();
 sg13g2_fill_2 FILLER_1_668 ();
 sg13g2_decap_4 FILLER_1_675 ();
 sg13g2_decap_8 FILLER_1_705 ();
 sg13g2_decap_8 FILLER_1_712 ();
 sg13g2_decap_4 FILLER_1_719 ();
 sg13g2_fill_1 FILLER_1_723 ();
 sg13g2_fill_2 FILLER_1_760 ();
 sg13g2_decap_4 FILLER_1_788 ();
 sg13g2_fill_2 FILLER_1_802 ();
 sg13g2_fill_2 FILLER_1_830 ();
 sg13g2_fill_1 FILLER_1_832 ();
 sg13g2_fill_2 FILLER_1_846 ();
 sg13g2_decap_8 FILLER_1_914 ();
 sg13g2_decap_8 FILLER_1_921 ();
 sg13g2_decap_4 FILLER_1_928 ();
 sg13g2_fill_2 FILLER_1_932 ();
 sg13g2_decap_8 FILLER_1_947 ();
 sg13g2_decap_8 FILLER_1_964 ();
 sg13g2_decap_8 FILLER_1_971 ();
 sg13g2_decap_8 FILLER_1_978 ();
 sg13g2_fill_1 FILLER_1_985 ();
 sg13g2_fill_2 FILLER_1_1026 ();
 sg13g2_fill_2 FILLER_1_1038 ();
 sg13g2_fill_1 FILLER_1_1040 ();
 sg13g2_decap_4 FILLER_1_1051 ();
 sg13g2_fill_2 FILLER_1_1081 ();
 sg13g2_fill_1 FILLER_1_1083 ();
 sg13g2_fill_2 FILLER_1_1094 ();
 sg13g2_decap_4 FILLER_1_1126 ();
 sg13g2_fill_2 FILLER_1_1130 ();
 sg13g2_decap_8 FILLER_1_1162 ();
 sg13g2_decap_8 FILLER_1_1195 ();
 sg13g2_fill_1 FILLER_1_1202 ();
 sg13g2_fill_2 FILLER_1_1241 ();
 sg13g2_fill_2 FILLER_1_1269 ();
 sg13g2_fill_1 FILLER_1_1276 ();
 sg13g2_fill_1 FILLER_1_1303 ();
 sg13g2_fill_2 FILLER_1_1376 ();
 sg13g2_fill_1 FILLER_1_1378 ();
 sg13g2_fill_1 FILLER_1_1412 ();
 sg13g2_decap_8 FILLER_1_1421 ();
 sg13g2_fill_1 FILLER_1_1428 ();
 sg13g2_decap_8 FILLER_1_1459 ();
 sg13g2_decap_8 FILLER_1_1466 ();
 sg13g2_decap_4 FILLER_1_1473 ();
 sg13g2_fill_2 FILLER_1_1477 ();
 sg13g2_fill_1 FILLER_1_1552 ();
 sg13g2_fill_1 FILLER_1_1587 ();
 sg13g2_decap_8 FILLER_1_1598 ();
 sg13g2_decap_4 FILLER_1_1657 ();
 sg13g2_fill_1 FILLER_1_1661 ();
 sg13g2_decap_8 FILLER_1_1670 ();
 sg13g2_decap_4 FILLER_1_1677 ();
 sg13g2_fill_1 FILLER_1_1681 ();
 sg13g2_fill_1 FILLER_1_1711 ();
 sg13g2_fill_1 FILLER_1_1716 ();
 sg13g2_fill_1 FILLER_1_1743 ();
 sg13g2_fill_1 FILLER_1_1748 ();
 sg13g2_fill_1 FILLER_1_1759 ();
 sg13g2_decap_8 FILLER_1_1770 ();
 sg13g2_decap_8 FILLER_1_1777 ();
 sg13g2_decap_8 FILLER_1_1784 ();
 sg13g2_fill_1 FILLER_1_1791 ();
 sg13g2_fill_2 FILLER_1_1818 ();
 sg13g2_fill_2 FILLER_1_1869 ();
 sg13g2_fill_2 FILLER_1_1927 ();
 sg13g2_fill_1 FILLER_1_1929 ();
 sg13g2_fill_1 FILLER_1_1956 ();
 sg13g2_decap_8 FILLER_1_1993 ();
 sg13g2_fill_1 FILLER_1_2000 ();
 sg13g2_decap_4 FILLER_1_2073 ();
 sg13g2_fill_2 FILLER_1_2107 ();
 sg13g2_decap_4 FILLER_1_2135 ();
 sg13g2_fill_2 FILLER_1_2139 ();
 sg13g2_fill_2 FILLER_1_2206 ();
 sg13g2_decap_4 FILLER_1_2248 ();
 sg13g2_fill_2 FILLER_1_2252 ();
 sg13g2_decap_8 FILLER_1_2290 ();
 sg13g2_fill_1 FILLER_1_2297 ();
 sg13g2_decap_4 FILLER_1_2324 ();
 sg13g2_fill_1 FILLER_1_2328 ();
 sg13g2_decap_4 FILLER_1_2355 ();
 sg13g2_decap_4 FILLER_1_2369 ();
 sg13g2_fill_2 FILLER_1_2373 ();
 sg13g2_decap_4 FILLER_1_2411 ();
 sg13g2_decap_8 FILLER_1_2419 ();
 sg13g2_decap_4 FILLER_1_2426 ();
 sg13g2_fill_1 FILLER_1_2430 ();
 sg13g2_decap_8 FILLER_1_2441 ();
 sg13g2_fill_2 FILLER_1_2448 ();
 sg13g2_fill_1 FILLER_1_2450 ();
 sg13g2_fill_1 FILLER_1_2495 ();
 sg13g2_decap_4 FILLER_1_2522 ();
 sg13g2_decap_8 FILLER_1_2530 ();
 sg13g2_fill_1 FILLER_1_2537 ();
 sg13g2_fill_1 FILLER_1_2564 ();
 sg13g2_decap_8 FILLER_1_2601 ();
 sg13g2_decap_8 FILLER_1_2608 ();
 sg13g2_decap_8 FILLER_1_2615 ();
 sg13g2_decap_8 FILLER_1_2622 ();
 sg13g2_decap_8 FILLER_1_2629 ();
 sg13g2_decap_8 FILLER_1_2636 ();
 sg13g2_decap_8 FILLER_1_2643 ();
 sg13g2_decap_8 FILLER_1_2650 ();
 sg13g2_decap_8 FILLER_1_2657 ();
 sg13g2_decap_4 FILLER_1_2664 ();
 sg13g2_fill_2 FILLER_1_2668 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_fill_2 FILLER_2_21 ();
 sg13g2_fill_1 FILLER_2_23 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_fill_2 FILLER_2_47 ();
 sg13g2_fill_1 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_92 ();
 sg13g2_decap_4 FILLER_2_99 ();
 sg13g2_fill_1 FILLER_2_103 ();
 sg13g2_decap_4 FILLER_2_130 ();
 sg13g2_fill_2 FILLER_2_134 ();
 sg13g2_fill_1 FILLER_2_166 ();
 sg13g2_fill_1 FILLER_2_171 ();
 sg13g2_fill_2 FILLER_2_219 ();
 sg13g2_fill_1 FILLER_2_221 ();
 sg13g2_fill_2 FILLER_2_278 ();
 sg13g2_fill_2 FILLER_2_326 ();
 sg13g2_fill_2 FILLER_2_370 ();
 sg13g2_fill_2 FILLER_2_385 ();
 sg13g2_fill_1 FILLER_2_395 ();
 sg13g2_fill_1 FILLER_2_422 ();
 sg13g2_fill_1 FILLER_2_449 ();
 sg13g2_decap_4 FILLER_2_455 ();
 sg13g2_fill_1 FILLER_2_473 ();
 sg13g2_fill_2 FILLER_2_500 ();
 sg13g2_fill_1 FILLER_2_511 ();
 sg13g2_fill_1 FILLER_2_521 ();
 sg13g2_fill_2 FILLER_2_526 ();
 sg13g2_fill_2 FILLER_2_552 ();
 sg13g2_fill_2 FILLER_2_573 ();
 sg13g2_fill_1 FILLER_2_665 ();
 sg13g2_fill_1 FILLER_2_671 ();
 sg13g2_fill_1 FILLER_2_677 ();
 sg13g2_fill_1 FILLER_2_683 ();
 sg13g2_decap_4 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_701 ();
 sg13g2_fill_1 FILLER_2_760 ();
 sg13g2_fill_1 FILLER_2_805 ();
 sg13g2_fill_1 FILLER_2_810 ();
 sg13g2_fill_1 FILLER_2_815 ();
 sg13g2_fill_1 FILLER_2_826 ();
 sg13g2_fill_2 FILLER_2_951 ();
 sg13g2_fill_1 FILLER_2_1013 ();
 sg13g2_fill_1 FILLER_2_1061 ();
 sg13g2_decap_8 FILLER_2_1066 ();
 sg13g2_decap_4 FILLER_2_1073 ();
 sg13g2_fill_1 FILLER_2_1077 ();
 sg13g2_fill_1 FILLER_2_1149 ();
 sg13g2_fill_1 FILLER_2_1160 ();
 sg13g2_fill_1 FILLER_2_1179 ();
 sg13g2_fill_2 FILLER_2_1224 ();
 sg13g2_fill_1 FILLER_2_1226 ();
 sg13g2_fill_1 FILLER_2_1253 ();
 sg13g2_fill_1 FILLER_2_1374 ();
 sg13g2_fill_1 FILLER_2_1391 ();
 sg13g2_fill_2 FILLER_2_1400 ();
 sg13g2_decap_4 FILLER_2_1423 ();
 sg13g2_fill_2 FILLER_2_1427 ();
 sg13g2_fill_1 FILLER_2_1433 ();
 sg13g2_decap_8 FILLER_2_1451 ();
 sg13g2_decap_4 FILLER_2_1458 ();
 sg13g2_fill_1 FILLER_2_1462 ();
 sg13g2_fill_1 FILLER_2_1563 ();
 sg13g2_fill_1 FILLER_2_1568 ();
 sg13g2_fill_1 FILLER_2_1595 ();
 sg13g2_fill_1 FILLER_2_1622 ();
 sg13g2_decap_8 FILLER_2_1627 ();
 sg13g2_fill_1 FILLER_2_1634 ();
 sg13g2_decap_4 FILLER_2_1639 ();
 sg13g2_fill_1 FILLER_2_1655 ();
 sg13g2_decap_8 FILLER_2_1692 ();
 sg13g2_fill_1 FILLER_2_1699 ();
 sg13g2_fill_2 FILLER_2_1835 ();
 sg13g2_fill_1 FILLER_2_1837 ();
 sg13g2_decap_4 FILLER_2_1890 ();
 sg13g2_fill_1 FILLER_2_1894 ();
 sg13g2_fill_2 FILLER_2_1899 ();
 sg13g2_fill_1 FILLER_2_1927 ();
 sg13g2_fill_1 FILLER_2_1964 ();
 sg13g2_decap_8 FILLER_2_1985 ();
 sg13g2_decap_8 FILLER_2_1992 ();
 sg13g2_decap_4 FILLER_2_1999 ();
 sg13g2_fill_2 FILLER_2_2003 ();
 sg13g2_fill_1 FILLER_2_2019 ();
 sg13g2_fill_1 FILLER_2_2030 ();
 sg13g2_decap_4 FILLER_2_2082 ();
 sg13g2_fill_1 FILLER_2_2086 ();
 sg13g2_fill_2 FILLER_2_2091 ();
 sg13g2_decap_4 FILLER_2_2103 ();
 sg13g2_fill_1 FILLER_2_2117 ();
 sg13g2_fill_2 FILLER_2_2122 ();
 sg13g2_fill_2 FILLER_2_2145 ();
 sg13g2_decap_4 FILLER_2_2253 ();
 sg13g2_fill_2 FILLER_2_2261 ();
 sg13g2_fill_1 FILLER_2_2351 ();
 sg13g2_fill_2 FILLER_2_2401 ();
 sg13g2_fill_1 FILLER_2_2403 ();
 sg13g2_decap_4 FILLER_2_2440 ();
 sg13g2_fill_2 FILLER_2_2448 ();
 sg13g2_fill_1 FILLER_2_2450 ();
 sg13g2_fill_1 FILLER_2_2481 ();
 sg13g2_fill_1 FILLER_2_2518 ();
 sg13g2_decap_8 FILLER_2_2605 ();
 sg13g2_decap_8 FILLER_2_2612 ();
 sg13g2_decap_8 FILLER_2_2619 ();
 sg13g2_decap_8 FILLER_2_2626 ();
 sg13g2_decap_8 FILLER_2_2633 ();
 sg13g2_decap_8 FILLER_2_2640 ();
 sg13g2_decap_8 FILLER_2_2647 ();
 sg13g2_decap_8 FILLER_2_2654 ();
 sg13g2_decap_8 FILLER_2_2661 ();
 sg13g2_fill_2 FILLER_2_2668 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_fill_2 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_93 ();
 sg13g2_fill_1 FILLER_3_100 ();
 sg13g2_decap_8 FILLER_3_127 ();
 sg13g2_decap_8 FILLER_3_134 ();
 sg13g2_fill_2 FILLER_3_141 ();
 sg13g2_fill_1 FILLER_3_143 ();
 sg13g2_fill_2 FILLER_3_160 ();
 sg13g2_fill_2 FILLER_3_185 ();
 sg13g2_decap_8 FILLER_3_200 ();
 sg13g2_fill_1 FILLER_3_207 ();
 sg13g2_fill_2 FILLER_3_251 ();
 sg13g2_fill_1 FILLER_3_253 ();
 sg13g2_fill_1 FILLER_3_258 ();
 sg13g2_fill_1 FILLER_3_297 ();
 sg13g2_fill_1 FILLER_3_311 ();
 sg13g2_decap_4 FILLER_3_326 ();
 sg13g2_fill_2 FILLER_3_359 ();
 sg13g2_fill_1 FILLER_3_361 ();
 sg13g2_fill_2 FILLER_3_378 ();
 sg13g2_fill_2 FILLER_3_388 ();
 sg13g2_fill_2 FILLER_3_395 ();
 sg13g2_fill_2 FILLER_3_410 ();
 sg13g2_fill_1 FILLER_3_412 ();
 sg13g2_decap_4 FILLER_3_422 ();
 sg13g2_fill_1 FILLER_3_426 ();
 sg13g2_fill_2 FILLER_3_431 ();
 sg13g2_fill_1 FILLER_3_433 ();
 sg13g2_fill_1 FILLER_3_449 ();
 sg13g2_decap_4 FILLER_3_486 ();
 sg13g2_fill_1 FILLER_3_503 ();
 sg13g2_fill_1 FILLER_3_514 ();
 sg13g2_fill_1 FILLER_3_530 ();
 sg13g2_fill_1 FILLER_3_557 ();
 sg13g2_fill_1 FILLER_3_568 ();
 sg13g2_fill_1 FILLER_3_592 ();
 sg13g2_fill_1 FILLER_3_619 ();
 sg13g2_decap_4 FILLER_3_624 ();
 sg13g2_decap_4 FILLER_3_654 ();
 sg13g2_fill_2 FILLER_3_668 ();
 sg13g2_fill_1 FILLER_3_670 ();
 sg13g2_fill_1 FILLER_3_675 ();
 sg13g2_fill_2 FILLER_3_721 ();
 sg13g2_fill_1 FILLER_3_723 ();
 sg13g2_fill_2 FILLER_3_771 ();
 sg13g2_fill_1 FILLER_3_773 ();
 sg13g2_fill_2 FILLER_3_821 ();
 sg13g2_decap_8 FILLER_3_884 ();
 sg13g2_decap_4 FILLER_3_926 ();
 sg13g2_fill_2 FILLER_3_930 ();
 sg13g2_fill_2 FILLER_3_966 ();
 sg13g2_decap_8 FILLER_3_972 ();
 sg13g2_decap_8 FILLER_3_979 ();
 sg13g2_fill_2 FILLER_3_1027 ();
 sg13g2_fill_2 FILLER_3_1039 ();
 sg13g2_fill_1 FILLER_3_1041 ();
 sg13g2_decap_8 FILLER_3_1085 ();
 sg13g2_decap_4 FILLER_3_1092 ();
 sg13g2_fill_1 FILLER_3_1096 ();
 sg13g2_decap_8 FILLER_3_1154 ();
 sg13g2_fill_2 FILLER_3_1161 ();
 sg13g2_fill_1 FILLER_3_1229 ();
 sg13g2_fill_1 FILLER_3_1234 ();
 sg13g2_fill_2 FILLER_3_1256 ();
 sg13g2_fill_2 FILLER_3_1330 ();
 sg13g2_fill_1 FILLER_3_1418 ();
 sg13g2_fill_2 FILLER_3_1424 ();
 sg13g2_decap_4 FILLER_3_1439 ();
 sg13g2_fill_2 FILLER_3_1443 ();
 sg13g2_decap_8 FILLER_3_1449 ();
 sg13g2_decap_4 FILLER_3_1456 ();
 sg13g2_fill_1 FILLER_3_1460 ();
 sg13g2_decap_8 FILLER_3_1509 ();
 sg13g2_fill_1 FILLER_3_1516 ();
 sg13g2_fill_1 FILLER_3_1527 ();
 sg13g2_decap_4 FILLER_3_1582 ();
 sg13g2_fill_1 FILLER_3_1586 ();
 sg13g2_fill_1 FILLER_3_1602 ();
 sg13g2_fill_1 FILLER_3_1613 ();
 sg13g2_fill_1 FILLER_3_1640 ();
 sg13g2_fill_1 FILLER_3_1645 ();
 sg13g2_fill_2 FILLER_3_1722 ();
 sg13g2_fill_2 FILLER_3_1745 ();
 sg13g2_fill_2 FILLER_3_1783 ();
 sg13g2_fill_2 FILLER_3_1829 ();
 sg13g2_decap_8 FILLER_3_1857 ();
 sg13g2_fill_1 FILLER_3_1864 ();
 sg13g2_fill_1 FILLER_3_1896 ();
 sg13g2_fill_1 FILLER_3_1923 ();
 sg13g2_fill_1 FILLER_3_1964 ();
 sg13g2_fill_2 FILLER_3_1969 ();
 sg13g2_fill_1 FILLER_3_2007 ();
 sg13g2_decap_8 FILLER_3_2072 ();
 sg13g2_decap_8 FILLER_3_2079 ();
 sg13g2_fill_2 FILLER_3_2086 ();
 sg13g2_fill_1 FILLER_3_2088 ();
 sg13g2_fill_2 FILLER_3_2161 ();
 sg13g2_fill_1 FILLER_3_2163 ();
 sg13g2_fill_1 FILLER_3_2168 ();
 sg13g2_decap_8 FILLER_3_2195 ();
 sg13g2_fill_2 FILLER_3_2202 ();
 sg13g2_fill_1 FILLER_3_2204 ();
 sg13g2_fill_2 FILLER_3_2215 ();
 sg13g2_fill_2 FILLER_3_2227 ();
 sg13g2_fill_1 FILLER_3_2233 ();
 sg13g2_fill_2 FILLER_3_2297 ();
 sg13g2_fill_2 FILLER_3_2307 ();
 sg13g2_fill_1 FILLER_3_2309 ();
 sg13g2_fill_1 FILLER_3_2314 ();
 sg13g2_fill_1 FILLER_3_2340 ();
 sg13g2_decap_8 FILLER_3_2345 ();
 sg13g2_fill_2 FILLER_3_2352 ();
 sg13g2_fill_1 FILLER_3_2354 ();
 sg13g2_fill_1 FILLER_3_2363 ();
 sg13g2_fill_2 FILLER_3_2394 ();
 sg13g2_decap_8 FILLER_3_2400 ();
 sg13g2_decap_4 FILLER_3_2407 ();
 sg13g2_decap_4 FILLER_3_2432 ();
 sg13g2_fill_2 FILLER_3_2436 ();
 sg13g2_fill_2 FILLER_3_2540 ();
 sg13g2_fill_1 FILLER_3_2552 ();
 sg13g2_fill_2 FILLER_3_2573 ();
 sg13g2_decap_8 FILLER_3_2601 ();
 sg13g2_decap_8 FILLER_3_2608 ();
 sg13g2_decap_8 FILLER_3_2615 ();
 sg13g2_decap_8 FILLER_3_2622 ();
 sg13g2_decap_8 FILLER_3_2629 ();
 sg13g2_decap_8 FILLER_3_2636 ();
 sg13g2_decap_8 FILLER_3_2643 ();
 sg13g2_decap_8 FILLER_3_2650 ();
 sg13g2_decap_8 FILLER_3_2657 ();
 sg13g2_decap_4 FILLER_3_2664 ();
 sg13g2_fill_2 FILLER_3_2668 ();
 sg13g2_decap_4 FILLER_4_0 ();
 sg13g2_fill_1 FILLER_4_4 ();
 sg13g2_fill_2 FILLER_4_36 ();
 sg13g2_fill_1 FILLER_4_44 ();
 sg13g2_fill_2 FILLER_4_50 ();
 sg13g2_fill_2 FILLER_4_67 ();
 sg13g2_fill_1 FILLER_4_69 ();
 sg13g2_fill_2 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_129 ();
 sg13g2_decap_8 FILLER_4_136 ();
 sg13g2_decap_8 FILLER_4_143 ();
 sg13g2_decap_4 FILLER_4_150 ();
 sg13g2_fill_1 FILLER_4_166 ();
 sg13g2_fill_2 FILLER_4_172 ();
 sg13g2_fill_1 FILLER_4_174 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_fill_1 FILLER_4_238 ();
 sg13g2_fill_2 FILLER_4_275 ();
 sg13g2_fill_1 FILLER_4_277 ();
 sg13g2_fill_2 FILLER_4_340 ();
 sg13g2_fill_1 FILLER_4_346 ();
 sg13g2_fill_2 FILLER_4_351 ();
 sg13g2_fill_2 FILLER_4_357 ();
 sg13g2_fill_2 FILLER_4_363 ();
 sg13g2_decap_8 FILLER_4_425 ();
 sg13g2_decap_8 FILLER_4_432 ();
 sg13g2_decap_8 FILLER_4_439 ();
 sg13g2_fill_1 FILLER_4_446 ();
 sg13g2_fill_2 FILLER_4_456 ();
 sg13g2_decap_4 FILLER_4_462 ();
 sg13g2_fill_2 FILLER_4_466 ();
 sg13g2_decap_4 FILLER_4_472 ();
 sg13g2_fill_2 FILLER_4_476 ();
 sg13g2_fill_1 FILLER_4_503 ();
 sg13g2_fill_1 FILLER_4_566 ();
 sg13g2_fill_2 FILLER_4_585 ();
 sg13g2_fill_2 FILLER_4_606 ();
 sg13g2_decap_8 FILLER_4_612 ();
 sg13g2_decap_8 FILLER_4_619 ();
 sg13g2_fill_2 FILLER_4_626 ();
 sg13g2_fill_2 FILLER_4_674 ();
 sg13g2_decap_4 FILLER_4_685 ();
 sg13g2_fill_1 FILLER_4_689 ();
 sg13g2_decap_8 FILLER_4_705 ();
 sg13g2_fill_2 FILLER_4_712 ();
 sg13g2_fill_1 FILLER_4_714 ();
 sg13g2_decap_4 FILLER_4_719 ();
 sg13g2_decap_4 FILLER_4_728 ();
 sg13g2_decap_4 FILLER_4_736 ();
 sg13g2_fill_1 FILLER_4_740 ();
 sg13g2_fill_2 FILLER_4_755 ();
 sg13g2_fill_1 FILLER_4_757 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_fill_2 FILLER_4_791 ();
 sg13g2_fill_1 FILLER_4_793 ();
 sg13g2_decap_4 FILLER_4_808 ();
 sg13g2_fill_1 FILLER_4_812 ();
 sg13g2_fill_2 FILLER_4_870 ();
 sg13g2_fill_1 FILLER_4_872 ();
 sg13g2_decap_8 FILLER_4_877 ();
 sg13g2_decap_8 FILLER_4_884 ();
 sg13g2_decap_8 FILLER_4_891 ();
 sg13g2_fill_2 FILLER_4_898 ();
 sg13g2_decap_8 FILLER_4_926 ();
 sg13g2_decap_8 FILLER_4_933 ();
 sg13g2_decap_4 FILLER_4_940 ();
 sg13g2_fill_2 FILLER_4_948 ();
 sg13g2_fill_1 FILLER_4_950 ();
 sg13g2_fill_2 FILLER_4_961 ();
 sg13g2_fill_1 FILLER_4_963 ();
 sg13g2_decap_8 FILLER_4_989 ();
 sg13g2_decap_4 FILLER_4_996 ();
 sg13g2_fill_2 FILLER_4_1055 ();
 sg13g2_decap_4 FILLER_4_1061 ();
 sg13g2_fill_2 FILLER_4_1065 ();
 sg13g2_decap_8 FILLER_4_1093 ();
 sg13g2_decap_8 FILLER_4_1100 ();
 sg13g2_decap_4 FILLER_4_1107 ();
 sg13g2_fill_2 FILLER_4_1111 ();
 sg13g2_decap_4 FILLER_4_1117 ();
 sg13g2_fill_1 FILLER_4_1141 ();
 sg13g2_fill_2 FILLER_4_1194 ();
 sg13g2_fill_1 FILLER_4_1196 ();
 sg13g2_fill_2 FILLER_4_1280 ();
 sg13g2_fill_1 FILLER_4_1302 ();
 sg13g2_fill_2 FILLER_4_1330 ();
 sg13g2_fill_2 FILLER_4_1342 ();
 sg13g2_fill_2 FILLER_4_1354 ();
 sg13g2_fill_1 FILLER_4_1356 ();
 sg13g2_decap_4 FILLER_4_1414 ();
 sg13g2_decap_4 FILLER_4_1448 ();
 sg13g2_fill_1 FILLER_4_1486 ();
 sg13g2_fill_2 FILLER_4_1501 ();
 sg13g2_decap_8 FILLER_4_1507 ();
 sg13g2_decap_4 FILLER_4_1514 ();
 sg13g2_fill_2 FILLER_4_1518 ();
 sg13g2_fill_2 FILLER_4_1582 ();
 sg13g2_decap_8 FILLER_4_1623 ();
 sg13g2_decap_4 FILLER_4_1630 ();
 sg13g2_decap_8 FILLER_4_1638 ();
 sg13g2_fill_1 FILLER_4_1645 ();
 sg13g2_fill_1 FILLER_4_1676 ();
 sg13g2_decap_8 FILLER_4_1698 ();
 sg13g2_decap_4 FILLER_4_1705 ();
 sg13g2_fill_1 FILLER_4_1749 ();
 sg13g2_fill_2 FILLER_4_1760 ();
 sg13g2_decap_8 FILLER_4_1787 ();
 sg13g2_fill_2 FILLER_4_1794 ();
 sg13g2_fill_1 FILLER_4_1796 ();
 sg13g2_fill_1 FILLER_4_1807 ();
 sg13g2_decap_4 FILLER_4_1843 ();
 sg13g2_fill_1 FILLER_4_1847 ();
 sg13g2_decap_8 FILLER_4_1869 ();
 sg13g2_decap_8 FILLER_4_1876 ();
 sg13g2_fill_2 FILLER_4_1883 ();
 sg13g2_fill_1 FILLER_4_1885 ();
 sg13g2_fill_1 FILLER_4_1906 ();
 sg13g2_decap_8 FILLER_4_1911 ();
 sg13g2_decap_8 FILLER_4_1918 ();
 sg13g2_decap_4 FILLER_4_1925 ();
 sg13g2_fill_1 FILLER_4_1929 ();
 sg13g2_fill_2 FILLER_4_1970 ();
 sg13g2_fill_1 FILLER_4_1976 ();
 sg13g2_fill_2 FILLER_4_1981 ();
 sg13g2_fill_2 FILLER_4_2009 ();
 sg13g2_fill_2 FILLER_4_2037 ();
 sg13g2_fill_1 FILLER_4_2039 ();
 sg13g2_decap_8 FILLER_4_2141 ();
 sg13g2_decap_8 FILLER_4_2148 ();
 sg13g2_decap_8 FILLER_4_2155 ();
 sg13g2_fill_1 FILLER_4_2162 ();
 sg13g2_fill_2 FILLER_4_2194 ();
 sg13g2_fill_1 FILLER_4_2196 ();
 sg13g2_fill_2 FILLER_4_2205 ();
 sg13g2_fill_1 FILLER_4_2207 ();
 sg13g2_fill_2 FILLER_4_2224 ();
 sg13g2_fill_1 FILLER_4_2226 ();
 sg13g2_fill_2 FILLER_4_2252 ();
 sg13g2_decap_8 FILLER_4_2316 ();
 sg13g2_fill_2 FILLER_4_2369 ();
 sg13g2_decap_8 FILLER_4_2436 ();
 sg13g2_decap_8 FILLER_4_2443 ();
 sg13g2_decap_4 FILLER_4_2450 ();
 sg13g2_fill_2 FILLER_4_2454 ();
 sg13g2_decap_8 FILLER_4_2481 ();
 sg13g2_fill_1 FILLER_4_2488 ();
 sg13g2_decap_4 FILLER_4_2493 ();
 sg13g2_fill_2 FILLER_4_2505 ();
 sg13g2_decap_8 FILLER_4_2528 ();
 sg13g2_decap_8 FILLER_4_2535 ();
 sg13g2_decap_4 FILLER_4_2542 ();
 sg13g2_fill_2 FILLER_4_2546 ();
 sg13g2_fill_2 FILLER_4_2560 ();
 sg13g2_fill_1 FILLER_4_2562 ();
 sg13g2_decap_4 FILLER_4_2576 ();
 sg13g2_fill_2 FILLER_4_2580 ();
 sg13g2_decap_8 FILLER_4_2586 ();
 sg13g2_decap_8 FILLER_4_2593 ();
 sg13g2_decap_8 FILLER_4_2600 ();
 sg13g2_decap_8 FILLER_4_2607 ();
 sg13g2_decap_8 FILLER_4_2614 ();
 sg13g2_decap_8 FILLER_4_2621 ();
 sg13g2_decap_8 FILLER_4_2628 ();
 sg13g2_decap_8 FILLER_4_2635 ();
 sg13g2_decap_8 FILLER_4_2642 ();
 sg13g2_decap_8 FILLER_4_2649 ();
 sg13g2_decap_8 FILLER_4_2656 ();
 sg13g2_decap_8 FILLER_4_2663 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_fill_2 FILLER_5_7 ();
 sg13g2_fill_1 FILLER_5_9 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_4 FILLER_5_70 ();
 sg13g2_fill_2 FILLER_5_84 ();
 sg13g2_fill_1 FILLER_5_86 ();
 sg13g2_fill_2 FILLER_5_92 ();
 sg13g2_fill_1 FILLER_5_94 ();
 sg13g2_decap_4 FILLER_5_105 ();
 sg13g2_fill_1 FILLER_5_113 ();
 sg13g2_decap_8 FILLER_5_118 ();
 sg13g2_fill_1 FILLER_5_125 ();
 sg13g2_decap_8 FILLER_5_152 ();
 sg13g2_decap_4 FILLER_5_159 ();
 sg13g2_fill_2 FILLER_5_163 ();
 sg13g2_fill_2 FILLER_5_178 ();
 sg13g2_fill_2 FILLER_5_206 ();
 sg13g2_fill_1 FILLER_5_208 ();
 sg13g2_fill_1 FILLER_5_213 ();
 sg13g2_decap_8 FILLER_5_240 ();
 sg13g2_fill_2 FILLER_5_247 ();
 sg13g2_fill_1 FILLER_5_269 ();
 sg13g2_fill_1 FILLER_5_274 ();
 sg13g2_fill_2 FILLER_5_286 ();
 sg13g2_fill_1 FILLER_5_288 ();
 sg13g2_fill_2 FILLER_5_324 ();
 sg13g2_fill_1 FILLER_5_340 ();
 sg13g2_decap_8 FILLER_5_345 ();
 sg13g2_decap_8 FILLER_5_352 ();
 sg13g2_fill_2 FILLER_5_359 ();
 sg13g2_fill_2 FILLER_5_404 ();
 sg13g2_fill_1 FILLER_5_406 ();
 sg13g2_decap_4 FILLER_5_421 ();
 sg13g2_fill_1 FILLER_5_425 ();
 sg13g2_fill_2 FILLER_5_431 ();
 sg13g2_decap_8 FILLER_5_437 ();
 sg13g2_fill_2 FILLER_5_448 ();
 sg13g2_fill_1 FILLER_5_450 ();
 sg13g2_decap_8 FILLER_5_477 ();
 sg13g2_decap_4 FILLER_5_484 ();
 sg13g2_fill_1 FILLER_5_498 ();
 sg13g2_fill_2 FILLER_5_504 ();
 sg13g2_fill_1 FILLER_5_514 ();
 sg13g2_decap_8 FILLER_5_524 ();
 sg13g2_decap_8 FILLER_5_531 ();
 sg13g2_decap_4 FILLER_5_538 ();
 sg13g2_fill_1 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_565 ();
 sg13g2_decap_4 FILLER_5_572 ();
 sg13g2_fill_1 FILLER_5_576 ();
 sg13g2_decap_8 FILLER_5_592 ();
 sg13g2_decap_4 FILLER_5_603 ();
 sg13g2_decap_8 FILLER_5_611 ();
 sg13g2_decap_8 FILLER_5_618 ();
 sg13g2_decap_4 FILLER_5_625 ();
 sg13g2_fill_1 FILLER_5_656 ();
 sg13g2_fill_1 FILLER_5_676 ();
 sg13g2_decap_8 FILLER_5_681 ();
 sg13g2_decap_4 FILLER_5_688 ();
 sg13g2_decap_8 FILLER_5_726 ();
 sg13g2_decap_8 FILLER_5_733 ();
 sg13g2_fill_2 FILLER_5_740 ();
 sg13g2_fill_1 FILLER_5_742 ();
 sg13g2_fill_2 FILLER_5_766 ();
 sg13g2_fill_1 FILLER_5_768 ();
 sg13g2_decap_8 FILLER_5_795 ();
 sg13g2_fill_1 FILLER_5_802 ();
 sg13g2_decap_4 FILLER_5_839 ();
 sg13g2_fill_1 FILLER_5_847 ();
 sg13g2_fill_2 FILLER_5_858 ();
 sg13g2_decap_8 FILLER_5_886 ();
 sg13g2_decap_8 FILLER_5_893 ();
 sg13g2_fill_2 FILLER_5_900 ();
 sg13g2_decap_8 FILLER_5_916 ();
 sg13g2_decap_8 FILLER_5_923 ();
 sg13g2_decap_8 FILLER_5_930 ();
 sg13g2_decap_8 FILLER_5_937 ();
 sg13g2_fill_1 FILLER_5_944 ();
 sg13g2_fill_2 FILLER_5_955 ();
 sg13g2_fill_1 FILLER_5_957 ();
 sg13g2_fill_1 FILLER_5_975 ();
 sg13g2_decap_8 FILLER_5_1012 ();
 sg13g2_decap_8 FILLER_5_1019 ();
 sg13g2_decap_8 FILLER_5_1026 ();
 sg13g2_fill_1 FILLER_5_1033 ();
 sg13g2_decap_8 FILLER_5_1056 ();
 sg13g2_fill_2 FILLER_5_1063 ();
 sg13g2_decap_8 FILLER_5_1101 ();
 sg13g2_decap_8 FILLER_5_1108 ();
 sg13g2_decap_4 FILLER_5_1115 ();
 sg13g2_fill_2 FILLER_5_1149 ();
 sg13g2_decap_4 FILLER_5_1191 ();
 sg13g2_fill_1 FILLER_5_1195 ();
 sg13g2_fill_1 FILLER_5_1204 ();
 sg13g2_fill_1 FILLER_5_1210 ();
 sg13g2_fill_2 FILLER_5_1237 ();
 sg13g2_fill_1 FILLER_5_1239 ();
 sg13g2_fill_1 FILLER_5_1271 ();
 sg13g2_decap_8 FILLER_5_1341 ();
 sg13g2_decap_8 FILLER_5_1348 ();
 sg13g2_decap_4 FILLER_5_1355 ();
 sg13g2_fill_2 FILLER_5_1363 ();
 sg13g2_fill_2 FILLER_5_1369 ();
 sg13g2_fill_1 FILLER_5_1397 ();
 sg13g2_fill_1 FILLER_5_1445 ();
 sg13g2_fill_2 FILLER_5_1450 ();
 sg13g2_fill_1 FILLER_5_1462 ();
 sg13g2_decap_8 FILLER_5_1477 ();
 sg13g2_decap_8 FILLER_5_1484 ();
 sg13g2_fill_1 FILLER_5_1491 ();
 sg13g2_fill_2 FILLER_5_1560 ();
 sg13g2_fill_1 FILLER_5_1562 ();
 sg13g2_decap_8 FILLER_5_1570 ();
 sg13g2_fill_2 FILLER_5_1577 ();
 sg13g2_fill_1 FILLER_5_1579 ();
 sg13g2_decap_8 FILLER_5_1665 ();
 sg13g2_fill_2 FILLER_5_1698 ();
 sg13g2_fill_1 FILLER_5_1700 ();
 sg13g2_decap_4 FILLER_5_1722 ();
 sg13g2_fill_2 FILLER_5_1726 ();
 sg13g2_decap_8 FILLER_5_1751 ();
 sg13g2_fill_2 FILLER_5_1758 ();
 sg13g2_decap_4 FILLER_5_1786 ();
 sg13g2_fill_2 FILLER_5_1790 ();
 sg13g2_decap_8 FILLER_5_1818 ();
 sg13g2_fill_2 FILLER_5_1830 ();
 sg13g2_decap_8 FILLER_5_1847 ();
 sg13g2_fill_2 FILLER_5_1854 ();
 sg13g2_decap_8 FILLER_5_1898 ();
 sg13g2_decap_8 FILLER_5_1905 ();
 sg13g2_decap_8 FILLER_5_1912 ();
 sg13g2_decap_4 FILLER_5_1919 ();
 sg13g2_fill_2 FILLER_5_1923 ();
 sg13g2_fill_1 FILLER_5_1952 ();
 sg13g2_fill_1 FILLER_5_1974 ();
 sg13g2_fill_1 FILLER_5_1996 ();
 sg13g2_fill_2 FILLER_5_2001 ();
 sg13g2_decap_4 FILLER_5_2013 ();
 sg13g2_decap_4 FILLER_5_2021 ();
 sg13g2_decap_4 FILLER_5_2035 ();
 sg13g2_fill_2 FILLER_5_2075 ();
 sg13g2_fill_1 FILLER_5_2087 ();
 sg13g2_fill_2 FILLER_5_2092 ();
 sg13g2_fill_1 FILLER_5_2094 ();
 sg13g2_fill_2 FILLER_5_2099 ();
 sg13g2_fill_1 FILLER_5_2101 ();
 sg13g2_fill_2 FILLER_5_2154 ();
 sg13g2_fill_1 FILLER_5_2156 ();
 sg13g2_decap_8 FILLER_5_2161 ();
 sg13g2_fill_2 FILLER_5_2178 ();
 sg13g2_fill_1 FILLER_5_2180 ();
 sg13g2_decap_8 FILLER_5_2240 ();
 sg13g2_decap_8 FILLER_5_2247 ();
 sg13g2_decap_8 FILLER_5_2254 ();
 sg13g2_decap_4 FILLER_5_2261 ();
 sg13g2_fill_2 FILLER_5_2286 ();
 sg13g2_fill_2 FILLER_5_2292 ();
 sg13g2_decap_8 FILLER_5_2320 ();
 sg13g2_fill_2 FILLER_5_2327 ();
 sg13g2_fill_1 FILLER_5_2329 ();
 sg13g2_decap_8 FILLER_5_2334 ();
 sg13g2_decap_8 FILLER_5_2341 ();
 sg13g2_decap_4 FILLER_5_2348 ();
 sg13g2_fill_2 FILLER_5_2352 ();
 sg13g2_decap_4 FILLER_5_2359 ();
 sg13g2_fill_1 FILLER_5_2363 ();
 sg13g2_decap_8 FILLER_5_2374 ();
 sg13g2_decap_8 FILLER_5_2381 ();
 sg13g2_fill_1 FILLER_5_2388 ();
 sg13g2_decap_4 FILLER_5_2393 ();
 sg13g2_fill_1 FILLER_5_2397 ();
 sg13g2_decap_8 FILLER_5_2442 ();
 sg13g2_fill_1 FILLER_5_2493 ();
 sg13g2_fill_2 FILLER_5_2506 ();
 sg13g2_fill_1 FILLER_5_2508 ();
 sg13g2_fill_2 FILLER_5_2519 ();
 sg13g2_fill_1 FILLER_5_2521 ();
 sg13g2_decap_8 FILLER_5_2532 ();
 sg13g2_decap_4 FILLER_5_2539 ();
 sg13g2_decap_8 FILLER_5_2564 ();
 sg13g2_fill_1 FILLER_5_2571 ();
 sg13g2_fill_1 FILLER_5_2582 ();
 sg13g2_decap_8 FILLER_5_2591 ();
 sg13g2_decap_8 FILLER_5_2598 ();
 sg13g2_decap_8 FILLER_5_2605 ();
 sg13g2_fill_2 FILLER_5_2612 ();
 sg13g2_fill_1 FILLER_5_2614 ();
 sg13g2_decap_8 FILLER_5_2619 ();
 sg13g2_decap_8 FILLER_5_2626 ();
 sg13g2_decap_8 FILLER_5_2633 ();
 sg13g2_decap_8 FILLER_5_2640 ();
 sg13g2_decap_8 FILLER_5_2647 ();
 sg13g2_decap_8 FILLER_5_2654 ();
 sg13g2_decap_8 FILLER_5_2661 ();
 sg13g2_fill_2 FILLER_5_2668 ();
 sg13g2_fill_2 FILLER_6_0 ();
 sg13g2_fill_2 FILLER_6_37 ();
 sg13g2_fill_1 FILLER_6_39 ();
 sg13g2_fill_2 FILLER_6_45 ();
 sg13g2_fill_2 FILLER_6_52 ();
 sg13g2_fill_1 FILLER_6_54 ();
 sg13g2_decap_4 FILLER_6_112 ();
 sg13g2_fill_1 FILLER_6_116 ();
 sg13g2_decap_4 FILLER_6_153 ();
 sg13g2_fill_1 FILLER_6_157 ();
 sg13g2_fill_1 FILLER_6_184 ();
 sg13g2_fill_2 FILLER_6_199 ();
 sg13g2_fill_1 FILLER_6_201 ();
 sg13g2_decap_8 FILLER_6_214 ();
 sg13g2_fill_1 FILLER_6_221 ();
 sg13g2_decap_8 FILLER_6_239 ();
 sg13g2_decap_8 FILLER_6_246 ();
 sg13g2_decap_8 FILLER_6_253 ();
 sg13g2_decap_8 FILLER_6_260 ();
 sg13g2_decap_8 FILLER_6_267 ();
 sg13g2_decap_8 FILLER_6_274 ();
 sg13g2_decap_4 FILLER_6_281 ();
 sg13g2_fill_1 FILLER_6_285 ();
 sg13g2_fill_1 FILLER_6_306 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_fill_1 FILLER_6_335 ();
 sg13g2_decap_8 FILLER_6_344 ();
 sg13g2_decap_8 FILLER_6_351 ();
 sg13g2_decap_4 FILLER_6_358 ();
 sg13g2_fill_1 FILLER_6_362 ();
 sg13g2_fill_2 FILLER_6_372 ();
 sg13g2_fill_2 FILLER_6_424 ();
 sg13g2_fill_1 FILLER_6_521 ();
 sg13g2_decap_8 FILLER_6_526 ();
 sg13g2_decap_8 FILLER_6_533 ();
 sg13g2_decap_8 FILLER_6_540 ();
 sg13g2_fill_2 FILLER_6_547 ();
 sg13g2_fill_1 FILLER_6_549 ();
 sg13g2_decap_8 FILLER_6_554 ();
 sg13g2_decap_8 FILLER_6_561 ();
 sg13g2_decap_8 FILLER_6_568 ();
 sg13g2_fill_1 FILLER_6_592 ();
 sg13g2_decap_8 FILLER_6_619 ();
 sg13g2_decap_4 FILLER_6_626 ();
 sg13g2_fill_1 FILLER_6_630 ();
 sg13g2_decap_4 FILLER_6_639 ();
 sg13g2_fill_2 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_688 ();
 sg13g2_decap_4 FILLER_6_695 ();
 sg13g2_fill_2 FILLER_6_703 ();
 sg13g2_fill_2 FILLER_6_731 ();
 sg13g2_decap_4 FILLER_6_759 ();
 sg13g2_fill_2 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_769 ();
 sg13g2_fill_1 FILLER_6_776 ();
 sg13g2_decap_8 FILLER_6_781 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_4 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_825 ();
 sg13g2_decap_8 FILLER_6_832 ();
 sg13g2_decap_8 FILLER_6_839 ();
 sg13g2_decap_4 FILLER_6_846 ();
 sg13g2_fill_2 FILLER_6_850 ();
 sg13g2_decap_4 FILLER_6_930 ();
 sg13g2_fill_1 FILLER_6_934 ();
 sg13g2_decap_4 FILLER_6_945 ();
 sg13g2_fill_2 FILLER_6_975 ();
 sg13g2_fill_1 FILLER_6_1003 ();
 sg13g2_decap_4 FILLER_6_1022 ();
 sg13g2_fill_1 FILLER_6_1046 ();
 sg13g2_fill_1 FILLER_6_1068 ();
 sg13g2_fill_2 FILLER_6_1079 ();
 sg13g2_fill_2 FILLER_6_1085 ();
 sg13g2_decap_4 FILLER_6_1113 ();
 sg13g2_fill_1 FILLER_6_1117 ();
 sg13g2_fill_1 FILLER_6_1144 ();
 sg13g2_decap_8 FILLER_6_1155 ();
 sg13g2_decap_8 FILLER_6_1162 ();
 sg13g2_fill_1 FILLER_6_1169 ();
 sg13g2_fill_2 FILLER_6_1174 ();
 sg13g2_fill_1 FILLER_6_1176 ();
 sg13g2_fill_2 FILLER_6_1197 ();
 sg13g2_decap_8 FILLER_6_1203 ();
 sg13g2_fill_1 FILLER_6_1215 ();
 sg13g2_decap_4 FILLER_6_1220 ();
 sg13g2_fill_2 FILLER_6_1224 ();
 sg13g2_decap_4 FILLER_6_1234 ();
 sg13g2_fill_2 FILLER_6_1238 ();
 sg13g2_decap_8 FILLER_6_1265 ();
 sg13g2_fill_1 FILLER_6_1272 ();
 sg13g2_fill_1 FILLER_6_1288 ();
 sg13g2_fill_1 FILLER_6_1353 ();
 sg13g2_decap_4 FILLER_6_1364 ();
 sg13g2_fill_1 FILLER_6_1368 ();
 sg13g2_fill_1 FILLER_6_1373 ();
 sg13g2_fill_1 FILLER_6_1382 ();
 sg13g2_fill_2 FILLER_6_1413 ();
 sg13g2_fill_1 FILLER_6_1415 ();
 sg13g2_fill_2 FILLER_6_1457 ();
 sg13g2_decap_8 FILLER_6_1485 ();
 sg13g2_decap_4 FILLER_6_1492 ();
 sg13g2_decap_8 FILLER_6_1566 ();
 sg13g2_decap_8 FILLER_6_1573 ();
 sg13g2_decap_8 FILLER_6_1580 ();
 sg13g2_decap_8 FILLER_6_1613 ();
 sg13g2_fill_1 FILLER_6_1620 ();
 sg13g2_decap_4 FILLER_6_1625 ();
 sg13g2_fill_2 FILLER_6_1644 ();
 sg13g2_fill_2 FILLER_6_1658 ();
 sg13g2_fill_1 FILLER_6_1660 ();
 sg13g2_decap_8 FILLER_6_1665 ();
 sg13g2_fill_1 FILLER_6_1672 ();
 sg13g2_fill_2 FILLER_6_1687 ();
 sg13g2_decap_8 FILLER_6_1725 ();
 sg13g2_decap_8 FILLER_6_1732 ();
 sg13g2_decap_8 FILLER_6_1739 ();
 sg13g2_decap_4 FILLER_6_1746 ();
 sg13g2_fill_2 FILLER_6_1750 ();
 sg13g2_decap_8 FILLER_6_1760 ();
 sg13g2_fill_1 FILLER_6_1767 ();
 sg13g2_decap_8 FILLER_6_1772 ();
 sg13g2_decap_8 FILLER_6_1779 ();
 sg13g2_decap_8 FILLER_6_1786 ();
 sg13g2_fill_1 FILLER_6_1802 ();
 sg13g2_fill_1 FILLER_6_1845 ();
 sg13g2_fill_2 FILLER_6_1851 ();
 sg13g2_decap_8 FILLER_6_1925 ();
 sg13g2_decap_4 FILLER_6_1932 ();
 sg13g2_fill_2 FILLER_6_1940 ();
 sg13g2_fill_1 FILLER_6_1942 ();
 sg13g2_decap_8 FILLER_6_1947 ();
 sg13g2_decap_8 FILLER_6_1954 ();
 sg13g2_fill_1 FILLER_6_1961 ();
 sg13g2_decap_8 FILLER_6_1966 ();
 sg13g2_decap_8 FILLER_6_1973 ();
 sg13g2_decap_4 FILLER_6_1980 ();
 sg13g2_fill_2 FILLER_6_1984 ();
 sg13g2_decap_8 FILLER_6_1996 ();
 sg13g2_decap_8 FILLER_6_2003 ();
 sg13g2_decap_8 FILLER_6_2010 ();
 sg13g2_fill_2 FILLER_6_2017 ();
 sg13g2_fill_1 FILLER_6_2019 ();
 sg13g2_decap_8 FILLER_6_2030 ();
 sg13g2_decap_4 FILLER_6_2037 ();
 sg13g2_decap_8 FILLER_6_2051 ();
 sg13g2_fill_2 FILLER_6_2058 ();
 sg13g2_decap_8 FILLER_6_2064 ();
 sg13g2_decap_8 FILLER_6_2071 ();
 sg13g2_fill_1 FILLER_6_2091 ();
 sg13g2_decap_4 FILLER_6_2106 ();
 sg13g2_fill_1 FILLER_6_2110 ();
 sg13g2_fill_2 FILLER_6_2121 ();
 sg13g2_fill_1 FILLER_6_2123 ();
 sg13g2_fill_2 FILLER_6_2134 ();
 sg13g2_fill_1 FILLER_6_2136 ();
 sg13g2_decap_8 FILLER_6_2141 ();
 sg13g2_fill_2 FILLER_6_2148 ();
 sg13g2_fill_1 FILLER_6_2150 ();
 sg13g2_decap_8 FILLER_6_2155 ();
 sg13g2_decap_8 FILLER_6_2162 ();
 sg13g2_fill_1 FILLER_6_2179 ();
 sg13g2_fill_1 FILLER_6_2190 ();
 sg13g2_fill_1 FILLER_6_2217 ();
 sg13g2_fill_2 FILLER_6_2244 ();
 sg13g2_fill_2 FILLER_6_2251 ();
 sg13g2_fill_1 FILLER_6_2253 ();
 sg13g2_decap_4 FILLER_6_2259 ();
 sg13g2_fill_1 FILLER_6_2263 ();
 sg13g2_decap_4 FILLER_6_2282 ();
 sg13g2_fill_1 FILLER_6_2312 ();
 sg13g2_decap_8 FILLER_6_2349 ();
 sg13g2_fill_1 FILLER_6_2356 ();
 sg13g2_fill_2 FILLER_6_2361 ();
 sg13g2_decap_4 FILLER_6_2399 ();
 sg13g2_fill_1 FILLER_6_2403 ();
 sg13g2_fill_2 FILLER_6_2439 ();
 sg13g2_fill_2 FILLER_6_2451 ();
 sg13g2_fill_2 FILLER_6_2457 ();
 sg13g2_fill_1 FILLER_6_2459 ();
 sg13g2_fill_2 FILLER_6_2489 ();
 sg13g2_decap_8 FILLER_6_2521 ();
 sg13g2_fill_2 FILLER_6_2528 ();
 sg13g2_decap_8 FILLER_6_2602 ();
 sg13g2_fill_2 FILLER_6_2609 ();
 sg13g2_decap_4 FILLER_6_2637 ();
 sg13g2_decap_8 FILLER_6_2645 ();
 sg13g2_decap_8 FILLER_6_2652 ();
 sg13g2_decap_8 FILLER_6_2659 ();
 sg13g2_decap_4 FILLER_6_2666 ();
 sg13g2_decap_4 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_4 ();
 sg13g2_decap_8 FILLER_7_10 ();
 sg13g2_fill_1 FILLER_7_17 ();
 sg13g2_fill_2 FILLER_7_21 ();
 sg13g2_fill_2 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_40 ();
 sg13g2_decap_4 FILLER_7_47 ();
 sg13g2_decap_4 FILLER_7_55 ();
 sg13g2_fill_2 FILLER_7_67 ();
 sg13g2_fill_2 FILLER_7_129 ();
 sg13g2_fill_1 FILLER_7_131 ();
 sg13g2_fill_2 FILLER_7_167 ();
 sg13g2_fill_1 FILLER_7_169 ();
 sg13g2_fill_2 FILLER_7_175 ();
 sg13g2_fill_1 FILLER_7_177 ();
 sg13g2_decap_4 FILLER_7_240 ();
 sg13g2_fill_1 FILLER_7_244 ();
 sg13g2_decap_4 FILLER_7_271 ();
 sg13g2_fill_1 FILLER_7_275 ();
 sg13g2_fill_2 FILLER_7_281 ();
 sg13g2_fill_1 FILLER_7_283 ();
 sg13g2_decap_4 FILLER_7_292 ();
 sg13g2_decap_8 FILLER_7_313 ();
 sg13g2_fill_2 FILLER_7_320 ();
 sg13g2_fill_1 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_352 ();
 sg13g2_fill_1 FILLER_7_359 ();
 sg13g2_fill_2 FILLER_7_394 ();
 sg13g2_decap_4 FILLER_7_401 ();
 sg13g2_decap_8 FILLER_7_409 ();
 sg13g2_decap_8 FILLER_7_416 ();
 sg13g2_fill_2 FILLER_7_423 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_fill_1 FILLER_7_440 ();
 sg13g2_fill_1 FILLER_7_451 ();
 sg13g2_fill_2 FILLER_7_457 ();
 sg13g2_fill_1 FILLER_7_463 ();
 sg13g2_decap_4 FILLER_7_488 ();
 sg13g2_decap_4 FILLER_7_496 ();
 sg13g2_fill_2 FILLER_7_500 ();
 sg13g2_fill_1 FILLER_7_517 ();
 sg13g2_fill_2 FILLER_7_537 ();
 sg13g2_fill_2 FILLER_7_573 ();
 sg13g2_fill_1 FILLER_7_593 ();
 sg13g2_decap_8 FILLER_7_638 ();
 sg13g2_fill_2 FILLER_7_659 ();
 sg13g2_fill_2 FILLER_7_673 ();
 sg13g2_fill_1 FILLER_7_675 ();
 sg13g2_fill_2 FILLER_7_681 ();
 sg13g2_fill_1 FILLER_7_683 ();
 sg13g2_fill_2 FILLER_7_689 ();
 sg13g2_fill_1 FILLER_7_691 ();
 sg13g2_fill_1 FILLER_7_706 ();
 sg13g2_fill_1 FILLER_7_721 ();
 sg13g2_fill_2 FILLER_7_727 ();
 sg13g2_fill_1 FILLER_7_733 ();
 sg13g2_decap_8 FILLER_7_769 ();
 sg13g2_decap_8 FILLER_7_776 ();
 sg13g2_decap_8 FILLER_7_783 ();
 sg13g2_decap_8 FILLER_7_790 ();
 sg13g2_decap_4 FILLER_7_797 ();
 sg13g2_fill_2 FILLER_7_801 ();
 sg13g2_decap_4 FILLER_7_817 ();
 sg13g2_fill_2 FILLER_7_821 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_fill_2 FILLER_7_859 ();
 sg13g2_decap_8 FILLER_7_901 ();
 sg13g2_decap_8 FILLER_7_912 ();
 sg13g2_fill_1 FILLER_7_919 ();
 sg13g2_decap_4 FILLER_7_1029 ();
 sg13g2_fill_1 FILLER_7_1033 ();
 sg13g2_decap_4 FILLER_7_1073 ();
 sg13g2_fill_1 FILLER_7_1077 ();
 sg13g2_decap_8 FILLER_7_1128 ();
 sg13g2_decap_8 FILLER_7_1135 ();
 sg13g2_decap_8 FILLER_7_1142 ();
 sg13g2_decap_8 FILLER_7_1149 ();
 sg13g2_decap_8 FILLER_7_1156 ();
 sg13g2_decap_8 FILLER_7_1163 ();
 sg13g2_fill_2 FILLER_7_1170 ();
 sg13g2_decap_4 FILLER_7_1176 ();
 sg13g2_decap_4 FILLER_7_1188 ();
 sg13g2_fill_1 FILLER_7_1192 ();
 sg13g2_decap_8 FILLER_7_1197 ();
 sg13g2_decap_4 FILLER_7_1208 ();
 sg13g2_fill_1 FILLER_7_1212 ();
 sg13g2_fill_2 FILLER_7_1217 ();
 sg13g2_decap_8 FILLER_7_1235 ();
 sg13g2_decap_8 FILLER_7_1242 ();
 sg13g2_fill_2 FILLER_7_1249 ();
 sg13g2_decap_4 FILLER_7_1264 ();
 sg13g2_fill_1 FILLER_7_1268 ();
 sg13g2_decap_8 FILLER_7_1350 ();
 sg13g2_decap_8 FILLER_7_1357 ();
 sg13g2_decap_8 FILLER_7_1364 ();
 sg13g2_decap_8 FILLER_7_1371 ();
 sg13g2_decap_4 FILLER_7_1378 ();
 sg13g2_fill_2 FILLER_7_1394 ();
 sg13g2_fill_1 FILLER_7_1396 ();
 sg13g2_decap_8 FILLER_7_1401 ();
 sg13g2_fill_2 FILLER_7_1408 ();
 sg13g2_fill_2 FILLER_7_1415 ();
 sg13g2_fill_2 FILLER_7_1456 ();
 sg13g2_fill_1 FILLER_7_1484 ();
 sg13g2_fill_1 FILLER_7_1489 ();
 sg13g2_fill_2 FILLER_7_1516 ();
 sg13g2_fill_2 FILLER_7_1528 ();
 sg13g2_fill_2 FILLER_7_1534 ();
 sg13g2_decap_4 FILLER_7_1576 ();
 sg13g2_fill_1 FILLER_7_1580 ();
 sg13g2_fill_2 FILLER_7_1601 ();
 sg13g2_fill_2 FILLER_7_1615 ();
 sg13g2_fill_2 FILLER_7_1627 ();
 sg13g2_fill_2 FILLER_7_1639 ();
 sg13g2_fill_1 FILLER_7_1641 ();
 sg13g2_decap_8 FILLER_7_1656 ();
 sg13g2_decap_8 FILLER_7_1663 ();
 sg13g2_decap_8 FILLER_7_1670 ();
 sg13g2_fill_2 FILLER_7_1677 ();
 sg13g2_decap_8 FILLER_7_1712 ();
 sg13g2_decap_8 FILLER_7_1719 ();
 sg13g2_decap_8 FILLER_7_1726 ();
 sg13g2_decap_8 FILLER_7_1733 ();
 sg13g2_decap_8 FILLER_7_1766 ();
 sg13g2_decap_4 FILLER_7_1773 ();
 sg13g2_fill_1 FILLER_7_1807 ();
 sg13g2_fill_1 FILLER_7_1825 ();
 sg13g2_fill_1 FILLER_7_1839 ();
 sg13g2_fill_2 FILLER_7_1866 ();
 sg13g2_fill_1 FILLER_7_1890 ();
 sg13g2_fill_1 FILLER_7_1917 ();
 sg13g2_fill_2 FILLER_7_1922 ();
 sg13g2_decap_8 FILLER_7_1928 ();
 sg13g2_fill_1 FILLER_7_1935 ();
 sg13g2_fill_1 FILLER_7_1944 ();
 sg13g2_fill_1 FILLER_7_1964 ();
 sg13g2_decap_8 FILLER_7_1974 ();
 sg13g2_decap_8 FILLER_7_1981 ();
 sg13g2_decap_8 FILLER_7_1988 ();
 sg13g2_decap_8 FILLER_7_1995 ();
 sg13g2_decap_8 FILLER_7_2002 ();
 sg13g2_fill_2 FILLER_7_2009 ();
 sg13g2_decap_8 FILLER_7_2021 ();
 sg13g2_fill_2 FILLER_7_2028 ();
 sg13g2_decap_4 FILLER_7_2060 ();
 sg13g2_fill_2 FILLER_7_2064 ();
 sg13g2_fill_1 FILLER_7_2084 ();
 sg13g2_decap_8 FILLER_7_2121 ();
 sg13g2_fill_2 FILLER_7_2128 ();
 sg13g2_fill_1 FILLER_7_2130 ();
 sg13g2_decap_8 FILLER_7_2135 ();
 sg13g2_decap_8 FILLER_7_2142 ();
 sg13g2_fill_2 FILLER_7_2149 ();
 sg13g2_decap_8 FILLER_7_2163 ();
 sg13g2_decap_4 FILLER_7_2170 ();
 sg13g2_fill_1 FILLER_7_2188 ();
 sg13g2_decap_4 FILLER_7_2238 ();
 sg13g2_decap_8 FILLER_7_2252 ();
 sg13g2_decap_4 FILLER_7_2259 ();
 sg13g2_fill_1 FILLER_7_2284 ();
 sg13g2_fill_1 FILLER_7_2295 ();
 sg13g2_decap_4 FILLER_7_2310 ();
 sg13g2_decap_4 FILLER_7_2335 ();
 sg13g2_fill_2 FILLER_7_2339 ();
 sg13g2_decap_4 FILLER_7_2345 ();
 sg13g2_fill_1 FILLER_7_2349 ();
 sg13g2_decap_4 FILLER_7_2386 ();
 sg13g2_fill_1 FILLER_7_2390 ();
 sg13g2_decap_4 FILLER_7_2404 ();
 sg13g2_fill_2 FILLER_7_2408 ();
 sg13g2_fill_2 FILLER_7_2420 ();
 sg13g2_fill_1 FILLER_7_2422 ();
 sg13g2_decap_4 FILLER_7_2520 ();
 sg13g2_fill_1 FILLER_7_2524 ();
 sg13g2_decap_8 FILLER_7_2659 ();
 sg13g2_decap_4 FILLER_7_2666 ();
 sg13g2_fill_2 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_34 ();
 sg13g2_fill_1 FILLER_8_45 ();
 sg13g2_fill_1 FILLER_8_50 ();
 sg13g2_fill_1 FILLER_8_56 ();
 sg13g2_fill_2 FILLER_8_62 ();
 sg13g2_fill_1 FILLER_8_64 ();
 sg13g2_fill_2 FILLER_8_79 ();
 sg13g2_fill_1 FILLER_8_81 ();
 sg13g2_fill_1 FILLER_8_90 ();
 sg13g2_decap_8 FILLER_8_127 ();
 sg13g2_fill_2 FILLER_8_134 ();
 sg13g2_fill_2 FILLER_8_140 ();
 sg13g2_fill_1 FILLER_8_142 ();
 sg13g2_fill_2 FILLER_8_147 ();
 sg13g2_fill_1 FILLER_8_149 ();
 sg13g2_decap_8 FILLER_8_167 ();
 sg13g2_fill_1 FILLER_8_187 ();
 sg13g2_fill_1 FILLER_8_192 ();
 sg13g2_fill_1 FILLER_8_219 ();
 sg13g2_fill_1 FILLER_8_250 ();
 sg13g2_fill_2 FILLER_8_255 ();
 sg13g2_fill_2 FILLER_8_283 ();
 sg13g2_fill_1 FILLER_8_293 ();
 sg13g2_fill_2 FILLER_8_302 ();
 sg13g2_fill_2 FILLER_8_312 ();
 sg13g2_fill_2 FILLER_8_319 ();
 sg13g2_decap_4 FILLER_8_351 ();
 sg13g2_fill_1 FILLER_8_355 ();
 sg13g2_fill_1 FILLER_8_362 ();
 sg13g2_fill_2 FILLER_8_366 ();
 sg13g2_fill_2 FILLER_8_373 ();
 sg13g2_fill_2 FILLER_8_379 ();
 sg13g2_fill_1 FILLER_8_381 ();
 sg13g2_decap_8 FILLER_8_397 ();
 sg13g2_decap_8 FILLER_8_404 ();
 sg13g2_fill_1 FILLER_8_411 ();
 sg13g2_decap_4 FILLER_8_452 ();
 sg13g2_fill_1 FILLER_8_456 ();
 sg13g2_fill_2 FILLER_8_461 ();
 sg13g2_fill_1 FILLER_8_463 ();
 sg13g2_fill_2 FILLER_8_469 ();
 sg13g2_fill_1 FILLER_8_471 ();
 sg13g2_decap_4 FILLER_8_477 ();
 sg13g2_fill_2 FILLER_8_486 ();
 sg13g2_decap_4 FILLER_8_493 ();
 sg13g2_fill_1 FILLER_8_497 ();
 sg13g2_fill_1 FILLER_8_514 ();
 sg13g2_decap_4 FILLER_8_577 ();
 sg13g2_decap_4 FILLER_8_601 ();
 sg13g2_fill_1 FILLER_8_605 ();
 sg13g2_decap_8 FILLER_8_610 ();
 sg13g2_decap_8 FILLER_8_617 ();
 sg13g2_decap_8 FILLER_8_624 ();
 sg13g2_decap_8 FILLER_8_631 ();
 sg13g2_fill_1 FILLER_8_638 ();
 sg13g2_fill_1 FILLER_8_665 ();
 sg13g2_fill_1 FILLER_8_702 ();
 sg13g2_fill_1 FILLER_8_712 ();
 sg13g2_fill_1 FILLER_8_722 ();
 sg13g2_fill_1 FILLER_8_728 ();
 sg13g2_fill_2 FILLER_8_752 ();
 sg13g2_decap_8 FILLER_8_764 ();
 sg13g2_fill_2 FILLER_8_771 ();
 sg13g2_decap_4 FILLER_8_797 ();
 sg13g2_decap_8 FILLER_8_857 ();
 sg13g2_decap_4 FILLER_8_864 ();
 sg13g2_fill_2 FILLER_8_868 ();
 sg13g2_fill_2 FILLER_8_883 ();
 sg13g2_fill_1 FILLER_8_885 ();
 sg13g2_fill_1 FILLER_8_890 ();
 sg13g2_fill_2 FILLER_8_927 ();
 sg13g2_fill_1 FILLER_8_929 ();
 sg13g2_decap_4 FILLER_8_977 ();
 sg13g2_fill_2 FILLER_8_1037 ();
 sg13g2_fill_2 FILLER_8_1043 ();
 sg13g2_fill_1 FILLER_8_1045 ();
 sg13g2_fill_2 FILLER_8_1072 ();
 sg13g2_fill_1 FILLER_8_1095 ();
 sg13g2_decap_4 FILLER_8_1100 ();
 sg13g2_fill_1 FILLER_8_1104 ();
 sg13g2_decap_8 FILLER_8_1109 ();
 sg13g2_decap_8 FILLER_8_1116 ();
 sg13g2_decap_8 FILLER_8_1123 ();
 sg13g2_decap_4 FILLER_8_1130 ();
 sg13g2_fill_2 FILLER_8_1134 ();
 sg13g2_fill_2 FILLER_8_1172 ();
 sg13g2_decap_4 FILLER_8_1227 ();
 sg13g2_fill_1 FILLER_8_1231 ();
 sg13g2_decap_4 FILLER_8_1242 ();
 sg13g2_fill_2 FILLER_8_1315 ();
 sg13g2_fill_2 FILLER_8_1343 ();
 sg13g2_fill_1 FILLER_8_1345 ();
 sg13g2_decap_8 FILLER_8_1350 ();
 sg13g2_decap_8 FILLER_8_1357 ();
 sg13g2_decap_8 FILLER_8_1364 ();
 sg13g2_fill_1 FILLER_8_1371 ();
 sg13g2_decap_4 FILLER_8_1377 ();
 sg13g2_fill_1 FILLER_8_1381 ();
 sg13g2_fill_1 FILLER_8_1386 ();
 sg13g2_fill_2 FILLER_8_1421 ();
 sg13g2_fill_2 FILLER_8_1427 ();
 sg13g2_fill_1 FILLER_8_1429 ();
 sg13g2_decap_4 FILLER_8_1434 ();
 sg13g2_fill_2 FILLER_8_1438 ();
 sg13g2_fill_2 FILLER_8_1466 ();
 sg13g2_fill_1 FILLER_8_1468 ();
 sg13g2_decap_4 FILLER_8_1473 ();
 sg13g2_fill_2 FILLER_8_1477 ();
 sg13g2_decap_4 FILLER_8_1532 ();
 sg13g2_fill_2 FILLER_8_1536 ();
 sg13g2_fill_2 FILLER_8_1610 ();
 sg13g2_decap_4 FILLER_8_1622 ();
 sg13g2_fill_1 FILLER_8_1626 ();
 sg13g2_decap_4 FILLER_8_1671 ();
 sg13g2_fill_2 FILLER_8_1675 ();
 sg13g2_fill_1 FILLER_8_1703 ();
 sg13g2_fill_2 FILLER_8_1714 ();
 sg13g2_fill_1 FILLER_8_1742 ();
 sg13g2_fill_2 FILLER_8_1769 ();
 sg13g2_decap_8 FILLER_8_1801 ();
 sg13g2_decap_8 FILLER_8_1808 ();
 sg13g2_decap_4 FILLER_8_1815 ();
 sg13g2_decap_8 FILLER_8_1863 ();
 sg13g2_decap_8 FILLER_8_1870 ();
 sg13g2_decap_4 FILLER_8_1877 ();
 sg13g2_fill_1 FILLER_8_1881 ();
 sg13g2_fill_1 FILLER_8_1897 ();
 sg13g2_decap_4 FILLER_8_1924 ();
 sg13g2_fill_2 FILLER_8_1928 ();
 sg13g2_fill_2 FILLER_8_1950 ();
 sg13g2_fill_1 FILLER_8_1952 ();
 sg13g2_fill_1 FILLER_8_1979 ();
 sg13g2_fill_1 FILLER_8_2006 ();
 sg13g2_fill_1 FILLER_8_2033 ();
 sg13g2_fill_1 FILLER_8_2038 ();
 sg13g2_decap_4 FILLER_8_2065 ();
 sg13g2_fill_1 FILLER_8_2121 ();
 sg13g2_fill_2 FILLER_8_2148 ();
 sg13g2_fill_1 FILLER_8_2150 ();
 sg13g2_fill_2 FILLER_8_2159 ();
 sg13g2_fill_1 FILLER_8_2165 ();
 sg13g2_fill_2 FILLER_8_2196 ();
 sg13g2_fill_1 FILLER_8_2198 ();
 sg13g2_fill_1 FILLER_8_2274 ();
 sg13g2_decap_4 FILLER_8_2301 ();
 sg13g2_decap_8 FILLER_8_2331 ();
 sg13g2_decap_8 FILLER_8_2338 ();
 sg13g2_fill_2 FILLER_8_2345 ();
 sg13g2_fill_1 FILLER_8_2347 ();
 sg13g2_decap_4 FILLER_8_2356 ();
 sg13g2_fill_1 FILLER_8_2360 ();
 sg13g2_fill_1 FILLER_8_2365 ();
 sg13g2_fill_2 FILLER_8_2392 ();
 sg13g2_fill_2 FILLER_8_2420 ();
 sg13g2_fill_2 FILLER_8_2493 ();
 sg13g2_fill_1 FILLER_8_2495 ();
 sg13g2_fill_2 FILLER_8_2536 ();
 sg13g2_fill_1 FILLER_8_2564 ();
 sg13g2_fill_2 FILLER_8_2569 ();
 sg13g2_fill_1 FILLER_8_2571 ();
 sg13g2_decap_4 FILLER_8_2622 ();
 sg13g2_decap_8 FILLER_8_2656 ();
 sg13g2_decap_8 FILLER_8_2663 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_4 FILLER_9_7 ();
 sg13g2_fill_1 FILLER_9_11 ();
 sg13g2_fill_2 FILLER_9_16 ();
 sg13g2_fill_1 FILLER_9_18 ();
 sg13g2_fill_1 FILLER_9_75 ();
 sg13g2_fill_2 FILLER_9_95 ();
 sg13g2_decap_8 FILLER_9_123 ();
 sg13g2_decap_8 FILLER_9_130 ();
 sg13g2_fill_1 FILLER_9_137 ();
 sg13g2_fill_1 FILLER_9_148 ();
 sg13g2_fill_1 FILLER_9_166 ();
 sg13g2_decap_8 FILLER_9_232 ();
 sg13g2_decap_4 FILLER_9_239 ();
 sg13g2_fill_2 FILLER_9_248 ();
 sg13g2_fill_1 FILLER_9_250 ();
 sg13g2_fill_2 FILLER_9_266 ();
 sg13g2_fill_1 FILLER_9_345 ();
 sg13g2_decap_4 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_398 ();
 sg13g2_decap_8 FILLER_9_405 ();
 sg13g2_decap_4 FILLER_9_412 ();
 sg13g2_fill_1 FILLER_9_416 ();
 sg13g2_fill_1 FILLER_9_492 ();
 sg13g2_fill_1 FILLER_9_497 ();
 sg13g2_fill_1 FILLER_9_524 ();
 sg13g2_fill_1 FILLER_9_556 ();
 sg13g2_fill_1 FILLER_9_561 ();
 sg13g2_fill_1 FILLER_9_572 ();
 sg13g2_decap_4 FILLER_9_582 ();
 sg13g2_fill_2 FILLER_9_616 ();
 sg13g2_fill_2 FILLER_9_622 ();
 sg13g2_fill_1 FILLER_9_624 ();
 sg13g2_fill_2 FILLER_9_630 ();
 sg13g2_fill_1 FILLER_9_663 ();
 sg13g2_fill_1 FILLER_9_669 ();
 sg13g2_fill_1 FILLER_9_675 ();
 sg13g2_decap_4 FILLER_9_695 ();
 sg13g2_fill_1 FILLER_9_699 ();
 sg13g2_fill_1 FILLER_9_730 ();
 sg13g2_fill_2 FILLER_9_740 ();
 sg13g2_fill_2 FILLER_9_751 ();
 sg13g2_decap_4 FILLER_9_770 ();
 sg13g2_fill_1 FILLER_9_800 ();
 sg13g2_fill_2 FILLER_9_827 ();
 sg13g2_fill_1 FILLER_9_829 ();
 sg13g2_decap_8 FILLER_9_891 ();
 sg13g2_fill_1 FILLER_9_908 ();
 sg13g2_decap_4 FILLER_9_943 ();
 sg13g2_fill_2 FILLER_9_952 ();
 sg13g2_fill_1 FILLER_9_954 ();
 sg13g2_decap_8 FILLER_9_969 ();
 sg13g2_decap_8 FILLER_9_976 ();
 sg13g2_fill_1 FILLER_9_983 ();
 sg13g2_fill_2 FILLER_9_1002 ();
 sg13g2_fill_1 FILLER_9_1014 ();
 sg13g2_fill_2 FILLER_9_1019 ();
 sg13g2_fill_2 FILLER_9_1031 ();
 sg13g2_fill_2 FILLER_9_1059 ();
 sg13g2_fill_1 FILLER_9_1061 ();
 sg13g2_fill_1 FILLER_9_1066 ();
 sg13g2_decap_8 FILLER_9_1077 ();
 sg13g2_decap_8 FILLER_9_1084 ();
 sg13g2_decap_8 FILLER_9_1091 ();
 sg13g2_fill_2 FILLER_9_1098 ();
 sg13g2_fill_1 FILLER_9_1100 ();
 sg13g2_decap_8 FILLER_9_1105 ();
 sg13g2_decap_8 FILLER_9_1112 ();
 sg13g2_decap_8 FILLER_9_1119 ();
 sg13g2_fill_2 FILLER_9_1126 ();
 sg13g2_decap_8 FILLER_9_1164 ();
 sg13g2_fill_1 FILLER_9_1197 ();
 sg13g2_decap_4 FILLER_9_1315 ();
 sg13g2_fill_2 FILLER_9_1319 ();
 sg13g2_decap_8 FILLER_9_1325 ();
 sg13g2_decap_8 FILLER_9_1332 ();
 sg13g2_decap_4 FILLER_9_1339 ();
 sg13g2_decap_8 FILLER_9_1373 ();
 sg13g2_decap_8 FILLER_9_1380 ();
 sg13g2_decap_4 FILLER_9_1387 ();
 sg13g2_fill_1 FILLER_9_1391 ();
 sg13g2_decap_8 FILLER_9_1423 ();
 sg13g2_decap_8 FILLER_9_1430 ();
 sg13g2_fill_2 FILLER_9_1437 ();
 sg13g2_decap_8 FILLER_9_1453 ();
 sg13g2_fill_2 FILLER_9_1460 ();
 sg13g2_fill_1 FILLER_9_1462 ();
 sg13g2_fill_2 FILLER_9_1473 ();
 sg13g2_fill_1 FILLER_9_1475 ();
 sg13g2_fill_2 FILLER_9_1596 ();
 sg13g2_fill_2 FILLER_9_1608 ();
 sg13g2_fill_1 FILLER_9_1610 ();
 sg13g2_fill_1 FILLER_9_1615 ();
 sg13g2_fill_2 FILLER_9_1642 ();
 sg13g2_fill_2 FILLER_9_1707 ();
 sg13g2_fill_1 FILLER_9_1796 ();
 sg13g2_fill_1 FILLER_9_1823 ();
 sg13g2_fill_1 FILLER_9_1839 ();
 sg13g2_fill_1 FILLER_9_1844 ();
 sg13g2_fill_2 FILLER_9_1866 ();
 sg13g2_fill_2 FILLER_9_1894 ();
 sg13g2_fill_2 FILLER_9_1900 ();
 sg13g2_fill_1 FILLER_9_1902 ();
 sg13g2_fill_1 FILLER_9_1907 ();
 sg13g2_fill_2 FILLER_9_1921 ();
 sg13g2_fill_1 FILLER_9_1923 ();
 sg13g2_fill_2 FILLER_9_1943 ();
 sg13g2_fill_1 FILLER_9_1971 ();
 sg13g2_fill_1 FILLER_9_1984 ();
 sg13g2_decap_4 FILLER_9_2011 ();
 sg13g2_fill_2 FILLER_9_2100 ();
 sg13g2_fill_1 FILLER_9_2102 ();
 sg13g2_decap_8 FILLER_9_2132 ();
 sg13g2_fill_1 FILLER_9_2139 ();
 sg13g2_fill_2 FILLER_9_2240 ();
 sg13g2_fill_1 FILLER_9_2259 ();
 sg13g2_fill_1 FILLER_9_2270 ();
 sg13g2_fill_2 FILLER_9_2297 ();
 sg13g2_decap_4 FILLER_9_2309 ();
 sg13g2_fill_1 FILLER_9_2313 ();
 sg13g2_decap_8 FILLER_9_2318 ();
 sg13g2_fill_2 FILLER_9_2325 ();
 sg13g2_decap_8 FILLER_9_2348 ();
 sg13g2_decap_4 FILLER_9_2355 ();
 sg13g2_fill_1 FILLER_9_2369 ();
 sg13g2_fill_2 FILLER_9_2399 ();
 sg13g2_fill_1 FILLER_9_2401 ();
 sg13g2_fill_2 FILLER_9_2431 ();
 sg13g2_fill_1 FILLER_9_2460 ();
 sg13g2_fill_2 FILLER_9_2492 ();
 sg13g2_fill_2 FILLER_9_2498 ();
 sg13g2_fill_1 FILLER_9_2500 ();
 sg13g2_fill_2 FILLER_9_2532 ();
 sg13g2_fill_1 FILLER_9_2534 ();
 sg13g2_decap_8 FILLER_9_2549 ();
 sg13g2_decap_8 FILLER_9_2556 ();
 sg13g2_decap_8 FILLER_9_2563 ();
 sg13g2_decap_4 FILLER_9_2570 ();
 sg13g2_fill_2 FILLER_9_2574 ();
 sg13g2_fill_2 FILLER_9_2614 ();
 sg13g2_decap_8 FILLER_9_2647 ();
 sg13g2_decap_8 FILLER_9_2654 ();
 sg13g2_decap_8 FILLER_9_2661 ();
 sg13g2_fill_2 FILLER_9_2668 ();
 sg13g2_decap_4 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_33 ();
 sg13g2_fill_1 FILLER_10_40 ();
 sg13g2_fill_2 FILLER_10_44 ();
 sg13g2_fill_2 FILLER_10_50 ();
 sg13g2_fill_2 FILLER_10_78 ();
 sg13g2_fill_1 FILLER_10_80 ();
 sg13g2_decap_8 FILLER_10_113 ();
 sg13g2_fill_1 FILLER_10_120 ();
 sg13g2_decap_8 FILLER_10_125 ();
 sg13g2_decap_8 FILLER_10_132 ();
 sg13g2_fill_1 FILLER_10_139 ();
 sg13g2_decap_4 FILLER_10_170 ();
 sg13g2_fill_1 FILLER_10_174 ();
 sg13g2_decap_8 FILLER_10_179 ();
 sg13g2_decap_8 FILLER_10_186 ();
 sg13g2_decap_8 FILLER_10_193 ();
 sg13g2_fill_1 FILLER_10_200 ();
 sg13g2_fill_2 FILLER_10_218 ();
 sg13g2_fill_1 FILLER_10_220 ();
 sg13g2_decap_8 FILLER_10_226 ();
 sg13g2_fill_2 FILLER_10_255 ();
 sg13g2_fill_2 FILLER_10_265 ();
 sg13g2_fill_2 FILLER_10_278 ();
 sg13g2_fill_2 FILLER_10_288 ();
 sg13g2_fill_1 FILLER_10_290 ();
 sg13g2_decap_4 FILLER_10_297 ();
 sg13g2_fill_1 FILLER_10_309 ();
 sg13g2_fill_1 FILLER_10_316 ();
 sg13g2_decap_4 FILLER_10_330 ();
 sg13g2_fill_2 FILLER_10_338 ();
 sg13g2_fill_1 FILLER_10_340 ();
 sg13g2_fill_2 FILLER_10_346 ();
 sg13g2_fill_1 FILLER_10_348 ();
 sg13g2_fill_1 FILLER_10_380 ();
 sg13g2_fill_1 FILLER_10_386 ();
 sg13g2_decap_8 FILLER_10_417 ();
 sg13g2_fill_2 FILLER_10_424 ();
 sg13g2_fill_1 FILLER_10_426 ();
 sg13g2_fill_2 FILLER_10_458 ();
 sg13g2_decap_8 FILLER_10_496 ();
 sg13g2_fill_2 FILLER_10_522 ();
 sg13g2_fill_1 FILLER_10_547 ();
 sg13g2_fill_1 FILLER_10_552 ();
 sg13g2_fill_2 FILLER_10_557 ();
 sg13g2_decap_8 FILLER_10_642 ();
 sg13g2_decap_4 FILLER_10_649 ();
 sg13g2_fill_2 FILLER_10_695 ();
 sg13g2_decap_4 FILLER_10_701 ();
 sg13g2_fill_2 FILLER_10_724 ();
 sg13g2_decap_4 FILLER_10_731 ();
 sg13g2_fill_1 FILLER_10_744 ();
 sg13g2_decap_8 FILLER_10_775 ();
 sg13g2_fill_1 FILLER_10_782 ();
 sg13g2_fill_1 FILLER_10_840 ();
 sg13g2_fill_2 FILLER_10_918 ();
 sg13g2_decap_4 FILLER_10_924 ();
 sg13g2_fill_1 FILLER_10_928 ();
 sg13g2_fill_2 FILLER_10_939 ();
 sg13g2_fill_2 FILLER_10_945 ();
 sg13g2_decap_8 FILLER_10_959 ();
 sg13g2_decap_8 FILLER_10_966 ();
 sg13g2_decap_8 FILLER_10_973 ();
 sg13g2_decap_8 FILLER_10_980 ();
 sg13g2_decap_8 FILLER_10_987 ();
 sg13g2_decap_8 FILLER_10_994 ();
 sg13g2_decap_8 FILLER_10_1001 ();
 sg13g2_decap_4 FILLER_10_1008 ();
 sg13g2_decap_4 FILLER_10_1056 ();
 sg13g2_fill_1 FILLER_10_1064 ();
 sg13g2_decap_4 FILLER_10_1117 ();
 sg13g2_decap_8 FILLER_10_1166 ();
 sg13g2_decap_4 FILLER_10_1173 ();
 sg13g2_fill_2 FILLER_10_1241 ();
 sg13g2_fill_2 FILLER_10_1278 ();
 sg13g2_fill_1 FILLER_10_1280 ();
 sg13g2_decap_8 FILLER_10_1317 ();
 sg13g2_fill_2 FILLER_10_1324 ();
 sg13g2_fill_1 FILLER_10_1326 ();
 sg13g2_fill_2 FILLER_10_1336 ();
 sg13g2_decap_4 FILLER_10_1343 ();
 sg13g2_decap_8 FILLER_10_1433 ();
 sg13g2_decap_8 FILLER_10_1440 ();
 sg13g2_fill_2 FILLER_10_1447 ();
 sg13g2_fill_2 FILLER_10_1453 ();
 sg13g2_fill_1 FILLER_10_1455 ();
 sg13g2_decap_8 FILLER_10_1482 ();
 sg13g2_decap_4 FILLER_10_1489 ();
 sg13g2_fill_1 FILLER_10_1493 ();
 sg13g2_decap_4 FILLER_10_1506 ();
 sg13g2_fill_2 FILLER_10_1510 ();
 sg13g2_fill_1 FILLER_10_1600 ();
 sg13g2_decap_4 FILLER_10_1631 ();
 sg13g2_fill_2 FILLER_10_1639 ();
 sg13g2_decap_8 FILLER_10_1661 ();
 sg13g2_decap_4 FILLER_10_1668 ();
 sg13g2_decap_4 FILLER_10_1682 ();
 sg13g2_fill_1 FILLER_10_1686 ();
 sg13g2_fill_2 FILLER_10_1691 ();
 sg13g2_fill_1 FILLER_10_1693 ();
 sg13g2_fill_1 FILLER_10_1718 ();
 sg13g2_fill_1 FILLER_10_1723 ();
 sg13g2_fill_1 FILLER_10_1728 ();
 sg13g2_decap_4 FILLER_10_1798 ();
 sg13g2_fill_2 FILLER_10_1802 ();
 sg13g2_decap_4 FILLER_10_1818 ();
 sg13g2_fill_2 FILLER_10_1822 ();
 sg13g2_decap_4 FILLER_10_1829 ();
 sg13g2_fill_1 FILLER_10_1833 ();
 sg13g2_fill_2 FILLER_10_1838 ();
 sg13g2_fill_1 FILLER_10_1840 ();
 sg13g2_fill_1 FILLER_10_1845 ();
 sg13g2_fill_1 FILLER_10_1894 ();
 sg13g2_decap_8 FILLER_10_1899 ();
 sg13g2_decap_4 FILLER_10_1906 ();
 sg13g2_fill_2 FILLER_10_1914 ();
 sg13g2_fill_1 FILLER_10_1916 ();
 sg13g2_fill_2 FILLER_10_1931 ();
 sg13g2_fill_1 FILLER_10_1943 ();
 sg13g2_fill_1 FILLER_10_1954 ();
 sg13g2_fill_2 FILLER_10_1959 ();
 sg13g2_decap_8 FILLER_10_1965 ();
 sg13g2_fill_2 FILLER_10_1982 ();
 sg13g2_fill_2 FILLER_10_1994 ();
 sg13g2_decap_8 FILLER_10_2000 ();
 sg13g2_decap_8 FILLER_10_2007 ();
 sg13g2_decap_8 FILLER_10_2014 ();
 sg13g2_fill_2 FILLER_10_2021 ();
 sg13g2_fill_2 FILLER_10_2033 ();
 sg13g2_fill_2 FILLER_10_2045 ();
 sg13g2_decap_8 FILLER_10_2051 ();
 sg13g2_decap_8 FILLER_10_2058 ();
 sg13g2_decap_4 FILLER_10_2065 ();
 sg13g2_fill_1 FILLER_10_2069 ();
 sg13g2_decap_8 FILLER_10_2074 ();
 sg13g2_decap_4 FILLER_10_2081 ();
 sg13g2_fill_2 FILLER_10_2085 ();
 sg13g2_fill_2 FILLER_10_2097 ();
 sg13g2_fill_2 FILLER_10_2103 ();
 sg13g2_fill_1 FILLER_10_2105 ();
 sg13g2_fill_1 FILLER_10_2116 ();
 sg13g2_fill_1 FILLER_10_2138 ();
 sg13g2_fill_1 FILLER_10_2165 ();
 sg13g2_fill_1 FILLER_10_2187 ();
 sg13g2_decap_4 FILLER_10_2196 ();
 sg13g2_decap_8 FILLER_10_2247 ();
 sg13g2_fill_1 FILLER_10_2254 ();
 sg13g2_fill_1 FILLER_10_2281 ();
 sg13g2_fill_1 FILLER_10_2286 ();
 sg13g2_fill_2 FILLER_10_2291 ();
 sg13g2_fill_1 FILLER_10_2293 ();
 sg13g2_fill_2 FILLER_10_2320 ();
 sg13g2_decap_4 FILLER_10_2348 ();
 sg13g2_fill_1 FILLER_10_2352 ();
 sg13g2_decap_8 FILLER_10_2376 ();
 sg13g2_decap_8 FILLER_10_2383 ();
 sg13g2_decap_8 FILLER_10_2390 ();
 sg13g2_decap_8 FILLER_10_2397 ();
 sg13g2_fill_2 FILLER_10_2404 ();
 sg13g2_fill_2 FILLER_10_2445 ();
 sg13g2_fill_1 FILLER_10_2460 ();
 sg13g2_decap_8 FILLER_10_2487 ();
 sg13g2_decap_8 FILLER_10_2494 ();
 sg13g2_fill_1 FILLER_10_2501 ();
 sg13g2_fill_1 FILLER_10_2506 ();
 sg13g2_fill_1 FILLER_10_2517 ();
 sg13g2_fill_2 FILLER_10_2544 ();
 sg13g2_fill_1 FILLER_10_2546 ();
 sg13g2_fill_1 FILLER_10_2603 ();
 sg13g2_decap_4 FILLER_10_2614 ();
 sg13g2_fill_2 FILLER_10_2618 ();
 sg13g2_decap_8 FILLER_10_2640 ();
 sg13g2_decap_8 FILLER_10_2647 ();
 sg13g2_decap_8 FILLER_10_2654 ();
 sg13g2_decap_8 FILLER_10_2661 ();
 sg13g2_fill_2 FILLER_10_2668 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_18 ();
 sg13g2_decap_8 FILLER_11_25 ();
 sg13g2_fill_1 FILLER_11_32 ();
 sg13g2_fill_1 FILLER_11_38 ();
 sg13g2_fill_1 FILLER_11_49 ();
 sg13g2_fill_1 FILLER_11_55 ();
 sg13g2_fill_1 FILLER_11_65 ();
 sg13g2_fill_1 FILLER_11_70 ();
 sg13g2_fill_1 FILLER_11_101 ();
 sg13g2_fill_1 FILLER_11_128 ();
 sg13g2_fill_2 FILLER_11_133 ();
 sg13g2_fill_1 FILLER_11_161 ();
 sg13g2_fill_1 FILLER_11_167 ();
 sg13g2_fill_1 FILLER_11_177 ();
 sg13g2_decap_4 FILLER_11_182 ();
 sg13g2_fill_2 FILLER_11_186 ();
 sg13g2_decap_8 FILLER_11_193 ();
 sg13g2_decap_8 FILLER_11_200 ();
 sg13g2_fill_2 FILLER_11_207 ();
 sg13g2_fill_1 FILLER_11_209 ();
 sg13g2_decap_4 FILLER_11_214 ();
 sg13g2_fill_1 FILLER_11_218 ();
 sg13g2_decap_4 FILLER_11_228 ();
 sg13g2_fill_2 FILLER_11_236 ();
 sg13g2_decap_8 FILLER_11_268 ();
 sg13g2_decap_8 FILLER_11_275 ();
 sg13g2_fill_2 FILLER_11_310 ();
 sg13g2_fill_1 FILLER_11_312 ();
 sg13g2_fill_2 FILLER_11_321 ();
 sg13g2_decap_4 FILLER_11_349 ();
 sg13g2_decap_4 FILLER_11_390 ();
 sg13g2_fill_1 FILLER_11_394 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_463 ();
 sg13g2_fill_1 FILLER_11_468 ();
 sg13g2_decap_8 FILLER_11_477 ();
 sg13g2_fill_2 FILLER_11_484 ();
 sg13g2_fill_2 FILLER_11_490 ();
 sg13g2_decap_8 FILLER_11_504 ();
 sg13g2_decap_4 FILLER_11_511 ();
 sg13g2_fill_1 FILLER_11_515 ();
 sg13g2_fill_1 FILLER_11_525 ();
 sg13g2_decap_4 FILLER_11_535 ();
 sg13g2_decap_8 FILLER_11_558 ();
 sg13g2_fill_1 FILLER_11_565 ();
 sg13g2_decap_8 FILLER_11_570 ();
 sg13g2_fill_1 FILLER_11_592 ();
 sg13g2_fill_2 FILLER_11_607 ();
 sg13g2_decap_8 FILLER_11_613 ();
 sg13g2_decap_4 FILLER_11_620 ();
 sg13g2_fill_1 FILLER_11_624 ();
 sg13g2_fill_2 FILLER_11_633 ();
 sg13g2_fill_1 FILLER_11_635 ();
 sg13g2_fill_2 FILLER_11_641 ();
 sg13g2_fill_1 FILLER_11_643 ();
 sg13g2_fill_1 FILLER_11_678 ();
 sg13g2_decap_8 FILLER_11_683 ();
 sg13g2_fill_2 FILLER_11_690 ();
 sg13g2_decap_4 FILLER_11_696 ();
 sg13g2_decap_8 FILLER_11_770 ();
 sg13g2_decap_8 FILLER_11_777 ();
 sg13g2_decap_8 FILLER_11_784 ();
 sg13g2_fill_2 FILLER_11_791 ();
 sg13g2_decap_8 FILLER_11_797 ();
 sg13g2_fill_2 FILLER_11_804 ();
 sg13g2_fill_1 FILLER_11_806 ();
 sg13g2_decap_8 FILLER_11_817 ();
 sg13g2_decap_8 FILLER_11_824 ();
 sg13g2_decap_4 FILLER_11_831 ();
 sg13g2_fill_2 FILLER_11_835 ();
 sg13g2_fill_2 FILLER_11_873 ();
 sg13g2_decap_8 FILLER_11_926 ();
 sg13g2_fill_1 FILLER_11_933 ();
 sg13g2_fill_2 FILLER_11_1000 ();
 sg13g2_decap_8 FILLER_11_1014 ();
 sg13g2_decap_8 FILLER_11_1021 ();
 sg13g2_fill_2 FILLER_11_1033 ();
 sg13g2_fill_1 FILLER_11_1035 ();
 sg13g2_fill_2 FILLER_11_1040 ();
 sg13g2_decap_8 FILLER_11_1046 ();
 sg13g2_decap_8 FILLER_11_1053 ();
 sg13g2_fill_1 FILLER_11_1060 ();
 sg13g2_decap_8 FILLER_11_1124 ();
 sg13g2_fill_2 FILLER_11_1135 ();
 sg13g2_fill_1 FILLER_11_1137 ();
 sg13g2_fill_2 FILLER_11_1173 ();
 sg13g2_fill_2 FILLER_11_1199 ();
 sg13g2_fill_2 FILLER_11_1209 ();
 sg13g2_fill_1 FILLER_11_1216 ();
 sg13g2_fill_2 FILLER_11_1222 ();
 sg13g2_fill_1 FILLER_11_1224 ();
 sg13g2_fill_2 FILLER_11_1229 ();
 sg13g2_fill_1 FILLER_11_1231 ();
 sg13g2_decap_8 FILLER_11_1244 ();
 sg13g2_fill_2 FILLER_11_1251 ();
 sg13g2_fill_2 FILLER_11_1267 ();
 sg13g2_decap_4 FILLER_11_1306 ();
 sg13g2_fill_1 FILLER_11_1310 ();
 sg13g2_decap_8 FILLER_11_1316 ();
 sg13g2_fill_1 FILLER_11_1323 ();
 sg13g2_fill_2 FILLER_11_1328 ();
 sg13g2_decap_4 FILLER_11_1339 ();
 sg13g2_fill_1 FILLER_11_1343 ();
 sg13g2_fill_2 FILLER_11_1349 ();
 sg13g2_fill_2 FILLER_11_1359 ();
 sg13g2_fill_1 FILLER_11_1361 ();
 sg13g2_fill_2 FILLER_11_1370 ();
 sg13g2_fill_1 FILLER_11_1372 ();
 sg13g2_fill_2 FILLER_11_1403 ();
 sg13g2_fill_2 FILLER_11_1419 ();
 sg13g2_fill_1 FILLER_11_1421 ();
 sg13g2_decap_8 FILLER_11_1468 ();
 sg13g2_decap_8 FILLER_11_1475 ();
 sg13g2_decap_4 FILLER_11_1482 ();
 sg13g2_fill_1 FILLER_11_1486 ();
 sg13g2_decap_4 FILLER_11_1497 ();
 sg13g2_fill_1 FILLER_11_1511 ();
 sg13g2_decap_8 FILLER_11_1524 ();
 sg13g2_fill_1 FILLER_11_1531 ();
 sg13g2_fill_2 FILLER_11_1558 ();
 sg13g2_fill_1 FILLER_11_1573 ();
 sg13g2_fill_2 FILLER_11_1584 ();
 sg13g2_fill_2 FILLER_11_1591 ();
 sg13g2_decap_8 FILLER_11_1633 ();
 sg13g2_decap_8 FILLER_11_1640 ();
 sg13g2_decap_8 FILLER_11_1647 ();
 sg13g2_decap_8 FILLER_11_1654 ();
 sg13g2_fill_1 FILLER_11_1661 ();
 sg13g2_fill_1 FILLER_11_1672 ();
 sg13g2_decap_8 FILLER_11_1710 ();
 sg13g2_fill_1 FILLER_11_1717 ();
 sg13g2_decap_8 FILLER_11_1722 ();
 sg13g2_fill_1 FILLER_11_1744 ();
 sg13g2_fill_2 FILLER_11_1754 ();
 sg13g2_fill_2 FILLER_11_1803 ();
 sg13g2_fill_1 FILLER_11_1805 ();
 sg13g2_fill_1 FILLER_11_1837 ();
 sg13g2_fill_1 FILLER_11_1843 ();
 sg13g2_fill_2 FILLER_11_1848 ();
 sg13g2_fill_1 FILLER_11_1850 ();
 sg13g2_fill_2 FILLER_11_1856 ();
 sg13g2_fill_1 FILLER_11_1858 ();
 sg13g2_fill_2 FILLER_11_1869 ();
 sg13g2_fill_2 FILLER_11_1875 ();
 sg13g2_decap_8 FILLER_11_1914 ();
 sg13g2_fill_1 FILLER_11_1921 ();
 sg13g2_decap_8 FILLER_11_1927 ();
 sg13g2_decap_8 FILLER_11_1934 ();
 sg13g2_decap_8 FILLER_11_1941 ();
 sg13g2_decap_4 FILLER_11_1948 ();
 sg13g2_decap_8 FILLER_11_1977 ();
 sg13g2_decap_4 FILLER_11_2010 ();
 sg13g2_fill_2 FILLER_11_2014 ();
 sg13g2_fill_2 FILLER_11_2021 ();
 sg13g2_fill_1 FILLER_11_2023 ();
 sg13g2_decap_8 FILLER_11_2034 ();
 sg13g2_fill_1 FILLER_11_2041 ();
 sg13g2_fill_2 FILLER_11_2068 ();
 sg13g2_decap_4 FILLER_11_2096 ();
 sg13g2_decap_4 FILLER_11_2110 ();
 sg13g2_decap_8 FILLER_11_2140 ();
 sg13g2_fill_2 FILLER_11_2147 ();
 sg13g2_fill_1 FILLER_11_2149 ();
 sg13g2_fill_2 FILLER_11_2160 ();
 sg13g2_fill_2 FILLER_11_2172 ();
 sg13g2_fill_2 FILLER_11_2200 ();
 sg13g2_decap_4 FILLER_11_2242 ();
 sg13g2_decap_8 FILLER_11_2256 ();
 sg13g2_fill_1 FILLER_11_2263 ();
 sg13g2_decap_8 FILLER_11_2268 ();
 sg13g2_fill_1 FILLER_11_2275 ();
 sg13g2_decap_4 FILLER_11_2286 ();
 sg13g2_fill_1 FILLER_11_2290 ();
 sg13g2_fill_1 FILLER_11_2305 ();
 sg13g2_fill_2 FILLER_11_2353 ();
 sg13g2_fill_1 FILLER_11_2355 ();
 sg13g2_decap_4 FILLER_11_2395 ();
 sg13g2_decap_8 FILLER_11_2404 ();
 sg13g2_fill_1 FILLER_11_2411 ();
 sg13g2_fill_1 FILLER_11_2448 ();
 sg13g2_decap_8 FILLER_11_2485 ();
 sg13g2_decap_8 FILLER_11_2492 ();
 sg13g2_decap_4 FILLER_11_2499 ();
 sg13g2_fill_1 FILLER_11_2529 ();
 sg13g2_fill_1 FILLER_11_2534 ();
 sg13g2_decap_8 FILLER_11_2594 ();
 sg13g2_fill_1 FILLER_11_2601 ();
 sg13g2_fill_1 FILLER_11_2628 ();
 sg13g2_decap_4 FILLER_11_2665 ();
 sg13g2_fill_1 FILLER_11_2669 ();
 sg13g2_fill_1 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_4 FILLER_12_49 ();
 sg13g2_fill_1 FILLER_12_53 ();
 sg13g2_decap_8 FILLER_12_58 ();
 sg13g2_decap_8 FILLER_12_65 ();
 sg13g2_decap_8 FILLER_12_72 ();
 sg13g2_fill_1 FILLER_12_87 ();
 sg13g2_fill_2 FILLER_12_92 ();
 sg13g2_fill_2 FILLER_12_98 ();
 sg13g2_fill_2 FILLER_12_104 ();
 sg13g2_fill_1 FILLER_12_106 ();
 sg13g2_decap_8 FILLER_12_153 ();
 sg13g2_fill_2 FILLER_12_160 ();
 sg13g2_decap_8 FILLER_12_192 ();
 sg13g2_decap_4 FILLER_12_199 ();
 sg13g2_fill_1 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_243 ();
 sg13g2_decap_4 FILLER_12_250 ();
 sg13g2_fill_1 FILLER_12_254 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_fill_2 FILLER_12_280 ();
 sg13g2_fill_1 FILLER_12_282 ();
 sg13g2_fill_1 FILLER_12_287 ();
 sg13g2_fill_2 FILLER_12_297 ();
 sg13g2_fill_1 FILLER_12_299 ();
 sg13g2_fill_1 FILLER_12_308 ();
 sg13g2_fill_1 FILLER_12_315 ();
 sg13g2_fill_2 FILLER_12_320 ();
 sg13g2_decap_8 FILLER_12_335 ();
 sg13g2_decap_8 FILLER_12_342 ();
 sg13g2_decap_8 FILLER_12_349 ();
 sg13g2_decap_4 FILLER_12_356 ();
 sg13g2_fill_2 FILLER_12_360 ();
 sg13g2_decap_8 FILLER_12_407 ();
 sg13g2_decap_4 FILLER_12_414 ();
 sg13g2_decap_8 FILLER_12_422 ();
 sg13g2_decap_4 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_12_437 ();
 sg13g2_decap_8 FILLER_12_444 ();
 sg13g2_decap_8 FILLER_12_451 ();
 sg13g2_fill_1 FILLER_12_458 ();
 sg13g2_decap_4 FILLER_12_468 ();
 sg13g2_fill_2 FILLER_12_472 ();
 sg13g2_decap_8 FILLER_12_516 ();
 sg13g2_decap_4 FILLER_12_523 ();
 sg13g2_fill_1 FILLER_12_576 ();
 sg13g2_fill_1 FILLER_12_587 ();
 sg13g2_decap_8 FILLER_12_615 ();
 sg13g2_decap_8 FILLER_12_622 ();
 sg13g2_decap_8 FILLER_12_629 ();
 sg13g2_decap_8 FILLER_12_636 ();
 sg13g2_decap_8 FILLER_12_643 ();
 sg13g2_decap_4 FILLER_12_663 ();
 sg13g2_decap_8 FILLER_12_677 ();
 sg13g2_decap_8 FILLER_12_684 ();
 sg13g2_fill_2 FILLER_12_691 ();
 sg13g2_fill_1 FILLER_12_693 ();
 sg13g2_decap_8 FILLER_12_698 ();
 sg13g2_decap_8 FILLER_12_705 ();
 sg13g2_fill_1 FILLER_12_712 ();
 sg13g2_decap_8 FILLER_12_717 ();
 sg13g2_fill_1 FILLER_12_724 ();
 sg13g2_fill_2 FILLER_12_730 ();
 sg13g2_fill_2 FILLER_12_737 ();
 sg13g2_fill_2 FILLER_12_753 ();
 sg13g2_decap_8 FILLER_12_759 ();
 sg13g2_fill_1 FILLER_12_766 ();
 sg13g2_decap_8 FILLER_12_776 ();
 sg13g2_decap_8 FILLER_12_783 ();
 sg13g2_fill_2 FILLER_12_790 ();
 sg13g2_fill_1 FILLER_12_792 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_4 FILLER_12_840 ();
 sg13g2_fill_1 FILLER_12_844 ();
 sg13g2_decap_4 FILLER_12_872 ();
 sg13g2_decap_4 FILLER_12_880 ();
 sg13g2_fill_1 FILLER_12_884 ();
 sg13g2_decap_8 FILLER_12_905 ();
 sg13g2_decap_8 FILLER_12_912 ();
 sg13g2_decap_8 FILLER_12_919 ();
 sg13g2_fill_2 FILLER_12_926 ();
 sg13g2_fill_1 FILLER_12_928 ();
 sg13g2_fill_2 FILLER_12_959 ();
 sg13g2_fill_1 FILLER_12_961 ();
 sg13g2_fill_2 FILLER_12_1011 ();
 sg13g2_fill_1 FILLER_12_1032 ();
 sg13g2_decap_4 FILLER_12_1059 ();
 sg13g2_fill_2 FILLER_12_1114 ();
 sg13g2_fill_1 FILLER_12_1116 ();
 sg13g2_fill_2 FILLER_12_1121 ();
 sg13g2_fill_1 FILLER_12_1123 ();
 sg13g2_fill_2 FILLER_12_1150 ();
 sg13g2_fill_1 FILLER_12_1152 ();
 sg13g2_fill_2 FILLER_12_1230 ();
 sg13g2_fill_2 FILLER_12_1265 ();
 sg13g2_fill_1 FILLER_12_1267 ();
 sg13g2_decap_4 FILLER_12_1282 ();
 sg13g2_fill_2 FILLER_12_1286 ();
 sg13g2_decap_8 FILLER_12_1296 ();
 sg13g2_decap_8 FILLER_12_1303 ();
 sg13g2_decap_4 FILLER_12_1310 ();
 sg13g2_fill_1 FILLER_12_1314 ();
 sg13g2_fill_2 FILLER_12_1358 ();
 sg13g2_fill_1 FILLER_12_1360 ();
 sg13g2_decap_8 FILLER_12_1365 ();
 sg13g2_decap_8 FILLER_12_1372 ();
 sg13g2_decap_4 FILLER_12_1379 ();
 sg13g2_decap_4 FILLER_12_1419 ();
 sg13g2_fill_1 FILLER_12_1423 ();
 sg13g2_fill_1 FILLER_12_1437 ();
 sg13g2_decap_8 FILLER_12_1442 ();
 sg13g2_fill_2 FILLER_12_1449 ();
 sg13g2_fill_1 FILLER_12_1451 ();
 sg13g2_fill_2 FILLER_12_1486 ();
 sg13g2_fill_1 FILLER_12_1488 ();
 sg13g2_fill_2 FILLER_12_1519 ();
 sg13g2_fill_1 FILLER_12_1521 ();
 sg13g2_fill_2 FILLER_12_1532 ();
 sg13g2_fill_2 FILLER_12_1544 ();
 sg13g2_fill_1 FILLER_12_1567 ();
 sg13g2_decap_4 FILLER_12_1598 ();
 sg13g2_fill_1 FILLER_12_1602 ();
 sg13g2_decap_8 FILLER_12_1629 ();
 sg13g2_decap_8 FILLER_12_1636 ();
 sg13g2_fill_2 FILLER_12_1643 ();
 sg13g2_fill_1 FILLER_12_1645 ();
 sg13g2_decap_4 FILLER_12_1698 ();
 sg13g2_fill_1 FILLER_12_1792 ();
 sg13g2_decap_4 FILLER_12_1838 ();
 sg13g2_fill_2 FILLER_12_1842 ();
 sg13g2_fill_2 FILLER_12_1864 ();
 sg13g2_fill_1 FILLER_12_1866 ();
 sg13g2_fill_1 FILLER_12_1887 ();
 sg13g2_decap_4 FILLER_12_1929 ();
 sg13g2_fill_2 FILLER_12_1933 ();
 sg13g2_fill_2 FILLER_12_1973 ();
 sg13g2_fill_1 FILLER_12_2015 ();
 sg13g2_fill_1 FILLER_12_2020 ();
 sg13g2_fill_1 FILLER_12_2047 ();
 sg13g2_fill_1 FILLER_12_2069 ();
 sg13g2_fill_1 FILLER_12_2074 ();
 sg13g2_decap_8 FILLER_12_2126 ();
 sg13g2_decap_8 FILLER_12_2133 ();
 sg13g2_decap_8 FILLER_12_2140 ();
 sg13g2_fill_2 FILLER_12_2147 ();
 sg13g2_fill_1 FILLER_12_2149 ();
 sg13g2_fill_1 FILLER_12_2163 ();
 sg13g2_fill_2 FILLER_12_2168 ();
 sg13g2_fill_1 FILLER_12_2170 ();
 sg13g2_fill_2 FILLER_12_2181 ();
 sg13g2_fill_1 FILLER_12_2183 ();
 sg13g2_decap_4 FILLER_12_2188 ();
 sg13g2_fill_2 FILLER_12_2192 ();
 sg13g2_decap_4 FILLER_12_2202 ();
 sg13g2_fill_2 FILLER_12_2206 ();
 sg13g2_fill_2 FILLER_12_2222 ();
 sg13g2_decap_8 FILLER_12_2247 ();
 sg13g2_decap_8 FILLER_12_2254 ();
 sg13g2_decap_8 FILLER_12_2261 ();
 sg13g2_fill_2 FILLER_12_2268 ();
 sg13g2_decap_8 FILLER_12_2291 ();
 sg13g2_decap_8 FILLER_12_2298 ();
 sg13g2_fill_2 FILLER_12_2305 ();
 sg13g2_fill_2 FILLER_12_2327 ();
 sg13g2_decap_8 FILLER_12_2333 ();
 sg13g2_decap_4 FILLER_12_2340 ();
 sg13g2_fill_2 FILLER_12_2344 ();
 sg13g2_decap_4 FILLER_12_2401 ();
 sg13g2_fill_2 FILLER_12_2405 ();
 sg13g2_fill_1 FILLER_12_2454 ();
 sg13g2_fill_1 FILLER_12_2465 ();
 sg13g2_decap_4 FILLER_12_2505 ();
 sg13g2_decap_4 FILLER_12_2513 ();
 sg13g2_fill_2 FILLER_12_2517 ();
 sg13g2_fill_2 FILLER_12_2529 ();
 sg13g2_fill_1 FILLER_12_2531 ();
 sg13g2_decap_8 FILLER_12_2537 ();
 sg13g2_fill_2 FILLER_12_2544 ();
 sg13g2_decap_4 FILLER_12_2576 ();
 sg13g2_fill_2 FILLER_12_2614 ();
 sg13g2_decap_8 FILLER_12_2652 ();
 sg13g2_decap_8 FILLER_12_2659 ();
 sg13g2_decap_4 FILLER_12_2666 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_37 ();
 sg13g2_decap_8 FILLER_13_44 ();
 sg13g2_fill_2 FILLER_13_51 ();
 sg13g2_fill_1 FILLER_13_92 ();
 sg13g2_fill_2 FILLER_13_123 ();
 sg13g2_decap_8 FILLER_13_129 ();
 sg13g2_fill_2 FILLER_13_140 ();
 sg13g2_fill_1 FILLER_13_142 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_fill_1 FILLER_13_166 ();
 sg13g2_fill_1 FILLER_13_173 ();
 sg13g2_fill_2 FILLER_13_193 ();
 sg13g2_decap_4 FILLER_13_246 ();
 sg13g2_fill_1 FILLER_13_250 ();
 sg13g2_fill_1 FILLER_13_255 ();
 sg13g2_fill_1 FILLER_13_282 ();
 sg13g2_fill_1 FILLER_13_309 ();
 sg13g2_fill_1 FILLER_13_341 ();
 sg13g2_fill_1 FILLER_13_347 ();
 sg13g2_fill_1 FILLER_13_352 ();
 sg13g2_fill_1 FILLER_13_357 ();
 sg13g2_decap_4 FILLER_13_380 ();
 sg13g2_decap_4 FILLER_13_388 ();
 sg13g2_fill_1 FILLER_13_392 ();
 sg13g2_fill_2 FILLER_13_437 ();
 sg13g2_fill_2 FILLER_13_449 ();
 sg13g2_fill_1 FILLER_13_451 ();
 sg13g2_fill_2 FILLER_13_456 ();
 sg13g2_fill_1 FILLER_13_458 ();
 sg13g2_decap_8 FILLER_13_463 ();
 sg13g2_fill_1 FILLER_13_470 ();
 sg13g2_decap_4 FILLER_13_485 ();
 sg13g2_decap_8 FILLER_13_523 ();
 sg13g2_fill_2 FILLER_13_530 ();
 sg13g2_fill_1 FILLER_13_532 ();
 sg13g2_decap_8 FILLER_13_636 ();
 sg13g2_fill_2 FILLER_13_643 ();
 sg13g2_fill_2 FILLER_13_649 ();
 sg13g2_fill_2 FILLER_13_682 ();
 sg13g2_fill_1 FILLER_13_684 ();
 sg13g2_decap_8 FILLER_13_711 ();
 sg13g2_decap_8 FILLER_13_718 ();
 sg13g2_decap_4 FILLER_13_725 ();
 sg13g2_fill_1 FILLER_13_729 ();
 sg13g2_fill_2 FILLER_13_752 ();
 sg13g2_fill_1 FILLER_13_754 ();
 sg13g2_decap_8 FILLER_13_786 ();
 sg13g2_decap_4 FILLER_13_793 ();
 sg13g2_fill_2 FILLER_13_797 ();
 sg13g2_fill_2 FILLER_13_846 ();
 sg13g2_decap_4 FILLER_13_862 ();
 sg13g2_fill_2 FILLER_13_866 ();
 sg13g2_decap_8 FILLER_13_878 ();
 sg13g2_decap_8 FILLER_13_921 ();
 sg13g2_decap_8 FILLER_13_928 ();
 sg13g2_fill_1 FILLER_13_935 ();
 sg13g2_decap_8 FILLER_13_946 ();
 sg13g2_fill_2 FILLER_13_953 ();
 sg13g2_fill_1 FILLER_13_955 ();
 sg13g2_fill_2 FILLER_13_998 ();
 sg13g2_fill_1 FILLER_13_1000 ();
 sg13g2_fill_1 FILLER_13_1069 ();
 sg13g2_decap_8 FILLER_13_1136 ();
 sg13g2_decap_4 FILLER_13_1143 ();
 sg13g2_fill_1 FILLER_13_1204 ();
 sg13g2_fill_1 FILLER_13_1273 ();
 sg13g2_fill_1 FILLER_13_1310 ();
 sg13g2_fill_1 FILLER_13_1329 ();
 sg13g2_decap_8 FILLER_13_1356 ();
 sg13g2_decap_4 FILLER_13_1363 ();
 sg13g2_decap_4 FILLER_13_1407 ();
 sg13g2_decap_8 FILLER_13_1467 ();
 sg13g2_fill_2 FILLER_13_1478 ();
 sg13g2_decap_4 FILLER_13_1524 ();
 sg13g2_fill_2 FILLER_13_1528 ();
 sg13g2_fill_2 FILLER_13_1552 ();
 sg13g2_fill_1 FILLER_13_1571 ();
 sg13g2_fill_1 FILLER_13_1576 ();
 sg13g2_fill_1 FILLER_13_1617 ();
 sg13g2_fill_1 FILLER_13_1656 ();
 sg13g2_fill_2 FILLER_13_1667 ();
 sg13g2_fill_1 FILLER_13_1673 ();
 sg13g2_fill_2 FILLER_13_1700 ();
 sg13g2_fill_1 FILLER_13_1702 ();
 sg13g2_fill_2 FILLER_13_1739 ();
 sg13g2_fill_2 FILLER_13_1745 ();
 sg13g2_fill_1 FILLER_13_1747 ();
 sg13g2_fill_1 FILLER_13_1813 ();
 sg13g2_fill_1 FILLER_13_1818 ();
 sg13g2_fill_1 FILLER_13_1840 ();
 sg13g2_decap_8 FILLER_13_1845 ();
 sg13g2_decap_4 FILLER_13_1852 ();
 sg13g2_fill_2 FILLER_13_1877 ();
 sg13g2_decap_4 FILLER_13_1918 ();
 sg13g2_fill_1 FILLER_13_1927 ();
 sg13g2_decap_4 FILLER_13_2001 ();
 sg13g2_fill_2 FILLER_13_2005 ();
 sg13g2_fill_2 FILLER_13_2051 ();
 sg13g2_decap_4 FILLER_13_2057 ();
 sg13g2_fill_1 FILLER_13_2094 ();
 sg13g2_decap_4 FILLER_13_2129 ();
 sg13g2_fill_2 FILLER_13_2141 ();
 sg13g2_fill_1 FILLER_13_2147 ();
 sg13g2_fill_1 FILLER_13_2162 ();
 sg13g2_fill_1 FILLER_13_2183 ();
 sg13g2_decap_8 FILLER_13_2188 ();
 sg13g2_decap_8 FILLER_13_2195 ();
 sg13g2_decap_8 FILLER_13_2212 ();
 sg13g2_decap_8 FILLER_13_2259 ();
 sg13g2_decap_4 FILLER_13_2266 ();
 sg13g2_fill_1 FILLER_13_2270 ();
 sg13g2_decap_4 FILLER_13_2275 ();
 sg13g2_fill_1 FILLER_13_2279 ();
 sg13g2_decap_8 FILLER_13_2301 ();
 sg13g2_decap_4 FILLER_13_2308 ();
 sg13g2_fill_1 FILLER_13_2312 ();
 sg13g2_decap_4 FILLER_13_2317 ();
 sg13g2_fill_2 FILLER_13_2321 ();
 sg13g2_fill_1 FILLER_13_2337 ();
 sg13g2_decap_4 FILLER_13_2402 ();
 sg13g2_decap_4 FILLER_13_2517 ();
 sg13g2_decap_8 FILLER_13_2531 ();
 sg13g2_decap_8 FILLER_13_2538 ();
 sg13g2_decap_8 FILLER_13_2545 ();
 sg13g2_fill_1 FILLER_13_2552 ();
 sg13g2_fill_2 FILLER_13_2557 ();
 sg13g2_fill_1 FILLER_13_2569 ();
 sg13g2_decap_8 FILLER_13_2591 ();
 sg13g2_decap_8 FILLER_13_2598 ();
 sg13g2_decap_8 FILLER_13_2605 ();
 sg13g2_decap_8 FILLER_13_2612 ();
 sg13g2_decap_4 FILLER_13_2666 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_7 ();
 sg13g2_fill_1 FILLER_14_52 ();
 sg13g2_fill_1 FILLER_14_102 ();
 sg13g2_decap_8 FILLER_14_120 ();
 sg13g2_decap_4 FILLER_14_127 ();
 sg13g2_fill_2 FILLER_14_131 ();
 sg13g2_decap_8 FILLER_14_137 ();
 sg13g2_fill_2 FILLER_14_144 ();
 sg13g2_fill_1 FILLER_14_146 ();
 sg13g2_fill_2 FILLER_14_173 ();
 sg13g2_fill_1 FILLER_14_175 ();
 sg13g2_fill_2 FILLER_14_186 ();
 sg13g2_fill_1 FILLER_14_188 ();
 sg13g2_fill_2 FILLER_14_220 ();
 sg13g2_decap_4 FILLER_14_230 ();
 sg13g2_fill_1 FILLER_14_234 ();
 sg13g2_fill_1 FILLER_14_241 ();
 sg13g2_fill_2 FILLER_14_278 ();
 sg13g2_fill_2 FILLER_14_297 ();
 sg13g2_fill_1 FILLER_14_321 ();
 sg13g2_fill_2 FILLER_14_329 ();
 sg13g2_fill_1 FILLER_14_339 ();
 sg13g2_fill_2 FILLER_14_396 ();
 sg13g2_decap_8 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_14_415 ();
 sg13g2_fill_2 FILLER_14_453 ();
 sg13g2_fill_1 FILLER_14_455 ();
 sg13g2_fill_1 FILLER_14_460 ();
 sg13g2_fill_1 FILLER_14_466 ();
 sg13g2_fill_2 FILLER_14_493 ();
 sg13g2_fill_1 FILLER_14_505 ();
 sg13g2_fill_2 FILLER_14_510 ();
 sg13g2_fill_1 FILLER_14_538 ();
 sg13g2_fill_2 FILLER_14_565 ();
 sg13g2_fill_2 FILLER_14_652 ();
 sg13g2_decap_8 FILLER_14_690 ();
 sg13g2_fill_1 FILLER_14_729 ();
 sg13g2_fill_2 FILLER_14_843 ();
 sg13g2_decap_4 FILLER_14_849 ();
 sg13g2_fill_2 FILLER_14_853 ();
 sg13g2_fill_1 FILLER_14_881 ();
 sg13g2_fill_2 FILLER_14_887 ();
 sg13g2_decap_4 FILLER_14_922 ();
 sg13g2_fill_2 FILLER_14_926 ();
 sg13g2_decap_4 FILLER_14_989 ();
 sg13g2_fill_1 FILLER_14_993 ();
 sg13g2_fill_2 FILLER_14_1030 ();
 sg13g2_fill_2 FILLER_14_1041 ();
 sg13g2_fill_2 FILLER_14_1079 ();
 sg13g2_decap_4 FILLER_14_1142 ();
 sg13g2_fill_2 FILLER_14_1150 ();
 sg13g2_fill_2 FILLER_14_1178 ();
 sg13g2_decap_4 FILLER_14_1184 ();
 sg13g2_decap_4 FILLER_14_1196 ();
 sg13g2_fill_2 FILLER_14_1205 ();
 sg13g2_decap_8 FILLER_14_1237 ();
 sg13g2_decap_4 FILLER_14_1244 ();
 sg13g2_fill_2 FILLER_14_1278 ();
 sg13g2_fill_1 FILLER_14_1280 ();
 sg13g2_decap_4 FILLER_14_1342 ();
 sg13g2_decap_8 FILLER_14_1389 ();
 sg13g2_fill_2 FILLER_14_1396 ();
 sg13g2_fill_1 FILLER_14_1398 ();
 sg13g2_decap_4 FILLER_14_1403 ();
 sg13g2_fill_1 FILLER_14_1407 ();
 sg13g2_decap_8 FILLER_14_1412 ();
 sg13g2_fill_2 FILLER_14_1419 ();
 sg13g2_fill_1 FILLER_14_1421 ();
 sg13g2_decap_8 FILLER_14_1435 ();
 sg13g2_decap_4 FILLER_14_1442 ();
 sg13g2_fill_1 FILLER_14_1446 ();
 sg13g2_fill_2 FILLER_14_1461 ();
 sg13g2_fill_1 FILLER_14_1473 ();
 sg13g2_fill_1 FILLER_14_1484 ();
 sg13g2_fill_2 FILLER_14_1511 ();
 sg13g2_fill_2 FILLER_14_1539 ();
 sg13g2_fill_1 FILLER_14_1545 ();
 sg13g2_fill_1 FILLER_14_1553 ();
 sg13g2_fill_1 FILLER_14_1559 ();
 sg13g2_fill_1 FILLER_14_1579 ();
 sg13g2_fill_2 FILLER_14_1638 ();
 sg13g2_decap_8 FILLER_14_1644 ();
 sg13g2_decap_4 FILLER_14_1651 ();
 sg13g2_fill_1 FILLER_14_1655 ();
 sg13g2_fill_2 FILLER_14_1660 ();
 sg13g2_fill_1 FILLER_14_1662 ();
 sg13g2_decap_4 FILLER_14_1673 ();
 sg13g2_fill_2 FILLER_14_1677 ();
 sg13g2_decap_8 FILLER_14_1689 ();
 sg13g2_decap_4 FILLER_14_1696 ();
 sg13g2_fill_1 FILLER_14_1700 ();
 sg13g2_fill_2 FILLER_14_1728 ();
 sg13g2_fill_1 FILLER_14_1730 ();
 sg13g2_fill_2 FILLER_14_1745 ();
 sg13g2_decap_8 FILLER_14_1760 ();
 sg13g2_fill_2 FILLER_14_1777 ();
 sg13g2_fill_1 FILLER_14_1779 ();
 sg13g2_fill_2 FILLER_14_1798 ();
 sg13g2_fill_1 FILLER_14_1800 ();
 sg13g2_fill_1 FILLER_14_1847 ();
 sg13g2_fill_2 FILLER_14_1854 ();
 sg13g2_fill_2 FILLER_14_1868 ();
 sg13g2_fill_1 FILLER_14_1876 ();
 sg13g2_fill_2 FILLER_14_1882 ();
 sg13g2_fill_1 FILLER_14_1884 ();
 sg13g2_fill_2 FILLER_14_1906 ();
 sg13g2_fill_1 FILLER_14_1908 ();
 sg13g2_decap_8 FILLER_14_1913 ();
 sg13g2_fill_2 FILLER_14_1920 ();
 sg13g2_fill_1 FILLER_14_1922 ();
 sg13g2_fill_2 FILLER_14_1951 ();
 sg13g2_fill_1 FILLER_14_1963 ();
 sg13g2_fill_2 FILLER_14_1968 ();
 sg13g2_fill_1 FILLER_14_1970 ();
 sg13g2_decap_8 FILLER_14_1975 ();
 sg13g2_fill_2 FILLER_14_1982 ();
 sg13g2_fill_1 FILLER_14_1984 ();
 sg13g2_decap_4 FILLER_14_2007 ();
 sg13g2_fill_2 FILLER_14_2011 ();
 sg13g2_decap_4 FILLER_14_2049 ();
 sg13g2_fill_1 FILLER_14_2053 ();
 sg13g2_decap_8 FILLER_14_2064 ();
 sg13g2_decap_8 FILLER_14_2071 ();
 sg13g2_fill_1 FILLER_14_2078 ();
 sg13g2_decap_8 FILLER_14_2092 ();
 sg13g2_decap_4 FILLER_14_2099 ();
 sg13g2_fill_1 FILLER_14_2103 ();
 sg13g2_fill_1 FILLER_14_2114 ();
 sg13g2_fill_1 FILLER_14_2141 ();
 sg13g2_fill_2 FILLER_14_2176 ();
 sg13g2_fill_2 FILLER_14_2204 ();
 sg13g2_fill_2 FILLER_14_2232 ();
 sg13g2_decap_4 FILLER_14_2260 ();
 sg13g2_fill_1 FILLER_14_2264 ();
 sg13g2_fill_2 FILLER_14_2288 ();
 sg13g2_decap_4 FILLER_14_2316 ();
 sg13g2_decap_8 FILLER_14_2346 ();
 sg13g2_decap_4 FILLER_14_2353 ();
 sg13g2_decap_8 FILLER_14_2393 ();
 sg13g2_fill_1 FILLER_14_2461 ();
 sg13g2_fill_2 FILLER_14_2495 ();
 sg13g2_fill_1 FILLER_14_2497 ();
 sg13g2_decap_8 FILLER_14_2502 ();
 sg13g2_decap_4 FILLER_14_2509 ();
 sg13g2_decap_4 FILLER_14_2539 ();
 sg13g2_fill_1 FILLER_14_2543 ();
 sg13g2_decap_8 FILLER_14_2548 ();
 sg13g2_decap_4 FILLER_14_2555 ();
 sg13g2_decap_8 FILLER_14_2580 ();
 sg13g2_fill_1 FILLER_14_2587 ();
 sg13g2_decap_8 FILLER_14_2604 ();
 sg13g2_decap_8 FILLER_14_2611 ();
 sg13g2_decap_8 FILLER_14_2618 ();
 sg13g2_decap_4 FILLER_14_2625 ();
 sg13g2_decap_4 FILLER_14_2643 ();
 sg13g2_fill_2 FILLER_14_2651 ();
 sg13g2_fill_1 FILLER_14_2653 ();
 sg13g2_decap_8 FILLER_14_2658 ();
 sg13g2_decap_4 FILLER_14_2665 ();
 sg13g2_fill_1 FILLER_14_2669 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_78 ();
 sg13g2_fill_2 FILLER_15_107 ();
 sg13g2_decap_8 FILLER_15_117 ();
 sg13g2_decap_4 FILLER_15_124 ();
 sg13g2_fill_2 FILLER_15_132 ();
 sg13g2_fill_1 FILLER_15_163 ();
 sg13g2_fill_2 FILLER_15_187 ();
 sg13g2_fill_1 FILLER_15_189 ();
 sg13g2_fill_2 FILLER_15_216 ();
 sg13g2_fill_1 FILLER_15_218 ();
 sg13g2_decap_4 FILLER_15_223 ();
 sg13g2_decap_8 FILLER_15_232 ();
 sg13g2_fill_1 FILLER_15_239 ();
 sg13g2_fill_1 FILLER_15_244 ();
 sg13g2_decap_4 FILLER_15_275 ();
 sg13g2_fill_2 FILLER_15_279 ();
 sg13g2_decap_4 FILLER_15_286 ();
 sg13g2_fill_2 FILLER_15_290 ();
 sg13g2_fill_1 FILLER_15_298 ();
 sg13g2_fill_1 FILLER_15_310 ();
 sg13g2_decap_4 FILLER_15_332 ();
 sg13g2_fill_2 FILLER_15_336 ();
 sg13g2_fill_1 FILLER_15_351 ();
 sg13g2_decap_4 FILLER_15_364 ();
 sg13g2_decap_4 FILLER_15_382 ();
 sg13g2_decap_8 FILLER_15_391 ();
 sg13g2_fill_1 FILLER_15_398 ();
 sg13g2_fill_2 FILLER_15_412 ();
 sg13g2_fill_2 FILLER_15_440 ();
 sg13g2_fill_1 FILLER_15_452 ();
 sg13g2_fill_2 FILLER_15_479 ();
 sg13g2_fill_2 FILLER_15_485 ();
 sg13g2_fill_2 FILLER_15_492 ();
 sg13g2_decap_4 FILLER_15_504 ();
 sg13g2_fill_2 FILLER_15_508 ();
 sg13g2_decap_4 FILLER_15_515 ();
 sg13g2_fill_1 FILLER_15_519 ();
 sg13g2_decap_8 FILLER_15_524 ();
 sg13g2_decap_4 FILLER_15_531 ();
 sg13g2_fill_2 FILLER_15_561 ();
 sg13g2_fill_2 FILLER_15_573 ();
 sg13g2_fill_1 FILLER_15_578 ();
 sg13g2_fill_2 FILLER_15_619 ();
 sg13g2_fill_1 FILLER_15_649 ();
 sg13g2_fill_2 FILLER_15_674 ();
 sg13g2_decap_8 FILLER_15_680 ();
 sg13g2_decap_8 FILLER_15_687 ();
 sg13g2_decap_8 FILLER_15_694 ();
 sg13g2_decap_4 FILLER_15_701 ();
 sg13g2_fill_1 FILLER_15_705 ();
 sg13g2_fill_1 FILLER_15_732 ();
 sg13g2_fill_1 FILLER_15_759 ();
 sg13g2_fill_1 FILLER_15_765 ();
 sg13g2_fill_1 FILLER_15_771 ();
 sg13g2_fill_1 FILLER_15_777 ();
 sg13g2_fill_2 FILLER_15_783 ();
 sg13g2_fill_2 FILLER_15_789 ();
 sg13g2_fill_2 FILLER_15_801 ();
 sg13g2_fill_1 FILLER_15_807 ();
 sg13g2_fill_2 FILLER_15_812 ();
 sg13g2_fill_1 FILLER_15_814 ();
 sg13g2_decap_8 FILLER_15_829 ();
 sg13g2_fill_2 FILLER_15_862 ();
 sg13g2_fill_2 FILLER_15_868 ();
 sg13g2_fill_2 FILLER_15_880 ();
 sg13g2_fill_1 FILLER_15_882 ();
 sg13g2_fill_1 FILLER_15_935 ();
 sg13g2_fill_1 FILLER_15_940 ();
 sg13g2_fill_2 FILLER_15_967 ();
 sg13g2_fill_1 FILLER_15_969 ();
 sg13g2_decap_8 FILLER_15_996 ();
 sg13g2_fill_2 FILLER_15_1003 ();
 sg13g2_fill_1 FILLER_15_1005 ();
 sg13g2_fill_2 FILLER_15_1081 ();
 sg13g2_fill_2 FILLER_15_1163 ();
 sg13g2_decap_8 FILLER_15_1169 ();
 sg13g2_decap_8 FILLER_15_1176 ();
 sg13g2_decap_8 FILLER_15_1183 ();
 sg13g2_fill_1 FILLER_15_1190 ();
 sg13g2_decap_8 FILLER_15_1195 ();
 sg13g2_decap_8 FILLER_15_1202 ();
 sg13g2_fill_2 FILLER_15_1209 ();
 sg13g2_fill_1 FILLER_15_1211 ();
 sg13g2_decap_8 FILLER_15_1220 ();
 sg13g2_decap_8 FILLER_15_1232 ();
 sg13g2_decap_8 FILLER_15_1331 ();
 sg13g2_decap_4 FILLER_15_1342 ();
 sg13g2_fill_1 FILLER_15_1346 ();
 sg13g2_fill_1 FILLER_15_1351 ();
 sg13g2_fill_1 FILLER_15_1357 ();
 sg13g2_decap_8 FILLER_15_1384 ();
 sg13g2_fill_2 FILLER_15_1427 ();
 sg13g2_decap_8 FILLER_15_1436 ();
 sg13g2_decap_8 FILLER_15_1443 ();
 sg13g2_fill_1 FILLER_15_1450 ();
 sg13g2_decap_4 FILLER_15_1485 ();
 sg13g2_fill_2 FILLER_15_1489 ();
 sg13g2_fill_2 FILLER_15_1498 ();
 sg13g2_fill_1 FILLER_15_1500 ();
 sg13g2_fill_2 FILLER_15_1514 ();
 sg13g2_fill_1 FILLER_15_1516 ();
 sg13g2_fill_2 FILLER_15_1521 ();
 sg13g2_decap_8 FILLER_15_1552 ();
 sg13g2_decap_4 FILLER_15_1559 ();
 sg13g2_fill_1 FILLER_15_1573 ();
 sg13g2_decap_4 FILLER_15_1577 ();
 sg13g2_fill_1 FILLER_15_1581 ();
 sg13g2_decap_8 FILLER_15_1586 ();
 sg13g2_fill_2 FILLER_15_1593 ();
 sg13g2_fill_1 FILLER_15_1595 ();
 sg13g2_fill_2 FILLER_15_1620 ();
 sg13g2_fill_2 FILLER_15_1648 ();
 sg13g2_fill_1 FILLER_15_1650 ();
 sg13g2_decap_8 FILLER_15_1713 ();
 sg13g2_decap_8 FILLER_15_1720 ();
 sg13g2_fill_2 FILLER_15_1731 ();
 sg13g2_fill_1 FILLER_15_1733 ();
 sg13g2_fill_1 FILLER_15_1781 ();
 sg13g2_decap_8 FILLER_15_1786 ();
 sg13g2_decap_4 FILLER_15_1793 ();
 sg13g2_decap_4 FILLER_15_1805 ();
 sg13g2_fill_1 FILLER_15_1809 ();
 sg13g2_decap_8 FILLER_15_1814 ();
 sg13g2_decap_8 FILLER_15_1821 ();
 sg13g2_decap_4 FILLER_15_1828 ();
 sg13g2_fill_1 FILLER_15_1832 ();
 sg13g2_decap_4 FILLER_15_1843 ();
 sg13g2_fill_2 FILLER_15_1847 ();
 sg13g2_decap_4 FILLER_15_1855 ();
 sg13g2_fill_1 FILLER_15_1859 ();
 sg13g2_decap_8 FILLER_15_1923 ();
 sg13g2_fill_1 FILLER_15_1930 ();
 sg13g2_fill_2 FILLER_15_1947 ();
 sg13g2_decap_8 FILLER_15_1975 ();
 sg13g2_decap_8 FILLER_15_1982 ();
 sg13g2_decap_4 FILLER_15_1989 ();
 sg13g2_fill_1 FILLER_15_1993 ();
 sg13g2_decap_4 FILLER_15_1998 ();
 sg13g2_decap_4 FILLER_15_2015 ();
 sg13g2_fill_2 FILLER_15_2019 ();
 sg13g2_decap_8 FILLER_15_2029 ();
 sg13g2_decap_8 FILLER_15_2036 ();
 sg13g2_fill_1 FILLER_15_2165 ();
 sg13g2_fill_1 FILLER_15_2195 ();
 sg13g2_fill_2 FILLER_15_2251 ();
 sg13g2_fill_1 FILLER_15_2315 ();
 sg13g2_decap_4 FILLER_15_2357 ();
 sg13g2_decap_8 FILLER_15_2365 ();
 sg13g2_fill_2 FILLER_15_2372 ();
 sg13g2_decap_8 FILLER_15_2378 ();
 sg13g2_decap_8 FILLER_15_2385 ();
 sg13g2_fill_1 FILLER_15_2392 ();
 sg13g2_fill_1 FILLER_15_2457 ();
 sg13g2_decap_8 FILLER_15_2497 ();
 sg13g2_decap_4 FILLER_15_2504 ();
 sg13g2_fill_1 FILLER_15_2508 ();
 sg13g2_decap_8 FILLER_15_2561 ();
 sg13g2_fill_2 FILLER_15_2568 ();
 sg13g2_fill_2 FILLER_15_2612 ();
 sg13g2_fill_2 FILLER_15_2618 ();
 sg13g2_fill_1 FILLER_15_2620 ();
 sg13g2_fill_2 FILLER_15_2668 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_4 FILLER_16_7 ();
 sg13g2_fill_1 FILLER_16_42 ();
 sg13g2_fill_1 FILLER_16_48 ();
 sg13g2_fill_1 FILLER_16_75 ();
 sg13g2_fill_2 FILLER_16_91 ();
 sg13g2_fill_2 FILLER_16_98 ();
 sg13g2_fill_1 FILLER_16_109 ();
 sg13g2_fill_2 FILLER_16_114 ();
 sg13g2_decap_8 FILLER_16_156 ();
 sg13g2_fill_1 FILLER_16_163 ();
 sg13g2_fill_2 FILLER_16_173 ();
 sg13g2_fill_2 FILLER_16_179 ();
 sg13g2_fill_2 FILLER_16_206 ();
 sg13g2_fill_1 FILLER_16_208 ();
 sg13g2_fill_2 FILLER_16_235 ();
 sg13g2_fill_2 FILLER_16_241 ();
 sg13g2_fill_1 FILLER_16_248 ();
 sg13g2_fill_1 FILLER_16_253 ();
 sg13g2_fill_2 FILLER_16_258 ();
 sg13g2_fill_2 FILLER_16_264 ();
 sg13g2_fill_2 FILLER_16_270 ();
 sg13g2_fill_2 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_fill_2 FILLER_16_294 ();
 sg13g2_fill_1 FILLER_16_304 ();
 sg13g2_fill_1 FILLER_16_325 ();
 sg13g2_fill_2 FILLER_16_335 ();
 sg13g2_decap_4 FILLER_16_346 ();
 sg13g2_fill_1 FILLER_16_350 ();
 sg13g2_fill_2 FILLER_16_357 ();
 sg13g2_fill_1 FILLER_16_364 ();
 sg13g2_fill_2 FILLER_16_396 ();
 sg13g2_fill_1 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_16_408 ();
 sg13g2_decap_4 FILLER_16_415 ();
 sg13g2_fill_2 FILLER_16_419 ();
 sg13g2_decap_4 FILLER_16_425 ();
 sg13g2_fill_2 FILLER_16_429 ();
 sg13g2_fill_1 FILLER_16_435 ();
 sg13g2_fill_1 FILLER_16_456 ();
 sg13g2_fill_2 FILLER_16_462 ();
 sg13g2_decap_4 FILLER_16_468 ();
 sg13g2_decap_4 FILLER_16_482 ();
 sg13g2_fill_1 FILLER_16_486 ();
 sg13g2_decap_8 FILLER_16_497 ();
 sg13g2_decap_8 FILLER_16_504 ();
 sg13g2_fill_1 FILLER_16_511 ();
 sg13g2_decap_4 FILLER_16_538 ();
 sg13g2_fill_1 FILLER_16_542 ();
 sg13g2_fill_2 FILLER_16_547 ();
 sg13g2_fill_2 FILLER_16_567 ();
 sg13g2_fill_2 FILLER_16_603 ();
 sg13g2_fill_1 FILLER_16_605 ();
 sg13g2_decap_8 FILLER_16_610 ();
 sg13g2_fill_1 FILLER_16_617 ();
 sg13g2_decap_8 FILLER_16_657 ();
 sg13g2_decap_8 FILLER_16_664 ();
 sg13g2_decap_8 FILLER_16_671 ();
 sg13g2_decap_8 FILLER_16_678 ();
 sg13g2_fill_1 FILLER_16_685 ();
 sg13g2_decap_8 FILLER_16_690 ();
 sg13g2_fill_1 FILLER_16_697 ();
 sg13g2_fill_2 FILLER_16_702 ();
 sg13g2_fill_2 FILLER_16_713 ();
 sg13g2_fill_1 FILLER_16_715 ();
 sg13g2_fill_2 FILLER_16_729 ();
 sg13g2_fill_1 FILLER_16_731 ();
 sg13g2_decap_8 FILLER_16_746 ();
 sg13g2_fill_1 FILLER_16_772 ();
 sg13g2_fill_1 FILLER_16_778 ();
 sg13g2_decap_8 FILLER_16_793 ();
 sg13g2_decap_8 FILLER_16_800 ();
 sg13g2_fill_1 FILLER_16_807 ();
 sg13g2_decap_4 FILLER_16_818 ();
 sg13g2_decap_8 FILLER_16_841 ();
 sg13g2_decap_4 FILLER_16_848 ();
 sg13g2_fill_1 FILLER_16_852 ();
 sg13g2_fill_1 FILLER_16_896 ();
 sg13g2_decap_8 FILLER_16_935 ();
 sg13g2_fill_2 FILLER_16_942 ();
 sg13g2_fill_1 FILLER_16_944 ();
 sg13g2_fill_1 FILLER_16_959 ();
 sg13g2_decap_4 FILLER_16_996 ();
 sg13g2_fill_1 FILLER_16_1000 ();
 sg13g2_fill_2 FILLER_16_1045 ();
 sg13g2_fill_2 FILLER_16_1147 ();
 sg13g2_fill_1 FILLER_16_1149 ();
 sg13g2_fill_1 FILLER_16_1176 ();
 sg13g2_fill_1 FILLER_16_1215 ();
 sg13g2_decap_4 FILLER_16_1224 ();
 sg13g2_decap_8 FILLER_16_1236 ();
 sg13g2_fill_1 FILLER_16_1243 ();
 sg13g2_decap_8 FILLER_16_1248 ();
 sg13g2_decap_4 FILLER_16_1255 ();
 sg13g2_fill_1 FILLER_16_1259 ();
 sg13g2_fill_2 FILLER_16_1264 ();
 sg13g2_fill_2 FILLER_16_1274 ();
 sg13g2_decap_4 FILLER_16_1301 ();
 sg13g2_fill_2 FILLER_16_1305 ();
 sg13g2_decap_4 FILLER_16_1315 ();
 sg13g2_fill_1 FILLER_16_1323 ();
 sg13g2_fill_1 FILLER_16_1345 ();
 sg13g2_fill_1 FILLER_16_1351 ();
 sg13g2_fill_1 FILLER_16_1360 ();
 sg13g2_fill_2 FILLER_16_1365 ();
 sg13g2_decap_8 FILLER_16_1371 ();
 sg13g2_fill_1 FILLER_16_1378 ();
 sg13g2_fill_1 FILLER_16_1431 ();
 sg13g2_fill_2 FILLER_16_1436 ();
 sg13g2_decap_4 FILLER_16_1472 ();
 sg13g2_fill_2 FILLER_16_1476 ();
 sg13g2_decap_8 FILLER_16_1488 ();
 sg13g2_fill_1 FILLER_16_1495 ();
 sg13g2_fill_2 FILLER_16_1508 ();
 sg13g2_fill_1 FILLER_16_1533 ();
 sg13g2_decap_8 FILLER_16_1539 ();
 sg13g2_decap_8 FILLER_16_1546 ();
 sg13g2_fill_2 FILLER_16_1592 ();
 sg13g2_decap_4 FILLER_16_1599 ();
 sg13g2_fill_1 FILLER_16_1603 ();
 sg13g2_decap_8 FILLER_16_1665 ();
 sg13g2_decap_8 FILLER_16_1676 ();
 sg13g2_decap_8 FILLER_16_1683 ();
 sg13g2_decap_4 FILLER_16_1690 ();
 sg13g2_fill_2 FILLER_16_1698 ();
 sg13g2_fill_1 FILLER_16_1700 ();
 sg13g2_decap_4 FILLER_16_1711 ();
 sg13g2_decap_8 FILLER_16_1719 ();
 sg13g2_decap_8 FILLER_16_1726 ();
 sg13g2_decap_4 FILLER_16_1733 ();
 sg13g2_decap_8 FILLER_16_1791 ();
 sg13g2_decap_8 FILLER_16_1798 ();
 sg13g2_fill_1 FILLER_16_1805 ();
 sg13g2_decap_4 FILLER_16_1811 ();
 sg13g2_fill_2 FILLER_16_1815 ();
 sg13g2_decap_8 FILLER_16_1831 ();
 sg13g2_fill_2 FILLER_16_1838 ();
 sg13g2_fill_1 FILLER_16_1861 ();
 sg13g2_decap_8 FILLER_16_1902 ();
 sg13g2_decap_8 FILLER_16_1909 ();
 sg13g2_decap_8 FILLER_16_1920 ();
 sg13g2_fill_2 FILLER_16_1941 ();
 sg13g2_decap_8 FILLER_16_1999 ();
 sg13g2_decap_8 FILLER_16_2006 ();
 sg13g2_fill_2 FILLER_16_2013 ();
 sg13g2_fill_1 FILLER_16_2101 ();
 sg13g2_fill_1 FILLER_16_2117 ();
 sg13g2_decap_4 FILLER_16_2122 ();
 sg13g2_fill_1 FILLER_16_2126 ();
 sg13g2_decap_8 FILLER_16_2131 ();
 sg13g2_fill_1 FILLER_16_2138 ();
 sg13g2_fill_2 FILLER_16_2143 ();
 sg13g2_fill_1 FILLER_16_2145 ();
 sg13g2_fill_2 FILLER_16_2221 ();
 sg13g2_decap_4 FILLER_16_2236 ();
 sg13g2_decap_4 FILLER_16_2261 ();
 sg13g2_fill_2 FILLER_16_2265 ();
 sg13g2_decap_4 FILLER_16_2311 ();
 sg13g2_fill_1 FILLER_16_2315 ();
 sg13g2_decap_8 FILLER_16_2341 ();
 sg13g2_decap_8 FILLER_16_2348 ();
 sg13g2_fill_2 FILLER_16_2355 ();
 sg13g2_fill_1 FILLER_16_2367 ();
 sg13g2_fill_1 FILLER_16_2377 ();
 sg13g2_fill_1 FILLER_16_2412 ();
 sg13g2_fill_1 FILLER_16_2465 ();
 sg13g2_fill_2 FILLER_16_2521 ();
 sg13g2_fill_1 FILLER_16_2523 ();
 sg13g2_fill_2 FILLER_16_2545 ();
 sg13g2_fill_1 FILLER_16_2547 ();
 sg13g2_decap_4 FILLER_16_2574 ();
 sg13g2_fill_2 FILLER_16_2578 ();
 sg13g2_fill_2 FILLER_16_2629 ();
 sg13g2_fill_1 FILLER_16_2631 ();
 sg13g2_fill_2 FILLER_16_2668 ();
 sg13g2_decap_4 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_46 ();
 sg13g2_fill_1 FILLER_17_48 ();
 sg13g2_fill_1 FILLER_17_64 ();
 sg13g2_fill_2 FILLER_17_138 ();
 sg13g2_fill_1 FILLER_17_140 ();
 sg13g2_fill_1 FILLER_17_156 ();
 sg13g2_decap_4 FILLER_17_183 ();
 sg13g2_decap_4 FILLER_17_191 ();
 sg13g2_fill_1 FILLER_17_195 ();
 sg13g2_decap_4 FILLER_17_205 ();
 sg13g2_fill_2 FILLER_17_209 ();
 sg13g2_fill_2 FILLER_17_218 ();
 sg13g2_fill_1 FILLER_17_252 ();
 sg13g2_fill_1 FILLER_17_278 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_4 FILLER_17_294 ();
 sg13g2_fill_2 FILLER_17_348 ();
 sg13g2_fill_1 FILLER_17_350 ();
 sg13g2_fill_2 FILLER_17_375 ();
 sg13g2_fill_1 FILLER_17_381 ();
 sg13g2_decap_8 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_17_415 ();
 sg13g2_decap_8 FILLER_17_422 ();
 sg13g2_fill_2 FILLER_17_429 ();
 sg13g2_fill_2 FILLER_17_455 ();
 sg13g2_fill_1 FILLER_17_457 ();
 sg13g2_fill_2 FILLER_17_474 ();
 sg13g2_fill_1 FILLER_17_476 ();
 sg13g2_decap_4 FILLER_17_481 ();
 sg13g2_fill_1 FILLER_17_485 ();
 sg13g2_decap_8 FILLER_17_490 ();
 sg13g2_decap_8 FILLER_17_497 ();
 sg13g2_fill_1 FILLER_17_504 ();
 sg13g2_fill_2 FILLER_17_513 ();
 sg13g2_fill_1 FILLER_17_515 ();
 sg13g2_fill_2 FILLER_17_527 ();
 sg13g2_fill_1 FILLER_17_529 ();
 sg13g2_fill_1 FILLER_17_547 ();
 sg13g2_fill_2 FILLER_17_556 ();
 sg13g2_fill_1 FILLER_17_595 ();
 sg13g2_decap_8 FILLER_17_607 ();
 sg13g2_decap_8 FILLER_17_614 ();
 sg13g2_fill_1 FILLER_17_625 ();
 sg13g2_fill_1 FILLER_17_633 ();
 sg13g2_fill_1 FILLER_17_659 ();
 sg13g2_fill_1 FILLER_17_666 ();
 sg13g2_fill_1 FILLER_17_673 ();
 sg13g2_fill_1 FILLER_17_678 ();
 sg13g2_fill_2 FILLER_17_684 ();
 sg13g2_decap_4 FILLER_17_722 ();
 sg13g2_fill_2 FILLER_17_736 ();
 sg13g2_fill_1 FILLER_17_738 ();
 sg13g2_decap_8 FILLER_17_744 ();
 sg13g2_decap_8 FILLER_17_751 ();
 sg13g2_fill_2 FILLER_17_758 ();
 sg13g2_decap_8 FILLER_17_805 ();
 sg13g2_decap_8 FILLER_17_812 ();
 sg13g2_decap_4 FILLER_17_819 ();
 sg13g2_fill_1 FILLER_17_859 ();
 sg13g2_decap_8 FILLER_17_889 ();
 sg13g2_fill_2 FILLER_17_896 ();
 sg13g2_fill_1 FILLER_17_929 ();
 sg13g2_decap_4 FILLER_17_956 ();
 sg13g2_decap_8 FILLER_17_970 ();
 sg13g2_fill_1 FILLER_17_977 ();
 sg13g2_decap_8 FILLER_17_986 ();
 sg13g2_decap_8 FILLER_17_993 ();
 sg13g2_fill_2 FILLER_17_1000 ();
 sg13g2_fill_2 FILLER_17_1048 ();
 sg13g2_fill_2 FILLER_17_1054 ();
 sg13g2_fill_1 FILLER_17_1082 ();
 sg13g2_fill_1 FILLER_17_1088 ();
 sg13g2_fill_1 FILLER_17_1123 ();
 sg13g2_decap_4 FILLER_17_1199 ();
 sg13g2_fill_1 FILLER_17_1203 ();
 sg13g2_decap_8 FILLER_17_1261 ();
 sg13g2_fill_2 FILLER_17_1268 ();
 sg13g2_fill_2 FILLER_17_1282 ();
 sg13g2_fill_1 FILLER_17_1284 ();
 sg13g2_fill_2 FILLER_17_1314 ();
 sg13g2_decap_4 FILLER_17_1320 ();
 sg13g2_fill_1 FILLER_17_1324 ();
 sg13g2_fill_1 FILLER_17_1341 ();
 sg13g2_fill_1 FILLER_17_1347 ();
 sg13g2_fill_2 FILLER_17_1374 ();
 sg13g2_fill_1 FILLER_17_1376 ();
 sg13g2_fill_2 FILLER_17_1413 ();
 sg13g2_fill_1 FILLER_17_1415 ();
 sg13g2_decap_8 FILLER_17_1420 ();
 sg13g2_fill_2 FILLER_17_1427 ();
 sg13g2_fill_1 FILLER_17_1429 ();
 sg13g2_decap_8 FILLER_17_1445 ();
 sg13g2_decap_4 FILLER_17_1452 ();
 sg13g2_fill_2 FILLER_17_1456 ();
 sg13g2_decap_4 FILLER_17_1484 ();
 sg13g2_fill_2 FILLER_17_1499 ();
 sg13g2_fill_1 FILLER_17_1533 ();
 sg13g2_decap_8 FILLER_17_1538 ();
 sg13g2_decap_8 FILLER_17_1545 ();
 sg13g2_decap_4 FILLER_17_1552 ();
 sg13g2_decap_4 FILLER_17_1560 ();
 sg13g2_fill_1 FILLER_17_1564 ();
 sg13g2_fill_1 FILLER_17_1570 ();
 sg13g2_fill_2 FILLER_17_1576 ();
 sg13g2_fill_2 FILLER_17_1588 ();
 sg13g2_fill_2 FILLER_17_1594 ();
 sg13g2_fill_1 FILLER_17_1596 ();
 sg13g2_fill_2 FILLER_17_1612 ();
 sg13g2_fill_2 FILLER_17_1632 ();
 sg13g2_fill_1 FILLER_17_1649 ();
 sg13g2_decap_8 FILLER_17_1658 ();
 sg13g2_decap_8 FILLER_17_1665 ();
 sg13g2_decap_4 FILLER_17_1672 ();
 sg13g2_fill_1 FILLER_17_1676 ();
 sg13g2_decap_4 FILLER_17_1772 ();
 sg13g2_decap_8 FILLER_17_1802 ();
 sg13g2_decap_8 FILLER_17_1809 ();
 sg13g2_decap_4 FILLER_17_1816 ();
 sg13g2_fill_1 FILLER_17_1820 ();
 sg13g2_fill_1 FILLER_17_1847 ();
 sg13g2_decap_8 FILLER_17_1891 ();
 sg13g2_decap_4 FILLER_17_1898 ();
 sg13g2_fill_1 FILLER_17_1902 ();
 sg13g2_decap_4 FILLER_17_1912 ();
 sg13g2_fill_2 FILLER_17_1916 ();
 sg13g2_fill_1 FILLER_17_1922 ();
 sg13g2_fill_2 FILLER_17_1933 ();
 sg13g2_fill_1 FILLER_17_1971 ();
 sg13g2_fill_2 FILLER_17_1976 ();
 sg13g2_decap_4 FILLER_17_2014 ();
 sg13g2_fill_2 FILLER_17_2022 ();
 sg13g2_fill_1 FILLER_17_2029 ();
 sg13g2_fill_1 FILLER_17_2034 ();
 sg13g2_fill_1 FILLER_17_2070 ();
 sg13g2_fill_2 FILLER_17_2075 ();
 sg13g2_fill_1 FILLER_17_2092 ();
 sg13g2_decap_8 FILLER_17_2118 ();
 sg13g2_decap_8 FILLER_17_2125 ();
 sg13g2_fill_2 FILLER_17_2132 ();
 sg13g2_fill_1 FILLER_17_2134 ();
 sg13g2_decap_8 FILLER_17_2143 ();
 sg13g2_fill_1 FILLER_17_2150 ();
 sg13g2_decap_4 FILLER_17_2155 ();
 sg13g2_fill_2 FILLER_17_2159 ();
 sg13g2_decap_8 FILLER_17_2166 ();
 sg13g2_decap_8 FILLER_17_2194 ();
 sg13g2_decap_4 FILLER_17_2217 ();
 sg13g2_fill_1 FILLER_17_2221 ();
 sg13g2_decap_8 FILLER_17_2243 ();
 sg13g2_decap_8 FILLER_17_2250 ();
 sg13g2_fill_2 FILLER_17_2257 ();
 sg13g2_fill_1 FILLER_17_2259 ();
 sg13g2_decap_4 FILLER_17_2300 ();
 sg13g2_fill_1 FILLER_17_2304 ();
 sg13g2_decap_8 FILLER_17_2341 ();
 sg13g2_decap_4 FILLER_17_2348 ();
 sg13g2_fill_2 FILLER_17_2352 ();
 sg13g2_fill_2 FILLER_17_2390 ();
 sg13g2_fill_1 FILLER_17_2475 ();
 sg13g2_decap_4 FILLER_17_2480 ();
 sg13g2_decap_4 FILLER_17_2488 ();
 sg13g2_fill_1 FILLER_17_2492 ();
 sg13g2_decap_4 FILLER_17_2503 ();
 sg13g2_fill_2 FILLER_17_2507 ();
 sg13g2_fill_2 FILLER_17_2519 ();
 sg13g2_fill_1 FILLER_17_2540 ();
 sg13g2_fill_1 FILLER_17_2551 ();
 sg13g2_fill_1 FILLER_17_2588 ();
 sg13g2_fill_2 FILLER_17_2655 ();
 sg13g2_decap_8 FILLER_17_2661 ();
 sg13g2_fill_2 FILLER_17_2668 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_fill_2 FILLER_18_41 ();
 sg13g2_fill_1 FILLER_18_43 ();
 sg13g2_fill_1 FILLER_18_89 ();
 sg13g2_fill_2 FILLER_18_119 ();
 sg13g2_fill_2 FILLER_18_128 ();
 sg13g2_fill_1 FILLER_18_138 ();
 sg13g2_fill_2 FILLER_18_144 ();
 sg13g2_fill_1 FILLER_18_146 ();
 sg13g2_decap_8 FILLER_18_151 ();
 sg13g2_decap_4 FILLER_18_158 ();
 sg13g2_fill_2 FILLER_18_162 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_fill_1 FILLER_18_189 ();
 sg13g2_fill_2 FILLER_18_194 ();
 sg13g2_decap_8 FILLER_18_222 ();
 sg13g2_fill_1 FILLER_18_234 ();
 sg13g2_fill_1 FILLER_18_238 ();
 sg13g2_fill_1 FILLER_18_266 ();
 sg13g2_fill_1 FILLER_18_303 ();
 sg13g2_decap_8 FILLER_18_342 ();
 sg13g2_decap_4 FILLER_18_349 ();
 sg13g2_fill_1 FILLER_18_353 ();
 sg13g2_fill_1 FILLER_18_370 ();
 sg13g2_fill_1 FILLER_18_375 ();
 sg13g2_fill_1 FILLER_18_380 ();
 sg13g2_fill_2 FILLER_18_390 ();
 sg13g2_fill_1 FILLER_18_392 ();
 sg13g2_fill_1 FILLER_18_397 ();
 sg13g2_decap_8 FILLER_18_402 ();
 sg13g2_decap_4 FILLER_18_409 ();
 sg13g2_fill_1 FILLER_18_413 ();
 sg13g2_fill_2 FILLER_18_440 ();
 sg13g2_fill_1 FILLER_18_442 ();
 sg13g2_fill_1 FILLER_18_453 ();
 sg13g2_fill_2 FILLER_18_506 ();
 sg13g2_fill_1 FILLER_18_508 ();
 sg13g2_fill_2 FILLER_18_522 ();
 sg13g2_fill_2 FILLER_18_530 ();
 sg13g2_fill_1 FILLER_18_558 ();
 sg13g2_fill_2 FILLER_18_608 ();
 sg13g2_fill_2 FILLER_18_650 ();
 sg13g2_fill_2 FILLER_18_658 ();
 sg13g2_fill_1 FILLER_18_660 ();
 sg13g2_fill_1 FILLER_18_667 ();
 sg13g2_fill_2 FILLER_18_699 ();
 sg13g2_fill_1 FILLER_18_701 ();
 sg13g2_decap_8 FILLER_18_707 ();
 sg13g2_decap_8 FILLER_18_714 ();
 sg13g2_decap_8 FILLER_18_721 ();
 sg13g2_fill_2 FILLER_18_728 ();
 sg13g2_fill_1 FILLER_18_730 ();
 sg13g2_decap_4 FILLER_18_739 ();
 sg13g2_decap_8 FILLER_18_749 ();
 sg13g2_fill_2 FILLER_18_756 ();
 sg13g2_decap_8 FILLER_18_762 ();
 sg13g2_decap_4 FILLER_18_769 ();
 sg13g2_fill_2 FILLER_18_773 ();
 sg13g2_decap_8 FILLER_18_829 ();
 sg13g2_decap_8 FILLER_18_836 ();
 sg13g2_fill_2 FILLER_18_843 ();
 sg13g2_fill_1 FILLER_18_845 ();
 sg13g2_fill_1 FILLER_18_872 ();
 sg13g2_decap_8 FILLER_18_883 ();
 sg13g2_decap_4 FILLER_18_890 ();
 sg13g2_decap_8 FILLER_18_904 ();
 sg13g2_decap_8 FILLER_18_911 ();
 sg13g2_decap_4 FILLER_18_918 ();
 sg13g2_fill_2 FILLER_18_922 ();
 sg13g2_decap_8 FILLER_18_960 ();
 sg13g2_fill_2 FILLER_18_967 ();
 sg13g2_fill_1 FILLER_18_969 ();
 sg13g2_decap_8 FILLER_18_974 ();
 sg13g2_fill_2 FILLER_18_981 ();
 sg13g2_fill_1 FILLER_18_993 ();
 sg13g2_fill_2 FILLER_18_1088 ();
 sg13g2_fill_1 FILLER_18_1103 ();
 sg13g2_fill_2 FILLER_18_1138 ();
 sg13g2_fill_2 FILLER_18_1162 ();
 sg13g2_fill_1 FILLER_18_1164 ();
 sg13g2_fill_1 FILLER_18_1170 ();
 sg13g2_fill_1 FILLER_18_1197 ();
 sg13g2_fill_2 FILLER_18_1206 ();
 sg13g2_decap_8 FILLER_18_1260 ();
 sg13g2_decap_4 FILLER_18_1267 ();
 sg13g2_fill_2 FILLER_18_1271 ();
 sg13g2_fill_2 FILLER_18_1277 ();
 sg13g2_fill_1 FILLER_18_1279 ();
 sg13g2_decap_8 FILLER_18_1366 ();
 sg13g2_fill_1 FILLER_18_1373 ();
 sg13g2_fill_1 FILLER_18_1388 ();
 sg13g2_decap_4 FILLER_18_1402 ();
 sg13g2_fill_2 FILLER_18_1420 ();
 sg13g2_fill_1 FILLER_18_1422 ();
 sg13g2_decap_8 FILLER_18_1438 ();
 sg13g2_decap_8 FILLER_18_1445 ();
 sg13g2_fill_1 FILLER_18_1452 ();
 sg13g2_fill_2 FILLER_18_1459 ();
 sg13g2_fill_1 FILLER_18_1485 ();
 sg13g2_fill_1 FILLER_18_1502 ();
 sg13g2_fill_1 FILLER_18_1508 ();
 sg13g2_fill_1 FILLER_18_1514 ();
 sg13g2_fill_1 FILLER_18_1520 ();
 sg13g2_fill_1 FILLER_18_1525 ();
 sg13g2_decap_4 FILLER_18_1535 ();
 sg13g2_fill_2 FILLER_18_1539 ();
 sg13g2_fill_1 FILLER_18_1545 ();
 sg13g2_decap_8 FILLER_18_1610 ();
 sg13g2_fill_1 FILLER_18_1640 ();
 sg13g2_fill_2 FILLER_18_1648 ();
 sg13g2_fill_2 FILLER_18_1660 ();
 sg13g2_decap_4 FILLER_18_1676 ();
 sg13g2_fill_2 FILLER_18_1690 ();
 sg13g2_decap_4 FILLER_18_1701 ();
 sg13g2_fill_2 FILLER_18_1755 ();
 sg13g2_decap_4 FILLER_18_1783 ();
 sg13g2_fill_2 FILLER_18_1787 ();
 sg13g2_fill_2 FILLER_18_1815 ();
 sg13g2_fill_1 FILLER_18_1883 ();
 sg13g2_decap_8 FILLER_18_1888 ();
 sg13g2_decap_8 FILLER_18_1895 ();
 sg13g2_decap_4 FILLER_18_1902 ();
 sg13g2_fill_2 FILLER_18_1906 ();
 sg13g2_fill_2 FILLER_18_1941 ();
 sg13g2_fill_2 FILLER_18_2035 ();
 sg13g2_decap_4 FILLER_18_2067 ();
 sg13g2_fill_1 FILLER_18_2071 ();
 sg13g2_decap_4 FILLER_18_2119 ();
 sg13g2_decap_8 FILLER_18_2127 ();
 sg13g2_decap_4 FILLER_18_2134 ();
 sg13g2_fill_1 FILLER_18_2138 ();
 sg13g2_fill_1 FILLER_18_2143 ();
 sg13g2_fill_2 FILLER_18_2148 ();
 sg13g2_decap_4 FILLER_18_2176 ();
 sg13g2_decap_8 FILLER_18_2190 ();
 sg13g2_decap_8 FILLER_18_2197 ();
 sg13g2_fill_1 FILLER_18_2204 ();
 sg13g2_fill_2 FILLER_18_2249 ();
 sg13g2_decap_8 FILLER_18_2261 ();
 sg13g2_fill_2 FILLER_18_2268 ();
 sg13g2_fill_2 FILLER_18_2306 ();
 sg13g2_decap_4 FILLER_18_2344 ();
 sg13g2_fill_1 FILLER_18_2400 ();
 sg13g2_fill_2 FILLER_18_2411 ();
 sg13g2_fill_1 FILLER_18_2427 ();
 sg13g2_fill_2 FILLER_18_2431 ();
 sg13g2_fill_1 FILLER_18_2436 ();
 sg13g2_fill_2 FILLER_18_2447 ();
 sg13g2_decap_4 FILLER_18_2498 ();
 sg13g2_fill_2 FILLER_18_2502 ();
 sg13g2_decap_8 FILLER_18_2508 ();
 sg13g2_decap_8 FILLER_18_2518 ();
 sg13g2_decap_8 FILLER_18_2525 ();
 sg13g2_decap_8 FILLER_18_2532 ();
 sg13g2_decap_8 FILLER_18_2539 ();
 sg13g2_fill_1 FILLER_18_2546 ();
 sg13g2_fill_1 FILLER_18_2561 ();
 sg13g2_fill_1 FILLER_18_2567 ();
 sg13g2_fill_1 FILLER_18_2572 ();
 sg13g2_fill_1 FILLER_18_2599 ();
 sg13g2_decap_4 FILLER_18_2607 ();
 sg13g2_decap_8 FILLER_18_2621 ();
 sg13g2_decap_4 FILLER_18_2628 ();
 sg13g2_fill_1 FILLER_18_2632 ();
 sg13g2_decap_8 FILLER_18_2637 ();
 sg13g2_decap_8 FILLER_18_2644 ();
 sg13g2_decap_8 FILLER_18_2651 ();
 sg13g2_decap_8 FILLER_18_2658 ();
 sg13g2_decap_4 FILLER_18_2665 ();
 sg13g2_fill_1 FILLER_18_2669 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_fill_1 FILLER_19_26 ();
 sg13g2_fill_2 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_148 ();
 sg13g2_fill_2 FILLER_19_155 ();
 sg13g2_decap_8 FILLER_19_192 ();
 sg13g2_decap_4 FILLER_19_199 ();
 sg13g2_fill_1 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_208 ();
 sg13g2_decap_8 FILLER_19_215 ();
 sg13g2_decap_8 FILLER_19_222 ();
 sg13g2_decap_4 FILLER_19_237 ();
 sg13g2_fill_2 FILLER_19_241 ();
 sg13g2_fill_1 FILLER_19_247 ();
 sg13g2_fill_1 FILLER_19_258 ();
 sg13g2_decap_4 FILLER_19_288 ();
 sg13g2_fill_2 FILLER_19_292 ();
 sg13g2_fill_2 FILLER_19_308 ();
 sg13g2_fill_1 FILLER_19_362 ();
 sg13g2_fill_2 FILLER_19_367 ();
 sg13g2_fill_1 FILLER_19_369 ();
 sg13g2_fill_1 FILLER_19_387 ();
 sg13g2_fill_1 FILLER_19_461 ();
 sg13g2_fill_1 FILLER_19_492 ();
 sg13g2_fill_1 FILLER_19_535 ();
 sg13g2_fill_2 FILLER_19_569 ();
 sg13g2_fill_2 FILLER_19_590 ();
 sg13g2_fill_1 FILLER_19_605 ();
 sg13g2_fill_1 FILLER_19_674 ();
 sg13g2_fill_1 FILLER_19_714 ();
 sg13g2_decap_4 FILLER_19_720 ();
 sg13g2_fill_1 FILLER_19_724 ();
 sg13g2_fill_1 FILLER_19_730 ();
 sg13g2_decap_8 FILLER_19_768 ();
 sg13g2_decap_4 FILLER_19_775 ();
 sg13g2_decap_4 FILLER_19_787 ();
 sg13g2_fill_2 FILLER_19_791 ();
 sg13g2_decap_8 FILLER_19_796 ();
 sg13g2_decap_8 FILLER_19_803 ();
 sg13g2_decap_8 FILLER_19_810 ();
 sg13g2_decap_8 FILLER_19_817 ();
 sg13g2_fill_2 FILLER_19_824 ();
 sg13g2_fill_2 FILLER_19_856 ();
 sg13g2_fill_1 FILLER_19_858 ();
 sg13g2_fill_1 FILLER_19_885 ();
 sg13g2_decap_8 FILLER_19_920 ();
 sg13g2_decap_4 FILLER_19_927 ();
 sg13g2_decap_8 FILLER_19_952 ();
 sg13g2_decap_4 FILLER_19_959 ();
 sg13g2_fill_1 FILLER_19_963 ();
 sg13g2_fill_2 FILLER_19_1000 ();
 sg13g2_fill_1 FILLER_19_1032 ();
 sg13g2_fill_1 FILLER_19_1219 ();
 sg13g2_fill_2 FILLER_19_1251 ();
 sg13g2_decap_4 FILLER_19_1300 ();
 sg13g2_decap_8 FILLER_19_1318 ();
 sg13g2_decap_4 FILLER_19_1325 ();
 sg13g2_decap_8 FILLER_19_1347 ();
 sg13g2_decap_8 FILLER_19_1354 ();
 sg13g2_fill_2 FILLER_19_1371 ();
 sg13g2_decap_8 FILLER_19_1377 ();
 sg13g2_fill_1 FILLER_19_1384 ();
 sg13g2_fill_2 FILLER_19_1389 ();
 sg13g2_decap_8 FILLER_19_1401 ();
 sg13g2_fill_2 FILLER_19_1408 ();
 sg13g2_fill_1 FILLER_19_1410 ();
 sg13g2_fill_2 FILLER_19_1421 ();
 sg13g2_fill_2 FILLER_19_1428 ();
 sg13g2_fill_1 FILLER_19_1430 ();
 sg13g2_decap_4 FILLER_19_1438 ();
 sg13g2_fill_1 FILLER_19_1442 ();
 sg13g2_fill_2 FILLER_19_1485 ();
 sg13g2_fill_2 FILLER_19_1509 ();
 sg13g2_fill_1 FILLER_19_1517 ();
 sg13g2_fill_1 FILLER_19_1528 ();
 sg13g2_decap_8 FILLER_19_1535 ();
 sg13g2_fill_2 FILLER_19_1542 ();
 sg13g2_fill_1 FILLER_19_1556 ();
 sg13g2_decap_4 FILLER_19_1585 ();
 sg13g2_fill_1 FILLER_19_1589 ();
 sg13g2_fill_2 FILLER_19_1600 ();
 sg13g2_fill_1 FILLER_19_1602 ();
 sg13g2_fill_1 FILLER_19_1608 ();
 sg13g2_fill_2 FILLER_19_1620 ();
 sg13g2_fill_2 FILLER_19_1653 ();
 sg13g2_fill_1 FILLER_19_1660 ();
 sg13g2_fill_2 FILLER_19_1677 ();
 sg13g2_fill_1 FILLER_19_1679 ();
 sg13g2_fill_2 FILLER_19_1690 ();
 sg13g2_fill_2 FILLER_19_1715 ();
 sg13g2_fill_2 FILLER_19_1743 ();
 sg13g2_fill_1 FILLER_19_1745 ();
 sg13g2_fill_2 FILLER_19_1759 ();
 sg13g2_fill_1 FILLER_19_1769 ();
 sg13g2_decap_4 FILLER_19_1780 ();
 sg13g2_fill_1 FILLER_19_1784 ();
 sg13g2_fill_1 FILLER_19_1795 ();
 sg13g2_decap_4 FILLER_19_1800 ();
 sg13g2_fill_2 FILLER_19_1823 ();
 sg13g2_fill_1 FILLER_19_1825 ();
 sg13g2_decap_8 FILLER_19_1872 ();
 sg13g2_decap_4 FILLER_19_1879 ();
 sg13g2_decap_8 FILLER_19_1888 ();
 sg13g2_fill_2 FILLER_19_1913 ();
 sg13g2_fill_1 FILLER_19_1919 ();
 sg13g2_decap_4 FILLER_19_1924 ();
 sg13g2_fill_1 FILLER_19_1928 ();
 sg13g2_fill_2 FILLER_19_1971 ();
 sg13g2_fill_2 FILLER_19_1983 ();
 sg13g2_fill_1 FILLER_19_1999 ();
 sg13g2_decap_8 FILLER_19_2010 ();
 sg13g2_fill_2 FILLER_19_2017 ();
 sg13g2_fill_1 FILLER_19_2019 ();
 sg13g2_decap_8 FILLER_19_2056 ();
 sg13g2_fill_2 FILLER_19_2063 ();
 sg13g2_fill_1 FILLER_19_2065 ();
 sg13g2_decap_4 FILLER_19_2076 ();
 sg13g2_fill_1 FILLER_19_2132 ();
 sg13g2_fill_1 FILLER_19_2159 ();
 sg13g2_fill_2 FILLER_19_2164 ();
 sg13g2_fill_1 FILLER_19_2232 ();
 sg13g2_fill_2 FILLER_19_2259 ();
 sg13g2_decap_8 FILLER_19_2287 ();
 sg13g2_fill_2 FILLER_19_2294 ();
 sg13g2_fill_2 FILLER_19_2306 ();
 sg13g2_decap_8 FILLER_19_2312 ();
 sg13g2_decap_4 FILLER_19_2319 ();
 sg13g2_fill_1 FILLER_19_2323 ();
 sg13g2_fill_1 FILLER_19_2344 ();
 sg13g2_fill_2 FILLER_19_2354 ();
 sg13g2_fill_1 FILLER_19_2356 ();
 sg13g2_fill_2 FILLER_19_2361 ();
 sg13g2_fill_1 FILLER_19_2363 ();
 sg13g2_fill_1 FILLER_19_2385 ();
 sg13g2_decap_4 FILLER_19_2412 ();
 sg13g2_fill_1 FILLER_19_2419 ();
 sg13g2_fill_1 FILLER_19_2436 ();
 sg13g2_fill_1 FILLER_19_2461 ();
 sg13g2_decap_8 FILLER_19_2531 ();
 sg13g2_fill_2 FILLER_19_2538 ();
 sg13g2_decap_8 FILLER_19_2550 ();
 sg13g2_decap_4 FILLER_19_2557 ();
 sg13g2_fill_2 FILLER_19_2561 ();
 sg13g2_fill_2 FILLER_19_2576 ();
 sg13g2_fill_1 FILLER_19_2578 ();
 sg13g2_fill_1 FILLER_19_2583 ();
 sg13g2_fill_2 FILLER_19_2622 ();
 sg13g2_fill_1 FILLER_19_2624 ();
 sg13g2_fill_1 FILLER_19_2635 ();
 sg13g2_decap_8 FILLER_19_2662 ();
 sg13g2_fill_1 FILLER_19_2669 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_28 ();
 sg13g2_decap_4 FILLER_20_44 ();
 sg13g2_decap_8 FILLER_20_52 ();
 sg13g2_decap_8 FILLER_20_59 ();
 sg13g2_fill_2 FILLER_20_86 ();
 sg13g2_fill_1 FILLER_20_102 ();
 sg13g2_fill_1 FILLER_20_112 ();
 sg13g2_fill_2 FILLER_20_118 ();
 sg13g2_fill_1 FILLER_20_134 ();
 sg13g2_fill_1 FILLER_20_148 ();
 sg13g2_decap_8 FILLER_20_159 ();
 sg13g2_decap_4 FILLER_20_166 ();
 sg13g2_fill_2 FILLER_20_180 ();
 sg13g2_decap_4 FILLER_20_215 ();
 sg13g2_fill_1 FILLER_20_219 ();
 sg13g2_fill_2 FILLER_20_229 ();
 sg13g2_fill_1 FILLER_20_231 ();
 sg13g2_fill_2 FILLER_20_236 ();
 sg13g2_fill_1 FILLER_20_238 ();
 sg13g2_fill_2 FILLER_20_265 ();
 sg13g2_fill_1 FILLER_20_267 ();
 sg13g2_fill_2 FILLER_20_285 ();
 sg13g2_fill_2 FILLER_20_293 ();
 sg13g2_fill_1 FILLER_20_295 ();
 sg13g2_decap_4 FILLER_20_308 ();
 sg13g2_fill_2 FILLER_20_312 ();
 sg13g2_decap_8 FILLER_20_323 ();
 sg13g2_decap_8 FILLER_20_330 ();
 sg13g2_decap_4 FILLER_20_345 ();
 sg13g2_fill_2 FILLER_20_359 ();
 sg13g2_fill_2 FILLER_20_393 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_decap_4 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_410 ();
 sg13g2_fill_1 FILLER_20_419 ();
 sg13g2_fill_2 FILLER_20_450 ();
 sg13g2_fill_1 FILLER_20_452 ();
 sg13g2_fill_1 FILLER_20_479 ();
 sg13g2_fill_1 FILLER_20_484 ();
 sg13g2_fill_1 FILLER_20_491 ();
 sg13g2_fill_1 FILLER_20_503 ();
 sg13g2_fill_1 FILLER_20_542 ();
 sg13g2_fill_1 FILLER_20_569 ();
 sg13g2_fill_1 FILLER_20_599 ();
 sg13g2_fill_1 FILLER_20_677 ();
 sg13g2_fill_1 FILLER_20_704 ();
 sg13g2_decap_4 FILLER_20_731 ();
 sg13g2_fill_1 FILLER_20_735 ();
 sg13g2_fill_1 FILLER_20_741 ();
 sg13g2_fill_1 FILLER_20_747 ();
 sg13g2_fill_2 FILLER_20_765 ();
 sg13g2_fill_2 FILLER_20_775 ();
 sg13g2_decap_8 FILLER_20_811 ();
 sg13g2_decap_8 FILLER_20_818 ();
 sg13g2_decap_8 FILLER_20_825 ();
 sg13g2_decap_4 FILLER_20_832 ();
 sg13g2_fill_1 FILLER_20_846 ();
 sg13g2_fill_1 FILLER_20_898 ();
 sg13g2_decap_4 FILLER_20_909 ();
 sg13g2_decap_4 FILLER_20_959 ();
 sg13g2_fill_2 FILLER_20_999 ();
 sg13g2_fill_1 FILLER_20_1001 ();
 sg13g2_decap_8 FILLER_20_1016 ();
 sg13g2_decap_8 FILLER_20_1027 ();
 sg13g2_fill_2 FILLER_20_1034 ();
 sg13g2_fill_1 FILLER_20_1036 ();
 sg13g2_decap_8 FILLER_20_1042 ();
 sg13g2_decap_4 FILLER_20_1049 ();
 sg13g2_fill_1 FILLER_20_1053 ();
 sg13g2_decap_4 FILLER_20_1059 ();
 sg13g2_fill_2 FILLER_20_1073 ();
 sg13g2_fill_2 FILLER_20_1128 ();
 sg13g2_fill_1 FILLER_20_1130 ();
 sg13g2_fill_2 FILLER_20_1153 ();
 sg13g2_fill_1 FILLER_20_1159 ();
 sg13g2_decap_4 FILLER_20_1172 ();
 sg13g2_fill_2 FILLER_20_1184 ();
 sg13g2_fill_2 FILLER_20_1194 ();
 sg13g2_fill_2 FILLER_20_1232 ();
 sg13g2_fill_1 FILLER_20_1238 ();
 sg13g2_fill_2 FILLER_20_1255 ();
 sg13g2_fill_1 FILLER_20_1309 ();
 sg13g2_fill_1 FILLER_20_1314 ();
 sg13g2_decap_8 FILLER_20_1319 ();
 sg13g2_decap_8 FILLER_20_1326 ();
 sg13g2_decap_4 FILLER_20_1333 ();
 sg13g2_decap_8 FILLER_20_1389 ();
 sg13g2_decap_4 FILLER_20_1396 ();
 sg13g2_fill_2 FILLER_20_1422 ();
 sg13g2_decap_4 FILLER_20_1429 ();
 sg13g2_decap_4 FILLER_20_1439 ();
 sg13g2_fill_2 FILLER_20_1448 ();
 sg13g2_fill_1 FILLER_20_1477 ();
 sg13g2_fill_1 FILLER_20_1489 ();
 sg13g2_fill_2 FILLER_20_1500 ();
 sg13g2_fill_1 FILLER_20_1502 ();
 sg13g2_fill_2 FILLER_20_1514 ();
 sg13g2_fill_1 FILLER_20_1524 ();
 sg13g2_decap_8 FILLER_20_1528 ();
 sg13g2_decap_8 FILLER_20_1535 ();
 sg13g2_fill_2 FILLER_20_1546 ();
 sg13g2_fill_1 FILLER_20_1548 ();
 sg13g2_fill_1 FILLER_20_1559 ();
 sg13g2_fill_2 FILLER_20_1565 ();
 sg13g2_fill_1 FILLER_20_1572 ();
 sg13g2_fill_2 FILLER_20_1583 ();
 sg13g2_fill_1 FILLER_20_1589 ();
 sg13g2_decap_4 FILLER_20_1602 ();
 sg13g2_fill_1 FILLER_20_1614 ();
 sg13g2_fill_1 FILLER_20_1619 ();
 sg13g2_fill_2 FILLER_20_1625 ();
 sg13g2_decap_4 FILLER_20_1637 ();
 sg13g2_fill_2 FILLER_20_1660 ();
 sg13g2_fill_2 FILLER_20_1694 ();
 sg13g2_fill_1 FILLER_20_1696 ();
 sg13g2_decap_4 FILLER_20_1707 ();
 sg13g2_fill_2 FILLER_20_1711 ();
 sg13g2_fill_2 FILLER_20_1723 ();
 sg13g2_decap_8 FILLER_20_1751 ();
 sg13g2_decap_8 FILLER_20_1758 ();
 sg13g2_decap_4 FILLER_20_1765 ();
 sg13g2_fill_1 FILLER_20_1769 ();
 sg13g2_fill_2 FILLER_20_1780 ();
 sg13g2_decap_8 FILLER_20_1808 ();
 sg13g2_fill_1 FILLER_20_1815 ();
 sg13g2_fill_2 FILLER_20_1825 ();
 sg13g2_fill_1 FILLER_20_1827 ();
 sg13g2_fill_1 FILLER_20_1838 ();
 sg13g2_decap_4 FILLER_20_1865 ();
 sg13g2_decap_8 FILLER_20_1878 ();
 sg13g2_decap_4 FILLER_20_1885 ();
 sg13g2_fill_1 FILLER_20_1889 ();
 sg13g2_decap_4 FILLER_20_1923 ();
 sg13g2_fill_2 FILLER_20_1927 ();
 sg13g2_fill_2 FILLER_20_1977 ();
 sg13g2_fill_2 FILLER_20_1991 ();
 sg13g2_fill_1 FILLER_20_1997 ();
 sg13g2_decap_8 FILLER_20_2021 ();
 sg13g2_decap_8 FILLER_20_2028 ();
 sg13g2_decap_8 FILLER_20_2039 ();
 sg13g2_decap_8 FILLER_20_2046 ();
 sg13g2_decap_8 FILLER_20_2053 ();
 sg13g2_decap_4 FILLER_20_2109 ();
 sg13g2_fill_1 FILLER_20_2113 ();
 sg13g2_fill_2 FILLER_20_2166 ();
 sg13g2_fill_2 FILLER_20_2195 ();
 sg13g2_decap_4 FILLER_20_2205 ();
 sg13g2_fill_2 FILLER_20_2209 ();
 sg13g2_fill_2 FILLER_20_2215 ();
 sg13g2_fill_1 FILLER_20_2217 ();
 sg13g2_fill_1 FILLER_20_2228 ();
 sg13g2_fill_2 FILLER_20_2271 ();
 sg13g2_fill_1 FILLER_20_2273 ();
 sg13g2_decap_8 FILLER_20_2277 ();
 sg13g2_fill_2 FILLER_20_2284 ();
 sg13g2_fill_1 FILLER_20_2286 ();
 sg13g2_fill_2 FILLER_20_2300 ();
 sg13g2_fill_1 FILLER_20_2328 ();
 sg13g2_fill_2 FILLER_20_2348 ();
 sg13g2_fill_1 FILLER_20_2360 ();
 sg13g2_fill_1 FILLER_20_2368 ();
 sg13g2_decap_4 FILLER_20_2379 ();
 sg13g2_decap_4 FILLER_20_2387 ();
 sg13g2_fill_1 FILLER_20_2391 ();
 sg13g2_decap_8 FILLER_20_2396 ();
 sg13g2_decap_8 FILLER_20_2403 ();
 sg13g2_fill_2 FILLER_20_2410 ();
 sg13g2_fill_1 FILLER_20_2412 ();
 sg13g2_fill_2 FILLER_20_2422 ();
 sg13g2_fill_1 FILLER_20_2427 ();
 sg13g2_fill_2 FILLER_20_2441 ();
 sg13g2_fill_2 FILLER_20_2473 ();
 sg13g2_fill_2 FILLER_20_2501 ();
 sg13g2_fill_2 FILLER_20_2631 ();
 sg13g2_decap_8 FILLER_20_2659 ();
 sg13g2_decap_4 FILLER_20_2666 ();
 sg13g2_fill_1 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_46 ();
 sg13g2_decap_8 FILLER_21_53 ();
 sg13g2_decap_4 FILLER_21_60 ();
 sg13g2_fill_2 FILLER_21_64 ();
 sg13g2_fill_1 FILLER_21_82 ();
 sg13g2_fill_2 FILLER_21_109 ();
 sg13g2_decap_8 FILLER_21_158 ();
 sg13g2_fill_1 FILLER_21_165 ();
 sg13g2_fill_1 FILLER_21_196 ();
 sg13g2_fill_1 FILLER_21_234 ();
 sg13g2_fill_2 FILLER_21_239 ();
 sg13g2_fill_2 FILLER_21_246 ();
 sg13g2_fill_2 FILLER_21_252 ();
 sg13g2_fill_1 FILLER_21_254 ();
 sg13g2_fill_1 FILLER_21_259 ();
 sg13g2_fill_2 FILLER_21_268 ();
 sg13g2_fill_2 FILLER_21_276 ();
 sg13g2_fill_2 FILLER_21_286 ();
 sg13g2_fill_1 FILLER_21_288 ();
 sg13g2_fill_1 FILLER_21_294 ();
 sg13g2_decap_4 FILLER_21_307 ();
 sg13g2_fill_2 FILLER_21_311 ();
 sg13g2_decap_8 FILLER_21_330 ();
 sg13g2_decap_4 FILLER_21_337 ();
 sg13g2_fill_1 FILLER_21_341 ();
 sg13g2_decap_4 FILLER_21_346 ();
 sg13g2_fill_2 FILLER_21_350 ();
 sg13g2_fill_1 FILLER_21_356 ();
 sg13g2_fill_1 FILLER_21_361 ();
 sg13g2_fill_2 FILLER_21_366 ();
 sg13g2_fill_2 FILLER_21_372 ();
 sg13g2_fill_2 FILLER_21_379 ();
 sg13g2_decap_4 FILLER_21_387 ();
 sg13g2_decap_8 FILLER_21_404 ();
 sg13g2_decap_8 FILLER_21_411 ();
 sg13g2_decap_4 FILLER_21_418 ();
 sg13g2_fill_1 FILLER_21_422 ();
 sg13g2_fill_2 FILLER_21_432 ();
 sg13g2_fill_1 FILLER_21_439 ();
 sg13g2_fill_1 FILLER_21_445 ();
 sg13g2_fill_2 FILLER_21_459 ();
 sg13g2_fill_1 FILLER_21_461 ();
 sg13g2_fill_2 FILLER_21_472 ();
 sg13g2_fill_2 FILLER_21_480 ();
 sg13g2_fill_1 FILLER_21_482 ();
 sg13g2_decap_4 FILLER_21_497 ();
 sg13g2_fill_1 FILLER_21_501 ();
 sg13g2_fill_1 FILLER_21_554 ();
 sg13g2_fill_1 FILLER_21_693 ();
 sg13g2_fill_1 FILLER_21_719 ();
 sg13g2_decap_8 FILLER_21_726 ();
 sg13g2_fill_1 FILLER_21_741 ();
 sg13g2_fill_1 FILLER_21_746 ();
 sg13g2_fill_1 FILLER_21_753 ();
 sg13g2_fill_1 FILLER_21_758 ();
 sg13g2_fill_1 FILLER_21_763 ();
 sg13g2_fill_2 FILLER_21_769 ();
 sg13g2_fill_2 FILLER_21_797 ();
 sg13g2_fill_1 FILLER_21_799 ();
 sg13g2_decap_8 FILLER_21_805 ();
 sg13g2_decap_4 FILLER_21_812 ();
 sg13g2_decap_4 FILLER_21_842 ();
 sg13g2_fill_2 FILLER_21_846 ();
 sg13g2_decap_8 FILLER_21_856 ();
 sg13g2_fill_2 FILLER_21_863 ();
 sg13g2_fill_1 FILLER_21_865 ();
 sg13g2_fill_2 FILLER_21_891 ();
 sg13g2_decap_4 FILLER_21_963 ();
 sg13g2_fill_1 FILLER_21_967 ();
 sg13g2_decap_8 FILLER_21_994 ();
 sg13g2_fill_1 FILLER_21_1001 ();
 sg13g2_fill_2 FILLER_21_1028 ();
 sg13g2_fill_1 FILLER_21_1030 ();
 sg13g2_fill_2 FILLER_21_1041 ();
 sg13g2_fill_2 FILLER_21_1171 ();
 sg13g2_fill_1 FILLER_21_1173 ();
 sg13g2_fill_2 FILLER_21_1214 ();
 sg13g2_fill_1 FILLER_21_1220 ();
 sg13g2_fill_2 FILLER_21_1229 ();
 sg13g2_fill_1 FILLER_21_1239 ();
 sg13g2_fill_1 FILLER_21_1244 ();
 sg13g2_fill_2 FILLER_21_1271 ();
 sg13g2_decap_8 FILLER_21_1334 ();
 sg13g2_decap_8 FILLER_21_1341 ();
 sg13g2_decap_8 FILLER_21_1348 ();
 sg13g2_decap_4 FILLER_21_1355 ();
 sg13g2_fill_2 FILLER_21_1359 ();
 sg13g2_decap_8 FILLER_21_1391 ();
 sg13g2_decap_4 FILLER_21_1398 ();
 sg13g2_decap_4 FILLER_21_1429 ();
 sg13g2_fill_1 FILLER_21_1433 ();
 sg13g2_fill_2 FILLER_21_1439 ();
 sg13g2_fill_2 FILLER_21_1449 ();
 sg13g2_decap_4 FILLER_21_1474 ();
 sg13g2_fill_2 FILLER_21_1491 ();
 sg13g2_decap_8 FILLER_21_1524 ();
 sg13g2_fill_1 FILLER_21_1531 ();
 sg13g2_fill_1 FILLER_21_1576 ();
 sg13g2_fill_1 FILLER_21_1583 ();
 sg13g2_fill_1 FILLER_21_1644 ();
 sg13g2_fill_1 FILLER_21_1650 ();
 sg13g2_fill_2 FILLER_21_1659 ();
 sg13g2_fill_1 FILLER_21_1679 ();
 sg13g2_decap_8 FILLER_21_1696 ();
 sg13g2_decap_4 FILLER_21_1703 ();
 sg13g2_decap_8 FILLER_21_1737 ();
 sg13g2_decap_4 FILLER_21_1744 ();
 sg13g2_fill_1 FILLER_21_1748 ();
 sg13g2_decap_4 FILLER_21_1759 ();
 sg13g2_decap_8 FILLER_21_1767 ();
 sg13g2_fill_2 FILLER_21_1774 ();
 sg13g2_decap_8 FILLER_21_1780 ();
 sg13g2_fill_2 FILLER_21_1787 ();
 sg13g2_decap_8 FILLER_21_1793 ();
 sg13g2_decap_8 FILLER_21_1800 ();
 sg13g2_decap_8 FILLER_21_1807 ();
 sg13g2_decap_8 FILLER_21_1814 ();
 sg13g2_fill_1 FILLER_21_1853 ();
 sg13g2_fill_1 FILLER_21_1868 ();
 sg13g2_fill_2 FILLER_21_1880 ();
 sg13g2_fill_1 FILLER_21_1882 ();
 sg13g2_fill_2 FILLER_21_1887 ();
 sg13g2_fill_1 FILLER_21_1901 ();
 sg13g2_decap_8 FILLER_21_1911 ();
 sg13g2_decap_4 FILLER_21_1918 ();
 sg13g2_fill_1 FILLER_21_1927 ();
 sg13g2_fill_1 FILLER_21_1973 ();
 sg13g2_fill_2 FILLER_21_2007 ();
 sg13g2_fill_2 FILLER_21_2016 ();
 sg13g2_decap_4 FILLER_21_2054 ();
 sg13g2_decap_8 FILLER_21_2084 ();
 sg13g2_decap_4 FILLER_21_2091 ();
 sg13g2_fill_1 FILLER_21_2095 ();
 sg13g2_decap_8 FILLER_21_2135 ();
 sg13g2_fill_2 FILLER_21_2142 ();
 sg13g2_fill_1 FILLER_21_2144 ();
 sg13g2_fill_1 FILLER_21_2149 ();
 sg13g2_fill_2 FILLER_21_2162 ();
 sg13g2_fill_1 FILLER_21_2164 ();
 sg13g2_decap_4 FILLER_21_2211 ();
 sg13g2_decap_4 FILLER_21_2225 ();
 sg13g2_decap_8 FILLER_21_2239 ();
 sg13g2_fill_2 FILLER_21_2246 ();
 sg13g2_fill_1 FILLER_21_2248 ();
 sg13g2_fill_1 FILLER_21_2264 ();
 sg13g2_fill_1 FILLER_21_2273 ();
 sg13g2_fill_2 FILLER_21_2286 ();
 sg13g2_fill_2 FILLER_21_2309 ();
 sg13g2_fill_1 FILLER_21_2311 ();
 sg13g2_fill_2 FILLER_21_2348 ();
 sg13g2_decap_8 FILLER_21_2392 ();
 sg13g2_decap_8 FILLER_21_2399 ();
 sg13g2_fill_1 FILLER_21_2406 ();
 sg13g2_fill_1 FILLER_21_2423 ();
 sg13g2_fill_2 FILLER_21_2430 ();
 sg13g2_fill_1 FILLER_21_2462 ();
 sg13g2_fill_1 FILLER_21_2468 ();
 sg13g2_fill_2 FILLER_21_2482 ();
 sg13g2_fill_2 FILLER_21_2520 ();
 sg13g2_fill_2 FILLER_21_2605 ();
 sg13g2_fill_1 FILLER_21_2632 ();
 sg13g2_decap_8 FILLER_21_2663 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_28 ();
 sg13g2_fill_1 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_54 ();
 sg13g2_decap_4 FILLER_22_61 ();
 sg13g2_fill_1 FILLER_22_65 ();
 sg13g2_fill_2 FILLER_22_125 ();
 sg13g2_decap_4 FILLER_22_167 ();
 sg13g2_fill_2 FILLER_22_171 ();
 sg13g2_fill_1 FILLER_22_232 ();
 sg13g2_fill_1 FILLER_22_237 ();
 sg13g2_fill_1 FILLER_22_264 ();
 sg13g2_fill_2 FILLER_22_291 ();
 sg13g2_fill_2 FILLER_22_344 ();
 sg13g2_fill_2 FILLER_22_350 ();
 sg13g2_fill_1 FILLER_22_377 ();
 sg13g2_decap_8 FILLER_22_412 ();
 sg13g2_decap_4 FILLER_22_419 ();
 sg13g2_fill_1 FILLER_22_423 ();
 sg13g2_decap_8 FILLER_22_432 ();
 sg13g2_decap_4 FILLER_22_439 ();
 sg13g2_decap_4 FILLER_22_453 ();
 sg13g2_decap_8 FILLER_22_466 ();
 sg13g2_decap_8 FILLER_22_473 ();
 sg13g2_decap_8 FILLER_22_480 ();
 sg13g2_decap_8 FILLER_22_487 ();
 sg13g2_decap_8 FILLER_22_494 ();
 sg13g2_decap_8 FILLER_22_501 ();
 sg13g2_decap_4 FILLER_22_508 ();
 sg13g2_fill_1 FILLER_22_527 ();
 sg13g2_fill_2 FILLER_22_604 ();
 sg13g2_fill_2 FILLER_22_632 ();
 sg13g2_fill_2 FILLER_22_654 ();
 sg13g2_decap_4 FILLER_22_705 ();
 sg13g2_fill_1 FILLER_22_709 ();
 sg13g2_fill_2 FILLER_22_770 ();
 sg13g2_fill_1 FILLER_22_785 ();
 sg13g2_fill_2 FILLER_22_791 ();
 sg13g2_fill_1 FILLER_22_814 ();
 sg13g2_decap_8 FILLER_22_855 ();
 sg13g2_decap_8 FILLER_22_862 ();
 sg13g2_decap_8 FILLER_22_869 ();
 sg13g2_decap_8 FILLER_22_905 ();
 sg13g2_fill_2 FILLER_22_912 ();
 sg13g2_decap_8 FILLER_22_961 ();
 sg13g2_decap_4 FILLER_22_968 ();
 sg13g2_fill_2 FILLER_22_972 ();
 sg13g2_fill_2 FILLER_22_978 ();
 sg13g2_fill_1 FILLER_22_980 ();
 sg13g2_decap_4 FILLER_22_985 ();
 sg13g2_decap_8 FILLER_22_1014 ();
 sg13g2_fill_2 FILLER_22_1021 ();
 sg13g2_decap_8 FILLER_22_1083 ();
 sg13g2_fill_2 FILLER_22_1109 ();
 sg13g2_fill_1 FILLER_22_1111 ();
 sg13g2_fill_1 FILLER_22_1164 ();
 sg13g2_fill_1 FILLER_22_1191 ();
 sg13g2_fill_2 FILLER_22_1206 ();
 sg13g2_fill_2 FILLER_22_1249 ();
 sg13g2_fill_1 FILLER_22_1260 ();
 sg13g2_fill_1 FILLER_22_1269 ();
 sg13g2_fill_2 FILLER_22_1275 ();
 sg13g2_decap_8 FILLER_22_1311 ();
 sg13g2_decap_8 FILLER_22_1322 ();
 sg13g2_decap_8 FILLER_22_1329 ();
 sg13g2_decap_4 FILLER_22_1336 ();
 sg13g2_fill_1 FILLER_22_1340 ();
 sg13g2_decap_4 FILLER_22_1377 ();
 sg13g2_fill_2 FILLER_22_1381 ();
 sg13g2_fill_1 FILLER_22_1420 ();
 sg13g2_fill_2 FILLER_22_1437 ();
 sg13g2_fill_1 FILLER_22_1439 ();
 sg13g2_fill_2 FILLER_22_1467 ();
 sg13g2_fill_1 FILLER_22_1469 ();
 sg13g2_fill_2 FILLER_22_1493 ();
 sg13g2_fill_2 FILLER_22_1501 ();
 sg13g2_decap_8 FILLER_22_1509 ();
 sg13g2_fill_1 FILLER_22_1521 ();
 sg13g2_decap_4 FILLER_22_1535 ();
 sg13g2_fill_2 FILLER_22_1539 ();
 sg13g2_fill_1 FILLER_22_1546 ();
 sg13g2_fill_1 FILLER_22_1566 ();
 sg13g2_decap_8 FILLER_22_1580 ();
 sg13g2_decap_4 FILLER_22_1597 ();
 sg13g2_fill_2 FILLER_22_1609 ();
 sg13g2_fill_1 FILLER_22_1618 ();
 sg13g2_fill_1 FILLER_22_1629 ();
 sg13g2_fill_2 FILLER_22_1725 ();
 sg13g2_decap_8 FILLER_22_1731 ();
 sg13g2_decap_8 FILLER_22_1738 ();
 sg13g2_decap_8 FILLER_22_1745 ();
 sg13g2_fill_1 FILLER_22_1752 ();
 sg13g2_decap_8 FILLER_22_1783 ();
 sg13g2_decap_8 FILLER_22_1790 ();
 sg13g2_fill_1 FILLER_22_1797 ();
 sg13g2_fill_2 FILLER_22_1802 ();
 sg13g2_fill_1 FILLER_22_1804 ();
 sg13g2_fill_2 FILLER_22_1809 ();
 sg13g2_fill_1 FILLER_22_1811 ();
 sg13g2_fill_1 FILLER_22_1817 ();
 sg13g2_decap_4 FILLER_22_1836 ();
 sg13g2_decap_4 FILLER_22_1871 ();
 sg13g2_fill_1 FILLER_22_1875 ();
 sg13g2_fill_2 FILLER_22_1888 ();
 sg13g2_fill_2 FILLER_22_1920 ();
 sg13g2_fill_2 FILLER_22_1930 ();
 sg13g2_fill_1 FILLER_22_2012 ();
 sg13g2_decap_8 FILLER_22_2025 ();
 sg13g2_decap_4 FILLER_22_2060 ();
 sg13g2_decap_8 FILLER_22_2068 ();
 sg13g2_decap_8 FILLER_22_2075 ();
 sg13g2_decap_4 FILLER_22_2082 ();
 sg13g2_fill_1 FILLER_22_2086 ();
 sg13g2_decap_8 FILLER_22_2091 ();
 sg13g2_decap_4 FILLER_22_2098 ();
 sg13g2_fill_1 FILLER_22_2102 ();
 sg13g2_decap_4 FILLER_22_2131 ();
 sg13g2_fill_2 FILLER_22_2135 ();
 sg13g2_fill_2 FILLER_22_2142 ();
 sg13g2_fill_1 FILLER_22_2144 ();
 sg13g2_fill_2 FILLER_22_2159 ();
 sg13g2_fill_2 FILLER_22_2182 ();
 sg13g2_fill_1 FILLER_22_2224 ();
 sg13g2_fill_1 FILLER_22_2251 ();
 sg13g2_fill_1 FILLER_22_2310 ();
 sg13g2_decap_8 FILLER_22_2316 ();
 sg13g2_fill_2 FILLER_22_2327 ();
 sg13g2_fill_1 FILLER_22_2506 ();
 sg13g2_fill_1 FILLER_22_2514 ();
 sg13g2_fill_2 FILLER_22_2567 ();
 sg13g2_fill_1 FILLER_22_2583 ();
 sg13g2_decap_8 FILLER_22_2623 ();
 sg13g2_fill_2 FILLER_22_2640 ();
 sg13g2_fill_1 FILLER_22_2642 ();
 sg13g2_fill_1 FILLER_22_2647 ();
 sg13g2_decap_8 FILLER_22_2652 ();
 sg13g2_decap_8 FILLER_22_2659 ();
 sg13g2_decap_4 FILLER_22_2666 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_13 ();
 sg13g2_decap_8 FILLER_23_20 ();
 sg13g2_fill_2 FILLER_23_27 ();
 sg13g2_fill_2 FILLER_23_33 ();
 sg13g2_decap_4 FILLER_23_41 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_fill_2 FILLER_23_63 ();
 sg13g2_fill_1 FILLER_23_65 ();
 sg13g2_decap_4 FILLER_23_128 ();
 sg13g2_fill_1 FILLER_23_132 ();
 sg13g2_decap_4 FILLER_23_137 ();
 sg13g2_decap_8 FILLER_23_155 ();
 sg13g2_decap_4 FILLER_23_162 ();
 sg13g2_decap_8 FILLER_23_171 ();
 sg13g2_fill_1 FILLER_23_178 ();
 sg13g2_fill_2 FILLER_23_214 ();
 sg13g2_decap_8 FILLER_23_230 ();
 sg13g2_decap_8 FILLER_23_237 ();
 sg13g2_decap_4 FILLER_23_248 ();
 sg13g2_fill_1 FILLER_23_257 ();
 sg13g2_fill_1 FILLER_23_270 ();
 sg13g2_fill_2 FILLER_23_298 ();
 sg13g2_fill_1 FILLER_23_300 ();
 sg13g2_fill_1 FILLER_23_350 ();
 sg13g2_fill_1 FILLER_23_356 ();
 sg13g2_decap_4 FILLER_23_383 ();
 sg13g2_fill_2 FILLER_23_391 ();
 sg13g2_decap_8 FILLER_23_397 ();
 sg13g2_decap_8 FILLER_23_404 ();
 sg13g2_decap_4 FILLER_23_411 ();
 sg13g2_fill_2 FILLER_23_415 ();
 sg13g2_fill_2 FILLER_23_443 ();
 sg13g2_fill_2 FILLER_23_449 ();
 sg13g2_fill_2 FILLER_23_457 ();
 sg13g2_decap_4 FILLER_23_494 ();
 sg13g2_fill_2 FILLER_23_504 ();
 sg13g2_fill_1 FILLER_23_506 ();
 sg13g2_decap_4 FILLER_23_513 ();
 sg13g2_fill_1 FILLER_23_521 ();
 sg13g2_fill_2 FILLER_23_527 ();
 sg13g2_fill_1 FILLER_23_547 ();
 sg13g2_fill_1 FILLER_23_592 ();
 sg13g2_fill_2 FILLER_23_599 ();
 sg13g2_fill_1 FILLER_23_610 ();
 sg13g2_fill_1 FILLER_23_628 ();
 sg13g2_fill_2 FILLER_23_663 ();
 sg13g2_decap_4 FILLER_23_691 ();
 sg13g2_fill_2 FILLER_23_695 ();
 sg13g2_fill_1 FILLER_23_701 ();
 sg13g2_fill_2 FILLER_23_733 ();
 sg13g2_fill_2 FILLER_23_749 ();
 sg13g2_fill_1 FILLER_23_756 ();
 sg13g2_fill_2 FILLER_23_761 ();
 sg13g2_decap_4 FILLER_23_814 ();
 sg13g2_fill_2 FILLER_23_818 ();
 sg13g2_decap_4 FILLER_23_858 ();
 sg13g2_fill_1 FILLER_23_862 ();
 sg13g2_decap_8 FILLER_23_889 ();
 sg13g2_decap_4 FILLER_23_896 ();
 sg13g2_fill_2 FILLER_23_900 ();
 sg13g2_fill_2 FILLER_23_944 ();
 sg13g2_fill_2 FILLER_23_977 ();
 sg13g2_fill_1 FILLER_23_979 ();
 sg13g2_decap_8 FILLER_23_1005 ();
 sg13g2_decap_8 FILLER_23_1012 ();
 sg13g2_decap_4 FILLER_23_1019 ();
 sg13g2_decap_8 FILLER_23_1036 ();
 sg13g2_decap_8 FILLER_23_1043 ();
 sg13g2_decap_4 FILLER_23_1050 ();
 sg13g2_decap_4 FILLER_23_1064 ();
 sg13g2_fill_1 FILLER_23_1068 ();
 sg13g2_decap_8 FILLER_23_1086 ();
 sg13g2_fill_1 FILLER_23_1093 ();
 sg13g2_decap_8 FILLER_23_1098 ();
 sg13g2_decap_8 FILLER_23_1105 ();
 sg13g2_fill_2 FILLER_23_1112 ();
 sg13g2_decap_8 FILLER_23_1124 ();
 sg13g2_decap_8 FILLER_23_1131 ();
 sg13g2_fill_2 FILLER_23_1138 ();
 sg13g2_decap_8 FILLER_23_1148 ();
 sg13g2_fill_1 FILLER_23_1165 ();
 sg13g2_fill_1 FILLER_23_1239 ();
 sg13g2_fill_1 FILLER_23_1255 ();
 sg13g2_fill_1 FILLER_23_1295 ();
 sg13g2_fill_1 FILLER_23_1300 ();
 sg13g2_decap_4 FILLER_23_1373 ();
 sg13g2_decap_4 FILLER_23_1413 ();
 sg13g2_fill_1 FILLER_23_1417 ();
 sg13g2_fill_2 FILLER_23_1431 ();
 sg13g2_fill_2 FILLER_23_1452 ();
 sg13g2_fill_1 FILLER_23_1454 ();
 sg13g2_fill_1 FILLER_23_1480 ();
 sg13g2_fill_2 FILLER_23_1493 ();
 sg13g2_fill_1 FILLER_23_1495 ();
 sg13g2_fill_2 FILLER_23_1505 ();
 sg13g2_fill_1 FILLER_23_1507 ();
 sg13g2_fill_1 FILLER_23_1513 ();
 sg13g2_decap_4 FILLER_23_1534 ();
 sg13g2_decap_4 FILLER_23_1578 ();
 sg13g2_fill_1 FILLER_23_1582 ();
 sg13g2_decap_8 FILLER_23_1589 ();
 sg13g2_fill_2 FILLER_23_1632 ();
 sg13g2_fill_1 FILLER_23_1634 ();
 sg13g2_decap_4 FILLER_23_1641 ();
 sg13g2_fill_1 FILLER_23_1645 ();
 sg13g2_fill_2 FILLER_23_1650 ();
 sg13g2_fill_1 FILLER_23_1666 ();
 sg13g2_fill_1 FILLER_23_1671 ();
 sg13g2_decap_4 FILLER_23_1678 ();
 sg13g2_fill_1 FILLER_23_1682 ();
 sg13g2_fill_2 FILLER_23_1686 ();
 sg13g2_fill_1 FILLER_23_1688 ();
 sg13g2_decap_4 FILLER_23_1738 ();
 sg13g2_fill_1 FILLER_23_1848 ();
 sg13g2_fill_2 FILLER_23_1854 ();
 sg13g2_decap_4 FILLER_23_1868 ();
 sg13g2_fill_1 FILLER_23_1872 ();
 sg13g2_fill_2 FILLER_23_1899 ();
 sg13g2_fill_1 FILLER_23_1901 ();
 sg13g2_fill_1 FILLER_23_1916 ();
 sg13g2_fill_2 FILLER_23_1931 ();
 sg13g2_fill_2 FILLER_23_1983 ();
 sg13g2_fill_2 FILLER_23_1995 ();
 sg13g2_fill_2 FILLER_23_2005 ();
 sg13g2_fill_2 FILLER_23_2041 ();
 sg13g2_fill_1 FILLER_23_2043 ();
 sg13g2_decap_4 FILLER_23_2070 ();
 sg13g2_fill_1 FILLER_23_2074 ();
 sg13g2_decap_4 FILLER_23_2096 ();
 sg13g2_fill_1 FILLER_23_2100 ();
 sg13g2_fill_1 FILLER_23_2115 ();
 sg13g2_decap_8 FILLER_23_2124 ();
 sg13g2_fill_2 FILLER_23_2131 ();
 sg13g2_decap_4 FILLER_23_2143 ();
 sg13g2_decap_8 FILLER_23_2199 ();
 sg13g2_decap_4 FILLER_23_2250 ();
 sg13g2_fill_1 FILLER_23_2254 ();
 sg13g2_decap_4 FILLER_23_2275 ();
 sg13g2_fill_1 FILLER_23_2279 ();
 sg13g2_decap_8 FILLER_23_2316 ();
 sg13g2_decap_4 FILLER_23_2328 ();
 sg13g2_fill_2 FILLER_23_2332 ();
 sg13g2_fill_2 FILLER_23_2360 ();
 sg13g2_fill_2 FILLER_23_2375 ();
 sg13g2_fill_2 FILLER_23_2382 ();
 sg13g2_fill_2 FILLER_23_2414 ();
 sg13g2_fill_1 FILLER_23_2419 ();
 sg13g2_fill_2 FILLER_23_2527 ();
 sg13g2_fill_1 FILLER_23_2533 ();
 sg13g2_fill_1 FILLER_23_2579 ();
 sg13g2_decap_4 FILLER_23_2619 ();
 sg13g2_fill_1 FILLER_23_2623 ();
 sg13g2_fill_2 FILLER_23_2660 ();
 sg13g2_decap_4 FILLER_23_2666 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_7 ();
 sg13g2_fill_1 FILLER_24_9 ();
 sg13g2_fill_1 FILLER_24_24 ();
 sg13g2_fill_2 FILLER_24_43 ();
 sg13g2_fill_1 FILLER_24_45 ();
 sg13g2_decap_4 FILLER_24_50 ();
 sg13g2_fill_1 FILLER_24_93 ();
 sg13g2_fill_1 FILLER_24_137 ();
 sg13g2_decap_4 FILLER_24_143 ();
 sg13g2_decap_8 FILLER_24_157 ();
 sg13g2_decap_8 FILLER_24_164 ();
 sg13g2_decap_8 FILLER_24_171 ();
 sg13g2_decap_8 FILLER_24_178 ();
 sg13g2_decap_4 FILLER_24_185 ();
 sg13g2_fill_1 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_194 ();
 sg13g2_fill_2 FILLER_24_201 ();
 sg13g2_fill_1 FILLER_24_203 ();
 sg13g2_fill_2 FILLER_24_212 ();
 sg13g2_fill_1 FILLER_24_214 ();
 sg13g2_decap_4 FILLER_24_220 ();
 sg13g2_fill_1 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_235 ();
 sg13g2_fill_1 FILLER_24_242 ();
 sg13g2_decap_4 FILLER_24_252 ();
 sg13g2_fill_2 FILLER_24_261 ();
 sg13g2_fill_1 FILLER_24_263 ();
 sg13g2_fill_2 FILLER_24_281 ();
 sg13g2_decap_4 FILLER_24_316 ();
 sg13g2_fill_2 FILLER_24_328 ();
 sg13g2_fill_1 FILLER_24_330 ();
 sg13g2_decap_8 FILLER_24_335 ();
 sg13g2_decap_8 FILLER_24_342 ();
 sg13g2_decap_8 FILLER_24_349 ();
 sg13g2_decap_4 FILLER_24_356 ();
 sg13g2_fill_2 FILLER_24_364 ();
 sg13g2_decap_4 FILLER_24_370 ();
 sg13g2_decap_8 FILLER_24_404 ();
 sg13g2_fill_2 FILLER_24_411 ();
 sg13g2_fill_1 FILLER_24_474 ();
 sg13g2_decap_8 FILLER_24_506 ();
 sg13g2_decap_4 FILLER_24_513 ();
 sg13g2_fill_2 FILLER_24_517 ();
 sg13g2_fill_2 FILLER_24_524 ();
 sg13g2_fill_1 FILLER_24_526 ();
 sg13g2_fill_2 FILLER_24_532 ();
 sg13g2_fill_1 FILLER_24_539 ();
 sg13g2_fill_1 FILLER_24_577 ();
 sg13g2_fill_1 FILLER_24_586 ();
 sg13g2_fill_2 FILLER_24_593 ();
 sg13g2_fill_2 FILLER_24_603 ();
 sg13g2_fill_1 FILLER_24_605 ();
 sg13g2_fill_1 FILLER_24_642 ();
 sg13g2_fill_1 FILLER_24_651 ();
 sg13g2_fill_2 FILLER_24_656 ();
 sg13g2_fill_1 FILLER_24_661 ();
 sg13g2_decap_8 FILLER_24_681 ();
 sg13g2_fill_1 FILLER_24_688 ();
 sg13g2_decap_4 FILLER_24_743 ();
 sg13g2_fill_1 FILLER_24_747 ();
 sg13g2_decap_8 FILLER_24_752 ();
 sg13g2_decap_8 FILLER_24_759 ();
 sg13g2_decap_8 FILLER_24_766 ();
 sg13g2_fill_2 FILLER_24_773 ();
 sg13g2_fill_1 FILLER_24_788 ();
 sg13g2_decap_8 FILLER_24_815 ();
 sg13g2_fill_1 FILLER_24_822 ();
 sg13g2_fill_1 FILLER_24_854 ();
 sg13g2_fill_2 FILLER_24_957 ();
 sg13g2_fill_1 FILLER_24_995 ();
 sg13g2_decap_8 FILLER_24_1006 ();
 sg13g2_decap_8 FILLER_24_1013 ();
 sg13g2_decap_4 FILLER_24_1020 ();
 sg13g2_fill_1 FILLER_24_1024 ();
 sg13g2_decap_4 FILLER_24_1061 ();
 sg13g2_fill_1 FILLER_24_1101 ();
 sg13g2_decap_8 FILLER_24_1112 ();
 sg13g2_decap_8 FILLER_24_1119 ();
 sg13g2_decap_4 FILLER_24_1126 ();
 sg13g2_fill_2 FILLER_24_1130 ();
 sg13g2_decap_8 FILLER_24_1142 ();
 sg13g2_decap_8 FILLER_24_1149 ();
 sg13g2_decap_8 FILLER_24_1156 ();
 sg13g2_fill_2 FILLER_24_1163 ();
 sg13g2_fill_2 FILLER_24_1170 ();
 sg13g2_fill_2 FILLER_24_1192 ();
 sg13g2_fill_1 FILLER_24_1220 ();
 sg13g2_fill_2 FILLER_24_1251 ();
 sg13g2_fill_2 FILLER_24_1291 ();
 sg13g2_fill_2 FILLER_24_1298 ();
 sg13g2_fill_2 FILLER_24_1336 ();
 sg13g2_fill_2 FILLER_24_1348 ();
 sg13g2_fill_1 FILLER_24_1350 ();
 sg13g2_fill_1 FILLER_24_1355 ();
 sg13g2_decap_8 FILLER_24_1360 ();
 sg13g2_fill_2 FILLER_24_1367 ();
 sg13g2_decap_8 FILLER_24_1374 ();
 sg13g2_decap_4 FILLER_24_1398 ();
 sg13g2_fill_2 FILLER_24_1402 ();
 sg13g2_fill_2 FILLER_24_1413 ();
 sg13g2_fill_2 FILLER_24_1420 ();
 sg13g2_fill_1 FILLER_24_1432 ();
 sg13g2_fill_2 FILLER_24_1439 ();
 sg13g2_fill_1 FILLER_24_1446 ();
 sg13g2_fill_1 FILLER_24_1456 ();
 sg13g2_decap_4 FILLER_24_1493 ();
 sg13g2_fill_2 FILLER_24_1509 ();
 sg13g2_fill_1 FILLER_24_1524 ();
 sg13g2_decap_4 FILLER_24_1530 ();
 sg13g2_fill_2 FILLER_24_1534 ();
 sg13g2_fill_1 FILLER_24_1551 ();
 sg13g2_fill_1 FILLER_24_1557 ();
 sg13g2_fill_1 FILLER_24_1568 ();
 sg13g2_fill_1 FILLER_24_1574 ();
 sg13g2_fill_2 FILLER_24_1581 ();
 sg13g2_fill_1 FILLER_24_1583 ();
 sg13g2_fill_2 FILLER_24_1588 ();
 sg13g2_fill_1 FILLER_24_1590 ();
 sg13g2_fill_2 FILLER_24_1613 ();
 sg13g2_decap_4 FILLER_24_1621 ();
 sg13g2_fill_2 FILLER_24_1625 ();
 sg13g2_fill_1 FILLER_24_1635 ();
 sg13g2_fill_1 FILLER_24_1670 ();
 sg13g2_fill_1 FILLER_24_1676 ();
 sg13g2_fill_2 FILLER_24_1696 ();
 sg13g2_fill_1 FILLER_24_1698 ();
 sg13g2_decap_8 FILLER_24_1761 ();
 sg13g2_fill_1 FILLER_24_1768 ();
 sg13g2_fill_2 FILLER_24_1809 ();
 sg13g2_fill_1 FILLER_24_1811 ();
 sg13g2_fill_2 FILLER_24_1838 ();
 sg13g2_fill_2 FILLER_24_1850 ();
 sg13g2_fill_2 FILLER_24_1856 ();
 sg13g2_fill_1 FILLER_24_1863 ();
 sg13g2_fill_1 FILLER_24_1869 ();
 sg13g2_fill_2 FILLER_24_1879 ();
 sg13g2_fill_2 FILLER_24_1888 ();
 sg13g2_fill_2 FILLER_24_1911 ();
 sg13g2_fill_1 FILLER_24_1923 ();
 sg13g2_fill_1 FILLER_24_1929 ();
 sg13g2_fill_1 FILLER_24_1935 ();
 sg13g2_fill_1 FILLER_24_1953 ();
 sg13g2_fill_2 FILLER_24_1984 ();
 sg13g2_fill_1 FILLER_24_2052 ();
 sg13g2_fill_1 FILLER_24_2073 ();
 sg13g2_fill_2 FILLER_24_2100 ();
 sg13g2_fill_2 FILLER_24_2179 ();
 sg13g2_fill_2 FILLER_24_2212 ();
 sg13g2_fill_2 FILLER_24_2250 ();
 sg13g2_fill_1 FILLER_24_2357 ();
 sg13g2_fill_2 FILLER_24_2408 ();
 sg13g2_fill_1 FILLER_24_2423 ();
 sg13g2_decap_4 FILLER_24_2463 ();
 sg13g2_fill_1 FILLER_24_2467 ();
 sg13g2_fill_1 FILLER_24_2515 ();
 sg13g2_fill_1 FILLER_24_2529 ();
 sg13g2_decap_8 FILLER_24_2663 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_33 ();
 sg13g2_decap_8 FILLER_25_47 ();
 sg13g2_decap_4 FILLER_25_54 ();
 sg13g2_fill_1 FILLER_25_58 ();
 sg13g2_fill_1 FILLER_25_63 ();
 sg13g2_fill_1 FILLER_25_68 ();
 sg13g2_fill_1 FILLER_25_79 ();
 sg13g2_fill_1 FILLER_25_90 ();
 sg13g2_fill_2 FILLER_25_119 ();
 sg13g2_fill_1 FILLER_25_121 ();
 sg13g2_fill_2 FILLER_25_135 ();
 sg13g2_decap_8 FILLER_25_167 ();
 sg13g2_decap_8 FILLER_25_174 ();
 sg13g2_decap_8 FILLER_25_181 ();
 sg13g2_decap_8 FILLER_25_188 ();
 sg13g2_decap_4 FILLER_25_195 ();
 sg13g2_fill_2 FILLER_25_259 ();
 sg13g2_fill_1 FILLER_25_261 ();
 sg13g2_decap_4 FILLER_25_286 ();
 sg13g2_fill_1 FILLER_25_323 ();
 sg13g2_decap_8 FILLER_25_338 ();
 sg13g2_fill_2 FILLER_25_345 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_decap_4 FILLER_25_406 ();
 sg13g2_fill_2 FILLER_25_410 ();
 sg13g2_fill_1 FILLER_25_436 ();
 sg13g2_fill_1 FILLER_25_474 ();
 sg13g2_fill_2 FILLER_25_541 ();
 sg13g2_fill_1 FILLER_25_577 ();
 sg13g2_fill_1 FILLER_25_583 ();
 sg13g2_fill_1 FILLER_25_588 ();
 sg13g2_fill_1 FILLER_25_594 ();
 sg13g2_fill_1 FILLER_25_600 ();
 sg13g2_fill_1 FILLER_25_627 ();
 sg13g2_decap_8 FILLER_25_641 ();
 sg13g2_decap_4 FILLER_25_648 ();
 sg13g2_fill_2 FILLER_25_652 ();
 sg13g2_fill_2 FILLER_25_659 ();
 sg13g2_decap_8 FILLER_25_669 ();
 sg13g2_decap_8 FILLER_25_676 ();
 sg13g2_fill_1 FILLER_25_697 ();
 sg13g2_fill_1 FILLER_25_707 ();
 sg13g2_decap_4 FILLER_25_722 ();
 sg13g2_fill_1 FILLER_25_731 ();
 sg13g2_fill_1 FILLER_25_775 ();
 sg13g2_fill_2 FILLER_25_788 ();
 sg13g2_fill_1 FILLER_25_795 ();
 sg13g2_fill_2 FILLER_25_800 ();
 sg13g2_fill_1 FILLER_25_802 ();
 sg13g2_fill_1 FILLER_25_808 ();
 sg13g2_fill_2 FILLER_25_814 ();
 sg13g2_fill_1 FILLER_25_816 ();
 sg13g2_fill_2 FILLER_25_847 ();
 sg13g2_fill_1 FILLER_25_849 ();
 sg13g2_fill_2 FILLER_25_854 ();
 sg13g2_fill_1 FILLER_25_856 ();
 sg13g2_decap_4 FILLER_25_881 ();
 sg13g2_fill_1 FILLER_25_885 ();
 sg13g2_fill_1 FILLER_25_926 ();
 sg13g2_fill_1 FILLER_25_941 ();
 sg13g2_fill_2 FILLER_25_952 ();
 sg13g2_fill_2 FILLER_25_964 ();
 sg13g2_fill_2 FILLER_25_970 ();
 sg13g2_fill_1 FILLER_25_972 ();
 sg13g2_fill_1 FILLER_25_1072 ();
 sg13g2_decap_4 FILLER_25_1120 ();
 sg13g2_fill_2 FILLER_25_1124 ();
 sg13g2_decap_8 FILLER_25_1156 ();
 sg13g2_decap_4 FILLER_25_1163 ();
 sg13g2_fill_1 FILLER_25_1167 ();
 sg13g2_fill_2 FILLER_25_1209 ();
 sg13g2_fill_2 FILLER_25_1221 ();
 sg13g2_fill_1 FILLER_25_1223 ();
 sg13g2_fill_1 FILLER_25_1228 ();
 sg13g2_fill_1 FILLER_25_1266 ();
 sg13g2_fill_2 FILLER_25_1278 ();
 sg13g2_fill_2 FILLER_25_1319 ();
 sg13g2_decap_8 FILLER_25_1325 ();
 sg13g2_decap_4 FILLER_25_1332 ();
 sg13g2_fill_1 FILLER_25_1336 ();
 sg13g2_decap_8 FILLER_25_1347 ();
 sg13g2_decap_8 FILLER_25_1354 ();
 sg13g2_decap_4 FILLER_25_1361 ();
 sg13g2_decap_4 FILLER_25_1405 ();
 sg13g2_decap_4 FILLER_25_1423 ();
 sg13g2_fill_2 FILLER_25_1427 ();
 sg13g2_decap_4 FILLER_25_1435 ();
 sg13g2_fill_2 FILLER_25_1474 ();
 sg13g2_decap_4 FILLER_25_1500 ();
 sg13g2_fill_1 FILLER_25_1504 ();
 sg13g2_fill_2 FILLER_25_1515 ();
 sg13g2_fill_1 FILLER_25_1517 ();
 sg13g2_decap_8 FILLER_25_1523 ();
 sg13g2_fill_1 FILLER_25_1530 ();
 sg13g2_fill_1 FILLER_25_1536 ();
 sg13g2_fill_2 FILLER_25_1543 ();
 sg13g2_fill_1 FILLER_25_1545 ();
 sg13g2_fill_1 FILLER_25_1552 ();
 sg13g2_decap_4 FILLER_25_1580 ();
 sg13g2_decap_8 FILLER_25_1588 ();
 sg13g2_decap_4 FILLER_25_1599 ();
 sg13g2_fill_2 FILLER_25_1603 ();
 sg13g2_decap_4 FILLER_25_1610 ();
 sg13g2_fill_2 FILLER_25_1614 ();
 sg13g2_fill_1 FILLER_25_1646 ();
 sg13g2_fill_1 FILLER_25_1669 ();
 sg13g2_decap_8 FILLER_25_1765 ();
 sg13g2_fill_1 FILLER_25_1772 ();
 sg13g2_decap_8 FILLER_25_1809 ();
 sg13g2_fill_2 FILLER_25_1816 ();
 sg13g2_fill_1 FILLER_25_1818 ();
 sg13g2_decap_8 FILLER_25_1823 ();
 sg13g2_fill_2 FILLER_25_1830 ();
 sg13g2_decap_8 FILLER_25_1841 ();
 sg13g2_fill_2 FILLER_25_1848 ();
 sg13g2_fill_1 FILLER_25_1850 ();
 sg13g2_fill_2 FILLER_25_1876 ();
 sg13g2_fill_2 FILLER_25_1884 ();
 sg13g2_fill_1 FILLER_25_1929 ();
 sg13g2_fill_2 FILLER_25_1939 ();
 sg13g2_fill_2 FILLER_25_1953 ();
 sg13g2_fill_1 FILLER_25_1962 ();
 sg13g2_fill_1 FILLER_25_1976 ();
 sg13g2_fill_2 FILLER_25_1980 ();
 sg13g2_decap_8 FILLER_25_2031 ();
 sg13g2_decap_8 FILLER_25_2038 ();
 sg13g2_decap_4 FILLER_25_2045 ();
 sg13g2_fill_2 FILLER_25_2059 ();
 sg13g2_fill_2 FILLER_25_2100 ();
 sg13g2_fill_2 FILLER_25_2128 ();
 sg13g2_fill_2 FILLER_25_2134 ();
 sg13g2_fill_1 FILLER_25_2136 ();
 sg13g2_decap_4 FILLER_25_2185 ();
 sg13g2_decap_4 FILLER_25_2206 ();
 sg13g2_fill_1 FILLER_25_2210 ();
 sg13g2_fill_2 FILLER_25_2247 ();
 sg13g2_fill_1 FILLER_25_2249 ();
 sg13g2_fill_1 FILLER_25_2264 ();
 sg13g2_fill_1 FILLER_25_2291 ();
 sg13g2_fill_2 FILLER_25_2347 ();
 sg13g2_fill_2 FILLER_25_2425 ();
 sg13g2_decap_4 FILLER_25_2451 ();
 sg13g2_decap_4 FILLER_25_2460 ();
 sg13g2_fill_1 FILLER_25_2464 ();
 sg13g2_decap_4 FILLER_25_2504 ();
 sg13g2_fill_2 FILLER_25_2544 ();
 sg13g2_decap_4 FILLER_25_2628 ();
 sg13g2_decap_8 FILLER_25_2658 ();
 sg13g2_decap_4 FILLER_25_2665 ();
 sg13g2_fill_1 FILLER_25_2669 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_4 FILLER_26_7 ();
 sg13g2_fill_1 FILLER_26_11 ();
 sg13g2_fill_2 FILLER_26_21 ();
 sg13g2_fill_1 FILLER_26_36 ();
 sg13g2_fill_1 FILLER_26_46 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_fill_2 FILLER_26_63 ();
 sg13g2_fill_1 FILLER_26_65 ();
 sg13g2_fill_1 FILLER_26_79 ();
 sg13g2_fill_1 FILLER_26_85 ();
 sg13g2_fill_2 FILLER_26_122 ();
 sg13g2_fill_2 FILLER_26_135 ();
 sg13g2_fill_1 FILLER_26_137 ();
 sg13g2_decap_8 FILLER_26_141 ();
 sg13g2_fill_2 FILLER_26_148 ();
 sg13g2_fill_2 FILLER_26_160 ();
 sg13g2_decap_4 FILLER_26_188 ();
 sg13g2_fill_1 FILLER_26_252 ();
 sg13g2_fill_2 FILLER_26_262 ();
 sg13g2_fill_1 FILLER_26_264 ();
 sg13g2_fill_2 FILLER_26_311 ();
 sg13g2_fill_2 FILLER_26_321 ();
 sg13g2_decap_8 FILLER_26_335 ();
 sg13g2_decap_8 FILLER_26_342 ();
 sg13g2_decap_4 FILLER_26_349 ();
 sg13g2_fill_2 FILLER_26_353 ();
 sg13g2_decap_4 FILLER_26_399 ();
 sg13g2_decap_4 FILLER_26_407 ();
 sg13g2_fill_1 FILLER_26_411 ();
 sg13g2_fill_2 FILLER_26_487 ();
 sg13g2_fill_1 FILLER_26_549 ();
 sg13g2_fill_1 FILLER_26_560 ();
 sg13g2_fill_1 FILLER_26_568 ();
 sg13g2_fill_1 FILLER_26_574 ();
 sg13g2_fill_2 FILLER_26_600 ();
 sg13g2_fill_1 FILLER_26_602 ();
 sg13g2_fill_1 FILLER_26_627 ();
 sg13g2_fill_1 FILLER_26_632 ();
 sg13g2_fill_1 FILLER_26_685 ();
 sg13g2_fill_2 FILLER_26_716 ();
 sg13g2_fill_1 FILLER_26_718 ();
 sg13g2_decap_8 FILLER_26_724 ();
 sg13g2_decap_4 FILLER_26_789 ();
 sg13g2_fill_2 FILLER_26_823 ();
 sg13g2_decap_4 FILLER_26_839 ();
 sg13g2_fill_2 FILLER_26_853 ();
 sg13g2_fill_1 FILLER_26_855 ();
 sg13g2_decap_8 FILLER_26_896 ();
 sg13g2_decap_8 FILLER_26_903 ();
 sg13g2_decap_8 FILLER_26_910 ();
 sg13g2_decap_8 FILLER_26_917 ();
 sg13g2_fill_1 FILLER_26_924 ();
 sg13g2_decap_8 FILLER_26_938 ();
 sg13g2_decap_8 FILLER_26_945 ();
 sg13g2_decap_8 FILLER_26_952 ();
 sg13g2_decap_8 FILLER_26_959 ();
 sg13g2_decap_8 FILLER_26_966 ();
 sg13g2_fill_1 FILLER_26_973 ();
 sg13g2_fill_1 FILLER_26_1019 ();
 sg13g2_decap_4 FILLER_26_1096 ();
 sg13g2_fill_1 FILLER_26_1100 ();
 sg13g2_fill_1 FILLER_26_1127 ();
 sg13g2_decap_4 FILLER_26_1179 ();
 sg13g2_decap_8 FILLER_26_1199 ();
 sg13g2_decap_8 FILLER_26_1206 ();
 sg13g2_decap_8 FILLER_26_1213 ();
 sg13g2_decap_8 FILLER_26_1220 ();
 sg13g2_decap_4 FILLER_26_1227 ();
 sg13g2_fill_1 FILLER_26_1231 ();
 sg13g2_fill_2 FILLER_26_1242 ();
 sg13g2_fill_1 FILLER_26_1244 ();
 sg13g2_fill_1 FILLER_26_1253 ();
 sg13g2_fill_2 FILLER_26_1284 ();
 sg13g2_decap_8 FILLER_26_1290 ();
 sg13g2_decap_4 FILLER_26_1297 ();
 sg13g2_fill_1 FILLER_26_1301 ();
 sg13g2_decap_4 FILLER_26_1309 ();
 sg13g2_fill_2 FILLER_26_1313 ();
 sg13g2_fill_1 FILLER_26_1320 ();
 sg13g2_decap_8 FILLER_26_1355 ();
 sg13g2_decap_8 FILLER_26_1362 ();
 sg13g2_decap_4 FILLER_26_1369 ();
 sg13g2_fill_2 FILLER_26_1373 ();
 sg13g2_decap_8 FILLER_26_1379 ();
 sg13g2_fill_1 FILLER_26_1386 ();
 sg13g2_decap_8 FILLER_26_1403 ();
 sg13g2_decap_8 FILLER_26_1410 ();
 sg13g2_decap_4 FILLER_26_1417 ();
 sg13g2_fill_1 FILLER_26_1421 ();
 sg13g2_fill_2 FILLER_26_1445 ();
 sg13g2_fill_1 FILLER_26_1470 ();
 sg13g2_fill_1 FILLER_26_1492 ();
 sg13g2_decap_4 FILLER_26_1505 ();
 sg13g2_fill_2 FILLER_26_1516 ();
 sg13g2_decap_8 FILLER_26_1536 ();
 sg13g2_decap_4 FILLER_26_1543 ();
 sg13g2_fill_2 FILLER_26_1547 ();
 sg13g2_decap_4 FILLER_26_1554 ();
 sg13g2_fill_2 FILLER_26_1558 ();
 sg13g2_decap_8 FILLER_26_1566 ();
 sg13g2_decap_8 FILLER_26_1573 ();
 sg13g2_fill_1 FILLER_26_1580 ();
 sg13g2_decap_8 FILLER_26_1598 ();
 sg13g2_decap_8 FILLER_26_1605 ();
 sg13g2_fill_2 FILLER_26_1612 ();
 sg13g2_fill_1 FILLER_26_1614 ();
 sg13g2_fill_1 FILLER_26_1620 ();
 sg13g2_decap_4 FILLER_26_1671 ();
 sg13g2_fill_2 FILLER_26_1712 ();
 sg13g2_fill_1 FILLER_26_1714 ();
 sg13g2_decap_8 FILLER_26_1758 ();
 sg13g2_fill_2 FILLER_26_1765 ();
 sg13g2_fill_1 FILLER_26_1767 ();
 sg13g2_decap_8 FILLER_26_1778 ();
 sg13g2_decap_8 FILLER_26_1785 ();
 sg13g2_decap_8 FILLER_26_1800 ();
 sg13g2_decap_8 FILLER_26_1807 ();
 sg13g2_decap_8 FILLER_26_1814 ();
 sg13g2_fill_1 FILLER_26_1821 ();
 sg13g2_fill_1 FILLER_26_1834 ();
 sg13g2_fill_1 FILLER_26_1848 ();
 sg13g2_fill_1 FILLER_26_1853 ();
 sg13g2_decap_4 FILLER_26_1873 ();
 sg13g2_fill_1 FILLER_26_1877 ();
 sg13g2_fill_2 FILLER_26_1888 ();
 sg13g2_fill_1 FILLER_26_1890 ();
 sg13g2_fill_1 FILLER_26_1895 ();
 sg13g2_decap_4 FILLER_26_1902 ();
 sg13g2_fill_2 FILLER_26_1906 ();
 sg13g2_decap_4 FILLER_26_1945 ();
 sg13g2_decap_8 FILLER_26_1952 ();
 sg13g2_fill_2 FILLER_26_1959 ();
 sg13g2_fill_2 FILLER_26_1998 ();
 sg13g2_decap_8 FILLER_26_2060 ();
 sg13g2_decap_8 FILLER_26_2067 ();
 sg13g2_fill_2 FILLER_26_2091 ();
 sg13g2_decap_8 FILLER_26_2124 ();
 sg13g2_decap_8 FILLER_26_2131 ();
 sg13g2_decap_4 FILLER_26_2138 ();
 sg13g2_fill_2 FILLER_26_2152 ();
 sg13g2_decap_8 FILLER_26_2192 ();
 sg13g2_fill_2 FILLER_26_2199 ();
 sg13g2_fill_2 FILLER_26_2227 ();
 sg13g2_fill_2 FILLER_26_2237 ();
 sg13g2_fill_1 FILLER_26_2239 ();
 sg13g2_fill_2 FILLER_26_2250 ();
 sg13g2_decap_4 FILLER_26_2278 ();
 sg13g2_fill_2 FILLER_26_2290 ();
 sg13g2_fill_1 FILLER_26_2352 ();
 sg13g2_fill_2 FILLER_26_2356 ();
 sg13g2_fill_1 FILLER_26_2373 ();
 sg13g2_fill_2 FILLER_26_2430 ();
 sg13g2_decap_4 FILLER_26_2439 ();
 sg13g2_fill_2 FILLER_26_2453 ();
 sg13g2_fill_1 FILLER_26_2455 ();
 sg13g2_fill_2 FILLER_26_2489 ();
 sg13g2_decap_4 FILLER_26_2517 ();
 sg13g2_fill_2 FILLER_26_2525 ();
 sg13g2_fill_2 FILLER_26_2540 ();
 sg13g2_fill_1 FILLER_26_2542 ();
 sg13g2_fill_1 FILLER_26_2575 ();
 sg13g2_decap_4 FILLER_26_2623 ();
 sg13g2_decap_8 FILLER_26_2663 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_32 ();
 sg13g2_fill_1 FILLER_27_34 ();
 sg13g2_decap_8 FILLER_27_54 ();
 sg13g2_fill_2 FILLER_27_91 ();
 sg13g2_fill_2 FILLER_27_111 ();
 sg13g2_fill_1 FILLER_27_113 ();
 sg13g2_fill_2 FILLER_27_168 ();
 sg13g2_decap_4 FILLER_27_178 ();
 sg13g2_fill_2 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_188 ();
 sg13g2_decap_4 FILLER_27_195 ();
 sg13g2_fill_1 FILLER_27_199 ();
 sg13g2_decap_4 FILLER_27_204 ();
 sg13g2_fill_2 FILLER_27_208 ();
 sg13g2_fill_2 FILLER_27_236 ();
 sg13g2_fill_1 FILLER_27_238 ();
 sg13g2_decap_8 FILLER_27_296 ();
 sg13g2_fill_1 FILLER_27_303 ();
 sg13g2_decap_4 FILLER_27_361 ();
 sg13g2_fill_1 FILLER_27_365 ();
 sg13g2_fill_2 FILLER_27_439 ();
 sg13g2_fill_2 FILLER_27_446 ();
 sg13g2_fill_2 FILLER_27_452 ();
 sg13g2_fill_1 FILLER_27_454 ();
 sg13g2_fill_2 FILLER_27_459 ();
 sg13g2_fill_1 FILLER_27_461 ();
 sg13g2_fill_2 FILLER_27_467 ();
 sg13g2_fill_1 FILLER_27_469 ();
 sg13g2_fill_1 FILLER_27_483 ();
 sg13g2_decap_4 FILLER_27_498 ();
 sg13g2_fill_1 FILLER_27_516 ();
 sg13g2_fill_1 FILLER_27_521 ();
 sg13g2_decap_4 FILLER_27_526 ();
 sg13g2_decap_4 FILLER_27_534 ();
 sg13g2_fill_2 FILLER_27_548 ();
 sg13g2_fill_2 FILLER_27_578 ();
 sg13g2_fill_2 FILLER_27_584 ();
 sg13g2_decap_8 FILLER_27_590 ();
 sg13g2_fill_2 FILLER_27_627 ();
 sg13g2_fill_1 FILLER_27_629 ();
 sg13g2_fill_1 FILLER_27_635 ();
 sg13g2_fill_1 FILLER_27_705 ();
 sg13g2_fill_2 FILLER_27_710 ();
 sg13g2_fill_1 FILLER_27_717 ();
 sg13g2_fill_2 FILLER_27_723 ();
 sg13g2_fill_1 FILLER_27_725 ();
 sg13g2_fill_2 FILLER_27_760 ();
 sg13g2_fill_1 FILLER_27_771 ();
 sg13g2_decap_8 FILLER_27_813 ();
 sg13g2_decap_8 FILLER_27_847 ();
 sg13g2_decap_8 FILLER_27_854 ();
 sg13g2_decap_4 FILLER_27_861 ();
 sg13g2_fill_2 FILLER_27_865 ();
 sg13g2_fill_1 FILLER_27_871 ();
 sg13g2_decap_8 FILLER_27_876 ();
 sg13g2_decap_4 FILLER_27_883 ();
 sg13g2_fill_2 FILLER_27_887 ();
 sg13g2_decap_8 FILLER_27_902 ();
 sg13g2_fill_2 FILLER_27_909 ();
 sg13g2_decap_8 FILLER_27_919 ();
 sg13g2_fill_1 FILLER_27_926 ();
 sg13g2_fill_1 FILLER_27_931 ();
 sg13g2_fill_1 FILLER_27_962 ();
 sg13g2_fill_1 FILLER_27_968 ();
 sg13g2_fill_2 FILLER_27_982 ();
 sg13g2_fill_1 FILLER_27_984 ();
 sg13g2_decap_8 FILLER_27_989 ();
 sg13g2_decap_8 FILLER_27_996 ();
 sg13g2_decap_8 FILLER_27_1003 ();
 sg13g2_decap_8 FILLER_27_1010 ();
 sg13g2_decap_8 FILLER_27_1017 ();
 sg13g2_decap_8 FILLER_27_1024 ();
 sg13g2_fill_2 FILLER_27_1041 ();
 sg13g2_decap_8 FILLER_27_1061 ();
 sg13g2_decap_8 FILLER_27_1068 ();
 sg13g2_decap_4 FILLER_27_1126 ();
 sg13g2_fill_1 FILLER_27_1130 ();
 sg13g2_fill_2 FILLER_27_1177 ();
 sg13g2_decap_4 FILLER_27_1184 ();
 sg13g2_fill_1 FILLER_27_1188 ();
 sg13g2_fill_2 FILLER_27_1215 ();
 sg13g2_fill_1 FILLER_27_1238 ();
 sg13g2_fill_1 FILLER_27_1265 ();
 sg13g2_decap_4 FILLER_27_1270 ();
 sg13g2_fill_2 FILLER_27_1274 ();
 sg13g2_fill_2 FILLER_27_1310 ();
 sg13g2_fill_1 FILLER_27_1312 ();
 sg13g2_decap_8 FILLER_27_1343 ();
 sg13g2_decap_8 FILLER_27_1350 ();
 sg13g2_decap_8 FILLER_27_1357 ();
 sg13g2_fill_2 FILLER_27_1394 ();
 sg13g2_fill_1 FILLER_27_1396 ();
 sg13g2_fill_2 FILLER_27_1401 ();
 sg13g2_fill_2 FILLER_27_1442 ();
 sg13g2_fill_1 FILLER_27_1444 ();
 sg13g2_fill_1 FILLER_27_1454 ();
 sg13g2_fill_2 FILLER_27_1461 ();
 sg13g2_fill_1 FILLER_27_1463 ();
 sg13g2_fill_2 FILLER_27_1479 ();
 sg13g2_decap_8 FILLER_27_1489 ();
 sg13g2_decap_8 FILLER_27_1496 ();
 sg13g2_decap_8 FILLER_27_1503 ();
 sg13g2_fill_2 FILLER_27_1510 ();
 sg13g2_fill_2 FILLER_27_1517 ();
 sg13g2_fill_1 FILLER_27_1519 ();
 sg13g2_decap_8 FILLER_27_1549 ();
 sg13g2_fill_2 FILLER_27_1556 ();
 sg13g2_fill_1 FILLER_27_1567 ();
 sg13g2_decap_8 FILLER_27_1579 ();
 sg13g2_fill_1 FILLER_27_1586 ();
 sg13g2_fill_2 FILLER_27_1649 ();
 sg13g2_decap_4 FILLER_27_1656 ();
 sg13g2_fill_2 FILLER_27_1670 ();
 sg13g2_fill_1 FILLER_27_1672 ();
 sg13g2_fill_2 FILLER_27_1722 ();
 sg13g2_fill_2 FILLER_27_1786 ();
 sg13g2_fill_1 FILLER_27_1814 ();
 sg13g2_decap_8 FILLER_27_1824 ();
 sg13g2_fill_1 FILLER_27_1831 ();
 sg13g2_fill_2 FILLER_27_1846 ();
 sg13g2_fill_1 FILLER_27_1874 ();
 sg13g2_fill_2 FILLER_27_1916 ();
 sg13g2_fill_1 FILLER_27_1918 ();
 sg13g2_fill_2 FILLER_27_1959 ();
 sg13g2_fill_1 FILLER_27_1961 ();
 sg13g2_fill_2 FILLER_27_1972 ();
 sg13g2_fill_2 FILLER_27_2023 ();
 sg13g2_decap_4 FILLER_27_2089 ();
 sg13g2_decap_8 FILLER_27_2106 ();
 sg13g2_decap_8 FILLER_27_2113 ();
 sg13g2_decap_8 FILLER_27_2120 ();
 sg13g2_decap_4 FILLER_27_2127 ();
 sg13g2_fill_2 FILLER_27_2131 ();
 sg13g2_decap_8 FILLER_27_2137 ();
 sg13g2_fill_1 FILLER_27_2144 ();
 sg13g2_decap_4 FILLER_27_2206 ();
 sg13g2_fill_1 FILLER_27_2210 ();
 sg13g2_fill_2 FILLER_27_2237 ();
 sg13g2_fill_1 FILLER_27_2254 ();
 sg13g2_fill_2 FILLER_27_2284 ();
 sg13g2_fill_1 FILLER_27_2299 ();
 sg13g2_fill_1 FILLER_27_2345 ();
 sg13g2_fill_2 FILLER_27_2362 ();
 sg13g2_fill_2 FILLER_27_2438 ();
 sg13g2_fill_1 FILLER_27_2476 ();
 sg13g2_fill_2 FILLER_27_2491 ();
 sg13g2_fill_1 FILLER_27_2493 ();
 sg13g2_decap_8 FILLER_27_2504 ();
 sg13g2_decap_4 FILLER_27_2511 ();
 sg13g2_fill_2 FILLER_27_2515 ();
 sg13g2_fill_1 FILLER_27_2548 ();
 sg13g2_fill_1 FILLER_27_2575 ();
 sg13g2_fill_1 FILLER_27_2586 ();
 sg13g2_fill_2 FILLER_27_2613 ();
 sg13g2_decap_8 FILLER_27_2629 ();
 sg13g2_fill_2 FILLER_27_2636 ();
 sg13g2_fill_1 FILLER_27_2638 ();
 sg13g2_decap_8 FILLER_27_2647 ();
 sg13g2_decap_8 FILLER_27_2654 ();
 sg13g2_decap_8 FILLER_27_2661 ();
 sg13g2_fill_2 FILLER_27_2668 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_7 ();
 sg13g2_fill_2 FILLER_28_11 ();
 sg13g2_fill_2 FILLER_28_17 ();
 sg13g2_fill_1 FILLER_28_45 ();
 sg13g2_fill_2 FILLER_28_50 ();
 sg13g2_fill_2 FILLER_28_78 ();
 sg13g2_fill_1 FILLER_28_126 ();
 sg13g2_fill_1 FILLER_28_148 ();
 sg13g2_fill_2 FILLER_28_158 ();
 sg13g2_fill_2 FILLER_28_190 ();
 sg13g2_decap_4 FILLER_28_200 ();
 sg13g2_decap_8 FILLER_28_208 ();
 sg13g2_fill_2 FILLER_28_215 ();
 sg13g2_fill_1 FILLER_28_221 ();
 sg13g2_fill_1 FILLER_28_253 ();
 sg13g2_fill_1 FILLER_28_258 ();
 sg13g2_fill_1 FILLER_28_263 ();
 sg13g2_fill_2 FILLER_28_278 ();
 sg13g2_decap_8 FILLER_28_292 ();
 sg13g2_decap_4 FILLER_28_299 ();
 sg13g2_fill_1 FILLER_28_303 ();
 sg13g2_decap_8 FILLER_28_329 ();
 sg13g2_fill_1 FILLER_28_336 ();
 sg13g2_decap_4 FILLER_28_373 ();
 sg13g2_fill_2 FILLER_28_377 ();
 sg13g2_fill_2 FILLER_28_387 ();
 sg13g2_fill_1 FILLER_28_389 ();
 sg13g2_decap_4 FILLER_28_420 ();
 sg13g2_decap_4 FILLER_28_434 ();
 sg13g2_fill_1 FILLER_28_453 ();
 sg13g2_decap_8 FILLER_28_472 ();
 sg13g2_decap_4 FILLER_28_479 ();
 sg13g2_fill_2 FILLER_28_483 ();
 sg13g2_fill_1 FILLER_28_515 ();
 sg13g2_decap_8 FILLER_28_525 ();
 sg13g2_decap_4 FILLER_28_532 ();
 sg13g2_fill_1 FILLER_28_542 ();
 sg13g2_fill_1 FILLER_28_608 ();
 sg13g2_fill_1 FILLER_28_620 ();
 sg13g2_fill_1 FILLER_28_630 ();
 sg13g2_decap_4 FILLER_28_703 ();
 sg13g2_fill_2 FILLER_28_748 ();
 sg13g2_fill_2 FILLER_28_767 ();
 sg13g2_fill_1 FILLER_28_789 ();
 sg13g2_fill_2 FILLER_28_816 ();
 sg13g2_decap_8 FILLER_28_858 ();
 sg13g2_decap_4 FILLER_28_865 ();
 sg13g2_fill_1 FILLER_28_869 ();
 sg13g2_fill_2 FILLER_28_874 ();
 sg13g2_fill_2 FILLER_28_886 ();
 sg13g2_fill_1 FILLER_28_888 ();
 sg13g2_fill_2 FILLER_28_910 ();
 sg13g2_fill_1 FILLER_28_912 ();
 sg13g2_fill_2 FILLER_28_949 ();
 sg13g2_decap_8 FILLER_28_961 ();
 sg13g2_fill_2 FILLER_28_968 ();
 sg13g2_decap_8 FILLER_28_1006 ();
 sg13g2_decap_8 FILLER_28_1013 ();
 sg13g2_decap_8 FILLER_28_1020 ();
 sg13g2_decap_8 FILLER_28_1027 ();
 sg13g2_decap_8 FILLER_28_1034 ();
 sg13g2_fill_2 FILLER_28_1041 ();
 sg13g2_fill_1 FILLER_28_1043 ();
 sg13g2_decap_8 FILLER_28_1070 ();
 sg13g2_fill_2 FILLER_28_1077 ();
 sg13g2_fill_1 FILLER_28_1079 ();
 sg13g2_fill_2 FILLER_28_1119 ();
 sg13g2_fill_1 FILLER_28_1121 ();
 sg13g2_fill_1 FILLER_28_1158 ();
 sg13g2_decap_8 FILLER_28_1181 ();
 sg13g2_fill_2 FILLER_28_1188 ();
 sg13g2_decap_8 FILLER_28_1230 ();
 sg13g2_fill_1 FILLER_28_1237 ();
 sg13g2_decap_8 FILLER_28_1259 ();
 sg13g2_fill_2 FILLER_28_1266 ();
 sg13g2_fill_1 FILLER_28_1273 ();
 sg13g2_fill_1 FILLER_28_1279 ();
 sg13g2_decap_4 FILLER_28_1318 ();
 sg13g2_fill_2 FILLER_28_1322 ();
 sg13g2_decap_4 FILLER_28_1328 ();
 sg13g2_fill_2 FILLER_28_1332 ();
 sg13g2_decap_8 FILLER_28_1344 ();
 sg13g2_decap_4 FILLER_28_1351 ();
 sg13g2_fill_1 FILLER_28_1355 ();
 sg13g2_fill_2 FILLER_28_1392 ();
 sg13g2_fill_1 FILLER_28_1404 ();
 sg13g2_fill_2 FILLER_28_1418 ();
 sg13g2_decap_8 FILLER_28_1424 ();
 sg13g2_fill_2 FILLER_28_1431 ();
 sg13g2_fill_1 FILLER_28_1446 ();
 sg13g2_fill_1 FILLER_28_1452 ();
 sg13g2_decap_4 FILLER_28_1463 ();
 sg13g2_fill_2 FILLER_28_1483 ();
 sg13g2_fill_2 FILLER_28_1490 ();
 sg13g2_fill_2 FILLER_28_1497 ();
 sg13g2_fill_1 FILLER_28_1499 ();
 sg13g2_fill_1 FILLER_28_1505 ();
 sg13g2_fill_2 FILLER_28_1528 ();
 sg13g2_fill_1 FILLER_28_1530 ();
 sg13g2_decap_4 FILLER_28_1535 ();
 sg13g2_fill_2 FILLER_28_1539 ();
 sg13g2_decap_8 FILLER_28_1546 ();
 sg13g2_decap_8 FILLER_28_1553 ();
 sg13g2_fill_2 FILLER_28_1560 ();
 sg13g2_fill_1 FILLER_28_1562 ();
 sg13g2_decap_4 FILLER_28_1568 ();
 sg13g2_fill_1 FILLER_28_1572 ();
 sg13g2_decap_4 FILLER_28_1578 ();
 sg13g2_fill_2 FILLER_28_1582 ();
 sg13g2_fill_1 FILLER_28_1631 ();
 sg13g2_fill_2 FILLER_28_1652 ();
 sg13g2_decap_8 FILLER_28_1661 ();
 sg13g2_decap_8 FILLER_28_1668 ();
 sg13g2_decap_8 FILLER_28_1675 ();
 sg13g2_decap_8 FILLER_28_1682 ();
 sg13g2_decap_4 FILLER_28_1689 ();
 sg13g2_fill_1 FILLER_28_1693 ();
 sg13g2_decap_8 FILLER_28_1759 ();
 sg13g2_fill_2 FILLER_28_1766 ();
 sg13g2_fill_1 FILLER_28_1768 ();
 sg13g2_fill_1 FILLER_28_1773 ();
 sg13g2_fill_1 FILLER_28_1800 ();
 sg13g2_fill_1 FILLER_28_1810 ();
 sg13g2_fill_1 FILLER_28_1845 ();
 sg13g2_fill_1 FILLER_28_1888 ();
 sg13g2_decap_8 FILLER_28_1933 ();
 sg13g2_fill_2 FILLER_28_1940 ();
 sg13g2_decap_4 FILLER_28_2001 ();
 sg13g2_fill_1 FILLER_28_2005 ();
 sg13g2_decap_8 FILLER_28_2015 ();
 sg13g2_decap_8 FILLER_28_2022 ();
 sg13g2_decap_8 FILLER_28_2029 ();
 sg13g2_decap_8 FILLER_28_2049 ();
 sg13g2_decap_8 FILLER_28_2123 ();
 sg13g2_decap_8 FILLER_28_2130 ();
 sg13g2_fill_1 FILLER_28_2155 ();
 sg13g2_fill_1 FILLER_28_2160 ();
 sg13g2_fill_2 FILLER_28_2186 ();
 sg13g2_fill_2 FILLER_28_2192 ();
 sg13g2_decap_8 FILLER_28_2237 ();
 sg13g2_decap_4 FILLER_28_2254 ();
 sg13g2_fill_1 FILLER_28_2352 ();
 sg13g2_fill_2 FILLER_28_2484 ();
 sg13g2_fill_1 FILLER_28_2486 ();
 sg13g2_fill_2 FILLER_28_2491 ();
 sg13g2_decap_8 FILLER_28_2533 ();
 sg13g2_fill_1 FILLER_28_2545 ();
 sg13g2_decap_4 FILLER_28_2560 ();
 sg13g2_fill_1 FILLER_28_2564 ();
 sg13g2_decap_8 FILLER_28_2582 ();
 sg13g2_fill_1 FILLER_28_2589 ();
 sg13g2_decap_4 FILLER_28_2597 ();
 sg13g2_fill_2 FILLER_28_2601 ();
 sg13g2_decap_8 FILLER_28_2616 ();
 sg13g2_decap_4 FILLER_28_2623 ();
 sg13g2_fill_2 FILLER_28_2627 ();
 sg13g2_decap_8 FILLER_28_2655 ();
 sg13g2_decap_8 FILLER_28_2662 ();
 sg13g2_fill_1 FILLER_28_2669 ();
 sg13g2_decap_4 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_4 ();
 sg13g2_decap_8 FILLER_29_9 ();
 sg13g2_fill_2 FILLER_29_31 ();
 sg13g2_fill_1 FILLER_29_48 ();
 sg13g2_decap_4 FILLER_29_106 ();
 sg13g2_fill_1 FILLER_29_110 ();
 sg13g2_fill_1 FILLER_29_121 ();
 sg13g2_fill_1 FILLER_29_127 ();
 sg13g2_fill_1 FILLER_29_133 ();
 sg13g2_fill_1 FILLER_29_143 ();
 sg13g2_fill_2 FILLER_29_162 ();
 sg13g2_fill_1 FILLER_29_164 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_decap_8 FILLER_29_182 ();
 sg13g2_fill_2 FILLER_29_189 ();
 sg13g2_fill_1 FILLER_29_191 ();
 sg13g2_fill_1 FILLER_29_199 ();
 sg13g2_decap_8 FILLER_29_226 ();
 sg13g2_fill_2 FILLER_29_233 ();
 sg13g2_fill_1 FILLER_29_235 ();
 sg13g2_decap_4 FILLER_29_240 ();
 sg13g2_decap_8 FILLER_29_248 ();
 sg13g2_decap_4 FILLER_29_255 ();
 sg13g2_decap_8 FILLER_29_282 ();
 sg13g2_fill_2 FILLER_29_289 ();
 sg13g2_decap_8 FILLER_29_295 ();
 sg13g2_decap_8 FILLER_29_302 ();
 sg13g2_decap_8 FILLER_29_309 ();
 sg13g2_decap_8 FILLER_29_332 ();
 sg13g2_fill_2 FILLER_29_339 ();
 sg13g2_fill_1 FILLER_29_341 ();
 sg13g2_decap_8 FILLER_29_346 ();
 sg13g2_fill_2 FILLER_29_353 ();
 sg13g2_fill_1 FILLER_29_355 ();
 sg13g2_decap_8 FILLER_29_360 ();
 sg13g2_decap_8 FILLER_29_367 ();
 sg13g2_decap_8 FILLER_29_374 ();
 sg13g2_decap_8 FILLER_29_381 ();
 sg13g2_decap_8 FILLER_29_388 ();
 sg13g2_decap_8 FILLER_29_395 ();
 sg13g2_fill_1 FILLER_29_402 ();
 sg13g2_decap_8 FILLER_29_471 ();
 sg13g2_decap_4 FILLER_29_478 ();
 sg13g2_fill_1 FILLER_29_482 ();
 sg13g2_fill_1 FILLER_29_493 ();
 sg13g2_fill_1 FILLER_29_500 ();
 sg13g2_fill_1 FILLER_29_506 ();
 sg13g2_fill_1 FILLER_29_517 ();
 sg13g2_decap_8 FILLER_29_524 ();
 sg13g2_decap_4 FILLER_29_531 ();
 sg13g2_decap_8 FILLER_29_560 ();
 sg13g2_decap_4 FILLER_29_567 ();
 sg13g2_fill_1 FILLER_29_571 ();
 sg13g2_decap_8 FILLER_29_580 ();
 sg13g2_decap_8 FILLER_29_587 ();
 sg13g2_decap_8 FILLER_29_594 ();
 sg13g2_fill_2 FILLER_29_601 ();
 sg13g2_fill_2 FILLER_29_621 ();
 sg13g2_fill_1 FILLER_29_623 ();
 sg13g2_decap_4 FILLER_29_650 ();
 sg13g2_fill_1 FILLER_29_654 ();
 sg13g2_decap_4 FILLER_29_660 ();
 sg13g2_fill_1 FILLER_29_664 ();
 sg13g2_fill_2 FILLER_29_669 ();
 sg13g2_fill_1 FILLER_29_671 ();
 sg13g2_fill_1 FILLER_29_676 ();
 sg13g2_fill_2 FILLER_29_685 ();
 sg13g2_fill_1 FILLER_29_687 ();
 sg13g2_decap_8 FILLER_29_693 ();
 sg13g2_decap_8 FILLER_29_700 ();
 sg13g2_fill_1 FILLER_29_707 ();
 sg13g2_fill_1 FILLER_29_712 ();
 sg13g2_decap_4 FILLER_29_716 ();
 sg13g2_fill_1 FILLER_29_727 ();
 sg13g2_decap_8 FILLER_29_734 ();
 sg13g2_decap_8 FILLER_29_741 ();
 sg13g2_fill_2 FILLER_29_748 ();
 sg13g2_fill_1 FILLER_29_750 ();
 sg13g2_fill_1 FILLER_29_804 ();
 sg13g2_decap_8 FILLER_29_809 ();
 sg13g2_decap_8 FILLER_29_816 ();
 sg13g2_fill_1 FILLER_29_823 ();
 sg13g2_fill_2 FILLER_29_860 ();
 sg13g2_fill_1 FILLER_29_862 ();
 sg13g2_fill_2 FILLER_29_915 ();
 sg13g2_decap_4 FILLER_29_943 ();
 sg13g2_fill_1 FILLER_29_993 ();
 sg13g2_fill_1 FILLER_29_998 ();
 sg13g2_decap_4 FILLER_29_1035 ();
 sg13g2_fill_1 FILLER_29_1039 ();
 sg13g2_decap_4 FILLER_29_1044 ();
 sg13g2_decap_8 FILLER_29_1058 ();
 sg13g2_fill_1 FILLER_29_1065 ();
 sg13g2_decap_4 FILLER_29_1076 ();
 sg13g2_fill_2 FILLER_29_1085 ();
 sg13g2_decap_4 FILLER_29_1113 ();
 sg13g2_fill_2 FILLER_29_1117 ();
 sg13g2_fill_2 FILLER_29_1205 ();
 sg13g2_fill_1 FILLER_29_1247 ();
 sg13g2_decap_8 FILLER_29_1252 ();
 sg13g2_decap_8 FILLER_29_1259 ();
 sg13g2_decap_4 FILLER_29_1266 ();
 sg13g2_fill_2 FILLER_29_1270 ();
 sg13g2_fill_1 FILLER_29_1333 ();
 sg13g2_fill_1 FILLER_29_1360 ();
 sg13g2_fill_1 FILLER_29_1387 ();
 sg13g2_fill_1 FILLER_29_1398 ();
 sg13g2_fill_2 FILLER_29_1409 ();
 sg13g2_fill_2 FILLER_29_1415 ();
 sg13g2_fill_1 FILLER_29_1417 ();
 sg13g2_decap_8 FILLER_29_1426 ();
 sg13g2_fill_2 FILLER_29_1433 ();
 sg13g2_decap_8 FILLER_29_1505 ();
 sg13g2_decap_4 FILLER_29_1512 ();
 sg13g2_fill_2 FILLER_29_1516 ();
 sg13g2_fill_2 FILLER_29_1523 ();
 sg13g2_fill_1 FILLER_29_1525 ();
 sg13g2_decap_8 FILLER_29_1537 ();
 sg13g2_fill_1 FILLER_29_1549 ();
 sg13g2_decap_8 FILLER_29_1555 ();
 sg13g2_fill_2 FILLER_29_1562 ();
 sg13g2_fill_1 FILLER_29_1564 ();
 sg13g2_decap_4 FILLER_29_1571 ();
 sg13g2_fill_2 FILLER_29_1575 ();
 sg13g2_fill_1 FILLER_29_1583 ();
 sg13g2_decap_8 FILLER_29_1670 ();
 sg13g2_fill_2 FILLER_29_1748 ();
 sg13g2_fill_1 FILLER_29_1750 ();
 sg13g2_fill_2 FILLER_29_1774 ();
 sg13g2_decap_4 FILLER_29_1798 ();
 sg13g2_decap_4 FILLER_29_1806 ();
 sg13g2_fill_2 FILLER_29_1815 ();
 sg13g2_fill_2 FILLER_29_1828 ();
 sg13g2_fill_2 FILLER_29_1842 ();
 sg13g2_decap_8 FILLER_29_1849 ();
 sg13g2_fill_2 FILLER_29_1856 ();
 sg13g2_fill_1 FILLER_29_1896 ();
 sg13g2_fill_1 FILLER_29_1913 ();
 sg13g2_decap_4 FILLER_29_1931 ();
 sg13g2_decap_4 FILLER_29_1970 ();
 sg13g2_fill_2 FILLER_29_1982 ();
 sg13g2_decap_4 FILLER_29_1993 ();
 sg13g2_fill_1 FILLER_29_1997 ();
 sg13g2_decap_8 FILLER_29_2024 ();
 sg13g2_decap_4 FILLER_29_2031 ();
 sg13g2_fill_1 FILLER_29_2079 ();
 sg13g2_fill_2 FILLER_29_2137 ();
 sg13g2_fill_1 FILLER_29_2165 ();
 sg13g2_fill_2 FILLER_29_2192 ();
 sg13g2_fill_1 FILLER_29_2208 ();
 sg13g2_fill_2 FILLER_29_2230 ();
 sg13g2_fill_2 FILLER_29_2236 ();
 sg13g2_decap_8 FILLER_29_2246 ();
 sg13g2_fill_1 FILLER_29_2253 ();
 sg13g2_fill_2 FILLER_29_2272 ();
 sg13g2_fill_1 FILLER_29_2274 ();
 sg13g2_fill_1 FILLER_29_2318 ();
 sg13g2_fill_2 FILLER_29_2332 ();
 sg13g2_fill_2 FILLER_29_2339 ();
 sg13g2_fill_1 FILLER_29_2386 ();
 sg13g2_fill_1 FILLER_29_2423 ();
 sg13g2_fill_1 FILLER_29_2450 ();
 sg13g2_fill_2 FILLER_29_2472 ();
 sg13g2_fill_2 FILLER_29_2563 ();
 sg13g2_decap_4 FILLER_29_2612 ();
 sg13g2_fill_1 FILLER_29_2616 ();
 sg13g2_decap_8 FILLER_29_2653 ();
 sg13g2_decap_8 FILLER_29_2660 ();
 sg13g2_fill_2 FILLER_29_2667 ();
 sg13g2_fill_1 FILLER_29_2669 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_38 ();
 sg13g2_fill_1 FILLER_30_40 ();
 sg13g2_fill_2 FILLER_30_46 ();
 sg13g2_fill_1 FILLER_30_48 ();
 sg13g2_decap_8 FILLER_30_53 ();
 sg13g2_fill_2 FILLER_30_70 ();
 sg13g2_fill_1 FILLER_30_72 ();
 sg13g2_fill_1 FILLER_30_77 ();
 sg13g2_decap_4 FILLER_30_100 ();
 sg13g2_fill_1 FILLER_30_104 ();
 sg13g2_fill_2 FILLER_30_119 ();
 sg13g2_fill_1 FILLER_30_133 ();
 sg13g2_fill_2 FILLER_30_139 ();
 sg13g2_fill_1 FILLER_30_141 ();
 sg13g2_fill_1 FILLER_30_155 ();
 sg13g2_fill_1 FILLER_30_164 ();
 sg13g2_fill_1 FILLER_30_175 ();
 sg13g2_fill_1 FILLER_30_180 ();
 sg13g2_fill_1 FILLER_30_191 ();
 sg13g2_fill_1 FILLER_30_202 ();
 sg13g2_fill_1 FILLER_30_211 ();
 sg13g2_decap_4 FILLER_30_216 ();
 sg13g2_decap_8 FILLER_30_233 ();
 sg13g2_decap_8 FILLER_30_240 ();
 sg13g2_decap_8 FILLER_30_247 ();
 sg13g2_fill_2 FILLER_30_254 ();
 sg13g2_fill_1 FILLER_30_270 ();
 sg13g2_fill_1 FILLER_30_280 ();
 sg13g2_decap_4 FILLER_30_287 ();
 sg13g2_fill_2 FILLER_30_300 ();
 sg13g2_fill_2 FILLER_30_316 ();
 sg13g2_decap_8 FILLER_30_335 ();
 sg13g2_decap_8 FILLER_30_342 ();
 sg13g2_fill_2 FILLER_30_349 ();
 sg13g2_decap_8 FILLER_30_360 ();
 sg13g2_decap_8 FILLER_30_367 ();
 sg13g2_decap_8 FILLER_30_374 ();
 sg13g2_decap_8 FILLER_30_381 ();
 sg13g2_decap_8 FILLER_30_388 ();
 sg13g2_decap_8 FILLER_30_395 ();
 sg13g2_decap_8 FILLER_30_402 ();
 sg13g2_decap_8 FILLER_30_409 ();
 sg13g2_fill_2 FILLER_30_416 ();
 sg13g2_fill_1 FILLER_30_418 ();
 sg13g2_decap_8 FILLER_30_423 ();
 sg13g2_fill_2 FILLER_30_430 ();
 sg13g2_fill_1 FILLER_30_464 ();
 sg13g2_fill_1 FILLER_30_496 ();
 sg13g2_decap_4 FILLER_30_537 ();
 sg13g2_fill_1 FILLER_30_541 ();
 sg13g2_decap_8 FILLER_30_553 ();
 sg13g2_fill_1 FILLER_30_560 ();
 sg13g2_decap_8 FILLER_30_579 ();
 sg13g2_decap_8 FILLER_30_586 ();
 sg13g2_fill_1 FILLER_30_593 ();
 sg13g2_decap_4 FILLER_30_603 ();
 sg13g2_fill_1 FILLER_30_607 ();
 sg13g2_decap_4 FILLER_30_613 ();
 sg13g2_fill_2 FILLER_30_617 ();
 sg13g2_decap_8 FILLER_30_624 ();
 sg13g2_decap_8 FILLER_30_635 ();
 sg13g2_fill_2 FILLER_30_642 ();
 sg13g2_fill_1 FILLER_30_644 ();
 sg13g2_decap_8 FILLER_30_649 ();
 sg13g2_decap_8 FILLER_30_656 ();
 sg13g2_decap_4 FILLER_30_663 ();
 sg13g2_fill_1 FILLER_30_667 ();
 sg13g2_decap_8 FILLER_30_673 ();
 sg13g2_fill_2 FILLER_30_680 ();
 sg13g2_fill_1 FILLER_30_682 ();
 sg13g2_fill_1 FILLER_30_719 ();
 sg13g2_fill_2 FILLER_30_727 ();
 sg13g2_decap_8 FILLER_30_737 ();
 sg13g2_decap_8 FILLER_30_744 ();
 sg13g2_decap_8 FILLER_30_751 ();
 sg13g2_decap_8 FILLER_30_758 ();
 sg13g2_decap_4 FILLER_30_765 ();
 sg13g2_decap_4 FILLER_30_774 ();
 sg13g2_fill_1 FILLER_30_778 ();
 sg13g2_decap_8 FILLER_30_783 ();
 sg13g2_decap_8 FILLER_30_790 ();
 sg13g2_decap_8 FILLER_30_797 ();
 sg13g2_decap_8 FILLER_30_804 ();
 sg13g2_decap_8 FILLER_30_811 ();
 sg13g2_decap_8 FILLER_30_818 ();
 sg13g2_fill_1 FILLER_30_825 ();
 sg13g2_fill_2 FILLER_30_862 ();
 sg13g2_fill_2 FILLER_30_885 ();
 sg13g2_fill_1 FILLER_30_887 ();
 sg13g2_fill_2 FILLER_30_945 ();
 sg13g2_fill_1 FILLER_30_947 ();
 sg13g2_fill_1 FILLER_30_974 ();
 sg13g2_decap_4 FILLER_30_1011 ();
 sg13g2_fill_2 FILLER_30_1041 ();
 sg13g2_fill_1 FILLER_30_1043 ();
 sg13g2_fill_2 FILLER_30_1070 ();
 sg13g2_decap_4 FILLER_30_1101 ();
 sg13g2_decap_4 FILLER_30_1109 ();
 sg13g2_fill_2 FILLER_30_1113 ();
 sg13g2_fill_1 FILLER_30_1127 ();
 sg13g2_fill_2 FILLER_30_1146 ();
 sg13g2_fill_2 FILLER_30_1173 ();
 sg13g2_fill_1 FILLER_30_1175 ();
 sg13g2_decap_8 FILLER_30_1202 ();
 sg13g2_decap_8 FILLER_30_1209 ();
 sg13g2_decap_8 FILLER_30_1216 ();
 sg13g2_decap_4 FILLER_30_1223 ();
 sg13g2_fill_1 FILLER_30_1227 ();
 sg13g2_fill_1 FILLER_30_1236 ();
 sg13g2_decap_8 FILLER_30_1242 ();
 sg13g2_decap_8 FILLER_30_1249 ();
 sg13g2_decap_4 FILLER_30_1256 ();
 sg13g2_fill_2 FILLER_30_1260 ();
 sg13g2_decap_4 FILLER_30_1272 ();
 sg13g2_decap_4 FILLER_30_1280 ();
 sg13g2_decap_4 FILLER_30_1320 ();
 sg13g2_fill_1 FILLER_30_1369 ();
 sg13g2_fill_2 FILLER_30_1390 ();
 sg13g2_fill_1 FILLER_30_1392 ();
 sg13g2_fill_1 FILLER_30_1406 ();
 sg13g2_fill_2 FILLER_30_1417 ();
 sg13g2_fill_2 FILLER_30_1424 ();
 sg13g2_fill_1 FILLER_30_1426 ();
 sg13g2_fill_1 FILLER_30_1434 ();
 sg13g2_fill_2 FILLER_30_1444 ();
 sg13g2_fill_1 FILLER_30_1460 ();
 sg13g2_fill_1 FILLER_30_1467 ();
 sg13g2_fill_1 FILLER_30_1500 ();
 sg13g2_decap_4 FILLER_30_1510 ();
 sg13g2_fill_1 FILLER_30_1514 ();
 sg13g2_fill_2 FILLER_30_1522 ();
 sg13g2_decap_8 FILLER_30_1536 ();
 sg13g2_fill_2 FILLER_30_1543 ();
 sg13g2_decap_8 FILLER_30_1555 ();
 sg13g2_decap_8 FILLER_30_1562 ();
 sg13g2_fill_2 FILLER_30_1569 ();
 sg13g2_fill_2 FILLER_30_1602 ();
 sg13g2_fill_2 FILLER_30_1617 ();
 sg13g2_fill_1 FILLER_30_1631 ();
 sg13g2_decap_4 FILLER_30_1668 ();
 sg13g2_fill_2 FILLER_30_1672 ();
 sg13g2_fill_2 FILLER_30_1684 ();
 sg13g2_fill_1 FILLER_30_1690 ();
 sg13g2_decap_8 FILLER_30_1724 ();
 sg13g2_decap_8 FILLER_30_1731 ();
 sg13g2_decap_4 FILLER_30_1738 ();
 sg13g2_fill_1 FILLER_30_1742 ();
 sg13g2_decap_8 FILLER_30_1784 ();
 sg13g2_decap_8 FILLER_30_1791 ();
 sg13g2_fill_1 FILLER_30_1798 ();
 sg13g2_fill_1 FILLER_30_1823 ();
 sg13g2_decap_4 FILLER_30_1839 ();
 sg13g2_decap_4 FILLER_30_1857 ();
 sg13g2_fill_2 FILLER_30_1861 ();
 sg13g2_decap_4 FILLER_30_1872 ();
 sg13g2_decap_8 FILLER_30_1889 ();
 sg13g2_fill_2 FILLER_30_1896 ();
 sg13g2_fill_1 FILLER_30_1898 ();
 sg13g2_fill_1 FILLER_30_1903 ();
 sg13g2_decap_4 FILLER_30_1909 ();
 sg13g2_fill_1 FILLER_30_1913 ();
 sg13g2_fill_1 FILLER_30_1920 ();
 sg13g2_decap_8 FILLER_30_1926 ();
 sg13g2_decap_8 FILLER_30_1933 ();
 sg13g2_fill_1 FILLER_30_1940 ();
 sg13g2_decap_8 FILLER_30_1981 ();
 sg13g2_decap_4 FILLER_30_2002 ();
 sg13g2_fill_1 FILLER_30_2006 ();
 sg13g2_decap_8 FILLER_30_2011 ();
 sg13g2_decap_8 FILLER_30_2018 ();
 sg13g2_decap_8 FILLER_30_2025 ();
 sg13g2_decap_8 FILLER_30_2032 ();
 sg13g2_decap_8 FILLER_30_2039 ();
 sg13g2_fill_1 FILLER_30_2079 ();
 sg13g2_fill_1 FILLER_30_2095 ();
 sg13g2_fill_2 FILLER_30_2110 ();
 sg13g2_fill_1 FILLER_30_2112 ();
 sg13g2_fill_2 FILLER_30_2134 ();
 sg13g2_fill_2 FILLER_30_2232 ();
 sg13g2_fill_1 FILLER_30_2234 ();
 sg13g2_decap_4 FILLER_30_2248 ();
 sg13g2_fill_2 FILLER_30_2252 ();
 sg13g2_fill_2 FILLER_30_2300 ();
 sg13g2_fill_1 FILLER_30_2302 ();
 sg13g2_fill_1 FILLER_30_2366 ();
 sg13g2_fill_2 FILLER_30_2371 ();
 sg13g2_decap_4 FILLER_30_2381 ();
 sg13g2_fill_1 FILLER_30_2415 ();
 sg13g2_fill_1 FILLER_30_2455 ();
 sg13g2_fill_1 FILLER_30_2499 ();
 sg13g2_decap_8 FILLER_30_2562 ();
 sg13g2_decap_8 FILLER_30_2569 ();
 sg13g2_fill_1 FILLER_30_2576 ();
 sg13g2_decap_8 FILLER_30_2580 ();
 sg13g2_decap_8 FILLER_30_2587 ();
 sg13g2_fill_2 FILLER_30_2594 ();
 sg13g2_fill_2 FILLER_30_2635 ();
 sg13g2_fill_1 FILLER_30_2637 ();
 sg13g2_decap_8 FILLER_30_2642 ();
 sg13g2_decap_8 FILLER_30_2649 ();
 sg13g2_decap_8 FILLER_30_2656 ();
 sg13g2_decap_8 FILLER_30_2663 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_13 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_87 ();
 sg13g2_decap_8 FILLER_31_94 ();
 sg13g2_decap_8 FILLER_31_101 ();
 sg13g2_decap_4 FILLER_31_108 ();
 sg13g2_fill_1 FILLER_31_112 ();
 sg13g2_decap_4 FILLER_31_135 ();
 sg13g2_decap_8 FILLER_31_149 ();
 sg13g2_fill_2 FILLER_31_156 ();
 sg13g2_fill_2 FILLER_31_182 ();
 sg13g2_fill_2 FILLER_31_241 ();
 sg13g2_fill_2 FILLER_31_262 ();
 sg13g2_fill_2 FILLER_31_274 ();
 sg13g2_fill_1 FILLER_31_276 ();
 sg13g2_fill_1 FILLER_31_309 ();
 sg13g2_fill_1 FILLER_31_336 ();
 sg13g2_fill_1 FILLER_31_341 ();
 sg13g2_fill_1 FILLER_31_347 ();
 sg13g2_fill_2 FILLER_31_388 ();
 sg13g2_fill_1 FILLER_31_390 ();
 sg13g2_fill_2 FILLER_31_395 ();
 sg13g2_fill_1 FILLER_31_427 ();
 sg13g2_fill_2 FILLER_31_438 ();
 sg13g2_fill_1 FILLER_31_445 ();
 sg13g2_fill_2 FILLER_31_450 ();
 sg13g2_fill_1 FILLER_31_470 ();
 sg13g2_fill_1 FILLER_31_476 ();
 sg13g2_decap_8 FILLER_31_485 ();
 sg13g2_decap_4 FILLER_31_492 ();
 sg13g2_fill_1 FILLER_31_496 ();
 sg13g2_fill_1 FILLER_31_503 ();
 sg13g2_fill_2 FILLER_31_539 ();
 sg13g2_fill_1 FILLER_31_586 ();
 sg13g2_fill_1 FILLER_31_601 ();
 sg13g2_fill_1 FILLER_31_607 ();
 sg13g2_fill_1 FILLER_31_612 ();
 sg13g2_decap_8 FILLER_31_617 ();
 sg13g2_fill_2 FILLER_31_624 ();
 sg13g2_fill_2 FILLER_31_630 ();
 sg13g2_fill_1 FILLER_31_632 ();
 sg13g2_fill_1 FILLER_31_638 ();
 sg13g2_fill_2 FILLER_31_645 ();
 sg13g2_fill_2 FILLER_31_651 ();
 sg13g2_fill_1 FILLER_31_665 ();
 sg13g2_fill_1 FILLER_31_675 ();
 sg13g2_fill_1 FILLER_31_695 ();
 sg13g2_fill_1 FILLER_31_765 ();
 sg13g2_decap_8 FILLER_31_770 ();
 sg13g2_decap_8 FILLER_31_791 ();
 sg13g2_decap_8 FILLER_31_798 ();
 sg13g2_decap_8 FILLER_31_805 ();
 sg13g2_decap_8 FILLER_31_812 ();
 sg13g2_decap_8 FILLER_31_819 ();
 sg13g2_decap_4 FILLER_31_826 ();
 sg13g2_fill_2 FILLER_31_838 ();
 sg13g2_fill_1 FILLER_31_840 ();
 sg13g2_fill_2 FILLER_31_871 ();
 sg13g2_fill_1 FILLER_31_873 ();
 sg13g2_fill_2 FILLER_31_910 ();
 sg13g2_fill_1 FILLER_31_916 ();
 sg13g2_decap_8 FILLER_31_934 ();
 sg13g2_fill_2 FILLER_31_941 ();
 sg13g2_fill_2 FILLER_31_950 ();
 sg13g2_fill_1 FILLER_31_967 ();
 sg13g2_fill_1 FILLER_31_994 ();
 sg13g2_decap_4 FILLER_31_1005 ();
 sg13g2_fill_2 FILLER_31_1019 ();
 sg13g2_fill_1 FILLER_31_1021 ();
 sg13g2_decap_4 FILLER_31_1026 ();
 sg13g2_fill_2 FILLER_31_1030 ();
 sg13g2_decap_4 FILLER_31_1045 ();
 sg13g2_fill_2 FILLER_31_1049 ();
 sg13g2_decap_4 FILLER_31_1055 ();
 sg13g2_fill_1 FILLER_31_1059 ();
 sg13g2_fill_2 FILLER_31_1111 ();
 sg13g2_fill_1 FILLER_31_1167 ();
 sg13g2_decap_4 FILLER_31_1211 ();
 sg13g2_decap_8 FILLER_31_1256 ();
 sg13g2_decap_4 FILLER_31_1263 ();
 sg13g2_decap_8 FILLER_31_1272 ();
 sg13g2_decap_8 FILLER_31_1279 ();
 sg13g2_decap_4 FILLER_31_1286 ();
 sg13g2_decap_4 FILLER_31_1294 ();
 sg13g2_fill_2 FILLER_31_1302 ();
 sg13g2_fill_2 FILLER_31_1314 ();
 sg13g2_fill_2 FILLER_31_1320 ();
 sg13g2_fill_1 FILLER_31_1352 ();
 sg13g2_fill_2 FILLER_31_1382 ();
 sg13g2_decap_4 FILLER_31_1394 ();
 sg13g2_fill_1 FILLER_31_1398 ();
 sg13g2_decap_4 FILLER_31_1412 ();
 sg13g2_fill_2 FILLER_31_1443 ();
 sg13g2_fill_2 FILLER_31_1450 ();
 sg13g2_fill_2 FILLER_31_1462 ();
 sg13g2_fill_2 FILLER_31_1483 ();
 sg13g2_fill_1 FILLER_31_1490 ();
 sg13g2_decap_8 FILLER_31_1496 ();
 sg13g2_decap_8 FILLER_31_1503 ();
 sg13g2_decap_8 FILLER_31_1510 ();
 sg13g2_fill_1 FILLER_31_1517 ();
 sg13g2_fill_1 FILLER_31_1553 ();
 sg13g2_fill_2 FILLER_31_1569 ();
 sg13g2_fill_2 FILLER_31_1619 ();
 sg13g2_fill_1 FILLER_31_1626 ();
 sg13g2_decap_4 FILLER_31_1635 ();
 sg13g2_fill_2 FILLER_31_1639 ();
 sg13g2_decap_4 FILLER_31_1646 ();
 sg13g2_fill_2 FILLER_31_1659 ();
 sg13g2_decap_8 FILLER_31_1667 ();
 sg13g2_fill_1 FILLER_31_1679 ();
 sg13g2_fill_2 FILLER_31_1685 ();
 sg13g2_fill_1 FILLER_31_1687 ();
 sg13g2_fill_2 FILLER_31_1706 ();
 sg13g2_fill_1 FILLER_31_1708 ();
 sg13g2_decap_8 FILLER_31_1719 ();
 sg13g2_decap_8 FILLER_31_1726 ();
 sg13g2_decap_8 FILLER_31_1733 ();
 sg13g2_fill_1 FILLER_31_1740 ();
 sg13g2_fill_2 FILLER_31_1755 ();
 sg13g2_fill_1 FILLER_31_1757 ();
 sg13g2_fill_2 FILLER_31_1789 ();
 sg13g2_decap_8 FILLER_31_1795 ();
 sg13g2_decap_4 FILLER_31_1802 ();
 sg13g2_fill_2 FILLER_31_1810 ();
 sg13g2_fill_2 FILLER_31_1815 ();
 sg13g2_fill_1 FILLER_31_1820 ();
 sg13g2_fill_2 FILLER_31_1848 ();
 sg13g2_fill_1 FILLER_31_1855 ();
 sg13g2_fill_2 FILLER_31_1861 ();
 sg13g2_fill_1 FILLER_31_1863 ();
 sg13g2_decap_8 FILLER_31_1874 ();
 sg13g2_fill_2 FILLER_31_1881 ();
 sg13g2_decap_4 FILLER_31_1913 ();
 sg13g2_fill_1 FILLER_31_1917 ();
 sg13g2_fill_2 FILLER_31_1926 ();
 sg13g2_decap_8 FILLER_31_1934 ();
 sg13g2_fill_1 FILLER_31_1993 ();
 sg13g2_fill_2 FILLER_31_2003 ();
 sg13g2_fill_1 FILLER_31_2005 ();
 sg13g2_fill_2 FILLER_31_2011 ();
 sg13g2_fill_1 FILLER_31_2013 ();
 sg13g2_fill_2 FILLER_31_2040 ();
 sg13g2_fill_2 FILLER_31_2046 ();
 sg13g2_fill_1 FILLER_31_2048 ();
 sg13g2_fill_2 FILLER_31_2098 ();
 sg13g2_fill_1 FILLER_31_2100 ();
 sg13g2_fill_2 FILLER_31_2127 ();
 sg13g2_decap_8 FILLER_31_2211 ();
 sg13g2_fill_2 FILLER_31_2218 ();
 sg13g2_fill_1 FILLER_31_2220 ();
 sg13g2_decap_4 FILLER_31_2255 ();
 sg13g2_decap_4 FILLER_31_2269 ();
 sg13g2_fill_2 FILLER_31_2273 ();
 sg13g2_decap_8 FILLER_31_2283 ();
 sg13g2_fill_1 FILLER_31_2290 ();
 sg13g2_fill_1 FILLER_31_2372 ();
 sg13g2_decap_8 FILLER_31_2397 ();
 sg13g2_decap_8 FILLER_31_2404 ();
 sg13g2_decap_4 FILLER_31_2411 ();
 sg13g2_fill_2 FILLER_31_2419 ();
 sg13g2_decap_4 FILLER_31_2424 ();
 sg13g2_fill_1 FILLER_31_2428 ();
 sg13g2_fill_2 FILLER_31_2435 ();
 sg13g2_fill_2 FILLER_31_2441 ();
 sg13g2_fill_2 FILLER_31_2468 ();
 sg13g2_fill_2 FILLER_31_2493 ();
 sg13g2_decap_8 FILLER_31_2616 ();
 sg13g2_decap_8 FILLER_31_2623 ();
 sg13g2_decap_8 FILLER_31_2630 ();
 sg13g2_decap_8 FILLER_31_2637 ();
 sg13g2_decap_8 FILLER_31_2644 ();
 sg13g2_decap_8 FILLER_31_2651 ();
 sg13g2_decap_8 FILLER_31_2658 ();
 sg13g2_decap_4 FILLER_31_2665 ();
 sg13g2_fill_1 FILLER_31_2669 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_13 ();
 sg13g2_fill_1 FILLER_32_36 ();
 sg13g2_fill_1 FILLER_32_53 ();
 sg13g2_decap_8 FILLER_32_58 ();
 sg13g2_decap_8 FILLER_32_65 ();
 sg13g2_decap_4 FILLER_32_72 ();
 sg13g2_decap_8 FILLER_32_81 ();
 sg13g2_decap_8 FILLER_32_97 ();
 sg13g2_fill_2 FILLER_32_104 ();
 sg13g2_fill_1 FILLER_32_106 ();
 sg13g2_fill_1 FILLER_32_129 ();
 sg13g2_decap_8 FILLER_32_134 ();
 sg13g2_fill_1 FILLER_32_141 ();
 sg13g2_decap_4 FILLER_32_146 ();
 sg13g2_fill_2 FILLER_32_150 ();
 sg13g2_fill_2 FILLER_32_165 ();
 sg13g2_decap_8 FILLER_32_197 ();
 sg13g2_decap_4 FILLER_32_204 ();
 sg13g2_fill_2 FILLER_32_208 ();
 sg13g2_fill_1 FILLER_32_217 ();
 sg13g2_fill_2 FILLER_32_248 ();
 sg13g2_fill_2 FILLER_32_253 ();
 sg13g2_fill_2 FILLER_32_264 ();
 sg13g2_fill_1 FILLER_32_266 ();
 sg13g2_fill_1 FILLER_32_282 ();
 sg13g2_fill_1 FILLER_32_293 ();
 sg13g2_fill_2 FILLER_32_298 ();
 sg13g2_fill_1 FILLER_32_310 ();
 sg13g2_fill_1 FILLER_32_338 ();
 sg13g2_fill_2 FILLER_32_374 ();
 sg13g2_fill_1 FILLER_32_376 ();
 sg13g2_fill_1 FILLER_32_414 ();
 sg13g2_decap_4 FILLER_32_450 ();
 sg13g2_fill_2 FILLER_32_454 ();
 sg13g2_fill_2 FILLER_32_474 ();
 sg13g2_fill_2 FILLER_32_481 ();
 sg13g2_fill_1 FILLER_32_483 ();
 sg13g2_decap_4 FILLER_32_510 ();
 sg13g2_fill_1 FILLER_32_514 ();
 sg13g2_decap_8 FILLER_32_523 ();
 sg13g2_decap_4 FILLER_32_530 ();
 sg13g2_decap_4 FILLER_32_538 ();
 sg13g2_fill_1 FILLER_32_542 ();
 sg13g2_fill_2 FILLER_32_547 ();
 sg13g2_fill_1 FILLER_32_562 ();
 sg13g2_decap_4 FILLER_32_593 ();
 sg13g2_fill_2 FILLER_32_597 ();
 sg13g2_decap_8 FILLER_32_604 ();
 sg13g2_fill_1 FILLER_32_611 ();
 sg13g2_fill_2 FILLER_32_659 ();
 sg13g2_fill_2 FILLER_32_731 ();
 sg13g2_fill_2 FILLER_32_785 ();
 sg13g2_fill_1 FILLER_32_793 ();
 sg13g2_fill_2 FILLER_32_798 ();
 sg13g2_fill_1 FILLER_32_800 ();
 sg13g2_decap_8 FILLER_32_831 ();
 sg13g2_decap_8 FILLER_32_838 ();
 sg13g2_decap_8 FILLER_32_871 ();
 sg13g2_decap_4 FILLER_32_878 ();
 sg13g2_decap_8 FILLER_32_896 ();
 sg13g2_decap_4 FILLER_32_903 ();
 sg13g2_decap_8 FILLER_32_911 ();
 sg13g2_decap_8 FILLER_32_918 ();
 sg13g2_fill_1 FILLER_32_925 ();
 sg13g2_decap_8 FILLER_32_948 ();
 sg13g2_fill_2 FILLER_32_955 ();
 sg13g2_fill_1 FILLER_32_957 ();
 sg13g2_decap_8 FILLER_32_965 ();
 sg13g2_fill_2 FILLER_32_972 ();
 sg13g2_decap_4 FILLER_32_996 ();
 sg13g2_decap_8 FILLER_32_1030 ();
 sg13g2_decap_8 FILLER_32_1037 ();
 sg13g2_fill_2 FILLER_32_1044 ();
 sg13g2_fill_2 FILLER_32_1082 ();
 sg13g2_fill_1 FILLER_32_1127 ();
 sg13g2_fill_1 FILLER_32_1160 ();
 sg13g2_fill_1 FILLER_32_1181 ();
 sg13g2_fill_1 FILLER_32_1209 ();
 sg13g2_fill_1 FILLER_32_1236 ();
 sg13g2_decap_4 FILLER_32_1263 ();
 sg13g2_fill_2 FILLER_32_1267 ();
 sg13g2_decap_8 FILLER_32_1273 ();
 sg13g2_decap_8 FILLER_32_1280 ();
 sg13g2_fill_2 FILLER_32_1359 ();
 sg13g2_fill_2 FILLER_32_1365 ();
 sg13g2_fill_1 FILLER_32_1367 ();
 sg13g2_fill_2 FILLER_32_1378 ();
 sg13g2_fill_1 FILLER_32_1380 ();
 sg13g2_fill_2 FILLER_32_1407 ();
 sg13g2_fill_1 FILLER_32_1427 ();
 sg13g2_fill_1 FILLER_32_1444 ();
 sg13g2_fill_2 FILLER_32_1450 ();
 sg13g2_fill_1 FILLER_32_1482 ();
 sg13g2_decap_4 FILLER_32_1499 ();
 sg13g2_decap_8 FILLER_32_1509 ();
 sg13g2_fill_2 FILLER_32_1516 ();
 sg13g2_fill_2 FILLER_32_1525 ();
 sg13g2_fill_2 FILLER_32_1532 ();
 sg13g2_fill_1 FILLER_32_1539 ();
 sg13g2_fill_1 FILLER_32_1557 ();
 sg13g2_decap_4 FILLER_32_1562 ();
 sg13g2_fill_1 FILLER_32_1566 ();
 sg13g2_fill_1 FILLER_32_1573 ();
 sg13g2_fill_2 FILLER_32_1624 ();
 sg13g2_fill_1 FILLER_32_1635 ();
 sg13g2_fill_2 FILLER_32_1646 ();
 sg13g2_fill_1 FILLER_32_1648 ();
 sg13g2_decap_4 FILLER_32_1685 ();
 sg13g2_fill_2 FILLER_32_1689 ();
 sg13g2_decap_8 FILLER_32_1704 ();
 sg13g2_fill_1 FILLER_32_1711 ();
 sg13g2_fill_1 FILLER_32_1778 ();
 sg13g2_fill_2 FILLER_32_1783 ();
 sg13g2_fill_1 FILLER_32_1785 ();
 sg13g2_fill_2 FILLER_32_1829 ();
 sg13g2_fill_2 FILLER_32_1857 ();
 sg13g2_fill_2 FILLER_32_1892 ();
 sg13g2_fill_2 FILLER_32_1903 ();
 sg13g2_fill_2 FILLER_32_1911 ();
 sg13g2_fill_1 FILLER_32_1913 ();
 sg13g2_fill_2 FILLER_32_1945 ();
 sg13g2_fill_2 FILLER_32_1953 ();
 sg13g2_fill_1 FILLER_32_1955 ();
 sg13g2_decap_4 FILLER_32_1960 ();
 sg13g2_fill_2 FILLER_32_1964 ();
 sg13g2_decap_8 FILLER_32_1975 ();
 sg13g2_decap_8 FILLER_32_1982 ();
 sg13g2_fill_2 FILLER_32_1993 ();
 sg13g2_fill_1 FILLER_32_1995 ();
 sg13g2_decap_8 FILLER_32_2032 ();
 sg13g2_decap_8 FILLER_32_2039 ();
 sg13g2_decap_4 FILLER_32_2046 ();
 sg13g2_fill_1 FILLER_32_2081 ();
 sg13g2_decap_8 FILLER_32_2116 ();
 sg13g2_fill_2 FILLER_32_2123 ();
 sg13g2_fill_2 FILLER_32_2128 ();
 sg13g2_fill_1 FILLER_32_2130 ();
 sg13g2_decap_4 FILLER_32_2135 ();
 sg13g2_fill_1 FILLER_32_2139 ();
 sg13g2_fill_1 FILLER_32_2148 ();
 sg13g2_fill_1 FILLER_32_2155 ();
 sg13g2_fill_1 FILLER_32_2164 ();
 sg13g2_fill_2 FILLER_32_2169 ();
 sg13g2_fill_1 FILLER_32_2175 ();
 sg13g2_decap_8 FILLER_32_2202 ();
 sg13g2_fill_2 FILLER_32_2209 ();
 sg13g2_fill_1 FILLER_32_2211 ();
 sg13g2_decap_4 FILLER_32_2216 ();
 sg13g2_decap_8 FILLER_32_2230 ();
 sg13g2_decap_4 FILLER_32_2237 ();
 sg13g2_fill_1 FILLER_32_2241 ();
 sg13g2_fill_2 FILLER_32_2294 ();
 sg13g2_decap_4 FILLER_32_2320 ();
 sg13g2_fill_1 FILLER_32_2324 ();
 sg13g2_fill_2 FILLER_32_2329 ();
 sg13g2_fill_2 FILLER_32_2349 ();
 sg13g2_fill_2 FILLER_32_2358 ();
 sg13g2_decap_8 FILLER_32_2394 ();
 sg13g2_decap_8 FILLER_32_2401 ();
 sg13g2_decap_8 FILLER_32_2408 ();
 sg13g2_decap_4 FILLER_32_2415 ();
 sg13g2_fill_1 FILLER_32_2419 ();
 sg13g2_fill_2 FILLER_32_2461 ();
 sg13g2_fill_1 FILLER_32_2463 ();
 sg13g2_fill_2 FILLER_32_2578 ();
 sg13g2_decap_8 FILLER_32_2642 ();
 sg13g2_decap_8 FILLER_32_2649 ();
 sg13g2_decap_8 FILLER_32_2656 ();
 sg13g2_decap_8 FILLER_32_2663 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_33 ();
 sg13g2_fill_2 FILLER_33_68 ();
 sg13g2_fill_1 FILLER_33_70 ();
 sg13g2_fill_1 FILLER_33_76 ();
 sg13g2_fill_2 FILLER_33_82 ();
 sg13g2_fill_2 FILLER_33_148 ();
 sg13g2_fill_1 FILLER_33_150 ();
 sg13g2_decap_4 FILLER_33_155 ();
 sg13g2_fill_2 FILLER_33_159 ();
 sg13g2_decap_4 FILLER_33_166 ();
 sg13g2_decap_4 FILLER_33_190 ();
 sg13g2_fill_1 FILLER_33_219 ();
 sg13g2_fill_2 FILLER_33_229 ();
 sg13g2_decap_4 FILLER_33_243 ();
 sg13g2_fill_2 FILLER_33_265 ();
 sg13g2_fill_1 FILLER_33_267 ();
 sg13g2_fill_1 FILLER_33_274 ();
 sg13g2_fill_1 FILLER_33_285 ();
 sg13g2_fill_1 FILLER_33_310 ();
 sg13g2_fill_2 FILLER_33_342 ();
 sg13g2_fill_1 FILLER_33_344 ();
 sg13g2_fill_1 FILLER_33_389 ();
 sg13g2_fill_1 FILLER_33_447 ();
 sg13g2_decap_8 FILLER_33_472 ();
 sg13g2_fill_2 FILLER_33_479 ();
 sg13g2_decap_8 FILLER_33_499 ();
 sg13g2_decap_4 FILLER_33_506 ();
 sg13g2_fill_2 FILLER_33_518 ();
 sg13g2_fill_1 FILLER_33_520 ();
 sg13g2_decap_8 FILLER_33_525 ();
 sg13g2_decap_8 FILLER_33_532 ();
 sg13g2_fill_2 FILLER_33_539 ();
 sg13g2_fill_1 FILLER_33_541 ();
 sg13g2_fill_2 FILLER_33_554 ();
 sg13g2_decap_8 FILLER_33_580 ();
 sg13g2_fill_1 FILLER_33_601 ();
 sg13g2_fill_2 FILLER_33_606 ();
 sg13g2_fill_1 FILLER_33_613 ();
 sg13g2_decap_4 FILLER_33_618 ();
 sg13g2_fill_2 FILLER_33_630 ();
 sg13g2_fill_1 FILLER_33_658 ();
 sg13g2_fill_1 FILLER_33_679 ();
 sg13g2_fill_1 FILLER_33_685 ();
 sg13g2_fill_1 FILLER_33_701 ();
 sg13g2_fill_1 FILLER_33_719 ();
 sg13g2_fill_1 FILLER_33_749 ();
 sg13g2_fill_2 FILLER_33_761 ();
 sg13g2_fill_1 FILLER_33_763 ();
 sg13g2_fill_1 FILLER_33_790 ();
 sg13g2_decap_8 FILLER_33_827 ();
 sg13g2_decap_8 FILLER_33_834 ();
 sg13g2_fill_2 FILLER_33_841 ();
 sg13g2_fill_2 FILLER_33_851 ();
 sg13g2_fill_1 FILLER_33_863 ();
 sg13g2_decap_8 FILLER_33_869 ();
 sg13g2_decap_4 FILLER_33_876 ();
 sg13g2_fill_1 FILLER_33_880 ();
 sg13g2_decap_4 FILLER_33_917 ();
 sg13g2_fill_2 FILLER_33_921 ();
 sg13g2_decap_8 FILLER_33_964 ();
 sg13g2_decap_8 FILLER_33_971 ();
 sg13g2_decap_4 FILLER_33_978 ();
 sg13g2_fill_1 FILLER_33_982 ();
 sg13g2_fill_1 FILLER_33_1004 ();
 sg13g2_decap_8 FILLER_33_1036 ();
 sg13g2_decap_8 FILLER_33_1043 ();
 sg13g2_fill_1 FILLER_33_1050 ();
 sg13g2_fill_1 FILLER_33_1072 ();
 sg13g2_fill_2 FILLER_33_1083 ();
 sg13g2_fill_2 FILLER_33_1090 ();
 sg13g2_decap_8 FILLER_33_1097 ();
 sg13g2_fill_2 FILLER_33_1104 ();
 sg13g2_fill_1 FILLER_33_1168 ();
 sg13g2_decap_8 FILLER_33_1287 ();
 sg13g2_decap_8 FILLER_33_1303 ();
 sg13g2_decap_4 FILLER_33_1314 ();
 sg13g2_fill_1 FILLER_33_1318 ();
 sg13g2_fill_2 FILLER_33_1324 ();
 sg13g2_fill_2 FILLER_33_1342 ();
 sg13g2_fill_2 FILLER_33_1354 ();
 sg13g2_fill_2 FILLER_33_1360 ();
 sg13g2_fill_2 FILLER_33_1388 ();
 sg13g2_decap_8 FILLER_33_1397 ();
 sg13g2_fill_2 FILLER_33_1404 ();
 sg13g2_fill_1 FILLER_33_1430 ();
 sg13g2_fill_2 FILLER_33_1443 ();
 sg13g2_fill_1 FILLER_33_1445 ();
 sg13g2_fill_1 FILLER_33_1451 ();
 sg13g2_fill_2 FILLER_33_1457 ();
 sg13g2_decap_8 FILLER_33_1468 ();
 sg13g2_fill_1 FILLER_33_1475 ();
 sg13g2_fill_2 FILLER_33_1481 ();
 sg13g2_fill_1 FILLER_33_1483 ();
 sg13g2_fill_1 FILLER_33_1504 ();
 sg13g2_decap_8 FILLER_33_1543 ();
 sg13g2_decap_8 FILLER_33_1550 ();
 sg13g2_decap_4 FILLER_33_1557 ();
 sg13g2_fill_2 FILLER_33_1561 ();
 sg13g2_fill_2 FILLER_33_1596 ();
 sg13g2_decap_8 FILLER_33_1627 ();
 sg13g2_decap_8 FILLER_33_1634 ();
 sg13g2_decap_4 FILLER_33_1641 ();
 sg13g2_fill_2 FILLER_33_1645 ();
 sg13g2_fill_2 FILLER_33_1670 ();
 sg13g2_fill_2 FILLER_33_1676 ();
 sg13g2_decap_8 FILLER_33_1696 ();
 sg13g2_decap_8 FILLER_33_1703 ();
 sg13g2_fill_2 FILLER_33_1746 ();
 sg13g2_decap_8 FILLER_33_1777 ();
 sg13g2_fill_2 FILLER_33_1798 ();
 sg13g2_fill_1 FILLER_33_1846 ();
 sg13g2_fill_2 FILLER_33_1851 ();
 sg13g2_fill_2 FILLER_33_1858 ();
 sg13g2_fill_2 FILLER_33_1866 ();
 sg13g2_decap_4 FILLER_33_1898 ();
 sg13g2_fill_1 FILLER_33_1915 ();
 sg13g2_decap_8 FILLER_33_1946 ();
 sg13g2_fill_1 FILLER_33_1957 ();
 sg13g2_fill_2 FILLER_33_1994 ();
 sg13g2_fill_2 FILLER_33_2052 ();
 sg13g2_fill_1 FILLER_33_2070 ();
 sg13g2_fill_1 FILLER_33_2096 ();
 sg13g2_fill_1 FILLER_33_2107 ();
 sg13g2_decap_4 FILLER_33_2144 ();
 sg13g2_decap_4 FILLER_33_2187 ();
 sg13g2_fill_1 FILLER_33_2199 ();
 sg13g2_fill_1 FILLER_33_2226 ();
 sg13g2_fill_2 FILLER_33_2263 ();
 sg13g2_fill_2 FILLER_33_2295 ();
 sg13g2_fill_1 FILLER_33_2297 ();
 sg13g2_decap_4 FILLER_33_2318 ();
 sg13g2_fill_2 FILLER_33_2322 ();
 sg13g2_decap_8 FILLER_33_2382 ();
 sg13g2_decap_8 FILLER_33_2389 ();
 sg13g2_fill_1 FILLER_33_2396 ();
 sg13g2_decap_8 FILLER_33_2407 ();
 sg13g2_fill_2 FILLER_33_2414 ();
 sg13g2_fill_2 FILLER_33_2462 ();
 sg13g2_fill_1 FILLER_33_2468 ();
 sg13g2_fill_1 FILLER_33_2507 ();
 sg13g2_decap_8 FILLER_33_2512 ();
 sg13g2_fill_1 FILLER_33_2519 ();
 sg13g2_fill_2 FILLER_33_2526 ();
 sg13g2_fill_2 FILLER_33_2542 ();
 sg13g2_fill_1 FILLER_33_2544 ();
 sg13g2_decap_4 FILLER_33_2620 ();
 sg13g2_decap_8 FILLER_33_2628 ();
 sg13g2_decap_8 FILLER_33_2635 ();
 sg13g2_decap_8 FILLER_33_2642 ();
 sg13g2_decap_8 FILLER_33_2649 ();
 sg13g2_decap_8 FILLER_33_2656 ();
 sg13g2_decap_8 FILLER_33_2663 ();
 sg13g2_fill_1 FILLER_34_29 ();
 sg13g2_decap_8 FILLER_34_62 ();
 sg13g2_fill_2 FILLER_34_69 ();
 sg13g2_fill_2 FILLER_34_100 ();
 sg13g2_fill_2 FILLER_34_120 ();
 sg13g2_fill_1 FILLER_34_127 ();
 sg13g2_fill_2 FILLER_34_132 ();
 sg13g2_fill_1 FILLER_34_138 ();
 sg13g2_fill_2 FILLER_34_143 ();
 sg13g2_fill_2 FILLER_34_150 ();
 sg13g2_fill_2 FILLER_34_185 ();
 sg13g2_fill_1 FILLER_34_187 ();
 sg13g2_fill_2 FILLER_34_198 ();
 sg13g2_fill_1 FILLER_34_226 ();
 sg13g2_fill_1 FILLER_34_236 ();
 sg13g2_fill_1 FILLER_34_259 ();
 sg13g2_fill_2 FILLER_34_275 ();
 sg13g2_fill_1 FILLER_34_326 ();
 sg13g2_decap_4 FILLER_34_339 ();
 sg13g2_fill_2 FILLER_34_347 ();
 sg13g2_fill_1 FILLER_34_364 ();
 sg13g2_decap_4 FILLER_34_369 ();
 sg13g2_fill_1 FILLER_34_384 ();
 sg13g2_fill_2 FILLER_34_433 ();
 sg13g2_fill_1 FILLER_34_435 ();
 sg13g2_fill_2 FILLER_34_441 ();
 sg13g2_fill_1 FILLER_34_443 ();
 sg13g2_fill_2 FILLER_34_496 ();
 sg13g2_fill_1 FILLER_34_498 ();
 sg13g2_fill_2 FILLER_34_543 ();
 sg13g2_fill_2 FILLER_34_550 ();
 sg13g2_fill_1 FILLER_34_552 ();
 sg13g2_decap_4 FILLER_34_596 ();
 sg13g2_fill_1 FILLER_34_600 ();
 sg13g2_fill_2 FILLER_34_610 ();
 sg13g2_fill_1 FILLER_34_612 ();
 sg13g2_fill_2 FILLER_34_622 ();
 sg13g2_decap_4 FILLER_34_628 ();
 sg13g2_fill_1 FILLER_34_632 ();
 sg13g2_fill_2 FILLER_34_646 ();
 sg13g2_fill_2 FILLER_34_653 ();
 sg13g2_fill_2 FILLER_34_668 ();
 sg13g2_fill_1 FILLER_34_684 ();
 sg13g2_fill_2 FILLER_34_721 ();
 sg13g2_fill_2 FILLER_34_726 ();
 sg13g2_fill_2 FILLER_34_776 ();
 sg13g2_decap_8 FILLER_34_787 ();
 sg13g2_decap_8 FILLER_34_794 ();
 sg13g2_decap_8 FILLER_34_827 ();
 sg13g2_fill_2 FILLER_34_834 ();
 sg13g2_decap_4 FILLER_34_883 ();
 sg13g2_fill_1 FILLER_34_887 ();
 sg13g2_fill_1 FILLER_34_898 ();
 sg13g2_fill_2 FILLER_34_925 ();
 sg13g2_fill_1 FILLER_34_973 ();
 sg13g2_decap_8 FILLER_34_978 ();
 sg13g2_fill_2 FILLER_34_985 ();
 sg13g2_decap_8 FILLER_34_1038 ();
 sg13g2_decap_8 FILLER_34_1045 ();
 sg13g2_fill_2 FILLER_34_1052 ();
 sg13g2_decap_8 FILLER_34_1084 ();
 sg13g2_fill_2 FILLER_34_1091 ();
 sg13g2_fill_1 FILLER_34_1133 ();
 sg13g2_decap_8 FILLER_34_1232 ();
 sg13g2_fill_2 FILLER_34_1239 ();
 sg13g2_fill_1 FILLER_34_1241 ();
 sg13g2_fill_1 FILLER_34_1278 ();
 sg13g2_decap_4 FILLER_34_1284 ();
 sg13g2_fill_1 FILLER_34_1288 ();
 sg13g2_decap_4 FILLER_34_1300 ();
 sg13g2_fill_1 FILLER_34_1304 ();
 sg13g2_fill_2 FILLER_34_1314 ();
 sg13g2_decap_4 FILLER_34_1348 ();
 sg13g2_fill_2 FILLER_34_1352 ();
 sg13g2_fill_1 FILLER_34_1393 ();
 sg13g2_fill_1 FILLER_34_1414 ();
 sg13g2_fill_1 FILLER_34_1429 ();
 sg13g2_fill_2 FILLER_34_1436 ();
 sg13g2_fill_2 FILLER_34_1453 ();
 sg13g2_fill_2 FILLER_34_1473 ();
 sg13g2_fill_1 FILLER_34_1479 ();
 sg13g2_fill_1 FILLER_34_1485 ();
 sg13g2_fill_1 FILLER_34_1495 ();
 sg13g2_fill_2 FILLER_34_1501 ();
 sg13g2_fill_1 FILLER_34_1503 ();
 sg13g2_fill_1 FILLER_34_1510 ();
 sg13g2_fill_1 FILLER_34_1533 ();
 sg13g2_fill_1 FILLER_34_1549 ();
 sg13g2_fill_1 FILLER_34_1569 ();
 sg13g2_fill_1 FILLER_34_1573 ();
 sg13g2_fill_2 FILLER_34_1587 ();
 sg13g2_fill_1 FILLER_34_1589 ();
 sg13g2_fill_2 FILLER_34_1620 ();
 sg13g2_fill_1 FILLER_34_1627 ();
 sg13g2_decap_4 FILLER_34_1700 ();
 sg13g2_decap_8 FILLER_34_1714 ();
 sg13g2_fill_1 FILLER_34_1721 ();
 sg13g2_fill_2 FILLER_34_1726 ();
 sg13g2_fill_2 FILLER_34_1742 ();
 sg13g2_fill_1 FILLER_34_1744 ();
 sg13g2_fill_1 FILLER_34_1778 ();
 sg13g2_decap_4 FILLER_34_1782 ();
 sg13g2_fill_1 FILLER_34_1820 ();
 sg13g2_decap_4 FILLER_34_1873 ();
 sg13g2_fill_2 FILLER_34_1887 ();
 sg13g2_fill_1 FILLER_34_1889 ();
 sg13g2_fill_1 FILLER_34_1896 ();
 sg13g2_fill_1 FILLER_34_1906 ();
 sg13g2_decap_8 FILLER_34_1932 ();
 sg13g2_decap_4 FILLER_34_1939 ();
 sg13g2_fill_1 FILLER_34_2011 ();
 sg13g2_fill_1 FILLER_34_2016 ();
 sg13g2_fill_1 FILLER_34_2042 ();
 sg13g2_fill_2 FILLER_34_2047 ();
 sg13g2_fill_1 FILLER_34_2049 ();
 sg13g2_fill_1 FILLER_34_2074 ();
 sg13g2_fill_1 FILLER_34_2081 ();
 sg13g2_decap_4 FILLER_34_2091 ();
 sg13g2_fill_2 FILLER_34_2128 ();
 sg13g2_decap_4 FILLER_34_2189 ();
 sg13g2_fill_2 FILLER_34_2193 ();
 sg13g2_fill_2 FILLER_34_2199 ();
 sg13g2_fill_1 FILLER_34_2206 ();
 sg13g2_fill_1 FILLER_34_2233 ();
 sg13g2_decap_8 FILLER_34_2238 ();
 sg13g2_decap_4 FILLER_34_2245 ();
 sg13g2_fill_2 FILLER_34_2249 ();
 sg13g2_decap_8 FILLER_34_2282 ();
 sg13g2_decap_8 FILLER_34_2289 ();
 sg13g2_fill_1 FILLER_34_2300 ();
 sg13g2_decap_4 FILLER_34_2345 ();
 sg13g2_fill_1 FILLER_34_2362 ();
 sg13g2_fill_2 FILLER_34_2367 ();
 sg13g2_fill_1 FILLER_34_2369 ();
 sg13g2_fill_1 FILLER_34_2380 ();
 sg13g2_fill_1 FILLER_34_2391 ();
 sg13g2_fill_2 FILLER_34_2401 ();
 sg13g2_fill_2 FILLER_34_2441 ();
 sg13g2_decap_8 FILLER_34_2469 ();
 sg13g2_decap_4 FILLER_34_2476 ();
 sg13g2_fill_2 FILLER_34_2492 ();
 sg13g2_fill_2 FILLER_34_2534 ();
 sg13g2_fill_1 FILLER_34_2573 ();
 sg13g2_fill_1 FILLER_34_2584 ();
 sg13g2_fill_2 FILLER_34_2598 ();
 sg13g2_decap_8 FILLER_34_2607 ();
 sg13g2_decap_8 FILLER_34_2614 ();
 sg13g2_decap_8 FILLER_34_2621 ();
 sg13g2_decap_8 FILLER_34_2628 ();
 sg13g2_decap_8 FILLER_34_2635 ();
 sg13g2_decap_8 FILLER_34_2642 ();
 sg13g2_decap_8 FILLER_34_2649 ();
 sg13g2_decap_8 FILLER_34_2656 ();
 sg13g2_decap_8 FILLER_34_2663 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_2 ();
 sg13g2_fill_1 FILLER_35_25 ();
 sg13g2_fill_2 FILLER_35_57 ();
 sg13g2_fill_1 FILLER_35_59 ();
 sg13g2_fill_1 FILLER_35_75 ();
 sg13g2_fill_2 FILLER_35_81 ();
 sg13g2_fill_1 FILLER_35_101 ();
 sg13g2_fill_2 FILLER_35_159 ();
 sg13g2_fill_2 FILLER_35_165 ();
 sg13g2_fill_1 FILLER_35_167 ();
 sg13g2_fill_2 FILLER_35_218 ();
 sg13g2_fill_2 FILLER_35_249 ();
 sg13g2_fill_1 FILLER_35_259 ();
 sg13g2_decap_4 FILLER_35_264 ();
 sg13g2_fill_2 FILLER_35_268 ();
 sg13g2_fill_2 FILLER_35_275 ();
 sg13g2_fill_1 FILLER_35_277 ();
 sg13g2_fill_1 FILLER_35_282 ();
 sg13g2_fill_1 FILLER_35_299 ();
 sg13g2_fill_1 FILLER_35_305 ();
 sg13g2_fill_2 FILLER_35_341 ();
 sg13g2_fill_1 FILLER_35_343 ();
 sg13g2_decap_4 FILLER_35_359 ();
 sg13g2_fill_1 FILLER_35_363 ();
 sg13g2_fill_2 FILLER_35_371 ();
 sg13g2_fill_2 FILLER_35_405 ();
 sg13g2_fill_2 FILLER_35_419 ();
 sg13g2_fill_2 FILLER_35_431 ();
 sg13g2_fill_2 FILLER_35_451 ();
 sg13g2_fill_1 FILLER_35_453 ();
 sg13g2_fill_2 FILLER_35_459 ();
 sg13g2_fill_1 FILLER_35_465 ();
 sg13g2_fill_1 FILLER_35_470 ();
 sg13g2_fill_2 FILLER_35_475 ();
 sg13g2_fill_2 FILLER_35_481 ();
 sg13g2_fill_1 FILLER_35_488 ();
 sg13g2_fill_1 FILLER_35_506 ();
 sg13g2_fill_2 FILLER_35_512 ();
 sg13g2_decap_4 FILLER_35_566 ();
 sg13g2_fill_1 FILLER_35_570 ();
 sg13g2_decap_4 FILLER_35_605 ();
 sg13g2_fill_1 FILLER_35_609 ();
 sg13g2_fill_2 FILLER_35_615 ();
 sg13g2_fill_1 FILLER_35_617 ();
 sg13g2_decap_4 FILLER_35_635 ();
 sg13g2_fill_1 FILLER_35_643 ();
 sg13g2_decap_4 FILLER_35_676 ();
 sg13g2_fill_1 FILLER_35_716 ();
 sg13g2_fill_1 FILLER_35_731 ();
 sg13g2_fill_1 FILLER_35_743 ();
 sg13g2_fill_1 FILLER_35_752 ();
 sg13g2_fill_2 FILLER_35_772 ();
 sg13g2_fill_1 FILLER_35_774 ();
 sg13g2_decap_8 FILLER_35_800 ();
 sg13g2_decap_8 FILLER_35_811 ();
 sg13g2_decap_8 FILLER_35_818 ();
 sg13g2_decap_8 FILLER_35_825 ();
 sg13g2_fill_2 FILLER_35_832 ();
 sg13g2_fill_2 FILLER_35_864 ();
 sg13g2_fill_1 FILLER_35_866 ();
 sg13g2_decap_4 FILLER_35_893 ();
 sg13g2_fill_1 FILLER_35_901 ();
 sg13g2_fill_2 FILLER_35_938 ();
 sg13g2_decap_4 FILLER_35_987 ();
 sg13g2_fill_2 FILLER_35_991 ();
 sg13g2_fill_1 FILLER_35_1008 ();
 sg13g2_decap_8 FILLER_35_1035 ();
 sg13g2_decap_4 FILLER_35_1089 ();
 sg13g2_fill_1 FILLER_35_1093 ();
 sg13g2_fill_2 FILLER_35_1123 ();
 sg13g2_fill_1 FILLER_35_1161 ();
 sg13g2_fill_2 FILLER_35_1168 ();
 sg13g2_fill_2 FILLER_35_1180 ();
 sg13g2_fill_2 FILLER_35_1192 ();
 sg13g2_decap_8 FILLER_35_1220 ();
 sg13g2_decap_4 FILLER_35_1227 ();
 sg13g2_fill_1 FILLER_35_1231 ();
 sg13g2_decap_8 FILLER_35_1236 ();
 sg13g2_decap_4 FILLER_35_1243 ();
 sg13g2_fill_2 FILLER_35_1273 ();
 sg13g2_fill_1 FILLER_35_1275 ();
 sg13g2_decap_8 FILLER_35_1320 ();
 sg13g2_decap_4 FILLER_35_1327 ();
 sg13g2_fill_2 FILLER_35_1331 ();
 sg13g2_decap_8 FILLER_35_1338 ();
 sg13g2_fill_1 FILLER_35_1345 ();
 sg13g2_decap_4 FILLER_35_1360 ();
 sg13g2_fill_2 FILLER_35_1406 ();
 sg13g2_fill_2 FILLER_35_1425 ();
 sg13g2_fill_1 FILLER_35_1427 ();
 sg13g2_fill_1 FILLER_35_1432 ();
 sg13g2_decap_8 FILLER_35_1447 ();
 sg13g2_fill_2 FILLER_35_1454 ();
 sg13g2_fill_1 FILLER_35_1461 ();
 sg13g2_fill_1 FILLER_35_1466 ();
 sg13g2_fill_1 FILLER_35_1472 ();
 sg13g2_fill_1 FILLER_35_1484 ();
 sg13g2_fill_1 FILLER_35_1488 ();
 sg13g2_fill_2 FILLER_35_1510 ();
 sg13g2_fill_2 FILLER_35_1542 ();
 sg13g2_fill_1 FILLER_35_1549 ();
 sg13g2_fill_2 FILLER_35_1554 ();
 sg13g2_fill_1 FILLER_35_1560 ();
 sg13g2_fill_1 FILLER_35_1617 ();
 sg13g2_decap_4 FILLER_35_1627 ();
 sg13g2_fill_1 FILLER_35_1631 ();
 sg13g2_fill_1 FILLER_35_1648 ();
 sg13g2_fill_1 FILLER_35_1654 ();
 sg13g2_fill_1 FILLER_35_1660 ();
 sg13g2_fill_2 FILLER_35_1666 ();
 sg13g2_fill_1 FILLER_35_1668 ();
 sg13g2_decap_4 FILLER_35_1692 ();
 sg13g2_fill_2 FILLER_35_1696 ();
 sg13g2_fill_2 FILLER_35_1702 ();
 sg13g2_fill_2 FILLER_35_1730 ();
 sg13g2_decap_4 FILLER_35_1766 ();
 sg13g2_fill_2 FILLER_35_1826 ();
 sg13g2_fill_2 FILLER_35_1840 ();
 sg13g2_fill_1 FILLER_35_1880 ();
 sg13g2_fill_1 FILLER_35_1886 ();
 sg13g2_fill_2 FILLER_35_1891 ();
 sg13g2_fill_2 FILLER_35_1911 ();
 sg13g2_fill_1 FILLER_35_1947 ();
 sg13g2_fill_1 FILLER_35_1958 ();
 sg13g2_fill_2 FILLER_35_1969 ();
 sg13g2_fill_1 FILLER_35_1971 ();
 sg13g2_decap_8 FILLER_35_1977 ();
 sg13g2_decap_8 FILLER_35_1984 ();
 sg13g2_fill_2 FILLER_35_1991 ();
 sg13g2_fill_1 FILLER_35_1993 ();
 sg13g2_decap_4 FILLER_35_2004 ();
 sg13g2_decap_4 FILLER_35_2024 ();
 sg13g2_fill_1 FILLER_35_2028 ();
 sg13g2_fill_1 FILLER_35_2045 ();
 sg13g2_fill_1 FILLER_35_2072 ();
 sg13g2_fill_2 FILLER_35_2099 ();
 sg13g2_fill_1 FILLER_35_2101 ();
 sg13g2_fill_1 FILLER_35_2106 ();
 sg13g2_fill_1 FILLER_35_2165 ();
 sg13g2_fill_2 FILLER_35_2182 ();
 sg13g2_fill_1 FILLER_35_2192 ();
 sg13g2_decap_8 FILLER_35_2234 ();
 sg13g2_fill_2 FILLER_35_2258 ();
 sg13g2_fill_1 FILLER_35_2260 ();
 sg13g2_fill_1 FILLER_35_2274 ();
 sg13g2_fill_1 FILLER_35_2280 ();
 sg13g2_decap_8 FILLER_35_2285 ();
 sg13g2_fill_1 FILLER_35_2292 ();
 sg13g2_fill_1 FILLER_35_2301 ();
 sg13g2_decap_8 FILLER_35_2306 ();
 sg13g2_fill_1 FILLER_35_2323 ();
 sg13g2_fill_1 FILLER_35_2350 ();
 sg13g2_fill_1 FILLER_35_2355 ();
 sg13g2_fill_1 FILLER_35_2382 ();
 sg13g2_fill_2 FILLER_35_2409 ();
 sg13g2_fill_1 FILLER_35_2477 ();
 sg13g2_fill_1 FILLER_35_2482 ();
 sg13g2_fill_1 FILLER_35_2550 ();
 sg13g2_fill_1 FILLER_35_2588 ();
 sg13g2_decap_8 FILLER_35_2625 ();
 sg13g2_decap_8 FILLER_35_2632 ();
 sg13g2_decap_8 FILLER_35_2639 ();
 sg13g2_decap_8 FILLER_35_2646 ();
 sg13g2_decap_8 FILLER_35_2653 ();
 sg13g2_decap_8 FILLER_35_2660 ();
 sg13g2_fill_2 FILLER_35_2667 ();
 sg13g2_fill_1 FILLER_35_2669 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_49 ();
 sg13g2_fill_2 FILLER_36_59 ();
 sg13g2_fill_2 FILLER_36_80 ();
 sg13g2_fill_2 FILLER_36_90 ();
 sg13g2_decap_8 FILLER_36_102 ();
 sg13g2_fill_2 FILLER_36_109 ();
 sg13g2_fill_1 FILLER_36_135 ();
 sg13g2_fill_1 FILLER_36_144 ();
 sg13g2_decap_4 FILLER_36_166 ();
 sg13g2_fill_2 FILLER_36_170 ();
 sg13g2_fill_1 FILLER_36_193 ();
 sg13g2_fill_1 FILLER_36_210 ();
 sg13g2_fill_1 FILLER_36_253 ();
 sg13g2_fill_1 FILLER_36_259 ();
 sg13g2_fill_1 FILLER_36_268 ();
 sg13g2_decap_4 FILLER_36_277 ();
 sg13g2_fill_2 FILLER_36_307 ();
 sg13g2_fill_1 FILLER_36_316 ();
 sg13g2_decap_4 FILLER_36_347 ();
 sg13g2_fill_2 FILLER_36_377 ();
 sg13g2_fill_2 FILLER_36_389 ();
 sg13g2_fill_1 FILLER_36_451 ();
 sg13g2_fill_2 FILLER_36_458 ();
 sg13g2_fill_1 FILLER_36_460 ();
 sg13g2_decap_4 FILLER_36_467 ();
 sg13g2_fill_2 FILLER_36_471 ();
 sg13g2_fill_1 FILLER_36_482 ();
 sg13g2_fill_1 FILLER_36_508 ();
 sg13g2_decap_8 FILLER_36_514 ();
 sg13g2_fill_2 FILLER_36_521 ();
 sg13g2_fill_1 FILLER_36_523 ();
 sg13g2_fill_1 FILLER_36_539 ();
 sg13g2_fill_1 FILLER_36_555 ();
 sg13g2_fill_2 FILLER_36_563 ();
 sg13g2_fill_2 FILLER_36_569 ();
 sg13g2_fill_1 FILLER_36_576 ();
 sg13g2_decap_4 FILLER_36_581 ();
 sg13g2_fill_1 FILLER_36_585 ();
 sg13g2_fill_1 FILLER_36_593 ();
 sg13g2_decap_8 FILLER_36_598 ();
 sg13g2_fill_2 FILLER_36_605 ();
 sg13g2_fill_1 FILLER_36_607 ();
 sg13g2_fill_2 FILLER_36_627 ();
 sg13g2_fill_2 FILLER_36_643 ();
 sg13g2_fill_1 FILLER_36_649 ();
 sg13g2_fill_1 FILLER_36_654 ();
 sg13g2_fill_2 FILLER_36_703 ();
 sg13g2_fill_1 FILLER_36_715 ();
 sg13g2_fill_1 FILLER_36_722 ();
 sg13g2_fill_2 FILLER_36_739 ();
 sg13g2_fill_1 FILLER_36_741 ();
 sg13g2_fill_2 FILLER_36_752 ();
 sg13g2_fill_2 FILLER_36_765 ();
 sg13g2_fill_1 FILLER_36_767 ();
 sg13g2_fill_1 FILLER_36_773 ();
 sg13g2_fill_1 FILLER_36_779 ();
 sg13g2_fill_2 FILLER_36_816 ();
 sg13g2_fill_1 FILLER_36_818 ();
 sg13g2_decap_8 FILLER_36_823 ();
 sg13g2_fill_2 FILLER_36_830 ();
 sg13g2_fill_1 FILLER_36_832 ();
 sg13g2_fill_2 FILLER_36_869 ();
 sg13g2_fill_2 FILLER_36_911 ();
 sg13g2_decap_8 FILLER_36_956 ();
 sg13g2_decap_4 FILLER_36_963 ();
 sg13g2_fill_2 FILLER_36_967 ();
 sg13g2_fill_1 FILLER_36_995 ();
 sg13g2_fill_2 FILLER_36_1011 ();
 sg13g2_fill_1 FILLER_36_1013 ();
 sg13g2_decap_4 FILLER_36_1028 ();
 sg13g2_fill_2 FILLER_36_1032 ();
 sg13g2_fill_2 FILLER_36_1124 ();
 sg13g2_fill_1 FILLER_36_1178 ();
 sg13g2_decap_4 FILLER_36_1210 ();
 sg13g2_fill_2 FILLER_36_1214 ();
 sg13g2_decap_8 FILLER_36_1223 ();
 sg13g2_fill_2 FILLER_36_1230 ();
 sg13g2_fill_1 FILLER_36_1232 ();
 sg13g2_decap_4 FILLER_36_1241 ();
 sg13g2_fill_2 FILLER_36_1245 ();
 sg13g2_fill_1 FILLER_36_1251 ();
 sg13g2_fill_1 FILLER_36_1256 ();
 sg13g2_fill_2 FILLER_36_1287 ();
 sg13g2_decap_8 FILLER_36_1292 ();
 sg13g2_fill_1 FILLER_36_1299 ();
 sg13g2_fill_2 FILLER_36_1304 ();
 sg13g2_fill_2 FILLER_36_1311 ();
 sg13g2_decap_8 FILLER_36_1317 ();
 sg13g2_decap_4 FILLER_36_1324 ();
 sg13g2_fill_2 FILLER_36_1332 ();
 sg13g2_fill_2 FILLER_36_1382 ();
 sg13g2_fill_1 FILLER_36_1407 ();
 sg13g2_fill_2 FILLER_36_1473 ();
 sg13g2_fill_1 FILLER_36_1475 ();
 sg13g2_fill_2 FILLER_36_1479 ();
 sg13g2_fill_2 FILLER_36_1512 ();
 sg13g2_fill_2 FILLER_36_1518 ();
 sg13g2_fill_2 FILLER_36_1529 ();
 sg13g2_fill_1 FILLER_36_1553 ();
 sg13g2_fill_2 FILLER_36_1580 ();
 sg13g2_decap_4 FILLER_36_1587 ();
 sg13g2_fill_2 FILLER_36_1599 ();
 sg13g2_fill_1 FILLER_36_1601 ();
 sg13g2_decap_4 FILLER_36_1612 ();
 sg13g2_fill_1 FILLER_36_1616 ();
 sg13g2_fill_1 FILLER_36_1635 ();
 sg13g2_decap_4 FILLER_36_1659 ();
 sg13g2_fill_1 FILLER_36_1663 ();
 sg13g2_decap_4 FILLER_36_1669 ();
 sg13g2_fill_2 FILLER_36_1673 ();
 sg13g2_fill_1 FILLER_36_1694 ();
 sg13g2_fill_1 FILLER_36_1705 ();
 sg13g2_decap_4 FILLER_36_1740 ();
 sg13g2_fill_1 FILLER_36_1744 ();
 sg13g2_fill_2 FILLER_36_1782 ();
 sg13g2_fill_1 FILLER_36_1793 ();
 sg13g2_fill_1 FILLER_36_1799 ();
 sg13g2_decap_8 FILLER_36_1828 ();
 sg13g2_decap_4 FILLER_36_1835 ();
 sg13g2_fill_2 FILLER_36_1839 ();
 sg13g2_decap_4 FILLER_36_1845 ();
 sg13g2_fill_1 FILLER_36_1849 ();
 sg13g2_fill_1 FILLER_36_1854 ();
 sg13g2_fill_1 FILLER_36_1859 ();
 sg13g2_fill_1 FILLER_36_1886 ();
 sg13g2_fill_1 FILLER_36_1913 ();
 sg13g2_decap_8 FILLER_36_1930 ();
 sg13g2_decap_4 FILLER_36_1937 ();
 sg13g2_fill_2 FILLER_36_1964 ();
 sg13g2_fill_1 FILLER_36_1966 ();
 sg13g2_decap_4 FILLER_36_1976 ();
 sg13g2_decap_4 FILLER_36_2000 ();
 sg13g2_decap_8 FILLER_36_2008 ();
 sg13g2_decap_8 FILLER_36_2015 ();
 sg13g2_decap_8 FILLER_36_2026 ();
 sg13g2_fill_2 FILLER_36_2033 ();
 sg13g2_fill_1 FILLER_36_2035 ();
 sg13g2_fill_2 FILLER_36_2047 ();
 sg13g2_decap_4 FILLER_36_2083 ();
 sg13g2_fill_2 FILLER_36_2126 ();
 sg13g2_fill_1 FILLER_36_2142 ();
 sg13g2_fill_1 FILLER_36_2172 ();
 sg13g2_fill_2 FILLER_36_2194 ();
 sg13g2_fill_2 FILLER_36_2217 ();
 sg13g2_fill_1 FILLER_36_2219 ();
 sg13g2_decap_8 FILLER_36_2234 ();
 sg13g2_fill_2 FILLER_36_2254 ();
 sg13g2_decap_4 FILLER_36_2292 ();
 sg13g2_fill_2 FILLER_36_2317 ();
 sg13g2_fill_1 FILLER_36_2319 ();
 sg13g2_fill_2 FILLER_36_2417 ();
 sg13g2_fill_2 FILLER_36_2445 ();
 sg13g2_fill_1 FILLER_36_2447 ();
 sg13g2_fill_2 FILLER_36_2474 ();
 sg13g2_fill_1 FILLER_36_2476 ();
 sg13g2_decap_4 FILLER_36_2481 ();
 sg13g2_fill_1 FILLER_36_2485 ();
 sg13g2_fill_2 FILLER_36_2496 ();
 sg13g2_fill_1 FILLER_36_2528 ();
 sg13g2_fill_1 FILLER_36_2539 ();
 sg13g2_fill_1 FILLER_36_2546 ();
 sg13g2_fill_2 FILLER_36_2581 ();
 sg13g2_decap_8 FILLER_36_2623 ();
 sg13g2_decap_8 FILLER_36_2630 ();
 sg13g2_decap_8 FILLER_36_2637 ();
 sg13g2_decap_8 FILLER_36_2644 ();
 sg13g2_decap_8 FILLER_36_2651 ();
 sg13g2_decap_8 FILLER_36_2658 ();
 sg13g2_decap_4 FILLER_36_2665 ();
 sg13g2_fill_1 FILLER_36_2669 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_4 FILLER_37_14 ();
 sg13g2_fill_2 FILLER_37_55 ();
 sg13g2_fill_1 FILLER_37_62 ();
 sg13g2_fill_1 FILLER_37_73 ();
 sg13g2_decap_8 FILLER_37_78 ();
 sg13g2_fill_2 FILLER_37_85 ();
 sg13g2_fill_1 FILLER_37_87 ();
 sg13g2_decap_4 FILLER_37_93 ();
 sg13g2_fill_1 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_172 ();
 sg13g2_fill_2 FILLER_37_179 ();
 sg13g2_fill_1 FILLER_37_181 ();
 sg13g2_fill_1 FILLER_37_213 ();
 sg13g2_fill_1 FILLER_37_240 ();
 sg13g2_decap_4 FILLER_37_272 ();
 sg13g2_fill_1 FILLER_37_276 ();
 sg13g2_fill_2 FILLER_37_286 ();
 sg13g2_fill_2 FILLER_37_350 ();
 sg13g2_fill_1 FILLER_37_365 ();
 sg13g2_fill_2 FILLER_37_376 ();
 sg13g2_fill_1 FILLER_37_395 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_2 FILLER_37_417 ();
 sg13g2_fill_2 FILLER_37_449 ();
 sg13g2_fill_1 FILLER_37_455 ();
 sg13g2_decap_8 FILLER_37_460 ();
 sg13g2_fill_2 FILLER_37_498 ();
 sg13g2_fill_1 FILLER_37_500 ();
 sg13g2_fill_2 FILLER_37_505 ();
 sg13g2_fill_1 FILLER_37_516 ();
 sg13g2_fill_1 FILLER_37_521 ();
 sg13g2_fill_1 FILLER_37_526 ();
 sg13g2_fill_2 FILLER_37_532 ();
 sg13g2_fill_1 FILLER_37_534 ();
 sg13g2_decap_4 FILLER_37_565 ();
 sg13g2_fill_2 FILLER_37_569 ();
 sg13g2_decap_4 FILLER_37_587 ();
 sg13g2_fill_1 FILLER_37_591 ();
 sg13g2_decap_4 FILLER_37_600 ();
 sg13g2_fill_1 FILLER_37_604 ();
 sg13g2_fill_2 FILLER_37_636 ();
 sg13g2_fill_2 FILLER_37_647 ();
 sg13g2_fill_1 FILLER_37_649 ();
 sg13g2_fill_1 FILLER_37_655 ();
 sg13g2_fill_2 FILLER_37_661 ();
 sg13g2_fill_2 FILLER_37_667 ();
 sg13g2_fill_1 FILLER_37_669 ();
 sg13g2_fill_2 FILLER_37_675 ();
 sg13g2_fill_1 FILLER_37_677 ();
 sg13g2_fill_1 FILLER_37_688 ();
 sg13g2_fill_1 FILLER_37_699 ();
 sg13g2_decap_8 FILLER_37_704 ();
 sg13g2_decap_8 FILLER_37_711 ();
 sg13g2_decap_4 FILLER_37_718 ();
 sg13g2_fill_2 FILLER_37_768 ();
 sg13g2_fill_1 FILLER_37_770 ();
 sg13g2_fill_1 FILLER_37_775 ();
 sg13g2_fill_1 FILLER_37_781 ();
 sg13g2_fill_2 FILLER_37_786 ();
 sg13g2_fill_2 FILLER_37_798 ();
 sg13g2_fill_2 FILLER_37_810 ();
 sg13g2_decap_8 FILLER_37_838 ();
 sg13g2_decap_4 FILLER_37_845 ();
 sg13g2_decap_4 FILLER_37_853 ();
 sg13g2_decap_8 FILLER_37_871 ();
 sg13g2_fill_1 FILLER_37_878 ();
 sg13g2_decap_8 FILLER_37_897 ();
 sg13g2_decap_4 FILLER_37_904 ();
 sg13g2_decap_8 FILLER_37_916 ();
 sg13g2_fill_2 FILLER_37_923 ();
 sg13g2_fill_1 FILLER_37_991 ();
 sg13g2_decap_8 FILLER_37_1018 ();
 sg13g2_fill_1 FILLER_37_1025 ();
 sg13g2_fill_1 FILLER_37_1171 ();
 sg13g2_fill_1 FILLER_37_1178 ();
 sg13g2_fill_2 FILLER_37_1219 ();
 sg13g2_decap_4 FILLER_37_1300 ();
 sg13g2_decap_8 FILLER_37_1330 ();
 sg13g2_fill_1 FILLER_37_1337 ();
 sg13g2_fill_2 FILLER_37_1374 ();
 sg13g2_fill_2 FILLER_37_1416 ();
 sg13g2_fill_2 FILLER_37_1438 ();
 sg13g2_fill_2 FILLER_37_1527 ();
 sg13g2_fill_2 FILLER_37_1578 ();
 sg13g2_fill_2 FILLER_37_1591 ();
 sg13g2_fill_1 FILLER_37_1593 ();
 sg13g2_decap_8 FILLER_37_1608 ();
 sg13g2_fill_2 FILLER_37_1615 ();
 sg13g2_fill_2 FILLER_37_1621 ();
 sg13g2_fill_1 FILLER_37_1633 ();
 sg13g2_fill_2 FILLER_37_1649 ();
 sg13g2_fill_1 FILLER_37_1651 ();
 sg13g2_fill_2 FILLER_37_1662 ();
 sg13g2_fill_1 FILLER_37_1669 ();
 sg13g2_decap_8 FILLER_37_1685 ();
 sg13g2_fill_2 FILLER_37_1692 ();
 sg13g2_fill_1 FILLER_37_1694 ();
 sg13g2_fill_2 FILLER_37_1705 ();
 sg13g2_fill_2 FILLER_37_1727 ();
 sg13g2_decap_4 FILLER_37_1758 ();
 sg13g2_fill_1 FILLER_37_1762 ();
 sg13g2_fill_1 FILLER_37_1778 ();
 sg13g2_decap_4 FILLER_37_1828 ();
 sg13g2_decap_4 FILLER_37_1889 ();
 sg13g2_fill_2 FILLER_37_1893 ();
 sg13g2_decap_4 FILLER_37_1899 ();
 sg13g2_fill_1 FILLER_37_1913 ();
 sg13g2_decap_8 FILLER_37_1932 ();
 sg13g2_decap_8 FILLER_37_1943 ();
 sg13g2_fill_2 FILLER_37_1950 ();
 sg13g2_fill_1 FILLER_37_1952 ();
 sg13g2_fill_1 FILLER_37_1983 ();
 sg13g2_decap_8 FILLER_37_2014 ();
 sg13g2_decap_8 FILLER_37_2021 ();
 sg13g2_decap_4 FILLER_37_2028 ();
 sg13g2_fill_2 FILLER_37_2072 ();
 sg13g2_fill_2 FILLER_37_2087 ();
 sg13g2_fill_2 FILLER_37_2115 ();
 sg13g2_fill_2 FILLER_37_2144 ();
 sg13g2_fill_2 FILLER_37_2155 ();
 sg13g2_decap_8 FILLER_37_2203 ();
 sg13g2_fill_2 FILLER_37_2210 ();
 sg13g2_decap_4 FILLER_37_2228 ();
 sg13g2_fill_2 FILLER_37_2232 ();
 sg13g2_decap_4 FILLER_37_2270 ();
 sg13g2_decap_4 FILLER_37_2314 ();
 sg13g2_fill_2 FILLER_37_2328 ();
 sg13g2_decap_4 FILLER_37_2369 ();
 sg13g2_decap_4 FILLER_37_2408 ();
 sg13g2_decap_8 FILLER_37_2459 ();
 sg13g2_fill_2 FILLER_37_2466 ();
 sg13g2_decap_4 FILLER_37_2488 ();
 sg13g2_fill_2 FILLER_37_2513 ();
 sg13g2_fill_2 FILLER_37_2530 ();
 sg13g2_fill_2 FILLER_37_2565 ();
 sg13g2_fill_2 FILLER_37_2598 ();
 sg13g2_decap_8 FILLER_37_2630 ();
 sg13g2_decap_8 FILLER_37_2637 ();
 sg13g2_decap_8 FILLER_37_2644 ();
 sg13g2_decap_8 FILLER_37_2651 ();
 sg13g2_decap_8 FILLER_37_2658 ();
 sg13g2_decap_4 FILLER_37_2665 ();
 sg13g2_fill_1 FILLER_37_2669 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_fill_1 FILLER_38_14 ();
 sg13g2_fill_1 FILLER_38_58 ();
 sg13g2_fill_2 FILLER_38_100 ();
 sg13g2_fill_2 FILLER_38_108 ();
 sg13g2_decap_8 FILLER_38_177 ();
 sg13g2_decap_8 FILLER_38_184 ();
 sg13g2_decap_4 FILLER_38_191 ();
 sg13g2_fill_1 FILLER_38_215 ();
 sg13g2_fill_1 FILLER_38_241 ();
 sg13g2_fill_1 FILLER_38_272 ();
 sg13g2_fill_1 FILLER_38_279 ();
 sg13g2_fill_1 FILLER_38_286 ();
 sg13g2_decap_4 FILLER_38_324 ();
 sg13g2_fill_1 FILLER_38_328 ();
 sg13g2_decap_8 FILLER_38_333 ();
 sg13g2_decap_8 FILLER_38_340 ();
 sg13g2_fill_2 FILLER_38_358 ();
 sg13g2_fill_2 FILLER_38_363 ();
 sg13g2_decap_4 FILLER_38_447 ();
 sg13g2_fill_1 FILLER_38_456 ();
 sg13g2_fill_1 FILLER_38_504 ();
 sg13g2_fill_1 FILLER_38_526 ();
 sg13g2_decap_4 FILLER_38_533 ();
 sg13g2_fill_2 FILLER_38_537 ();
 sg13g2_fill_1 FILLER_38_543 ();
 sg13g2_fill_1 FILLER_38_554 ();
 sg13g2_fill_1 FILLER_38_570 ();
 sg13g2_decap_8 FILLER_38_585 ();
 sg13g2_decap_4 FILLER_38_592 ();
 sg13g2_fill_2 FILLER_38_596 ();
 sg13g2_fill_2 FILLER_38_624 ();
 sg13g2_fill_1 FILLER_38_626 ();
 sg13g2_fill_1 FILLER_38_637 ();
 sg13g2_fill_1 FILLER_38_687 ();
 sg13g2_decap_4 FILLER_38_719 ();
 sg13g2_fill_2 FILLER_38_723 ();
 sg13g2_fill_1 FILLER_38_729 ();
 sg13g2_fill_1 FILLER_38_808 ();
 sg13g2_decap_8 FILLER_38_835 ();
 sg13g2_decap_8 FILLER_38_842 ();
 sg13g2_fill_1 FILLER_38_849 ();
 sg13g2_fill_1 FILLER_38_854 ();
 sg13g2_fill_2 FILLER_38_859 ();
 sg13g2_decap_8 FILLER_38_865 ();
 sg13g2_decap_8 FILLER_38_872 ();
 sg13g2_decap_8 FILLER_38_879 ();
 sg13g2_decap_4 FILLER_38_896 ();
 sg13g2_decap_4 FILLER_38_934 ();
 sg13g2_fill_2 FILLER_38_942 ();
 sg13g2_fill_2 FILLER_38_957 ();
 sg13g2_fill_2 FILLER_38_1000 ();
 sg13g2_decap_8 FILLER_38_1006 ();
 sg13g2_fill_2 FILLER_38_1013 ();
 sg13g2_decap_8 FILLER_38_1019 ();
 sg13g2_decap_8 FILLER_38_1026 ();
 sg13g2_decap_8 FILLER_38_1033 ();
 sg13g2_decap_4 FILLER_38_1040 ();
 sg13g2_fill_1 FILLER_38_1044 ();
 sg13g2_decap_8 FILLER_38_1076 ();
 sg13g2_fill_2 FILLER_38_1083 ();
 sg13g2_fill_1 FILLER_38_1085 ();
 sg13g2_fill_2 FILLER_38_1090 ();
 sg13g2_fill_1 FILLER_38_1092 ();
 sg13g2_fill_1 FILLER_38_1100 ();
 sg13g2_fill_1 FILLER_38_1105 ();
 sg13g2_fill_2 FILLER_38_1154 ();
 sg13g2_fill_1 FILLER_38_1195 ();
 sg13g2_fill_1 FILLER_38_1222 ();
 sg13g2_fill_1 FILLER_38_1226 ();
 sg13g2_fill_1 FILLER_38_1270 ();
 sg13g2_fill_1 FILLER_38_1275 ();
 sg13g2_fill_1 FILLER_38_1338 ();
 sg13g2_fill_1 FILLER_38_1343 ();
 sg13g2_fill_1 FILLER_38_1348 ();
 sg13g2_fill_1 FILLER_38_1375 ();
 sg13g2_fill_2 FILLER_38_1423 ();
 sg13g2_fill_1 FILLER_38_1437 ();
 sg13g2_fill_1 FILLER_38_1445 ();
 sg13g2_fill_2 FILLER_38_1470 ();
 sg13g2_fill_2 FILLER_38_1476 ();
 sg13g2_fill_2 FILLER_38_1490 ();
 sg13g2_fill_1 FILLER_38_1549 ();
 sg13g2_fill_1 FILLER_38_1568 ();
 sg13g2_decap_8 FILLER_38_1582 ();
 sg13g2_decap_8 FILLER_38_1589 ();
 sg13g2_decap_8 FILLER_38_1596 ();
 sg13g2_decap_8 FILLER_38_1672 ();
 sg13g2_fill_2 FILLER_38_1679 ();
 sg13g2_fill_1 FILLER_38_1686 ();
 sg13g2_decap_4 FILLER_38_1695 ();
 sg13g2_fill_1 FILLER_38_1699 ();
 sg13g2_fill_1 FILLER_38_1726 ();
 sg13g2_decap_4 FILLER_38_1753 ();
 sg13g2_fill_2 FILLER_38_1757 ();
 sg13g2_fill_1 FILLER_38_1799 ();
 sg13g2_fill_2 FILLER_38_1825 ();
 sg13g2_decap_8 FILLER_38_1831 ();
 sg13g2_decap_4 FILLER_38_1878 ();
 sg13g2_fill_1 FILLER_38_1891 ();
 sg13g2_fill_1 FILLER_38_1931 ();
 sg13g2_fill_2 FILLER_38_1941 ();
 sg13g2_fill_1 FILLER_38_1975 ();
 sg13g2_fill_1 FILLER_38_1980 ();
 sg13g2_fill_1 FILLER_38_2050 ();
 sg13g2_fill_2 FILLER_38_2056 ();
 sg13g2_decap_4 FILLER_38_2062 ();
 sg13g2_fill_1 FILLER_38_2071 ();
 sg13g2_fill_2 FILLER_38_2108 ();
 sg13g2_fill_1 FILLER_38_2136 ();
 sg13g2_fill_2 FILLER_38_2184 ();
 sg13g2_fill_1 FILLER_38_2221 ();
 sg13g2_fill_1 FILLER_38_2234 ();
 sg13g2_fill_2 FILLER_38_2287 ();
 sg13g2_fill_1 FILLER_38_2289 ();
 sg13g2_fill_2 FILLER_38_2342 ();
 sg13g2_decap_4 FILLER_38_2354 ();
 sg13g2_decap_4 FILLER_38_2362 ();
 sg13g2_fill_2 FILLER_38_2376 ();
 sg13g2_fill_1 FILLER_38_2378 ();
 sg13g2_decap_4 FILLER_38_2410 ();
 sg13g2_fill_1 FILLER_38_2427 ();
 sg13g2_decap_4 FILLER_38_2454 ();
 sg13g2_fill_1 FILLER_38_2458 ();
 sg13g2_fill_2 FILLER_38_2489 ();
 sg13g2_decap_8 FILLER_38_2501 ();
 sg13g2_decap_8 FILLER_38_2589 ();
 sg13g2_decap_4 FILLER_38_2596 ();
 sg13g2_fill_2 FILLER_38_2600 ();
 sg13g2_decap_8 FILLER_38_2606 ();
 sg13g2_decap_8 FILLER_38_2613 ();
 sg13g2_decap_8 FILLER_38_2620 ();
 sg13g2_decap_8 FILLER_38_2627 ();
 sg13g2_decap_8 FILLER_38_2634 ();
 sg13g2_decap_8 FILLER_38_2641 ();
 sg13g2_decap_8 FILLER_38_2648 ();
 sg13g2_decap_8 FILLER_38_2655 ();
 sg13g2_decap_8 FILLER_38_2662 ();
 sg13g2_fill_1 FILLER_38_2669 ();
 sg13g2_fill_2 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_56 ();
 sg13g2_fill_1 FILLER_39_58 ();
 sg13g2_fill_1 FILLER_39_68 ();
 sg13g2_decap_4 FILLER_39_80 ();
 sg13g2_fill_1 FILLER_39_98 ();
 sg13g2_fill_1 FILLER_39_150 ();
 sg13g2_fill_2 FILLER_39_161 ();
 sg13g2_fill_1 FILLER_39_211 ();
 sg13g2_fill_2 FILLER_39_219 ();
 sg13g2_fill_2 FILLER_39_226 ();
 sg13g2_decap_8 FILLER_39_234 ();
 sg13g2_decap_8 FILLER_39_241 ();
 sg13g2_decap_4 FILLER_39_248 ();
 sg13g2_fill_2 FILLER_39_252 ();
 sg13g2_fill_1 FILLER_39_258 ();
 sg13g2_decap_8 FILLER_39_263 ();
 sg13g2_fill_2 FILLER_39_276 ();
 sg13g2_fill_1 FILLER_39_295 ();
 sg13g2_decap_8 FILLER_39_300 ();
 sg13g2_decap_8 FILLER_39_307 ();
 sg13g2_decap_8 FILLER_39_314 ();
 sg13g2_decap_8 FILLER_39_321 ();
 sg13g2_fill_2 FILLER_39_409 ();
 sg13g2_fill_2 FILLER_39_425 ();
 sg13g2_fill_2 FILLER_39_445 ();
 sg13g2_decap_4 FILLER_39_532 ();
 sg13g2_fill_1 FILLER_39_536 ();
 sg13g2_decap_4 FILLER_39_543 ();
 sg13g2_fill_2 FILLER_39_547 ();
 sg13g2_fill_2 FILLER_39_552 ();
 sg13g2_fill_2 FILLER_39_562 ();
 sg13g2_fill_1 FILLER_39_564 ();
 sg13g2_decap_4 FILLER_39_596 ();
 sg13g2_fill_1 FILLER_39_605 ();
 sg13g2_fill_2 FILLER_39_637 ();
 sg13g2_fill_1 FILLER_39_639 ();
 sg13g2_decap_4 FILLER_39_679 ();
 sg13g2_fill_1 FILLER_39_683 ();
 sg13g2_fill_2 FILLER_39_703 ();
 sg13g2_decap_8 FILLER_39_709 ();
 sg13g2_fill_1 FILLER_39_716 ();
 sg13g2_fill_1 FILLER_39_721 ();
 sg13g2_fill_1 FILLER_39_769 ();
 sg13g2_fill_2 FILLER_39_774 ();
 sg13g2_fill_2 FILLER_39_781 ();
 sg13g2_fill_1 FILLER_39_783 ();
 sg13g2_fill_2 FILLER_39_794 ();
 sg13g2_decap_8 FILLER_39_835 ();
 sg13g2_fill_2 FILLER_39_873 ();
 sg13g2_fill_1 FILLER_39_875 ();
 sg13g2_fill_1 FILLER_39_895 ();
 sg13g2_fill_1 FILLER_39_906 ();
 sg13g2_decap_4 FILLER_39_944 ();
 sg13g2_decap_8 FILLER_39_952 ();
 sg13g2_fill_1 FILLER_39_959 ();
 sg13g2_decap_8 FILLER_39_965 ();
 sg13g2_decap_4 FILLER_39_972 ();
 sg13g2_fill_2 FILLER_39_976 ();
 sg13g2_decap_8 FILLER_39_982 ();
 sg13g2_decap_8 FILLER_39_989 ();
 sg13g2_decap_4 FILLER_39_996 ();
 sg13g2_decap_4 FILLER_39_1015 ();
 sg13g2_fill_2 FILLER_39_1019 ();
 sg13g2_decap_8 FILLER_39_1025 ();
 sg13g2_decap_8 FILLER_39_1032 ();
 sg13g2_fill_1 FILLER_39_1039 ();
 sg13g2_decap_4 FILLER_39_1051 ();
 sg13g2_fill_2 FILLER_39_1059 ();
 sg13g2_fill_1 FILLER_39_1061 ();
 sg13g2_decap_4 FILLER_39_1076 ();
 sg13g2_fill_2 FILLER_39_1080 ();
 sg13g2_decap_4 FILLER_39_1086 ();
 sg13g2_fill_1 FILLER_39_1090 ();
 sg13g2_fill_1 FILLER_39_1118 ();
 sg13g2_fill_1 FILLER_39_1135 ();
 sg13g2_fill_2 FILLER_39_1156 ();
 sg13g2_fill_1 FILLER_39_1161 ();
 sg13g2_fill_1 FILLER_39_1176 ();
 sg13g2_fill_2 FILLER_39_1218 ();
 sg13g2_decap_8 FILLER_39_1258 ();
 sg13g2_decap_8 FILLER_39_1265 ();
 sg13g2_decap_4 FILLER_39_1272 ();
 sg13g2_fill_1 FILLER_39_1276 ();
 sg13g2_decap_4 FILLER_39_1316 ();
 sg13g2_fill_1 FILLER_39_1320 ();
 sg13g2_decap_8 FILLER_39_1325 ();
 sg13g2_decap_8 FILLER_39_1332 ();
 sg13g2_decap_8 FILLER_39_1339 ();
 sg13g2_fill_2 FILLER_39_1346 ();
 sg13g2_fill_2 FILLER_39_1362 ();
 sg13g2_fill_1 FILLER_39_1364 ();
 sg13g2_decap_8 FILLER_39_1391 ();
 sg13g2_fill_1 FILLER_39_1398 ();
 sg13g2_decap_8 FILLER_39_1474 ();
 sg13g2_fill_1 FILLER_39_1496 ();
 sg13g2_fill_2 FILLER_39_1501 ();
 sg13g2_fill_2 FILLER_39_1532 ();
 sg13g2_fill_1 FILLER_39_1558 ();
 sg13g2_fill_1 FILLER_39_1564 ();
 sg13g2_decap_4 FILLER_39_1568 ();
 sg13g2_decap_8 FILLER_39_1577 ();
 sg13g2_decap_4 FILLER_39_1598 ();
 sg13g2_fill_2 FILLER_39_1602 ();
 sg13g2_fill_1 FILLER_39_1636 ();
 sg13g2_fill_2 FILLER_39_1660 ();
 sg13g2_fill_2 FILLER_39_1671 ();
 sg13g2_fill_1 FILLER_39_1673 ();
 sg13g2_fill_2 FILLER_39_1714 ();
 sg13g2_fill_2 FILLER_39_1742 ();
 sg13g2_fill_1 FILLER_39_1744 ();
 sg13g2_decap_8 FILLER_39_1749 ();
 sg13g2_decap_8 FILLER_39_1763 ();
 sg13g2_decap_8 FILLER_39_1770 ();
 sg13g2_decap_8 FILLER_39_1832 ();
 sg13g2_decap_4 FILLER_39_1839 ();
 sg13g2_fill_1 FILLER_39_1843 ();
 sg13g2_fill_1 FILLER_39_1852 ();
 sg13g2_decap_4 FILLER_39_1886 ();
 sg13g2_fill_2 FILLER_39_1909 ();
 sg13g2_fill_1 FILLER_39_1911 ();
 sg13g2_fill_2 FILLER_39_1920 ();
 sg13g2_fill_1 FILLER_39_1926 ();
 sg13g2_fill_1 FILLER_39_1943 ();
 sg13g2_fill_1 FILLER_39_1950 ();
 sg13g2_fill_1 FILLER_39_1956 ();
 sg13g2_fill_1 FILLER_39_1983 ();
 sg13g2_fill_2 FILLER_39_1989 ();
 sg13g2_fill_1 FILLER_39_1999 ();
 sg13g2_fill_1 FILLER_39_2004 ();
 sg13g2_fill_1 FILLER_39_2035 ();
 sg13g2_fill_1 FILLER_39_2041 ();
 sg13g2_fill_2 FILLER_39_2046 ();
 sg13g2_decap_8 FILLER_39_2053 ();
 sg13g2_decap_8 FILLER_39_2060 ();
 sg13g2_decap_8 FILLER_39_2067 ();
 sg13g2_fill_2 FILLER_39_2074 ();
 sg13g2_fill_1 FILLER_39_2076 ();
 sg13g2_fill_2 FILLER_39_2085 ();
 sg13g2_fill_2 FILLER_39_2117 ();
 sg13g2_fill_1 FILLER_39_2272 ();
 sg13g2_decap_4 FILLER_39_2318 ();
 sg13g2_fill_1 FILLER_39_2322 ();
 sg13g2_decap_8 FILLER_39_2327 ();
 sg13g2_decap_8 FILLER_39_2338 ();
 sg13g2_decap_4 FILLER_39_2345 ();
 sg13g2_fill_2 FILLER_39_2349 ();
 sg13g2_fill_1 FILLER_39_2377 ();
 sg13g2_fill_2 FILLER_39_2388 ();
 sg13g2_fill_2 FILLER_39_2421 ();
 sg13g2_fill_1 FILLER_39_2423 ();
 sg13g2_fill_2 FILLER_39_2445 ();
 sg13g2_fill_1 FILLER_39_2447 ();
 sg13g2_fill_2 FILLER_39_2465 ();
 sg13g2_fill_1 FILLER_39_2467 ();
 sg13g2_fill_2 FILLER_39_2494 ();
 sg13g2_fill_2 FILLER_39_2541 ();
 sg13g2_fill_2 FILLER_39_2546 ();
 sg13g2_fill_1 FILLER_39_2592 ();
 sg13g2_decap_8 FILLER_39_2597 ();
 sg13g2_decap_8 FILLER_39_2604 ();
 sg13g2_decap_8 FILLER_39_2611 ();
 sg13g2_decap_8 FILLER_39_2618 ();
 sg13g2_decap_8 FILLER_39_2625 ();
 sg13g2_decap_8 FILLER_39_2632 ();
 sg13g2_decap_8 FILLER_39_2639 ();
 sg13g2_decap_8 FILLER_39_2646 ();
 sg13g2_decap_8 FILLER_39_2653 ();
 sg13g2_decap_8 FILLER_39_2660 ();
 sg13g2_fill_2 FILLER_39_2667 ();
 sg13g2_fill_1 FILLER_39_2669 ();
 sg13g2_fill_1 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_6 ();
 sg13g2_fill_1 FILLER_40_12 ();
 sg13g2_fill_1 FILLER_40_17 ();
 sg13g2_fill_1 FILLER_40_23 ();
 sg13g2_fill_1 FILLER_40_29 ();
 sg13g2_fill_2 FILLER_40_34 ();
 sg13g2_fill_1 FILLER_40_46 ();
 sg13g2_fill_2 FILLER_40_56 ();
 sg13g2_fill_1 FILLER_40_58 ();
 sg13g2_fill_1 FILLER_40_82 ();
 sg13g2_decap_4 FILLER_40_88 ();
 sg13g2_fill_1 FILLER_40_105 ();
 sg13g2_fill_2 FILLER_40_110 ();
 sg13g2_fill_1 FILLER_40_112 ();
 sg13g2_fill_2 FILLER_40_117 ();
 sg13g2_fill_1 FILLER_40_119 ();
 sg13g2_fill_1 FILLER_40_156 ();
 sg13g2_fill_2 FILLER_40_171 ();
 sg13g2_fill_1 FILLER_40_173 ();
 sg13g2_decap_8 FILLER_40_190 ();
 sg13g2_decap_8 FILLER_40_197 ();
 sg13g2_fill_1 FILLER_40_204 ();
 sg13g2_fill_2 FILLER_40_249 ();
 sg13g2_decap_8 FILLER_40_288 ();
 sg13g2_fill_1 FILLER_40_295 ();
 sg13g2_fill_2 FILLER_40_328 ();
 sg13g2_fill_2 FILLER_40_334 ();
 sg13g2_fill_1 FILLER_40_372 ();
 sg13g2_fill_2 FILLER_40_396 ();
 sg13g2_fill_1 FILLER_40_406 ();
 sg13g2_fill_2 FILLER_40_422 ();
 sg13g2_fill_1 FILLER_40_433 ();
 sg13g2_fill_2 FILLER_40_441 ();
 sg13g2_fill_2 FILLER_40_477 ();
 sg13g2_decap_8 FILLER_40_483 ();
 sg13g2_fill_2 FILLER_40_495 ();
 sg13g2_fill_1 FILLER_40_506 ();
 sg13g2_decap_4 FILLER_40_533 ();
 sg13g2_fill_2 FILLER_40_537 ();
 sg13g2_fill_1 FILLER_40_543 ();
 sg13g2_fill_1 FILLER_40_548 ();
 sg13g2_fill_2 FILLER_40_553 ();
 sg13g2_fill_1 FILLER_40_555 ();
 sg13g2_fill_2 FILLER_40_573 ();
 sg13g2_decap_4 FILLER_40_592 ();
 sg13g2_fill_1 FILLER_40_596 ();
 sg13g2_fill_1 FILLER_40_602 ();
 sg13g2_fill_2 FILLER_40_660 ();
 sg13g2_fill_1 FILLER_40_662 ();
 sg13g2_fill_2 FILLER_40_668 ();
 sg13g2_fill_1 FILLER_40_670 ();
 sg13g2_fill_2 FILLER_40_676 ();
 sg13g2_fill_1 FILLER_40_678 ();
 sg13g2_fill_1 FILLER_40_693 ();
 sg13g2_fill_1 FILLER_40_724 ();
 sg13g2_fill_1 FILLER_40_730 ();
 sg13g2_fill_1 FILLER_40_746 ();
 sg13g2_fill_1 FILLER_40_751 ();
 sg13g2_decap_4 FILLER_40_757 ();
 sg13g2_decap_8 FILLER_40_771 ();
 sg13g2_decap_8 FILLER_40_778 ();
 sg13g2_decap_8 FILLER_40_785 ();
 sg13g2_fill_1 FILLER_40_802 ();
 sg13g2_decap_8 FILLER_40_814 ();
 sg13g2_fill_1 FILLER_40_821 ();
 sg13g2_decap_8 FILLER_40_826 ();
 sg13g2_fill_2 FILLER_40_843 ();
 sg13g2_fill_1 FILLER_40_855 ();
 sg13g2_fill_2 FILLER_40_866 ();
 sg13g2_decap_8 FILLER_40_949 ();
 sg13g2_decap_8 FILLER_40_956 ();
 sg13g2_fill_2 FILLER_40_963 ();
 sg13g2_fill_1 FILLER_40_965 ();
 sg13g2_decap_8 FILLER_40_970 ();
 sg13g2_fill_2 FILLER_40_977 ();
 sg13g2_decap_8 FILLER_40_993 ();
 sg13g2_fill_1 FILLER_40_1000 ();
 sg13g2_decap_8 FILLER_40_1040 ();
 sg13g2_fill_1 FILLER_40_1047 ();
 sg13g2_fill_1 FILLER_40_1051 ();
 sg13g2_decap_8 FILLER_40_1078 ();
 sg13g2_fill_2 FILLER_40_1085 ();
 sg13g2_fill_1 FILLER_40_1087 ();
 sg13g2_fill_2 FILLER_40_1166 ();
 sg13g2_fill_1 FILLER_40_1182 ();
 sg13g2_decap_8 FILLER_40_1187 ();
 sg13g2_fill_1 FILLER_40_1224 ();
 sg13g2_decap_4 FILLER_40_1230 ();
 sg13g2_fill_1 FILLER_40_1234 ();
 sg13g2_fill_2 FILLER_40_1239 ();
 sg13g2_fill_2 FILLER_40_1262 ();
 sg13g2_fill_1 FILLER_40_1264 ();
 sg13g2_decap_4 FILLER_40_1273 ();
 sg13g2_fill_1 FILLER_40_1277 ();
 sg13g2_fill_1 FILLER_40_1286 ();
 sg13g2_fill_2 FILLER_40_1291 ();
 sg13g2_decap_4 FILLER_40_1301 ();
 sg13g2_fill_2 FILLER_40_1314 ();
 sg13g2_fill_1 FILLER_40_1316 ();
 sg13g2_decap_8 FILLER_40_1329 ();
 sg13g2_decap_8 FILLER_40_1336 ();
 sg13g2_decap_8 FILLER_40_1343 ();
 sg13g2_fill_2 FILLER_40_1350 ();
 sg13g2_decap_8 FILLER_40_1362 ();
 sg13g2_decap_4 FILLER_40_1369 ();
 sg13g2_fill_1 FILLER_40_1373 ();
 sg13g2_decap_4 FILLER_40_1378 ();
 sg13g2_decap_8 FILLER_40_1386 ();
 sg13g2_decap_4 FILLER_40_1393 ();
 sg13g2_fill_2 FILLER_40_1407 ();
 sg13g2_decap_8 FILLER_40_1455 ();
 sg13g2_decap_8 FILLER_40_1462 ();
 sg13g2_decap_8 FILLER_40_1469 ();
 sg13g2_decap_4 FILLER_40_1476 ();
 sg13g2_fill_1 FILLER_40_1480 ();
 sg13g2_fill_2 FILLER_40_1489 ();
 sg13g2_fill_1 FILLER_40_1491 ();
 sg13g2_fill_2 FILLER_40_1504 ();
 sg13g2_fill_1 FILLER_40_1515 ();
 sg13g2_fill_1 FILLER_40_1520 ();
 sg13g2_decap_4 FILLER_40_1552 ();
 sg13g2_decap_8 FILLER_40_1569 ();
 sg13g2_decap_8 FILLER_40_1576 ();
 sg13g2_decap_4 FILLER_40_1583 ();
 sg13g2_fill_2 FILLER_40_1587 ();
 sg13g2_decap_4 FILLER_40_1599 ();
 sg13g2_fill_2 FILLER_40_1603 ();
 sg13g2_decap_8 FILLER_40_1611 ();
 sg13g2_decap_4 FILLER_40_1674 ();
 sg13g2_fill_2 FILLER_40_1678 ();
 sg13g2_decap_4 FILLER_40_1684 ();
 sg13g2_fill_2 FILLER_40_1691 ();
 sg13g2_fill_1 FILLER_40_1693 ();
 sg13g2_fill_2 FILLER_40_1704 ();
 sg13g2_fill_1 FILLER_40_1706 ();
 sg13g2_decap_4 FILLER_40_1712 ();
 sg13g2_fill_1 FILLER_40_1716 ();
 sg13g2_decap_4 FILLER_40_1727 ();
 sg13g2_fill_2 FILLER_40_1731 ();
 sg13g2_fill_2 FILLER_40_1784 ();
 sg13g2_fill_1 FILLER_40_1802 ();
 sg13g2_fill_2 FILLER_40_1820 ();
 sg13g2_fill_1 FILLER_40_1826 ();
 sg13g2_decap_8 FILLER_40_1843 ();
 sg13g2_fill_2 FILLER_40_1850 ();
 sg13g2_fill_1 FILLER_40_1852 ();
 sg13g2_decap_4 FILLER_40_1867 ();
 sg13g2_fill_1 FILLER_40_1892 ();
 sg13g2_decap_4 FILLER_40_1898 ();
 sg13g2_fill_1 FILLER_40_1916 ();
 sg13g2_fill_1 FILLER_40_1953 ();
 sg13g2_decap_4 FILLER_40_1959 ();
 sg13g2_fill_1 FILLER_40_1963 ();
 sg13g2_fill_1 FILLER_40_1968 ();
 sg13g2_decap_8 FILLER_40_1980 ();
 sg13g2_decap_4 FILLER_40_1987 ();
 sg13g2_fill_2 FILLER_40_1991 ();
 sg13g2_fill_1 FILLER_40_1997 ();
 sg13g2_fill_2 FILLER_40_2019 ();
 sg13g2_fill_1 FILLER_40_2021 ();
 sg13g2_fill_1 FILLER_40_2027 ();
 sg13g2_fill_1 FILLER_40_2039 ();
 sg13g2_decap_4 FILLER_40_2092 ();
 sg13g2_fill_1 FILLER_40_2110 ();
 sg13g2_fill_1 FILLER_40_2149 ();
 sg13g2_decap_8 FILLER_40_2192 ();
 sg13g2_fill_1 FILLER_40_2199 ();
 sg13g2_fill_2 FILLER_40_2204 ();
 sg13g2_fill_1 FILLER_40_2215 ();
 sg13g2_fill_2 FILLER_40_2230 ();
 sg13g2_fill_2 FILLER_40_2239 ();
 sg13g2_fill_1 FILLER_40_2268 ();
 sg13g2_fill_1 FILLER_40_2277 ();
 sg13g2_fill_1 FILLER_40_2296 ();
 sg13g2_decap_8 FILLER_40_2333 ();
 sg13g2_decap_8 FILLER_40_2340 ();
 sg13g2_decap_8 FILLER_40_2347 ();
 sg13g2_fill_2 FILLER_40_2354 ();
 sg13g2_fill_1 FILLER_40_2356 ();
 sg13g2_decap_4 FILLER_40_2387 ();
 sg13g2_fill_2 FILLER_40_2417 ();
 sg13g2_decap_4 FILLER_40_2429 ();
 sg13g2_fill_2 FILLER_40_2433 ();
 sg13g2_fill_1 FILLER_40_2479 ();
 sg13g2_decap_4 FILLER_40_2485 ();
 sg13g2_fill_1 FILLER_40_2489 ();
 sg13g2_fill_1 FILLER_40_2500 ();
 sg13g2_decap_8 FILLER_40_2505 ();
 sg13g2_fill_2 FILLER_40_2512 ();
 sg13g2_decap_8 FILLER_40_2576 ();
 sg13g2_decap_8 FILLER_40_2609 ();
 sg13g2_decap_8 FILLER_40_2616 ();
 sg13g2_decap_8 FILLER_40_2623 ();
 sg13g2_decap_8 FILLER_40_2630 ();
 sg13g2_decap_8 FILLER_40_2637 ();
 sg13g2_decap_8 FILLER_40_2644 ();
 sg13g2_decap_8 FILLER_40_2651 ();
 sg13g2_decap_8 FILLER_40_2658 ();
 sg13g2_decap_4 FILLER_40_2665 ();
 sg13g2_fill_1 FILLER_40_2669 ();
 sg13g2_fill_2 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_32 ();
 sg13g2_fill_1 FILLER_41_34 ();
 sg13g2_fill_1 FILLER_41_50 ();
 sg13g2_fill_1 FILLER_41_56 ();
 sg13g2_decap_4 FILLER_41_69 ();
 sg13g2_decap_8 FILLER_41_83 ();
 sg13g2_fill_2 FILLER_41_153 ();
 sg13g2_fill_1 FILLER_41_169 ();
 sg13g2_decap_8 FILLER_41_196 ();
 sg13g2_decap_8 FILLER_41_203 ();
 sg13g2_decap_4 FILLER_41_210 ();
 sg13g2_fill_2 FILLER_41_214 ();
 sg13g2_fill_1 FILLER_41_221 ();
 sg13g2_fill_1 FILLER_41_226 ();
 sg13g2_fill_2 FILLER_41_231 ();
 sg13g2_fill_2 FILLER_41_242 ();
 sg13g2_decap_4 FILLER_41_249 ();
 sg13g2_fill_1 FILLER_41_253 ();
 sg13g2_fill_2 FILLER_41_298 ();
 sg13g2_fill_1 FILLER_41_317 ();
 sg13g2_fill_2 FILLER_41_321 ();
 sg13g2_fill_1 FILLER_41_338 ();
 sg13g2_fill_2 FILLER_41_363 ();
 sg13g2_fill_2 FILLER_41_408 ();
 sg13g2_fill_1 FILLER_41_417 ();
 sg13g2_fill_2 FILLER_41_428 ();
 sg13g2_fill_1 FILLER_41_447 ();
 sg13g2_decap_8 FILLER_41_474 ();
 sg13g2_decap_8 FILLER_41_481 ();
 sg13g2_fill_2 FILLER_41_488 ();
 sg13g2_fill_1 FILLER_41_490 ();
 sg13g2_fill_1 FILLER_41_500 ();
 sg13g2_decap_8 FILLER_41_515 ();
 sg13g2_fill_1 FILLER_41_522 ();
 sg13g2_fill_2 FILLER_41_549 ();
 sg13g2_decap_8 FILLER_41_566 ();
 sg13g2_decap_8 FILLER_41_573 ();
 sg13g2_decap_4 FILLER_41_580 ();
 sg13g2_decap_8 FILLER_41_589 ();
 sg13g2_decap_8 FILLER_41_596 ();
 sg13g2_decap_8 FILLER_41_607 ();
 sg13g2_fill_1 FILLER_41_614 ();
 sg13g2_decap_8 FILLER_41_619 ();
 sg13g2_decap_4 FILLER_41_626 ();
 sg13g2_fill_2 FILLER_41_635 ();
 sg13g2_fill_1 FILLER_41_643 ();
 sg13g2_fill_2 FILLER_41_649 ();
 sg13g2_fill_2 FILLER_41_656 ();
 sg13g2_fill_2 FILLER_41_663 ();
 sg13g2_fill_1 FILLER_41_665 ();
 sg13g2_decap_4 FILLER_41_686 ();
 sg13g2_fill_1 FILLER_41_721 ();
 sg13g2_fill_1 FILLER_41_736 ();
 sg13g2_fill_2 FILLER_41_763 ();
 sg13g2_fill_2 FILLER_41_826 ();
 sg13g2_fill_1 FILLER_41_828 ();
 sg13g2_fill_2 FILLER_41_881 ();
 sg13g2_fill_2 FILLER_41_914 ();
 sg13g2_fill_1 FILLER_41_916 ();
 sg13g2_fill_2 FILLER_41_1019 ();
 sg13g2_fill_1 FILLER_41_1053 ();
 sg13g2_fill_2 FILLER_41_1069 ();
 sg13g2_fill_2 FILLER_41_1080 ();
 sg13g2_fill_2 FILLER_41_1092 ();
 sg13g2_fill_2 FILLER_41_1149 ();
 sg13g2_decap_8 FILLER_41_1194 ();
 sg13g2_decap_4 FILLER_41_1201 ();
 sg13g2_decap_4 FILLER_41_1211 ();
 sg13g2_fill_1 FILLER_41_1215 ();
 sg13g2_fill_2 FILLER_41_1220 ();
 sg13g2_fill_1 FILLER_41_1222 ();
 sg13g2_fill_1 FILLER_41_1243 ();
 sg13g2_decap_4 FILLER_41_1275 ();
 sg13g2_decap_8 FILLER_41_1283 ();
 sg13g2_decap_4 FILLER_41_1290 ();
 sg13g2_fill_2 FILLER_41_1309 ();
 sg13g2_decap_8 FILLER_41_1337 ();
 sg13g2_decap_8 FILLER_41_1344 ();
 sg13g2_decap_8 FILLER_41_1351 ();
 sg13g2_decap_4 FILLER_41_1358 ();
 sg13g2_fill_1 FILLER_41_1362 ();
 sg13g2_decap_8 FILLER_41_1366 ();
 sg13g2_fill_2 FILLER_41_1373 ();
 sg13g2_fill_2 FILLER_41_1401 ();
 sg13g2_fill_2 FILLER_41_1461 ();
 sg13g2_fill_2 FILLER_41_1476 ();
 sg13g2_fill_1 FILLER_41_1478 ();
 sg13g2_fill_1 FILLER_41_1505 ();
 sg13g2_fill_2 FILLER_41_1514 ();
 sg13g2_fill_1 FILLER_41_1516 ();
 sg13g2_fill_1 FILLER_41_1526 ();
 sg13g2_fill_2 FILLER_41_1534 ();
 sg13g2_fill_1 FILLER_41_1584 ();
 sg13g2_decap_8 FILLER_41_1589 ();
 sg13g2_fill_2 FILLER_41_1596 ();
 sg13g2_fill_1 FILLER_41_1598 ();
 sg13g2_decap_8 FILLER_41_1603 ();
 sg13g2_decap_8 FILLER_41_1610 ();
 sg13g2_fill_2 FILLER_41_1617 ();
 sg13g2_fill_1 FILLER_41_1622 ();
 sg13g2_fill_1 FILLER_41_1627 ();
 sg13g2_fill_1 FILLER_41_1633 ();
 sg13g2_fill_2 FILLER_41_1644 ();
 sg13g2_fill_1 FILLER_41_1674 ();
 sg13g2_decap_4 FILLER_41_1715 ();
 sg13g2_fill_1 FILLER_41_1719 ();
 sg13g2_fill_1 FILLER_41_1750 ();
 sg13g2_fill_1 FILLER_41_1786 ();
 sg13g2_fill_1 FILLER_41_1798 ();
 sg13g2_fill_1 FILLER_41_1804 ();
 sg13g2_fill_2 FILLER_41_1882 ();
 sg13g2_fill_1 FILLER_41_1884 ();
 sg13g2_fill_2 FILLER_41_1933 ();
 sg13g2_fill_1 FILLER_41_1977 ();
 sg13g2_fill_1 FILLER_41_1982 ();
 sg13g2_fill_1 FILLER_41_1987 ();
 sg13g2_fill_1 FILLER_41_1993 ();
 sg13g2_fill_1 FILLER_41_1998 ();
 sg13g2_fill_1 FILLER_41_2004 ();
 sg13g2_fill_1 FILLER_41_2010 ();
 sg13g2_fill_1 FILLER_41_2017 ();
 sg13g2_fill_1 FILLER_41_2030 ();
 sg13g2_fill_2 FILLER_41_2035 ();
 sg13g2_fill_1 FILLER_41_2037 ();
 sg13g2_decap_8 FILLER_41_2096 ();
 sg13g2_fill_2 FILLER_41_2103 ();
 sg13g2_fill_1 FILLER_41_2105 ();
 sg13g2_fill_1 FILLER_41_2126 ();
 sg13g2_fill_2 FILLER_41_2144 ();
 sg13g2_fill_1 FILLER_41_2156 ();
 sg13g2_fill_2 FILLER_41_2162 ();
 sg13g2_fill_1 FILLER_41_2182 ();
 sg13g2_decap_8 FILLER_41_2186 ();
 sg13g2_decap_8 FILLER_41_2193 ();
 sg13g2_decap_8 FILLER_41_2287 ();
 sg13g2_decap_8 FILLER_41_2294 ();
 sg13g2_decap_4 FILLER_41_2301 ();
 sg13g2_fill_1 FILLER_41_2305 ();
 sg13g2_decap_8 FILLER_41_2309 ();
 sg13g2_decap_8 FILLER_41_2316 ();
 sg13g2_decap_8 FILLER_41_2323 ();
 sg13g2_decap_8 FILLER_41_2330 ();
 sg13g2_decap_8 FILLER_41_2337 ();
 sg13g2_decap_8 FILLER_41_2344 ();
 sg13g2_decap_8 FILLER_41_2351 ();
 sg13g2_decap_4 FILLER_41_2358 ();
 sg13g2_fill_1 FILLER_41_2362 ();
 sg13g2_fill_2 FILLER_41_2371 ();
 sg13g2_fill_2 FILLER_41_2399 ();
 sg13g2_fill_1 FILLER_41_2401 ();
 sg13g2_fill_1 FILLER_41_2420 ();
 sg13g2_decap_8 FILLER_41_2431 ();
 sg13g2_fill_2 FILLER_41_2438 ();
 sg13g2_decap_8 FILLER_41_2444 ();
 sg13g2_decap_8 FILLER_41_2451 ();
 sg13g2_fill_2 FILLER_41_2458 ();
 sg13g2_fill_1 FILLER_41_2460 ();
 sg13g2_decap_8 FILLER_41_2487 ();
 sg13g2_decap_4 FILLER_41_2494 ();
 sg13g2_fill_1 FILLER_41_2498 ();
 sg13g2_fill_2 FILLER_41_2538 ();
 sg13g2_fill_2 FILLER_41_2567 ();
 sg13g2_decap_8 FILLER_41_2579 ();
 sg13g2_fill_2 FILLER_41_2586 ();
 sg13g2_decap_8 FILLER_41_2592 ();
 sg13g2_decap_8 FILLER_41_2599 ();
 sg13g2_decap_8 FILLER_41_2606 ();
 sg13g2_decap_8 FILLER_41_2613 ();
 sg13g2_decap_8 FILLER_41_2620 ();
 sg13g2_decap_8 FILLER_41_2627 ();
 sg13g2_decap_8 FILLER_41_2634 ();
 sg13g2_decap_8 FILLER_41_2641 ();
 sg13g2_decap_8 FILLER_41_2648 ();
 sg13g2_decap_8 FILLER_41_2655 ();
 sg13g2_decap_8 FILLER_41_2662 ();
 sg13g2_fill_1 FILLER_41_2669 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_13 ();
 sg13g2_fill_2 FILLER_42_32 ();
 sg13g2_fill_1 FILLER_42_34 ();
 sg13g2_fill_2 FILLER_42_39 ();
 sg13g2_fill_1 FILLER_42_41 ();
 sg13g2_fill_2 FILLER_42_73 ();
 sg13g2_decap_4 FILLER_42_88 ();
 sg13g2_fill_1 FILLER_42_92 ();
 sg13g2_decap_4 FILLER_42_192 ();
 sg13g2_decap_8 FILLER_42_213 ();
 sg13g2_decap_4 FILLER_42_220 ();
 sg13g2_fill_2 FILLER_42_224 ();
 sg13g2_fill_1 FILLER_42_273 ();
 sg13g2_fill_1 FILLER_42_279 ();
 sg13g2_fill_2 FILLER_42_285 ();
 sg13g2_fill_1 FILLER_42_291 ();
 sg13g2_fill_1 FILLER_42_298 ();
 sg13g2_fill_2 FILLER_42_314 ();
 sg13g2_fill_1 FILLER_42_344 ();
 sg13g2_fill_2 FILLER_42_363 ();
 sg13g2_fill_1 FILLER_42_407 ();
 sg13g2_fill_1 FILLER_42_416 ();
 sg13g2_fill_2 FILLER_42_453 ();
 sg13g2_fill_1 FILLER_42_459 ();
 sg13g2_decap_8 FILLER_42_469 ();
 sg13g2_decap_8 FILLER_42_476 ();
 sg13g2_fill_2 FILLER_42_483 ();
 sg13g2_decap_8 FILLER_42_506 ();
 sg13g2_fill_1 FILLER_42_513 ();
 sg13g2_fill_2 FILLER_42_556 ();
 sg13g2_fill_1 FILLER_42_572 ();
 sg13g2_fill_1 FILLER_42_582 ();
 sg13g2_fill_1 FILLER_42_587 ();
 sg13g2_fill_1 FILLER_42_608 ();
 sg13g2_decap_8 FILLER_42_614 ();
 sg13g2_fill_1 FILLER_42_657 ();
 sg13g2_fill_2 FILLER_42_663 ();
 sg13g2_decap_4 FILLER_42_670 ();
 sg13g2_fill_2 FILLER_42_674 ();
 sg13g2_fill_1 FILLER_42_727 ();
 sg13g2_fill_1 FILLER_42_765 ();
 sg13g2_decap_4 FILLER_42_788 ();
 sg13g2_decap_8 FILLER_42_802 ();
 sg13g2_decap_8 FILLER_42_809 ();
 sg13g2_decap_8 FILLER_42_816 ();
 sg13g2_decap_8 FILLER_42_823 ();
 sg13g2_fill_2 FILLER_42_830 ();
 sg13g2_fill_1 FILLER_42_832 ();
 sg13g2_fill_2 FILLER_42_837 ();
 sg13g2_decap_8 FILLER_42_850 ();
 sg13g2_decap_4 FILLER_42_857 ();
 sg13g2_fill_1 FILLER_42_861 ();
 sg13g2_fill_2 FILLER_42_891 ();
 sg13g2_decap_4 FILLER_42_903 ();
 sg13g2_fill_1 FILLER_42_907 ();
 sg13g2_fill_1 FILLER_42_928 ();
 sg13g2_decap_8 FILLER_42_933 ();
 sg13g2_decap_4 FILLER_42_950 ();
 sg13g2_fill_2 FILLER_42_954 ();
 sg13g2_fill_1 FILLER_42_960 ();
 sg13g2_fill_1 FILLER_42_975 ();
 sg13g2_fill_1 FILLER_42_1038 ();
 sg13g2_fill_1 FILLER_42_1060 ();
 sg13g2_fill_1 FILLER_42_1066 ();
 sg13g2_fill_1 FILLER_42_1088 ();
 sg13g2_fill_2 FILLER_42_1114 ();
 sg13g2_fill_2 FILLER_42_1155 ();
 sg13g2_fill_1 FILLER_42_1181 ();
 sg13g2_fill_1 FILLER_42_1187 ();
 sg13g2_decap_4 FILLER_42_1193 ();
 sg13g2_fill_1 FILLER_42_1204 ();
 sg13g2_fill_2 FILLER_42_1211 ();
 sg13g2_fill_1 FILLER_42_1213 ();
 sg13g2_fill_2 FILLER_42_1227 ();
 sg13g2_fill_1 FILLER_42_1283 ();
 sg13g2_fill_1 FILLER_42_1306 ();
 sg13g2_fill_1 FILLER_42_1320 ();
 sg13g2_fill_2 FILLER_42_1325 ();
 sg13g2_fill_1 FILLER_42_1327 ();
 sg13g2_fill_2 FILLER_42_1354 ();
 sg13g2_fill_1 FILLER_42_1356 ();
 sg13g2_fill_2 FILLER_42_1361 ();
 sg13g2_decap_8 FILLER_42_1392 ();
 sg13g2_fill_1 FILLER_42_1399 ();
 sg13g2_decap_4 FILLER_42_1409 ();
 sg13g2_fill_1 FILLER_42_1413 ();
 sg13g2_fill_1 FILLER_42_1443 ();
 sg13g2_fill_2 FILLER_42_1464 ();
 sg13g2_decap_4 FILLER_42_1475 ();
 sg13g2_fill_2 FILLER_42_1479 ();
 sg13g2_fill_2 FILLER_42_1489 ();
 sg13g2_fill_1 FILLER_42_1496 ();
 sg13g2_fill_1 FILLER_42_1502 ();
 sg13g2_fill_2 FILLER_42_1516 ();
 sg13g2_fill_1 FILLER_42_1518 ();
 sg13g2_decap_4 FILLER_42_1536 ();
 sg13g2_decap_4 FILLER_42_1545 ();
 sg13g2_fill_2 FILLER_42_1575 ();
 sg13g2_fill_2 FILLER_42_1580 ();
 sg13g2_decap_8 FILLER_42_1594 ();
 sg13g2_decap_8 FILLER_42_1601 ();
 sg13g2_decap_8 FILLER_42_1608 ();
 sg13g2_decap_4 FILLER_42_1615 ();
 sg13g2_decap_8 FILLER_42_1625 ();
 sg13g2_decap_4 FILLER_42_1632 ();
 sg13g2_fill_2 FILLER_42_1636 ();
 sg13g2_fill_2 FILLER_42_1665 ();
 sg13g2_fill_1 FILLER_42_1667 ();
 sg13g2_decap_8 FILLER_42_1686 ();
 sg13g2_decap_8 FILLER_42_1693 ();
 sg13g2_fill_2 FILLER_42_1700 ();
 sg13g2_fill_1 FILLER_42_1702 ();
 sg13g2_decap_4 FILLER_42_1739 ();
 sg13g2_fill_2 FILLER_42_1747 ();
 sg13g2_fill_1 FILLER_42_1749 ();
 sg13g2_decap_8 FILLER_42_1754 ();
 sg13g2_fill_2 FILLER_42_1761 ();
 sg13g2_fill_2 FILLER_42_1767 ();
 sg13g2_fill_1 FILLER_42_1769 ();
 sg13g2_fill_1 FILLER_42_1792 ();
 sg13g2_fill_1 FILLER_42_1802 ();
 sg13g2_fill_1 FILLER_42_1808 ();
 sg13g2_fill_2 FILLER_42_1828 ();
 sg13g2_fill_1 FILLER_42_1856 ();
 sg13g2_fill_1 FILLER_42_1862 ();
 sg13g2_fill_2 FILLER_42_1871 ();
 sg13g2_fill_1 FILLER_42_1873 ();
 sg13g2_fill_1 FILLER_42_1904 ();
 sg13g2_fill_2 FILLER_42_1952 ();
 sg13g2_fill_1 FILLER_42_1959 ();
 sg13g2_fill_1 FILLER_42_1969 ();
 sg13g2_decap_4 FILLER_42_1996 ();
 sg13g2_decap_4 FILLER_42_2005 ();
 sg13g2_fill_1 FILLER_42_2009 ();
 sg13g2_decap_4 FILLER_42_2070 ();
 sg13g2_fill_2 FILLER_42_2078 ();
 sg13g2_fill_1 FILLER_42_2080 ();
 sg13g2_decap_8 FILLER_42_2085 ();
 sg13g2_decap_8 FILLER_42_2092 ();
 sg13g2_fill_2 FILLER_42_2099 ();
 sg13g2_fill_1 FILLER_42_2186 ();
 sg13g2_decap_4 FILLER_42_2222 ();
 sg13g2_fill_2 FILLER_42_2226 ();
 sg13g2_fill_2 FILLER_42_2238 ();
 sg13g2_fill_1 FILLER_42_2261 ();
 sg13g2_decap_4 FILLER_42_2354 ();
 sg13g2_fill_2 FILLER_42_2358 ();
 sg13g2_decap_8 FILLER_42_2377 ();
 sg13g2_decap_8 FILLER_42_2384 ();
 sg13g2_fill_1 FILLER_42_2391 ();
 sg13g2_fill_1 FILLER_42_2396 ();
 sg13g2_fill_2 FILLER_42_2427 ();
 sg13g2_fill_1 FILLER_42_2429 ();
 sg13g2_decap_8 FILLER_42_2492 ();
 sg13g2_decap_8 FILLER_42_2499 ();
 sg13g2_decap_8 FILLER_42_2506 ();
 sg13g2_decap_4 FILLER_42_2513 ();
 sg13g2_fill_2 FILLER_42_2517 ();
 sg13g2_decap_8 FILLER_42_2527 ();
 sg13g2_decap_8 FILLER_42_2534 ();
 sg13g2_decap_8 FILLER_42_2541 ();
 sg13g2_decap_8 FILLER_42_2548 ();
 sg13g2_decap_4 FILLER_42_2555 ();
 sg13g2_decap_8 FILLER_42_2563 ();
 sg13g2_decap_8 FILLER_42_2570 ();
 sg13g2_decap_8 FILLER_42_2577 ();
 sg13g2_decap_8 FILLER_42_2584 ();
 sg13g2_decap_8 FILLER_42_2591 ();
 sg13g2_decap_8 FILLER_42_2598 ();
 sg13g2_decap_8 FILLER_42_2605 ();
 sg13g2_decap_8 FILLER_42_2612 ();
 sg13g2_decap_8 FILLER_42_2619 ();
 sg13g2_decap_8 FILLER_42_2626 ();
 sg13g2_decap_8 FILLER_42_2633 ();
 sg13g2_decap_8 FILLER_42_2640 ();
 sg13g2_decap_8 FILLER_42_2647 ();
 sg13g2_decap_8 FILLER_42_2654 ();
 sg13g2_decap_8 FILLER_42_2661 ();
 sg13g2_fill_2 FILLER_42_2668 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_4 FILLER_43_11 ();
 sg13g2_decap_8 FILLER_43_41 ();
 sg13g2_fill_1 FILLER_43_48 ();
 sg13g2_fill_1 FILLER_43_128 ();
 sg13g2_fill_2 FILLER_43_147 ();
 sg13g2_decap_8 FILLER_43_153 ();
 sg13g2_fill_1 FILLER_43_160 ();
 sg13g2_fill_1 FILLER_43_201 ();
 sg13g2_fill_1 FILLER_43_219 ();
 sg13g2_decap_4 FILLER_43_224 ();
 sg13g2_decap_8 FILLER_43_252 ();
 sg13g2_fill_1 FILLER_43_259 ();
 sg13g2_fill_1 FILLER_43_276 ();
 sg13g2_fill_1 FILLER_43_337 ();
 sg13g2_fill_1 FILLER_43_358 ();
 sg13g2_fill_2 FILLER_43_378 ();
 sg13g2_fill_1 FILLER_43_394 ();
 sg13g2_fill_2 FILLER_43_418 ();
 sg13g2_decap_4 FILLER_43_459 ();
 sg13g2_fill_2 FILLER_43_463 ();
 sg13g2_fill_1 FILLER_43_474 ();
 sg13g2_fill_1 FILLER_43_485 ();
 sg13g2_fill_2 FILLER_43_507 ();
 sg13g2_fill_2 FILLER_43_520 ();
 sg13g2_fill_1 FILLER_43_522 ();
 sg13g2_fill_1 FILLER_43_574 ();
 sg13g2_fill_2 FILLER_43_581 ();
 sg13g2_fill_1 FILLER_43_594 ();
 sg13g2_fill_2 FILLER_43_605 ();
 sg13g2_decap_8 FILLER_43_616 ();
 sg13g2_decap_4 FILLER_43_623 ();
 sg13g2_fill_1 FILLER_43_627 ();
 sg13g2_fill_1 FILLER_43_684 ();
 sg13g2_fill_1 FILLER_43_713 ();
 sg13g2_fill_1 FILLER_43_720 ();
 sg13g2_fill_1 FILLER_43_735 ();
 sg13g2_fill_1 FILLER_43_741 ();
 sg13g2_fill_1 FILLER_43_746 ();
 sg13g2_fill_1 FILLER_43_757 ();
 sg13g2_fill_2 FILLER_43_764 ();
 sg13g2_fill_2 FILLER_43_771 ();
 sg13g2_decap_8 FILLER_43_795 ();
 sg13g2_decap_8 FILLER_43_802 ();
 sg13g2_fill_2 FILLER_43_809 ();
 sg13g2_fill_1 FILLER_43_811 ();
 sg13g2_decap_4 FILLER_43_822 ();
 sg13g2_fill_1 FILLER_43_852 ();
 sg13g2_fill_1 FILLER_43_867 ();
 sg13g2_decap_4 FILLER_43_885 ();
 sg13g2_fill_1 FILLER_43_893 ();
 sg13g2_decap_8 FILLER_43_921 ();
 sg13g2_fill_1 FILLER_43_928 ();
 sg13g2_decap_8 FILLER_43_934 ();
 sg13g2_fill_1 FILLER_43_941 ();
 sg13g2_decap_8 FILLER_43_950 ();
 sg13g2_fill_2 FILLER_43_957 ();
 sg13g2_fill_1 FILLER_43_959 ();
 sg13g2_fill_2 FILLER_43_969 ();
 sg13g2_fill_2 FILLER_43_1041 ();
 sg13g2_fill_1 FILLER_43_1054 ();
 sg13g2_fill_1 FILLER_43_1078 ();
 sg13g2_fill_1 FILLER_43_1092 ();
 sg13g2_fill_1 FILLER_43_1126 ();
 sg13g2_fill_2 FILLER_43_1139 ();
 sg13g2_fill_2 FILLER_43_1145 ();
 sg13g2_decap_8 FILLER_43_1180 ();
 sg13g2_fill_2 FILLER_43_1202 ();
 sg13g2_fill_1 FILLER_43_1204 ();
 sg13g2_decap_4 FILLER_43_1221 ();
 sg13g2_fill_2 FILLER_43_1225 ();
 sg13g2_fill_2 FILLER_43_1231 ();
 sg13g2_decap_4 FILLER_43_1254 ();
 sg13g2_fill_1 FILLER_43_1292 ();
 sg13g2_fill_1 FILLER_43_1299 ();
 sg13g2_decap_4 FILLER_43_1303 ();
 sg13g2_fill_1 FILLER_43_1307 ();
 sg13g2_fill_2 FILLER_43_1312 ();
 sg13g2_fill_1 FILLER_43_1326 ();
 sg13g2_fill_2 FILLER_43_1344 ();
 sg13g2_fill_1 FILLER_43_1355 ();
 sg13g2_fill_2 FILLER_43_1370 ();
 sg13g2_fill_1 FILLER_43_1387 ();
 sg13g2_fill_2 FILLER_43_1422 ();
 sg13g2_fill_1 FILLER_43_1458 ();
 sg13g2_decap_4 FILLER_43_1467 ();
 sg13g2_fill_1 FILLER_43_1471 ();
 sg13g2_decap_4 FILLER_43_1507 ();
 sg13g2_fill_2 FILLER_43_1560 ();
 sg13g2_fill_1 FILLER_43_1562 ();
 sg13g2_fill_1 FILLER_43_1567 ();
 sg13g2_fill_2 FILLER_43_1572 ();
 sg13g2_decap_8 FILLER_43_1592 ();
 sg13g2_decap_8 FILLER_43_1607 ();
 sg13g2_decap_8 FILLER_43_1614 ();
 sg13g2_decap_8 FILLER_43_1621 ();
 sg13g2_decap_8 FILLER_43_1628 ();
 sg13g2_decap_4 FILLER_43_1635 ();
 sg13g2_fill_2 FILLER_43_1639 ();
 sg13g2_fill_2 FILLER_43_1647 ();
 sg13g2_fill_2 FILLER_43_1658 ();
 sg13g2_fill_2 FILLER_43_1668 ();
 sg13g2_fill_1 FILLER_43_1670 ();
 sg13g2_decap_8 FILLER_43_1689 ();
 sg13g2_decap_8 FILLER_43_1696 ();
 sg13g2_decap_8 FILLER_43_1703 ();
 sg13g2_decap_8 FILLER_43_1710 ();
 sg13g2_fill_2 FILLER_43_1717 ();
 sg13g2_fill_1 FILLER_43_1719 ();
 sg13g2_decap_8 FILLER_43_1724 ();
 sg13g2_decap_8 FILLER_43_1731 ();
 sg13g2_decap_8 FILLER_43_1738 ();
 sg13g2_decap_8 FILLER_43_1745 ();
 sg13g2_fill_2 FILLER_43_1752 ();
 sg13g2_fill_2 FILLER_43_1767 ();
 sg13g2_fill_1 FILLER_43_1769 ();
 sg13g2_fill_2 FILLER_43_1782 ();
 sg13g2_fill_1 FILLER_43_1810 ();
 sg13g2_fill_1 FILLER_43_1816 ();
 sg13g2_fill_1 FILLER_43_1926 ();
 sg13g2_fill_2 FILLER_43_1940 ();
 sg13g2_fill_2 FILLER_43_1953 ();
 sg13g2_fill_2 FILLER_43_1968 ();
 sg13g2_decap_8 FILLER_43_2013 ();
 sg13g2_decap_4 FILLER_43_2024 ();
 sg13g2_fill_2 FILLER_43_2028 ();
 sg13g2_decap_4 FILLER_43_2039 ();
 sg13g2_fill_1 FILLER_43_2048 ();
 sg13g2_fill_2 FILLER_43_2057 ();
 sg13g2_fill_1 FILLER_43_2059 ();
 sg13g2_decap_8 FILLER_43_2064 ();
 sg13g2_decap_8 FILLER_43_2071 ();
 sg13g2_decap_8 FILLER_43_2078 ();
 sg13g2_decap_8 FILLER_43_2085 ();
 sg13g2_fill_2 FILLER_43_2092 ();
 sg13g2_fill_2 FILLER_43_2175 ();
 sg13g2_fill_1 FILLER_43_2296 ();
 sg13g2_fill_1 FILLER_43_2309 ();
 sg13g2_fill_1 FILLER_43_2336 ();
 sg13g2_decap_8 FILLER_43_2363 ();
 sg13g2_decap_4 FILLER_43_2370 ();
 sg13g2_fill_1 FILLER_43_2374 ();
 sg13g2_decap_8 FILLER_43_2378 ();
 sg13g2_fill_2 FILLER_43_2415 ();
 sg13g2_fill_1 FILLER_43_2417 ();
 sg13g2_fill_2 FILLER_43_2448 ();
 sg13g2_fill_2 FILLER_43_2489 ();
 sg13g2_decap_8 FILLER_43_2504 ();
 sg13g2_decap_8 FILLER_43_2511 ();
 sg13g2_decap_8 FILLER_43_2518 ();
 sg13g2_decap_8 FILLER_43_2525 ();
 sg13g2_decap_8 FILLER_43_2532 ();
 sg13g2_decap_8 FILLER_43_2539 ();
 sg13g2_decap_8 FILLER_43_2546 ();
 sg13g2_decap_8 FILLER_43_2553 ();
 sg13g2_decap_8 FILLER_43_2560 ();
 sg13g2_decap_8 FILLER_43_2567 ();
 sg13g2_decap_8 FILLER_43_2574 ();
 sg13g2_decap_8 FILLER_43_2581 ();
 sg13g2_decap_8 FILLER_43_2588 ();
 sg13g2_decap_8 FILLER_43_2595 ();
 sg13g2_decap_8 FILLER_43_2602 ();
 sg13g2_decap_8 FILLER_43_2609 ();
 sg13g2_decap_8 FILLER_43_2616 ();
 sg13g2_decap_8 FILLER_43_2623 ();
 sg13g2_decap_8 FILLER_43_2630 ();
 sg13g2_decap_8 FILLER_43_2637 ();
 sg13g2_decap_8 FILLER_43_2644 ();
 sg13g2_decap_8 FILLER_43_2651 ();
 sg13g2_decap_8 FILLER_43_2658 ();
 sg13g2_decap_4 FILLER_43_2665 ();
 sg13g2_fill_1 FILLER_43_2669 ();
 sg13g2_fill_1 FILLER_44_0 ();
 sg13g2_decap_4 FILLER_44_32 ();
 sg13g2_decap_8 FILLER_44_41 ();
 sg13g2_decap_8 FILLER_44_48 ();
 sg13g2_fill_2 FILLER_44_55 ();
 sg13g2_fill_1 FILLER_44_57 ();
 sg13g2_fill_1 FILLER_44_70 ();
 sg13g2_decap_4 FILLER_44_75 ();
 sg13g2_fill_1 FILLER_44_79 ();
 sg13g2_decap_4 FILLER_44_90 ();
 sg13g2_fill_2 FILLER_44_94 ();
 sg13g2_fill_2 FILLER_44_126 ();
 sg13g2_fill_2 FILLER_44_132 ();
 sg13g2_decap_8 FILLER_44_139 ();
 sg13g2_decap_8 FILLER_44_146 ();
 sg13g2_fill_2 FILLER_44_153 ();
 sg13g2_decap_8 FILLER_44_159 ();
 sg13g2_decap_4 FILLER_44_166 ();
 sg13g2_fill_2 FILLER_44_170 ();
 sg13g2_fill_1 FILLER_44_212 ();
 sg13g2_fill_1 FILLER_44_218 ();
 sg13g2_decap_8 FILLER_44_223 ();
 sg13g2_decap_4 FILLER_44_239 ();
 sg13g2_decap_8 FILLER_44_251 ();
 sg13g2_fill_2 FILLER_44_258 ();
 sg13g2_fill_2 FILLER_44_276 ();
 sg13g2_fill_2 FILLER_44_283 ();
 sg13g2_fill_2 FILLER_44_332 ();
 sg13g2_fill_1 FILLER_44_344 ();
 sg13g2_fill_1 FILLER_44_371 ();
 sg13g2_fill_1 FILLER_44_377 ();
 sg13g2_fill_2 FILLER_44_412 ();
 sg13g2_decap_8 FILLER_44_499 ();
 sg13g2_decap_8 FILLER_44_506 ();
 sg13g2_decap_8 FILLER_44_513 ();
 sg13g2_decap_8 FILLER_44_520 ();
 sg13g2_decap_8 FILLER_44_527 ();
 sg13g2_fill_2 FILLER_44_534 ();
 sg13g2_fill_1 FILLER_44_536 ();
 sg13g2_fill_2 FILLER_44_565 ();
 sg13g2_fill_2 FILLER_44_602 ();
 sg13g2_decap_8 FILLER_44_616 ();
 sg13g2_decap_8 FILLER_44_623 ();
 sg13g2_decap_8 FILLER_44_630 ();
 sg13g2_fill_2 FILLER_44_658 ();
 sg13g2_decap_8 FILLER_44_668 ();
 sg13g2_fill_2 FILLER_44_675 ();
 sg13g2_decap_8 FILLER_44_695 ();
 sg13g2_fill_2 FILLER_44_702 ();
 sg13g2_fill_1 FILLER_44_704 ();
 sg13g2_decap_4 FILLER_44_709 ();
 sg13g2_fill_1 FILLER_44_713 ();
 sg13g2_decap_4 FILLER_44_720 ();
 sg13g2_fill_1 FILLER_44_734 ();
 sg13g2_fill_2 FILLER_44_761 ();
 sg13g2_fill_2 FILLER_44_773 ();
 sg13g2_fill_2 FILLER_44_801 ();
 sg13g2_fill_2 FILLER_44_813 ();
 sg13g2_fill_1 FILLER_44_815 ();
 sg13g2_fill_1 FILLER_44_842 ();
 sg13g2_fill_2 FILLER_44_853 ();
 sg13g2_fill_1 FILLER_44_855 ();
 sg13g2_decap_8 FILLER_44_887 ();
 sg13g2_decap_4 FILLER_44_894 ();
 sg13g2_fill_1 FILLER_44_898 ();
 sg13g2_decap_8 FILLER_44_904 ();
 sg13g2_decap_8 FILLER_44_911 ();
 sg13g2_fill_1 FILLER_44_918 ();
 sg13g2_decap_8 FILLER_44_945 ();
 sg13g2_decap_4 FILLER_44_952 ();
 sg13g2_fill_1 FILLER_44_956 ();
 sg13g2_fill_1 FILLER_44_987 ();
 sg13g2_fill_1 FILLER_44_995 ();
 sg13g2_fill_2 FILLER_44_1070 ();
 sg13g2_fill_1 FILLER_44_1104 ();
 sg13g2_fill_2 FILLER_44_1162 ();
 sg13g2_fill_1 FILLER_44_1183 ();
 sg13g2_fill_2 FILLER_44_1206 ();
 sg13g2_fill_1 FILLER_44_1208 ();
 sg13g2_decap_8 FILLER_44_1223 ();
 sg13g2_fill_2 FILLER_44_1230 ();
 sg13g2_decap_8 FILLER_44_1241 ();
 sg13g2_decap_4 FILLER_44_1268 ();
 sg13g2_fill_1 FILLER_44_1310 ();
 sg13g2_fill_2 FILLER_44_1340 ();
 sg13g2_fill_1 FILLER_44_1342 ();
 sg13g2_decap_8 FILLER_44_1353 ();
 sg13g2_decap_4 FILLER_44_1360 ();
 sg13g2_fill_2 FILLER_44_1372 ();
 sg13g2_decap_4 FILLER_44_1378 ();
 sg13g2_fill_1 FILLER_44_1382 ();
 sg13g2_fill_2 FILLER_44_1419 ();
 sg13g2_fill_1 FILLER_44_1433 ();
 sg13g2_decap_8 FILLER_44_1455 ();
 sg13g2_decap_8 FILLER_44_1462 ();
 sg13g2_decap_4 FILLER_44_1469 ();
 sg13g2_fill_2 FILLER_44_1473 ();
 sg13g2_decap_4 FILLER_44_1505 ();
 sg13g2_fill_1 FILLER_44_1509 ();
 sg13g2_fill_2 FILLER_44_1527 ();
 sg13g2_fill_1 FILLER_44_1551 ();
 sg13g2_decap_4 FILLER_44_1579 ();
 sg13g2_fill_1 FILLER_44_1583 ();
 sg13g2_decap_8 FILLER_44_1588 ();
 sg13g2_decap_8 FILLER_44_1630 ();
 sg13g2_decap_4 FILLER_44_1637 ();
 sg13g2_decap_8 FILLER_44_1674 ();
 sg13g2_decap_8 FILLER_44_1681 ();
 sg13g2_decap_8 FILLER_44_1688 ();
 sg13g2_decap_8 FILLER_44_1695 ();
 sg13g2_fill_2 FILLER_44_1702 ();
 sg13g2_fill_1 FILLER_44_1704 ();
 sg13g2_decap_8 FILLER_44_1718 ();
 sg13g2_fill_2 FILLER_44_1725 ();
 sg13g2_fill_1 FILLER_44_1727 ();
 sg13g2_fill_1 FILLER_44_1732 ();
 sg13g2_fill_2 FILLER_44_1737 ();
 sg13g2_decap_8 FILLER_44_1743 ();
 sg13g2_fill_1 FILLER_44_1759 ();
 sg13g2_fill_1 FILLER_44_1777 ();
 sg13g2_fill_2 FILLER_44_1793 ();
 sg13g2_fill_2 FILLER_44_1800 ();
 sg13g2_fill_2 FILLER_44_1807 ();
 sg13g2_fill_1 FILLER_44_1809 ();
 sg13g2_fill_1 FILLER_44_1815 ();
 sg13g2_fill_1 FILLER_44_1831 ();
 sg13g2_fill_1 FILLER_44_1837 ();
 sg13g2_fill_2 FILLER_44_1842 ();
 sg13g2_fill_2 FILLER_44_1888 ();
 sg13g2_fill_1 FILLER_44_1890 ();
 sg13g2_fill_1 FILLER_44_1937 ();
 sg13g2_fill_2 FILLER_44_1943 ();
 sg13g2_fill_1 FILLER_44_1963 ();
 sg13g2_fill_1 FILLER_44_1969 ();
 sg13g2_fill_1 FILLER_44_1976 ();
 sg13g2_fill_1 FILLER_44_1981 ();
 sg13g2_fill_2 FILLER_44_1988 ();
 sg13g2_fill_2 FILLER_44_2011 ();
 sg13g2_fill_1 FILLER_44_2013 ();
 sg13g2_fill_1 FILLER_44_2027 ();
 sg13g2_fill_1 FILLER_44_2041 ();
 sg13g2_decap_8 FILLER_44_2055 ();
 sg13g2_fill_2 FILLER_44_2062 ();
 sg13g2_fill_1 FILLER_44_2064 ();
 sg13g2_fill_1 FILLER_44_2112 ();
 sg13g2_fill_2 FILLER_44_2132 ();
 sg13g2_fill_2 FILLER_44_2164 ();
 sg13g2_fill_1 FILLER_44_2173 ();
 sg13g2_fill_1 FILLER_44_2200 ();
 sg13g2_decap_4 FILLER_44_2230 ();
 sg13g2_fill_2 FILLER_44_2242 ();
 sg13g2_decap_4 FILLER_44_2336 ();
 sg13g2_fill_1 FILLER_44_2340 ();
 sg13g2_fill_1 FILLER_44_2346 ();
 sg13g2_fill_2 FILLER_44_2373 ();
 sg13g2_decap_8 FILLER_44_2404 ();
 sg13g2_decap_4 FILLER_44_2411 ();
 sg13g2_fill_2 FILLER_44_2415 ();
 sg13g2_fill_1 FILLER_44_2423 ();
 sg13g2_decap_8 FILLER_44_2514 ();
 sg13g2_decap_8 FILLER_44_2521 ();
 sg13g2_decap_8 FILLER_44_2528 ();
 sg13g2_decap_8 FILLER_44_2535 ();
 sg13g2_decap_8 FILLER_44_2542 ();
 sg13g2_decap_8 FILLER_44_2549 ();
 sg13g2_decap_8 FILLER_44_2556 ();
 sg13g2_decap_8 FILLER_44_2563 ();
 sg13g2_decap_8 FILLER_44_2570 ();
 sg13g2_decap_8 FILLER_44_2577 ();
 sg13g2_decap_8 FILLER_44_2584 ();
 sg13g2_decap_8 FILLER_44_2591 ();
 sg13g2_decap_8 FILLER_44_2598 ();
 sg13g2_decap_8 FILLER_44_2605 ();
 sg13g2_decap_8 FILLER_44_2612 ();
 sg13g2_decap_8 FILLER_44_2619 ();
 sg13g2_decap_8 FILLER_44_2626 ();
 sg13g2_decap_8 FILLER_44_2633 ();
 sg13g2_decap_8 FILLER_44_2640 ();
 sg13g2_decap_8 FILLER_44_2647 ();
 sg13g2_decap_8 FILLER_44_2654 ();
 sg13g2_decap_8 FILLER_44_2661 ();
 sg13g2_fill_2 FILLER_44_2668 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_7 ();
 sg13g2_fill_1 FILLER_45_31 ();
 sg13g2_decap_8 FILLER_45_40 ();
 sg13g2_decap_8 FILLER_45_47 ();
 sg13g2_decap_8 FILLER_45_54 ();
 sg13g2_decap_8 FILLER_45_61 ();
 sg13g2_decap_8 FILLER_45_68 ();
 sg13g2_decap_8 FILLER_45_75 ();
 sg13g2_decap_8 FILLER_45_82 ();
 sg13g2_fill_2 FILLER_45_89 ();
 sg13g2_fill_1 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_96 ();
 sg13g2_decap_4 FILLER_45_103 ();
 sg13g2_fill_2 FILLER_45_107 ();
 sg13g2_fill_2 FILLER_45_122 ();
 sg13g2_fill_1 FILLER_45_159 ();
 sg13g2_decap_8 FILLER_45_164 ();
 sg13g2_decap_8 FILLER_45_171 ();
 sg13g2_fill_1 FILLER_45_182 ();
 sg13g2_fill_2 FILLER_45_214 ();
 sg13g2_fill_2 FILLER_45_242 ();
 sg13g2_fill_1 FILLER_45_302 ();
 sg13g2_fill_1 FILLER_45_306 ();
 sg13g2_fill_1 FILLER_45_373 ();
 sg13g2_fill_1 FILLER_45_405 ();
 sg13g2_fill_1 FILLER_45_409 ();
 sg13g2_fill_2 FILLER_45_436 ();
 sg13g2_decap_8 FILLER_45_499 ();
 sg13g2_decap_8 FILLER_45_506 ();
 sg13g2_decap_8 FILLER_45_519 ();
 sg13g2_decap_8 FILLER_45_526 ();
 sg13g2_decap_4 FILLER_45_542 ();
 sg13g2_fill_1 FILLER_45_546 ();
 sg13g2_fill_2 FILLER_45_553 ();
 sg13g2_fill_2 FILLER_45_616 ();
 sg13g2_fill_2 FILLER_45_622 ();
 sg13g2_fill_2 FILLER_45_628 ();
 sg13g2_fill_1 FILLER_45_630 ();
 sg13g2_fill_2 FILLER_45_654 ();
 sg13g2_decap_8 FILLER_45_662 ();
 sg13g2_fill_2 FILLER_45_669 ();
 sg13g2_fill_1 FILLER_45_671 ();
 sg13g2_decap_8 FILLER_45_676 ();
 sg13g2_decap_8 FILLER_45_683 ();
 sg13g2_decap_8 FILLER_45_690 ();
 sg13g2_fill_2 FILLER_45_697 ();
 sg13g2_fill_1 FILLER_45_699 ();
 sg13g2_fill_1 FILLER_45_704 ();
 sg13g2_fill_1 FILLER_45_714 ();
 sg13g2_fill_2 FILLER_45_720 ();
 sg13g2_decap_8 FILLER_45_727 ();
 sg13g2_decap_4 FILLER_45_734 ();
 sg13g2_fill_2 FILLER_45_754 ();
 sg13g2_fill_1 FILLER_45_766 ();
 sg13g2_fill_1 FILLER_45_777 ();
 sg13g2_fill_1 FILLER_45_781 ();
 sg13g2_fill_2 FILLER_45_792 ();
 sg13g2_fill_1 FILLER_45_856 ();
 sg13g2_fill_1 FILLER_45_883 ();
 sg13g2_fill_2 FILLER_45_910 ();
 sg13g2_fill_1 FILLER_45_912 ();
 sg13g2_fill_1 FILLER_45_923 ();
 sg13g2_fill_2 FILLER_45_987 ();
 sg13g2_fill_1 FILLER_45_1015 ();
 sg13g2_fill_1 FILLER_45_1087 ();
 sg13g2_fill_1 FILLER_45_1118 ();
 sg13g2_fill_1 FILLER_45_1185 ();
 sg13g2_fill_1 FILLER_45_1203 ();
 sg13g2_decap_8 FILLER_45_1225 ();
 sg13g2_decap_8 FILLER_45_1232 ();
 sg13g2_decap_8 FILLER_45_1239 ();
 sg13g2_decap_4 FILLER_45_1246 ();
 sg13g2_fill_1 FILLER_45_1250 ();
 sg13g2_decap_4 FILLER_45_1256 ();
 sg13g2_fill_2 FILLER_45_1260 ();
 sg13g2_decap_4 FILLER_45_1267 ();
 sg13g2_fill_2 FILLER_45_1271 ();
 sg13g2_decap_8 FILLER_45_1278 ();
 sg13g2_fill_2 FILLER_45_1285 ();
 sg13g2_fill_1 FILLER_45_1292 ();
 sg13g2_fill_1 FILLER_45_1301 ();
 sg13g2_fill_1 FILLER_45_1312 ();
 sg13g2_fill_2 FILLER_45_1324 ();
 sg13g2_decap_8 FILLER_45_1333 ();
 sg13g2_fill_1 FILLER_45_1343 ();
 sg13g2_fill_2 FILLER_45_1348 ();
 sg13g2_fill_1 FILLER_45_1350 ();
 sg13g2_decap_8 FILLER_45_1356 ();
 sg13g2_decap_8 FILLER_45_1363 ();
 sg13g2_decap_4 FILLER_45_1370 ();
 sg13g2_decap_8 FILLER_45_1379 ();
 sg13g2_fill_2 FILLER_45_1386 ();
 sg13g2_fill_1 FILLER_45_1388 ();
 sg13g2_fill_2 FILLER_45_1402 ();
 sg13g2_decap_8 FILLER_45_1408 ();
 sg13g2_fill_1 FILLER_45_1423 ();
 sg13g2_fill_2 FILLER_45_1475 ();
 sg13g2_fill_1 FILLER_45_1477 ();
 sg13g2_fill_2 FILLER_45_1484 ();
 sg13g2_decap_8 FILLER_45_1490 ();
 sg13g2_fill_2 FILLER_45_1497 ();
 sg13g2_decap_8 FILLER_45_1502 ();
 sg13g2_decap_8 FILLER_45_1509 ();
 sg13g2_fill_1 FILLER_45_1516 ();
 sg13g2_decap_4 FILLER_45_1521 ();
 sg13g2_fill_2 FILLER_45_1538 ();
 sg13g2_fill_1 FILLER_45_1540 ();
 sg13g2_fill_2 FILLER_45_1551 ();
 sg13g2_fill_2 FILLER_45_1574 ();
 sg13g2_fill_1 FILLER_45_1576 ();
 sg13g2_decap_4 FILLER_45_1586 ();
 sg13g2_fill_2 FILLER_45_1604 ();
 sg13g2_decap_4 FILLER_45_1619 ();
 sg13g2_fill_1 FILLER_45_1623 ();
 sg13g2_fill_1 FILLER_45_1645 ();
 sg13g2_fill_1 FILLER_45_1651 ();
 sg13g2_decap_4 FILLER_45_1660 ();
 sg13g2_fill_2 FILLER_45_1664 ();
 sg13g2_fill_2 FILLER_45_1671 ();
 sg13g2_fill_2 FILLER_45_1740 ();
 sg13g2_decap_4 FILLER_45_1779 ();
 sg13g2_decap_8 FILLER_45_1801 ();
 sg13g2_decap_4 FILLER_45_1808 ();
 sg13g2_decap_8 FILLER_45_1816 ();
 sg13g2_fill_1 FILLER_45_1823 ();
 sg13g2_fill_2 FILLER_45_1855 ();
 sg13g2_fill_1 FILLER_45_1892 ();
 sg13g2_decap_4 FILLER_45_1902 ();
 sg13g2_fill_1 FILLER_45_1951 ();
 sg13g2_decap_8 FILLER_45_2043 ();
 sg13g2_fill_1 FILLER_45_2050 ();
 sg13g2_fill_1 FILLER_45_2085 ();
 sg13g2_fill_2 FILLER_45_2107 ();
 sg13g2_fill_2 FILLER_45_2140 ();
 sg13g2_fill_2 FILLER_45_2278 ();
 sg13g2_decap_4 FILLER_45_2332 ();
 sg13g2_fill_1 FILLER_45_2405 ();
 sg13g2_fill_1 FILLER_45_2419 ();
 sg13g2_fill_2 FILLER_45_2444 ();
 sg13g2_fill_1 FILLER_45_2459 ();
 sg13g2_fill_2 FILLER_45_2506 ();
 sg13g2_decap_8 FILLER_45_2512 ();
 sg13g2_decap_8 FILLER_45_2519 ();
 sg13g2_decap_8 FILLER_45_2526 ();
 sg13g2_decap_8 FILLER_45_2533 ();
 sg13g2_decap_8 FILLER_45_2540 ();
 sg13g2_decap_8 FILLER_45_2547 ();
 sg13g2_decap_8 FILLER_45_2554 ();
 sg13g2_decap_8 FILLER_45_2561 ();
 sg13g2_decap_8 FILLER_45_2568 ();
 sg13g2_decap_8 FILLER_45_2575 ();
 sg13g2_decap_8 FILLER_45_2582 ();
 sg13g2_decap_8 FILLER_45_2589 ();
 sg13g2_decap_8 FILLER_45_2596 ();
 sg13g2_decap_8 FILLER_45_2603 ();
 sg13g2_decap_8 FILLER_45_2610 ();
 sg13g2_decap_8 FILLER_45_2617 ();
 sg13g2_decap_8 FILLER_45_2624 ();
 sg13g2_decap_8 FILLER_45_2631 ();
 sg13g2_decap_8 FILLER_45_2638 ();
 sg13g2_decap_8 FILLER_45_2645 ();
 sg13g2_decap_8 FILLER_45_2652 ();
 sg13g2_decap_8 FILLER_45_2659 ();
 sg13g2_decap_4 FILLER_45_2666 ();
 sg13g2_decap_4 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_4 ();
 sg13g2_decap_8 FILLER_46_39 ();
 sg13g2_decap_8 FILLER_46_46 ();
 sg13g2_decap_4 FILLER_46_83 ();
 sg13g2_fill_1 FILLER_46_87 ();
 sg13g2_fill_1 FILLER_46_124 ();
 sg13g2_fill_2 FILLER_46_128 ();
 sg13g2_fill_1 FILLER_46_130 ();
 sg13g2_fill_1 FILLER_46_175 ();
 sg13g2_fill_1 FILLER_46_199 ();
 sg13g2_fill_1 FILLER_46_238 ();
 sg13g2_fill_1 FILLER_46_269 ();
 sg13g2_fill_1 FILLER_46_274 ();
 sg13g2_fill_1 FILLER_46_289 ();
 sg13g2_fill_1 FILLER_46_307 ();
 sg13g2_fill_1 FILLER_46_333 ();
 sg13g2_fill_1 FILLER_46_362 ();
 sg13g2_fill_2 FILLER_46_374 ();
 sg13g2_fill_1 FILLER_46_386 ();
 sg13g2_fill_2 FILLER_46_435 ();
 sg13g2_fill_1 FILLER_46_474 ();
 sg13g2_decap_4 FILLER_46_527 ();
 sg13g2_decap_8 FILLER_46_535 ();
 sg13g2_fill_1 FILLER_46_542 ();
 sg13g2_fill_1 FILLER_46_547 ();
 sg13g2_fill_2 FILLER_46_579 ();
 sg13g2_fill_2 FILLER_46_619 ();
 sg13g2_decap_8 FILLER_46_648 ();
 sg13g2_decap_8 FILLER_46_655 ();
 sg13g2_fill_1 FILLER_46_662 ();
 sg13g2_decap_8 FILLER_46_689 ();
 sg13g2_fill_2 FILLER_46_696 ();
 sg13g2_fill_1 FILLER_46_698 ();
 sg13g2_decap_8 FILLER_46_735 ();
 sg13g2_fill_1 FILLER_46_742 ();
 sg13g2_fill_2 FILLER_46_748 ();
 sg13g2_decap_8 FILLER_46_759 ();
 sg13g2_decap_8 FILLER_46_813 ();
 sg13g2_decap_4 FILLER_46_820 ();
 sg13g2_decap_4 FILLER_46_833 ();
 sg13g2_fill_2 FILLER_46_851 ();
 sg13g2_fill_2 FILLER_46_913 ();
 sg13g2_fill_2 FILLER_46_968 ();
 sg13g2_fill_1 FILLER_46_1014 ();
 sg13g2_fill_2 FILLER_46_1025 ();
 sg13g2_fill_2 FILLER_46_1056 ();
 sg13g2_fill_1 FILLER_46_1076 ();
 sg13g2_fill_1 FILLER_46_1105 ();
 sg13g2_fill_1 FILLER_46_1137 ();
 sg13g2_fill_2 FILLER_46_1150 ();
 sg13g2_decap_4 FILLER_46_1182 ();
 sg13g2_fill_2 FILLER_46_1186 ();
 sg13g2_fill_2 FILLER_46_1230 ();
 sg13g2_fill_1 FILLER_46_1252 ();
 sg13g2_fill_1 FILLER_46_1261 ();
 sg13g2_fill_1 FILLER_46_1266 ();
 sg13g2_fill_1 FILLER_46_1272 ();
 sg13g2_fill_1 FILLER_46_1278 ();
 sg13g2_fill_1 FILLER_46_1287 ();
 sg13g2_decap_8 FILLER_46_1292 ();
 sg13g2_decap_4 FILLER_46_1299 ();
 sg13g2_fill_2 FILLER_46_1303 ();
 sg13g2_fill_1 FILLER_46_1335 ();
 sg13g2_decap_4 FILLER_46_1366 ();
 sg13g2_decap_8 FILLER_46_1379 ();
 sg13g2_decap_8 FILLER_46_1386 ();
 sg13g2_decap_8 FILLER_46_1393 ();
 sg13g2_decap_8 FILLER_46_1400 ();
 sg13g2_decap_4 FILLER_46_1407 ();
 sg13g2_fill_1 FILLER_46_1411 ();
 sg13g2_fill_1 FILLER_46_1420 ();
 sg13g2_fill_1 FILLER_46_1424 ();
 sg13g2_fill_2 FILLER_46_1432 ();
 sg13g2_fill_2 FILLER_46_1442 ();
 sg13g2_decap_4 FILLER_46_1448 ();
 sg13g2_fill_2 FILLER_46_1452 ();
 sg13g2_decap_8 FILLER_46_1458 ();
 sg13g2_decap_8 FILLER_46_1465 ();
 sg13g2_fill_2 FILLER_46_1472 ();
 sg13g2_fill_1 FILLER_46_1474 ();
 sg13g2_fill_1 FILLER_46_1485 ();
 sg13g2_decap_4 FILLER_46_1490 ();
 sg13g2_fill_2 FILLER_46_1494 ();
 sg13g2_fill_2 FILLER_46_1507 ();
 sg13g2_fill_2 FILLER_46_1519 ();
 sg13g2_fill_1 FILLER_46_1531 ();
 sg13g2_fill_1 FILLER_46_1536 ();
 sg13g2_fill_1 FILLER_46_1555 ();
 sg13g2_fill_2 FILLER_46_1569 ();
 sg13g2_fill_1 FILLER_46_1571 ();
 sg13g2_fill_1 FILLER_46_1577 ();
 sg13g2_fill_1 FILLER_46_1586 ();
 sg13g2_fill_2 FILLER_46_1595 ();
 sg13g2_fill_2 FILLER_46_1603 ();
 sg13g2_fill_2 FILLER_46_1671 ();
 sg13g2_fill_1 FILLER_46_1673 ();
 sg13g2_fill_1 FILLER_46_1678 ();
 sg13g2_fill_2 FILLER_46_1683 ();
 sg13g2_fill_1 FILLER_46_1689 ();
 sg13g2_decap_4 FILLER_46_1759 ();
 sg13g2_fill_2 FILLER_46_1763 ();
 sg13g2_decap_4 FILLER_46_1773 ();
 sg13g2_fill_1 FILLER_46_1777 ();
 sg13g2_decap_4 FILLER_46_1783 ();
 sg13g2_fill_1 FILLER_46_1787 ();
 sg13g2_decap_4 FILLER_46_1808 ();
 sg13g2_fill_1 FILLER_46_1812 ();
 sg13g2_decap_8 FILLER_46_1821 ();
 sg13g2_fill_1 FILLER_46_1828 ();
 sg13g2_fill_1 FILLER_46_1837 ();
 sg13g2_fill_1 FILLER_46_1883 ();
 sg13g2_fill_1 FILLER_46_1905 ();
 sg13g2_fill_1 FILLER_46_1927 ();
 sg13g2_fill_1 FILLER_46_1977 ();
 sg13g2_decap_8 FILLER_46_2008 ();
 sg13g2_decap_4 FILLER_46_2015 ();
 sg13g2_decap_8 FILLER_46_2023 ();
 sg13g2_fill_1 FILLER_46_2030 ();
 sg13g2_decap_4 FILLER_46_2037 ();
 sg13g2_fill_1 FILLER_46_2041 ();
 sg13g2_fill_1 FILLER_46_2075 ();
 sg13g2_fill_1 FILLER_46_2079 ();
 sg13g2_fill_1 FILLER_46_2106 ();
 sg13g2_fill_2 FILLER_46_2159 ();
 sg13g2_fill_2 FILLER_46_2166 ();
 sg13g2_fill_1 FILLER_46_2229 ();
 sg13g2_fill_1 FILLER_46_2252 ();
 sg13g2_fill_2 FILLER_46_2280 ();
 sg13g2_fill_1 FILLER_46_2317 ();
 sg13g2_fill_1 FILLER_46_2325 ();
 sg13g2_fill_2 FILLER_46_2335 ();
 sg13g2_fill_2 FILLER_46_2347 ();
 sg13g2_fill_2 FILLER_46_2359 ();
 sg13g2_fill_1 FILLER_46_2390 ();
 sg13g2_decap_4 FILLER_46_2414 ();
 sg13g2_fill_2 FILLER_46_2426 ();
 sg13g2_fill_1 FILLER_46_2436 ();
 sg13g2_fill_1 FILLER_46_2483 ();
 sg13g2_decap_8 FILLER_46_2529 ();
 sg13g2_decap_8 FILLER_46_2536 ();
 sg13g2_decap_8 FILLER_46_2543 ();
 sg13g2_decap_8 FILLER_46_2550 ();
 sg13g2_decap_8 FILLER_46_2557 ();
 sg13g2_decap_8 FILLER_46_2564 ();
 sg13g2_decap_8 FILLER_46_2571 ();
 sg13g2_decap_8 FILLER_46_2578 ();
 sg13g2_decap_8 FILLER_46_2585 ();
 sg13g2_decap_8 FILLER_46_2592 ();
 sg13g2_decap_8 FILLER_46_2599 ();
 sg13g2_decap_8 FILLER_46_2606 ();
 sg13g2_decap_8 FILLER_46_2613 ();
 sg13g2_decap_8 FILLER_46_2620 ();
 sg13g2_decap_8 FILLER_46_2627 ();
 sg13g2_decap_8 FILLER_46_2634 ();
 sg13g2_decap_8 FILLER_46_2641 ();
 sg13g2_decap_8 FILLER_46_2648 ();
 sg13g2_decap_8 FILLER_46_2655 ();
 sg13g2_decap_8 FILLER_46_2662 ();
 sg13g2_fill_1 FILLER_46_2669 ();
 sg13g2_fill_2 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_2 ();
 sg13g2_decap_4 FILLER_47_33 ();
 sg13g2_fill_2 FILLER_47_37 ();
 sg13g2_fill_1 FILLER_47_43 ();
 sg13g2_fill_2 FILLER_47_57 ();
 sg13g2_fill_1 FILLER_47_67 ();
 sg13g2_decap_4 FILLER_47_71 ();
 sg13g2_fill_1 FILLER_47_80 ();
 sg13g2_fill_2 FILLER_47_85 ();
 sg13g2_fill_1 FILLER_47_87 ();
 sg13g2_decap_4 FILLER_47_92 ();
 sg13g2_fill_1 FILLER_47_96 ();
 sg13g2_fill_1 FILLER_47_131 ();
 sg13g2_fill_1 FILLER_47_145 ();
 sg13g2_fill_2 FILLER_47_172 ();
 sg13g2_fill_1 FILLER_47_174 ();
 sg13g2_decap_8 FILLER_47_178 ();
 sg13g2_fill_2 FILLER_47_193 ();
 sg13g2_fill_1 FILLER_47_195 ();
 sg13g2_fill_2 FILLER_47_210 ();
 sg13g2_fill_1 FILLER_47_262 ();
 sg13g2_fill_1 FILLER_47_274 ();
 sg13g2_fill_2 FILLER_47_285 ();
 sg13g2_fill_2 FILLER_47_304 ();
 sg13g2_fill_1 FILLER_47_310 ();
 sg13g2_fill_2 FILLER_47_322 ();
 sg13g2_fill_1 FILLER_47_356 ();
 sg13g2_fill_2 FILLER_47_361 ();
 sg13g2_fill_1 FILLER_47_371 ();
 sg13g2_fill_1 FILLER_47_391 ();
 sg13g2_fill_2 FILLER_47_404 ();
 sg13g2_fill_1 FILLER_47_414 ();
 sg13g2_fill_2 FILLER_47_431 ();
 sg13g2_fill_1 FILLER_47_453 ();
 sg13g2_fill_2 FILLER_47_468 ();
 sg13g2_fill_1 FILLER_47_470 ();
 sg13g2_fill_2 FILLER_47_484 ();
 sg13g2_decap_4 FILLER_47_500 ();
 sg13g2_fill_2 FILLER_47_514 ();
 sg13g2_decap_4 FILLER_47_521 ();
 sg13g2_fill_1 FILLER_47_525 ();
 sg13g2_decap_8 FILLER_47_531 ();
 sg13g2_fill_1 FILLER_47_538 ();
 sg13g2_fill_2 FILLER_47_585 ();
 sg13g2_fill_1 FILLER_47_598 ();
 sg13g2_fill_1 FILLER_47_655 ();
 sg13g2_decap_4 FILLER_47_691 ();
 sg13g2_fill_2 FILLER_47_699 ();
 sg13g2_decap_4 FILLER_47_755 ();
 sg13g2_fill_2 FILLER_47_764 ();
 sg13g2_fill_2 FILLER_47_771 ();
 sg13g2_fill_1 FILLER_47_777 ();
 sg13g2_fill_2 FILLER_47_788 ();
 sg13g2_fill_2 FILLER_47_794 ();
 sg13g2_fill_2 FILLER_47_801 ();
 sg13g2_decap_8 FILLER_47_807 ();
 sg13g2_decap_8 FILLER_47_814 ();
 sg13g2_decap_8 FILLER_47_821 ();
 sg13g2_decap_8 FILLER_47_828 ();
 sg13g2_decap_4 FILLER_47_845 ();
 sg13g2_fill_2 FILLER_47_849 ();
 sg13g2_fill_2 FILLER_47_877 ();
 sg13g2_fill_2 FILLER_47_889 ();
 sg13g2_fill_1 FILLER_47_895 ();
 sg13g2_fill_2 FILLER_47_901 ();
 sg13g2_fill_2 FILLER_47_924 ();
 sg13g2_fill_1 FILLER_47_926 ();
 sg13g2_fill_1 FILLER_47_931 ();
 sg13g2_decap_4 FILLER_47_936 ();
 sg13g2_fill_2 FILLER_47_940 ();
 sg13g2_fill_2 FILLER_47_973 ();
 sg13g2_fill_2 FILLER_47_979 ();
 sg13g2_fill_2 FILLER_47_985 ();
 sg13g2_fill_1 FILLER_47_1000 ();
 sg13g2_fill_1 FILLER_47_1060 ();
 sg13g2_fill_2 FILLER_47_1064 ();
 sg13g2_fill_1 FILLER_47_1098 ();
 sg13g2_fill_1 FILLER_47_1124 ();
 sg13g2_fill_1 FILLER_47_1134 ();
 sg13g2_fill_1 FILLER_47_1192 ();
 sg13g2_fill_1 FILLER_47_1200 ();
 sg13g2_fill_1 FILLER_47_1209 ();
 sg13g2_fill_1 FILLER_47_1222 ();
 sg13g2_fill_2 FILLER_47_1228 ();
 sg13g2_fill_2 FILLER_47_1249 ();
 sg13g2_fill_2 FILLER_47_1268 ();
 sg13g2_fill_1 FILLER_47_1292 ();
 sg13g2_decap_4 FILLER_47_1301 ();
 sg13g2_fill_2 FILLER_47_1305 ();
 sg13g2_fill_1 FILLER_47_1339 ();
 sg13g2_decap_4 FILLER_47_1349 ();
 sg13g2_fill_1 FILLER_47_1353 ();
 sg13g2_decap_8 FILLER_47_1374 ();
 sg13g2_fill_2 FILLER_47_1406 ();
 sg13g2_fill_1 FILLER_47_1408 ();
 sg13g2_fill_2 FILLER_47_1417 ();
 sg13g2_decap_4 FILLER_47_1435 ();
 sg13g2_fill_2 FILLER_47_1439 ();
 sg13g2_decap_8 FILLER_47_1446 ();
 sg13g2_decap_8 FILLER_47_1453 ();
 sg13g2_fill_1 FILLER_47_1460 ();
 sg13g2_fill_2 FILLER_47_1486 ();
 sg13g2_fill_1 FILLER_47_1488 ();
 sg13g2_fill_1 FILLER_47_1500 ();
 sg13g2_fill_1 FILLER_47_1517 ();
 sg13g2_decap_4 FILLER_47_1527 ();
 sg13g2_fill_1 FILLER_47_1531 ();
 sg13g2_fill_1 FILLER_47_1542 ();
 sg13g2_decap_4 FILLER_47_1579 ();
 sg13g2_fill_2 FILLER_47_1597 ();
 sg13g2_fill_2 FILLER_47_1603 ();
 sg13g2_fill_2 FILLER_47_1610 ();
 sg13g2_fill_2 FILLER_47_1617 ();
 sg13g2_fill_1 FILLER_47_1619 ();
 sg13g2_fill_2 FILLER_47_1668 ();
 sg13g2_fill_1 FILLER_47_1670 ();
 sg13g2_decap_4 FILLER_47_1706 ();
 sg13g2_decap_4 FILLER_47_1715 ();
 sg13g2_fill_1 FILLER_47_1719 ();
 sg13g2_fill_2 FILLER_47_1724 ();
 sg13g2_decap_4 FILLER_47_1730 ();
 sg13g2_fill_1 FILLER_47_1734 ();
 sg13g2_fill_2 FILLER_47_1740 ();
 sg13g2_fill_1 FILLER_47_1742 ();
 sg13g2_decap_8 FILLER_47_1769 ();
 sg13g2_decap_8 FILLER_47_1776 ();
 sg13g2_decap_8 FILLER_47_1783 ();
 sg13g2_decap_4 FILLER_47_1790 ();
 sg13g2_fill_2 FILLER_47_1794 ();
 sg13g2_fill_2 FILLER_47_1822 ();
 sg13g2_fill_1 FILLER_47_1824 ();
 sg13g2_fill_1 FILLER_47_1853 ();
 sg13g2_fill_1 FILLER_47_1859 ();
 sg13g2_fill_1 FILLER_47_1894 ();
 sg13g2_fill_1 FILLER_47_1928 ();
 sg13g2_fill_2 FILLER_47_1955 ();
 sg13g2_decap_8 FILLER_47_2000 ();
 sg13g2_decap_8 FILLER_47_2007 ();
 sg13g2_decap_8 FILLER_47_2014 ();
 sg13g2_fill_2 FILLER_47_2021 ();
 sg13g2_fill_2 FILLER_47_2034 ();
 sg13g2_fill_2 FILLER_47_2046 ();
 sg13g2_fill_1 FILLER_47_2079 ();
 sg13g2_fill_1 FILLER_47_2130 ();
 sg13g2_fill_2 FILLER_47_2199 ();
 sg13g2_decap_4 FILLER_47_2305 ();
 sg13g2_fill_2 FILLER_47_2309 ();
 sg13g2_decap_8 FILLER_47_2355 ();
 sg13g2_decap_8 FILLER_47_2514 ();
 sg13g2_decap_8 FILLER_47_2521 ();
 sg13g2_decap_8 FILLER_47_2528 ();
 sg13g2_decap_8 FILLER_47_2535 ();
 sg13g2_decap_8 FILLER_47_2542 ();
 sg13g2_decap_8 FILLER_47_2549 ();
 sg13g2_decap_8 FILLER_47_2556 ();
 sg13g2_decap_8 FILLER_47_2563 ();
 sg13g2_decap_8 FILLER_47_2570 ();
 sg13g2_decap_8 FILLER_47_2577 ();
 sg13g2_decap_8 FILLER_47_2584 ();
 sg13g2_decap_8 FILLER_47_2591 ();
 sg13g2_decap_8 FILLER_47_2598 ();
 sg13g2_decap_8 FILLER_47_2605 ();
 sg13g2_decap_8 FILLER_47_2612 ();
 sg13g2_decap_8 FILLER_47_2619 ();
 sg13g2_decap_8 FILLER_47_2626 ();
 sg13g2_decap_8 FILLER_47_2633 ();
 sg13g2_decap_8 FILLER_47_2640 ();
 sg13g2_decap_8 FILLER_47_2647 ();
 sg13g2_decap_8 FILLER_47_2654 ();
 sg13g2_decap_8 FILLER_47_2661 ();
 sg13g2_fill_2 FILLER_47_2668 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_fill_2 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_20 ();
 sg13g2_fill_1 FILLER_48_66 ();
 sg13g2_fill_1 FILLER_48_82 ();
 sg13g2_fill_2 FILLER_48_106 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_fill_2 FILLER_48_152 ();
 sg13g2_fill_2 FILLER_48_158 ();
 sg13g2_decap_4 FILLER_48_164 ();
 sg13g2_fill_1 FILLER_48_168 ();
 sg13g2_decap_8 FILLER_48_174 ();
 sg13g2_decap_8 FILLER_48_181 ();
 sg13g2_fill_2 FILLER_48_188 ();
 sg13g2_fill_1 FILLER_48_190 ();
 sg13g2_fill_2 FILLER_48_221 ();
 sg13g2_fill_2 FILLER_48_306 ();
 sg13g2_fill_2 FILLER_48_316 ();
 sg13g2_fill_1 FILLER_48_322 ();
 sg13g2_fill_2 FILLER_48_328 ();
 sg13g2_fill_2 FILLER_48_346 ();
 sg13g2_fill_2 FILLER_48_369 ();
 sg13g2_fill_2 FILLER_48_385 ();
 sg13g2_fill_1 FILLER_48_460 ();
 sg13g2_decap_4 FILLER_48_466 ();
 sg13g2_fill_1 FILLER_48_470 ();
 sg13g2_fill_1 FILLER_48_475 ();
 sg13g2_fill_1 FILLER_48_502 ();
 sg13g2_fill_1 FILLER_48_508 ();
 sg13g2_decap_8 FILLER_48_513 ();
 sg13g2_decap_8 FILLER_48_520 ();
 sg13g2_fill_1 FILLER_48_527 ();
 sg13g2_fill_1 FILLER_48_567 ();
 sg13g2_fill_1 FILLER_48_619 ();
 sg13g2_fill_2 FILLER_48_625 ();
 sg13g2_fill_2 FILLER_48_653 ();
 sg13g2_fill_2 FILLER_48_660 ();
 sg13g2_fill_1 FILLER_48_696 ();
 sg13g2_fill_2 FILLER_48_732 ();
 sg13g2_fill_2 FILLER_48_760 ();
 sg13g2_fill_1 FILLER_48_762 ();
 sg13g2_fill_1 FILLER_48_767 ();
 sg13g2_fill_1 FILLER_48_804 ();
 sg13g2_fill_2 FILLER_48_834 ();
 sg13g2_fill_1 FILLER_48_836 ();
 sg13g2_decap_4 FILLER_48_863 ();
 sg13g2_fill_1 FILLER_48_867 ();
 sg13g2_decap_8 FILLER_48_881 ();
 sg13g2_fill_1 FILLER_48_888 ();
 sg13g2_fill_1 FILLER_48_899 ();
 sg13g2_fill_1 FILLER_48_924 ();
 sg13g2_fill_1 FILLER_48_957 ();
 sg13g2_fill_1 FILLER_48_1007 ();
 sg13g2_fill_1 FILLER_48_1028 ();
 sg13g2_fill_1 FILLER_48_1056 ();
 sg13g2_fill_1 FILLER_48_1069 ();
 sg13g2_fill_1 FILLER_48_1095 ();
 sg13g2_fill_2 FILLER_48_1119 ();
 sg13g2_fill_1 FILLER_48_1149 ();
 sg13g2_decap_4 FILLER_48_1166 ();
 sg13g2_fill_1 FILLER_48_1170 ();
 sg13g2_fill_2 FILLER_48_1175 ();
 sg13g2_fill_1 FILLER_48_1177 ();
 sg13g2_decap_8 FILLER_48_1183 ();
 sg13g2_fill_1 FILLER_48_1190 ();
 sg13g2_fill_1 FILLER_48_1194 ();
 sg13g2_fill_2 FILLER_48_1234 ();
 sg13g2_decap_4 FILLER_48_1244 ();
 sg13g2_fill_1 FILLER_48_1258 ();
 sg13g2_fill_1 FILLER_48_1263 ();
 sg13g2_fill_1 FILLER_48_1312 ();
 sg13g2_fill_1 FILLER_48_1332 ();
 sg13g2_fill_2 FILLER_48_1339 ();
 sg13g2_decap_4 FILLER_48_1354 ();
 sg13g2_decap_4 FILLER_48_1371 ();
 sg13g2_decap_4 FILLER_48_1379 ();
 sg13g2_decap_4 FILLER_48_1407 ();
 sg13g2_fill_2 FILLER_48_1411 ();
 sg13g2_fill_1 FILLER_48_1418 ();
 sg13g2_fill_2 FILLER_48_1442 ();
 sg13g2_fill_1 FILLER_48_1444 ();
 sg13g2_decap_8 FILLER_48_1456 ();
 sg13g2_decap_8 FILLER_48_1463 ();
 sg13g2_decap_4 FILLER_48_1470 ();
 sg13g2_fill_1 FILLER_48_1474 ();
 sg13g2_fill_2 FILLER_48_1484 ();
 sg13g2_fill_2 FILLER_48_1534 ();
 sg13g2_fill_2 FILLER_48_1541 ();
 sg13g2_fill_1 FILLER_48_1564 ();
 sg13g2_fill_2 FILLER_48_1593 ();
 sg13g2_fill_1 FILLER_48_1595 ();
 sg13g2_decap_4 FILLER_48_1606 ();
 sg13g2_fill_1 FILLER_48_1610 ();
 sg13g2_fill_2 FILLER_48_1618 ();
 sg13g2_fill_2 FILLER_48_1625 ();
 sg13g2_fill_1 FILLER_48_1627 ();
 sg13g2_fill_1 FILLER_48_1654 ();
 sg13g2_fill_2 FILLER_48_1667 ();
 sg13g2_fill_1 FILLER_48_1669 ();
 sg13g2_decap_8 FILLER_48_1702 ();
 sg13g2_decap_8 FILLER_48_1709 ();
 sg13g2_decap_8 FILLER_48_1716 ();
 sg13g2_decap_8 FILLER_48_1723 ();
 sg13g2_decap_8 FILLER_48_1730 ();
 sg13g2_decap_8 FILLER_48_1737 ();
 sg13g2_decap_4 FILLER_48_1744 ();
 sg13g2_fill_2 FILLER_48_1748 ();
 sg13g2_decap_8 FILLER_48_1758 ();
 sg13g2_decap_8 FILLER_48_1765 ();
 sg13g2_decap_8 FILLER_48_1772 ();
 sg13g2_fill_2 FILLER_48_1779 ();
 sg13g2_decap_8 FILLER_48_1785 ();
 sg13g2_fill_2 FILLER_48_1792 ();
 sg13g2_fill_1 FILLER_48_1794 ();
 sg13g2_fill_2 FILLER_48_1808 ();
 sg13g2_fill_2 FILLER_48_1818 ();
 sg13g2_fill_1 FILLER_48_1820 ();
 sg13g2_fill_1 FILLER_48_1845 ();
 sg13g2_fill_2 FILLER_48_1859 ();
 sg13g2_fill_2 FILLER_48_1887 ();
 sg13g2_fill_1 FILLER_48_1893 ();
 sg13g2_fill_2 FILLER_48_1898 ();
 sg13g2_fill_1 FILLER_48_1926 ();
 sg13g2_fill_2 FILLER_48_1953 ();
 sg13g2_fill_1 FILLER_48_1989 ();
 sg13g2_decap_8 FILLER_48_1994 ();
 sg13g2_decap_4 FILLER_48_2001 ();
 sg13g2_fill_2 FILLER_48_2009 ();
 sg13g2_fill_1 FILLER_48_2011 ();
 sg13g2_fill_1 FILLER_48_2047 ();
 sg13g2_decap_8 FILLER_48_2074 ();
 sg13g2_decap_4 FILLER_48_2081 ();
 sg13g2_fill_1 FILLER_48_2085 ();
 sg13g2_fill_2 FILLER_48_2103 ();
 sg13g2_fill_1 FILLER_48_2117 ();
 sg13g2_fill_1 FILLER_48_2122 ();
 sg13g2_fill_2 FILLER_48_2133 ();
 sg13g2_fill_2 FILLER_48_2197 ();
 sg13g2_fill_1 FILLER_48_2229 ();
 sg13g2_fill_2 FILLER_48_2236 ();
 sg13g2_decap_4 FILLER_48_2397 ();
 sg13g2_fill_2 FILLER_48_2401 ();
 sg13g2_fill_1 FILLER_48_2413 ();
 sg13g2_fill_1 FILLER_48_2424 ();
 sg13g2_fill_1 FILLER_48_2467 ();
 sg13g2_fill_2 FILLER_48_2507 ();
 sg13g2_decap_8 FILLER_48_2513 ();
 sg13g2_decap_8 FILLER_48_2520 ();
 sg13g2_decap_8 FILLER_48_2527 ();
 sg13g2_decap_8 FILLER_48_2534 ();
 sg13g2_decap_8 FILLER_48_2541 ();
 sg13g2_decap_8 FILLER_48_2548 ();
 sg13g2_decap_8 FILLER_48_2555 ();
 sg13g2_decap_8 FILLER_48_2562 ();
 sg13g2_decap_8 FILLER_48_2569 ();
 sg13g2_decap_8 FILLER_48_2576 ();
 sg13g2_decap_8 FILLER_48_2583 ();
 sg13g2_decap_8 FILLER_48_2590 ();
 sg13g2_decap_8 FILLER_48_2597 ();
 sg13g2_decap_8 FILLER_48_2604 ();
 sg13g2_decap_8 FILLER_48_2611 ();
 sg13g2_decap_8 FILLER_48_2618 ();
 sg13g2_decap_8 FILLER_48_2625 ();
 sg13g2_decap_8 FILLER_48_2632 ();
 sg13g2_decap_8 FILLER_48_2639 ();
 sg13g2_decap_8 FILLER_48_2646 ();
 sg13g2_decap_8 FILLER_48_2653 ();
 sg13g2_decap_8 FILLER_48_2660 ();
 sg13g2_fill_2 FILLER_48_2667 ();
 sg13g2_fill_1 FILLER_48_2669 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_fill_2 FILLER_49_21 ();
 sg13g2_fill_1 FILLER_49_23 ();
 sg13g2_fill_2 FILLER_49_54 ();
 sg13g2_fill_1 FILLER_49_85 ();
 sg13g2_fill_1 FILLER_49_91 ();
 sg13g2_fill_1 FILLER_49_97 ();
 sg13g2_fill_1 FILLER_49_107 ();
 sg13g2_fill_1 FILLER_49_113 ();
 sg13g2_decap_8 FILLER_49_117 ();
 sg13g2_decap_4 FILLER_49_124 ();
 sg13g2_decap_8 FILLER_49_131 ();
 sg13g2_decap_8 FILLER_49_138 ();
 sg13g2_decap_8 FILLER_49_145 ();
 sg13g2_decap_4 FILLER_49_152 ();
 sg13g2_fill_1 FILLER_49_156 ();
 sg13g2_fill_1 FILLER_49_166 ();
 sg13g2_fill_1 FILLER_49_171 ();
 sg13g2_fill_2 FILLER_49_191 ();
 sg13g2_fill_1 FILLER_49_210 ();
 sg13g2_fill_1 FILLER_49_227 ();
 sg13g2_fill_1 FILLER_49_314 ();
 sg13g2_fill_1 FILLER_49_366 ();
 sg13g2_fill_1 FILLER_49_392 ();
 sg13g2_fill_1 FILLER_49_409 ();
 sg13g2_fill_1 FILLER_49_424 ();
 sg13g2_fill_1 FILLER_49_471 ();
 sg13g2_fill_1 FILLER_49_477 ();
 sg13g2_fill_1 FILLER_49_482 ();
 sg13g2_fill_1 FILLER_49_487 ();
 sg13g2_decap_8 FILLER_49_503 ();
 sg13g2_fill_1 FILLER_49_510 ();
 sg13g2_decap_8 FILLER_49_521 ();
 sg13g2_fill_1 FILLER_49_528 ();
 sg13g2_fill_1 FILLER_49_543 ();
 sg13g2_decap_8 FILLER_49_625 ();
 sg13g2_fill_2 FILLER_49_632 ();
 sg13g2_fill_1 FILLER_49_634 ();
 sg13g2_decap_4 FILLER_49_644 ();
 sg13g2_fill_2 FILLER_49_648 ();
 sg13g2_fill_2 FILLER_49_672 ();
 sg13g2_decap_4 FILLER_49_682 ();
 sg13g2_fill_1 FILLER_49_686 ();
 sg13g2_fill_2 FILLER_49_700 ();
 sg13g2_fill_2 FILLER_49_728 ();
 sg13g2_decap_8 FILLER_49_775 ();
 sg13g2_decap_8 FILLER_49_782 ();
 sg13g2_decap_4 FILLER_49_789 ();
 sg13g2_fill_1 FILLER_49_849 ();
 sg13g2_decap_8 FILLER_49_886 ();
 sg13g2_fill_2 FILLER_49_893 ();
 sg13g2_fill_1 FILLER_49_895 ();
 sg13g2_fill_2 FILLER_49_900 ();
 sg13g2_decap_8 FILLER_49_906 ();
 sg13g2_decap_8 FILLER_49_913 ();
 sg13g2_fill_2 FILLER_49_920 ();
 sg13g2_decap_4 FILLER_49_932 ();
 sg13g2_fill_2 FILLER_49_936 ();
 sg13g2_fill_2 FILLER_49_942 ();
 sg13g2_fill_1 FILLER_49_944 ();
 sg13g2_fill_2 FILLER_49_1016 ();
 sg13g2_fill_2 FILLER_49_1038 ();
 sg13g2_fill_2 FILLER_49_1067 ();
 sg13g2_fill_1 FILLER_49_1077 ();
 sg13g2_fill_1 FILLER_49_1087 ();
 sg13g2_fill_2 FILLER_49_1156 ();
 sg13g2_fill_1 FILLER_49_1158 ();
 sg13g2_decap_8 FILLER_49_1166 ();
 sg13g2_decap_4 FILLER_49_1173 ();
 sg13g2_fill_2 FILLER_49_1182 ();
 sg13g2_fill_1 FILLER_49_1184 ();
 sg13g2_fill_2 FILLER_49_1189 ();
 sg13g2_fill_2 FILLER_49_1199 ();
 sg13g2_fill_1 FILLER_49_1201 ();
 sg13g2_fill_2 FILLER_49_1219 ();
 sg13g2_fill_1 FILLER_49_1233 ();
 sg13g2_decap_4 FILLER_49_1242 ();
 sg13g2_decap_8 FILLER_49_1250 ();
 sg13g2_fill_1 FILLER_49_1257 ();
 sg13g2_fill_2 FILLER_49_1262 ();
 sg13g2_fill_2 FILLER_49_1269 ();
 sg13g2_fill_1 FILLER_49_1275 ();
 sg13g2_fill_2 FILLER_49_1279 ();
 sg13g2_fill_1 FILLER_49_1281 ();
 sg13g2_fill_2 FILLER_49_1286 ();
 sg13g2_decap_4 FILLER_49_1300 ();
 sg13g2_decap_8 FILLER_49_1316 ();
 sg13g2_fill_2 FILLER_49_1348 ();
 sg13g2_decap_4 FILLER_49_1367 ();
 sg13g2_fill_2 FILLER_49_1371 ();
 sg13g2_decap_8 FILLER_49_1378 ();
 sg13g2_decap_4 FILLER_49_1394 ();
 sg13g2_fill_2 FILLER_49_1398 ();
 sg13g2_fill_2 FILLER_49_1408 ();
 sg13g2_fill_1 FILLER_49_1410 ();
 sg13g2_fill_1 FILLER_49_1416 ();
 sg13g2_decap_8 FILLER_49_1421 ();
 sg13g2_fill_2 FILLER_49_1428 ();
 sg13g2_decap_8 FILLER_49_1450 ();
 sg13g2_fill_1 FILLER_49_1457 ();
 sg13g2_decap_4 FILLER_49_1468 ();
 sg13g2_fill_1 FILLER_49_1472 ();
 sg13g2_fill_2 FILLER_49_1502 ();
 sg13g2_decap_4 FILLER_49_1512 ();
 sg13g2_fill_1 FILLER_49_1516 ();
 sg13g2_fill_2 FILLER_49_1521 ();
 sg13g2_decap_8 FILLER_49_1526 ();
 sg13g2_fill_1 FILLER_49_1549 ();
 sg13g2_fill_1 FILLER_49_1563 ();
 sg13g2_decap_8 FILLER_49_1585 ();
 sg13g2_decap_8 FILLER_49_1592 ();
 sg13g2_fill_2 FILLER_49_1599 ();
 sg13g2_fill_1 FILLER_49_1601 ();
 sg13g2_decap_8 FILLER_49_1610 ();
 sg13g2_fill_2 FILLER_49_1617 ();
 sg13g2_fill_1 FILLER_49_1619 ();
 sg13g2_decap_8 FILLER_49_1638 ();
 sg13g2_fill_2 FILLER_49_1645 ();
 sg13g2_decap_8 FILLER_49_1655 ();
 sg13g2_fill_2 FILLER_49_1662 ();
 sg13g2_decap_8 FILLER_49_1669 ();
 sg13g2_decap_8 FILLER_49_1676 ();
 sg13g2_fill_2 FILLER_49_1696 ();
 sg13g2_decap_4 FILLER_49_1739 ();
 sg13g2_fill_1 FILLER_49_1743 ();
 sg13g2_fill_1 FILLER_49_1800 ();
 sg13g2_fill_2 FILLER_49_1841 ();
 sg13g2_fill_2 FILLER_49_1859 ();
 sg13g2_fill_1 FILLER_49_1872 ();
 sg13g2_decap_8 FILLER_49_1877 ();
 sg13g2_fill_2 FILLER_49_1884 ();
 sg13g2_fill_1 FILLER_49_1886 ();
 sg13g2_decap_4 FILLER_49_1943 ();
 sg13g2_fill_1 FILLER_49_1947 ();
 sg13g2_decap_4 FILLER_49_1978 ();
 sg13g2_decap_8 FILLER_49_1986 ();
 sg13g2_decap_8 FILLER_49_1993 ();
 sg13g2_fill_2 FILLER_49_2000 ();
 sg13g2_fill_1 FILLER_49_2002 ();
 sg13g2_decap_4 FILLER_49_2027 ();
 sg13g2_fill_2 FILLER_49_2031 ();
 sg13g2_fill_2 FILLER_49_2060 ();
 sg13g2_decap_8 FILLER_49_2072 ();
 sg13g2_decap_4 FILLER_49_2079 ();
 sg13g2_fill_1 FILLER_49_2083 ();
 sg13g2_fill_1 FILLER_49_2088 ();
 sg13g2_fill_2 FILLER_49_2103 ();
 sg13g2_fill_2 FILLER_49_2112 ();
 sg13g2_fill_2 FILLER_49_2117 ();
 sg13g2_fill_1 FILLER_49_2132 ();
 sg13g2_fill_2 FILLER_49_2166 ();
 sg13g2_fill_2 FILLER_49_2270 ();
 sg13g2_fill_2 FILLER_49_2305 ();
 sg13g2_fill_1 FILLER_49_2307 ();
 sg13g2_decap_4 FILLER_49_2318 ();
 sg13g2_fill_2 FILLER_49_2322 ();
 sg13g2_fill_1 FILLER_49_2383 ();
 sg13g2_decap_4 FILLER_49_2390 ();
 sg13g2_fill_1 FILLER_49_2394 ();
 sg13g2_fill_1 FILLER_49_2405 ();
 sg13g2_fill_2 FILLER_49_2410 ();
 sg13g2_fill_1 FILLER_49_2416 ();
 sg13g2_fill_1 FILLER_49_2443 ();
 sg13g2_fill_1 FILLER_49_2448 ();
 sg13g2_fill_1 FILLER_49_2459 ();
 sg13g2_fill_1 FILLER_49_2500 ();
 sg13g2_fill_2 FILLER_49_2531 ();
 sg13g2_fill_1 FILLER_49_2533 ();
 sg13g2_decap_8 FILLER_49_2560 ();
 sg13g2_decap_8 FILLER_49_2567 ();
 sg13g2_decap_8 FILLER_49_2574 ();
 sg13g2_decap_8 FILLER_49_2581 ();
 sg13g2_decap_8 FILLER_49_2588 ();
 sg13g2_decap_8 FILLER_49_2595 ();
 sg13g2_decap_8 FILLER_49_2602 ();
 sg13g2_decap_8 FILLER_49_2609 ();
 sg13g2_decap_8 FILLER_49_2616 ();
 sg13g2_decap_8 FILLER_49_2623 ();
 sg13g2_decap_8 FILLER_49_2630 ();
 sg13g2_decap_8 FILLER_49_2637 ();
 sg13g2_decap_8 FILLER_49_2644 ();
 sg13g2_decap_8 FILLER_49_2651 ();
 sg13g2_decap_8 FILLER_49_2658 ();
 sg13g2_decap_4 FILLER_49_2665 ();
 sg13g2_fill_1 FILLER_49_2669 ();
 sg13g2_fill_2 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_41 ();
 sg13g2_decap_4 FILLER_50_48 ();
 sg13g2_fill_2 FILLER_50_52 ();
 sg13g2_fill_1 FILLER_50_82 ();
 sg13g2_fill_1 FILLER_50_92 ();
 sg13g2_fill_1 FILLER_50_110 ();
 sg13g2_fill_2 FILLER_50_130 ();
 sg13g2_fill_2 FILLER_50_137 ();
 sg13g2_fill_1 FILLER_50_145 ();
 sg13g2_fill_1 FILLER_50_150 ();
 sg13g2_fill_1 FILLER_50_158 ();
 sg13g2_fill_1 FILLER_50_164 ();
 sg13g2_fill_2 FILLER_50_176 ();
 sg13g2_fill_2 FILLER_50_243 ();
 sg13g2_fill_1 FILLER_50_245 ();
 sg13g2_fill_2 FILLER_50_250 ();
 sg13g2_fill_1 FILLER_50_261 ();
 sg13g2_fill_1 FILLER_50_277 ();
 sg13g2_fill_1 FILLER_50_310 ();
 sg13g2_fill_1 FILLER_50_346 ();
 sg13g2_fill_1 FILLER_50_358 ();
 sg13g2_fill_1 FILLER_50_364 ();
 sg13g2_fill_1 FILLER_50_373 ();
 sg13g2_fill_2 FILLER_50_379 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_fill_2 FILLER_50_446 ();
 sg13g2_fill_2 FILLER_50_453 ();
 sg13g2_fill_1 FILLER_50_465 ();
 sg13g2_fill_1 FILLER_50_492 ();
 sg13g2_fill_1 FILLER_50_497 ();
 sg13g2_fill_1 FILLER_50_536 ();
 sg13g2_fill_1 FILLER_50_542 ();
 sg13g2_fill_1 FILLER_50_548 ();
 sg13g2_fill_1 FILLER_50_554 ();
 sg13g2_fill_2 FILLER_50_560 ();
 sg13g2_fill_1 FILLER_50_580 ();
 sg13g2_decap_8 FILLER_50_614 ();
 sg13g2_decap_8 FILLER_50_621 ();
 sg13g2_fill_1 FILLER_50_628 ();
 sg13g2_decap_8 FILLER_50_637 ();
 sg13g2_fill_2 FILLER_50_644 ();
 sg13g2_fill_2 FILLER_50_668 ();
 sg13g2_fill_1 FILLER_50_670 ();
 sg13g2_decap_8 FILLER_50_681 ();
 sg13g2_decap_8 FILLER_50_688 ();
 sg13g2_decap_8 FILLER_50_695 ();
 sg13g2_fill_1 FILLER_50_728 ();
 sg13g2_fill_2 FILLER_50_761 ();
 sg13g2_fill_1 FILLER_50_763 ();
 sg13g2_decap_4 FILLER_50_790 ();
 sg13g2_fill_1 FILLER_50_794 ();
 sg13g2_fill_1 FILLER_50_799 ();
 sg13g2_fill_1 FILLER_50_835 ();
 sg13g2_fill_1 FILLER_50_840 ();
 sg13g2_fill_2 FILLER_50_844 ();
 sg13g2_fill_2 FILLER_50_853 ();
 sg13g2_fill_1 FILLER_50_855 ();
 sg13g2_decap_4 FILLER_50_860 ();
 sg13g2_fill_1 FILLER_50_875 ();
 sg13g2_fill_2 FILLER_50_880 ();
 sg13g2_fill_1 FILLER_50_882 ();
 sg13g2_decap_4 FILLER_50_916 ();
 sg13g2_fill_2 FILLER_50_920 ();
 sg13g2_fill_2 FILLER_50_961 ();
 sg13g2_fill_2 FILLER_50_982 ();
 sg13g2_fill_2 FILLER_50_992 ();
 sg13g2_fill_2 FILLER_50_1005 ();
 sg13g2_fill_1 FILLER_50_1045 ();
 sg13g2_fill_1 FILLER_50_1068 ();
 sg13g2_fill_1 FILLER_50_1107 ();
 sg13g2_fill_2 FILLER_50_1147 ();
 sg13g2_fill_1 FILLER_50_1162 ();
 sg13g2_fill_2 FILLER_50_1175 ();
 sg13g2_fill_1 FILLER_50_1177 ();
 sg13g2_decap_8 FILLER_50_1187 ();
 sg13g2_decap_4 FILLER_50_1194 ();
 sg13g2_fill_1 FILLER_50_1198 ();
 sg13g2_decap_4 FILLER_50_1202 ();
 sg13g2_fill_2 FILLER_50_1211 ();
 sg13g2_fill_1 FILLER_50_1220 ();
 sg13g2_decap_4 FILLER_50_1225 ();
 sg13g2_decap_4 FILLER_50_1238 ();
 sg13g2_fill_2 FILLER_50_1250 ();
 sg13g2_fill_1 FILLER_50_1252 ();
 sg13g2_fill_1 FILLER_50_1265 ();
 sg13g2_decap_8 FILLER_50_1271 ();
 sg13g2_decap_4 FILLER_50_1278 ();
 sg13g2_decap_4 FILLER_50_1292 ();
 sg13g2_decap_4 FILLER_50_1312 ();
 sg13g2_fill_2 FILLER_50_1316 ();
 sg13g2_fill_2 FILLER_50_1328 ();
 sg13g2_fill_2 FILLER_50_1343 ();
 sg13g2_fill_1 FILLER_50_1345 ();
 sg13g2_fill_1 FILLER_50_1356 ();
 sg13g2_fill_1 FILLER_50_1382 ();
 sg13g2_fill_2 FILLER_50_1388 ();
 sg13g2_fill_1 FILLER_50_1390 ();
 sg13g2_fill_2 FILLER_50_1395 ();
 sg13g2_fill_2 FILLER_50_1405 ();
 sg13g2_fill_1 FILLER_50_1417 ();
 sg13g2_fill_2 FILLER_50_1427 ();
 sg13g2_fill_1 FILLER_50_1429 ();
 sg13g2_decap_4 FILLER_50_1435 ();
 sg13g2_decap_4 FILLER_50_1447 ();
 sg13g2_decap_4 FILLER_50_1455 ();
 sg13g2_fill_2 FILLER_50_1471 ();
 sg13g2_fill_1 FILLER_50_1490 ();
 sg13g2_fill_1 FILLER_50_1498 ();
 sg13g2_fill_2 FILLER_50_1521 ();
 sg13g2_fill_1 FILLER_50_1526 ();
 sg13g2_decap_8 FILLER_50_1539 ();
 sg13g2_fill_1 FILLER_50_1558 ();
 sg13g2_fill_2 FILLER_50_1564 ();
 sg13g2_fill_2 FILLER_50_1579 ();
 sg13g2_fill_2 FILLER_50_1607 ();
 sg13g2_fill_1 FILLER_50_1609 ();
 sg13g2_decap_8 FILLER_50_1636 ();
 sg13g2_fill_1 FILLER_50_1643 ();
 sg13g2_fill_2 FILLER_50_1648 ();
 sg13g2_decap_8 FILLER_50_1686 ();
 sg13g2_decap_4 FILLER_50_1723 ();
 sg13g2_decap_8 FILLER_50_1753 ();
 sg13g2_fill_2 FILLER_50_1760 ();
 sg13g2_fill_1 FILLER_50_1762 ();
 sg13g2_decap_8 FILLER_50_1793 ();
 sg13g2_decap_8 FILLER_50_1800 ();
 sg13g2_decap_4 FILLER_50_1807 ();
 sg13g2_fill_2 FILLER_50_1811 ();
 sg13g2_decap_8 FILLER_50_1848 ();
 sg13g2_fill_1 FILLER_50_1855 ();
 sg13g2_decap_8 FILLER_50_1865 ();
 sg13g2_decap_8 FILLER_50_1872 ();
 sg13g2_fill_2 FILLER_50_1879 ();
 sg13g2_fill_1 FILLER_50_1881 ();
 sg13g2_decap_8 FILLER_50_1886 ();
 sg13g2_decap_8 FILLER_50_1897 ();
 sg13g2_decap_4 FILLER_50_1904 ();
 sg13g2_fill_1 FILLER_50_1908 ();
 sg13g2_decap_8 FILLER_50_1913 ();
 sg13g2_decap_4 FILLER_50_1920 ();
 sg13g2_fill_2 FILLER_50_1932 ();
 sg13g2_fill_1 FILLER_50_1934 ();
 sg13g2_decap_8 FILLER_50_1939 ();
 sg13g2_decap_8 FILLER_50_1946 ();
 sg13g2_decap_4 FILLER_50_1953 ();
 sg13g2_fill_1 FILLER_50_1957 ();
 sg13g2_decap_8 FILLER_50_1962 ();
 sg13g2_decap_8 FILLER_50_1969 ();
 sg13g2_decap_8 FILLER_50_1976 ();
 sg13g2_fill_2 FILLER_50_1983 ();
 sg13g2_fill_1 FILLER_50_1985 ();
 sg13g2_decap_8 FILLER_50_2017 ();
 sg13g2_fill_2 FILLER_50_2024 ();
 sg13g2_fill_2 FILLER_50_2062 ();
 sg13g2_fill_1 FILLER_50_2068 ();
 sg13g2_fill_2 FILLER_50_2130 ();
 sg13g2_fill_1 FILLER_50_2136 ();
 sg13g2_fill_1 FILLER_50_2140 ();
 sg13g2_fill_1 FILLER_50_2226 ();
 sg13g2_fill_1 FILLER_50_2249 ();
 sg13g2_fill_1 FILLER_50_2260 ();
 sg13g2_fill_2 FILLER_50_2287 ();
 sg13g2_fill_2 FILLER_50_2315 ();
 sg13g2_fill_2 FILLER_50_2327 ();
 sg13g2_fill_1 FILLER_50_2329 ();
 sg13g2_decap_4 FILLER_50_2334 ();
 sg13g2_decap_4 FILLER_50_2378 ();
 sg13g2_fill_1 FILLER_50_2450 ();
 sg13g2_fill_2 FILLER_50_2497 ();
 sg13g2_decap_4 FILLER_50_2522 ();
 sg13g2_fill_2 FILLER_50_2526 ();
 sg13g2_decap_8 FILLER_50_2564 ();
 sg13g2_decap_8 FILLER_50_2571 ();
 sg13g2_decap_8 FILLER_50_2578 ();
 sg13g2_decap_8 FILLER_50_2585 ();
 sg13g2_decap_8 FILLER_50_2592 ();
 sg13g2_decap_8 FILLER_50_2599 ();
 sg13g2_decap_8 FILLER_50_2606 ();
 sg13g2_decap_8 FILLER_50_2613 ();
 sg13g2_decap_8 FILLER_50_2620 ();
 sg13g2_decap_8 FILLER_50_2627 ();
 sg13g2_decap_8 FILLER_50_2634 ();
 sg13g2_decap_8 FILLER_50_2641 ();
 sg13g2_decap_8 FILLER_50_2648 ();
 sg13g2_decap_8 FILLER_50_2655 ();
 sg13g2_decap_8 FILLER_50_2662 ();
 sg13g2_fill_1 FILLER_50_2669 ();
 sg13g2_fill_1 FILLER_51_0 ();
 sg13g2_fill_2 FILLER_51_31 ();
 sg13g2_fill_1 FILLER_51_38 ();
 sg13g2_fill_2 FILLER_51_42 ();
 sg13g2_fill_1 FILLER_51_44 ();
 sg13g2_decap_4 FILLER_51_54 ();
 sg13g2_fill_1 FILLER_51_58 ();
 sg13g2_fill_2 FILLER_51_79 ();
 sg13g2_fill_1 FILLER_51_81 ();
 sg13g2_fill_2 FILLER_51_87 ();
 sg13g2_fill_1 FILLER_51_94 ();
 sg13g2_fill_1 FILLER_51_110 ();
 sg13g2_fill_2 FILLER_51_119 ();
 sg13g2_fill_1 FILLER_51_138 ();
 sg13g2_fill_1 FILLER_51_144 ();
 sg13g2_fill_1 FILLER_51_171 ();
 sg13g2_decap_4 FILLER_51_206 ();
 sg13g2_decap_4 FILLER_51_214 ();
 sg13g2_decap_8 FILLER_51_223 ();
 sg13g2_fill_2 FILLER_51_230 ();
 sg13g2_fill_2 FILLER_51_246 ();
 sg13g2_fill_2 FILLER_51_256 ();
 sg13g2_fill_2 FILLER_51_261 ();
 sg13g2_fill_1 FILLER_51_323 ();
 sg13g2_fill_2 FILLER_51_360 ();
 sg13g2_fill_2 FILLER_51_377 ();
 sg13g2_fill_2 FILLER_51_383 ();
 sg13g2_fill_2 FILLER_51_413 ();
 sg13g2_fill_2 FILLER_51_452 ();
 sg13g2_fill_1 FILLER_51_458 ();
 sg13g2_fill_2 FILLER_51_464 ();
 sg13g2_fill_1 FILLER_51_471 ();
 sg13g2_decap_8 FILLER_51_479 ();
 sg13g2_decap_8 FILLER_51_486 ();
 sg13g2_fill_1 FILLER_51_493 ();
 sg13g2_fill_2 FILLER_51_508 ();
 sg13g2_fill_1 FILLER_51_510 ();
 sg13g2_fill_2 FILLER_51_524 ();
 sg13g2_fill_1 FILLER_51_542 ();
 sg13g2_fill_1 FILLER_51_563 ();
 sg13g2_fill_2 FILLER_51_569 ();
 sg13g2_fill_1 FILLER_51_579 ();
 sg13g2_fill_2 FILLER_51_585 ();
 sg13g2_fill_2 FILLER_51_600 ();
 sg13g2_decap_8 FILLER_51_615 ();
 sg13g2_decap_4 FILLER_51_622 ();
 sg13g2_fill_2 FILLER_51_626 ();
 sg13g2_fill_2 FILLER_51_637 ();
 sg13g2_decap_8 FILLER_51_691 ();
 sg13g2_fill_2 FILLER_51_698 ();
 sg13g2_fill_1 FILLER_51_704 ();
 sg13g2_decap_4 FILLER_51_741 ();
 sg13g2_decap_4 FILLER_51_767 ();
 sg13g2_fill_2 FILLER_51_771 ();
 sg13g2_decap_4 FILLER_51_777 ();
 sg13g2_fill_2 FILLER_51_781 ();
 sg13g2_decap_4 FILLER_51_836 ();
 sg13g2_fill_1 FILLER_51_840 ();
 sg13g2_fill_1 FILLER_51_844 ();
 sg13g2_decap_4 FILLER_51_850 ();
 sg13g2_fill_2 FILLER_51_854 ();
 sg13g2_fill_2 FILLER_51_960 ();
 sg13g2_fill_2 FILLER_51_1024 ();
 sg13g2_fill_2 FILLER_51_1042 ();
 sg13g2_fill_2 FILLER_51_1049 ();
 sg13g2_fill_1 FILLER_51_1066 ();
 sg13g2_fill_1 FILLER_51_1099 ();
 sg13g2_fill_1 FILLER_51_1115 ();
 sg13g2_fill_1 FILLER_51_1120 ();
 sg13g2_fill_1 FILLER_51_1130 ();
 sg13g2_fill_1 FILLER_51_1145 ();
 sg13g2_fill_1 FILLER_51_1151 ();
 sg13g2_decap_8 FILLER_51_1178 ();
 sg13g2_fill_2 FILLER_51_1185 ();
 sg13g2_decap_4 FILLER_51_1206 ();
 sg13g2_decap_4 FILLER_51_1214 ();
 sg13g2_decap_8 FILLER_51_1246 ();
 sg13g2_decap_4 FILLER_51_1253 ();
 sg13g2_fill_2 FILLER_51_1274 ();
 sg13g2_fill_1 FILLER_51_1276 ();
 sg13g2_fill_2 FILLER_51_1281 ();
 sg13g2_fill_1 FILLER_51_1283 ();
 sg13g2_fill_1 FILLER_51_1294 ();
 sg13g2_fill_1 FILLER_51_1300 ();
 sg13g2_fill_2 FILLER_51_1306 ();
 sg13g2_fill_1 FILLER_51_1314 ();
 sg13g2_fill_1 FILLER_51_1320 ();
 sg13g2_decap_4 FILLER_51_1332 ();
 sg13g2_fill_1 FILLER_51_1336 ();
 sg13g2_fill_2 FILLER_51_1342 ();
 sg13g2_fill_1 FILLER_51_1358 ();
 sg13g2_fill_1 FILLER_51_1366 ();
 sg13g2_fill_1 FILLER_51_1398 ();
 sg13g2_decap_8 FILLER_51_1408 ();
 sg13g2_fill_1 FILLER_51_1415 ();
 sg13g2_decap_8 FILLER_51_1429 ();
 sg13g2_fill_1 FILLER_51_1436 ();
 sg13g2_fill_2 FILLER_51_1449 ();
 sg13g2_fill_2 FILLER_51_1456 ();
 sg13g2_fill_1 FILLER_51_1458 ();
 sg13g2_fill_2 FILLER_51_1475 ();
 sg13g2_fill_1 FILLER_51_1477 ();
 sg13g2_fill_1 FILLER_51_1490 ();
 sg13g2_fill_2 FILLER_51_1506 ();
 sg13g2_fill_1 FILLER_51_1523 ();
 sg13g2_fill_2 FILLER_51_1553 ();
 sg13g2_fill_2 FILLER_51_1563 ();
 sg13g2_fill_2 FILLER_51_1570 ();
 sg13g2_fill_1 FILLER_51_1572 ();
 sg13g2_fill_2 FILLER_51_1587 ();
 sg13g2_fill_2 FILLER_51_1596 ();
 sg13g2_fill_1 FILLER_51_1606 ();
 sg13g2_fill_2 FILLER_51_1612 ();
 sg13g2_fill_1 FILLER_51_1614 ();
 sg13g2_decap_4 FILLER_51_1619 ();
 sg13g2_fill_2 FILLER_51_1623 ();
 sg13g2_decap_4 FILLER_51_1724 ();
 sg13g2_decap_8 FILLER_51_1751 ();
 sg13g2_fill_2 FILLER_51_1758 ();
 sg13g2_decap_8 FILLER_51_1774 ();
 sg13g2_decap_8 FILLER_51_1781 ();
 sg13g2_decap_4 FILLER_51_1788 ();
 sg13g2_fill_2 FILLER_51_1792 ();
 sg13g2_fill_2 FILLER_51_1817 ();
 sg13g2_decap_8 FILLER_51_1827 ();
 sg13g2_decap_8 FILLER_51_1834 ();
 sg13g2_decap_8 FILLER_51_1845 ();
 sg13g2_decap_8 FILLER_51_1852 ();
 sg13g2_decap_4 FILLER_51_1859 ();
 sg13g2_fill_2 FILLER_51_1863 ();
 sg13g2_decap_8 FILLER_51_1895 ();
 sg13g2_decap_8 FILLER_51_1902 ();
 sg13g2_fill_2 FILLER_51_1909 ();
 sg13g2_fill_1 FILLER_51_1911 ();
 sg13g2_decap_8 FILLER_51_1917 ();
 sg13g2_decap_4 FILLER_51_1924 ();
 sg13g2_fill_2 FILLER_51_1928 ();
 sg13g2_decap_8 FILLER_51_1943 ();
 sg13g2_decap_8 FILLER_51_1950 ();
 sg13g2_decap_4 FILLER_51_1957 ();
 sg13g2_fill_1 FILLER_51_1961 ();
 sg13g2_decap_8 FILLER_51_1979 ();
 sg13g2_fill_2 FILLER_51_1986 ();
 sg13g2_decap_4 FILLER_51_2027 ();
 sg13g2_fill_1 FILLER_51_2031 ();
 sg13g2_fill_1 FILLER_51_2037 ();
 sg13g2_decap_8 FILLER_51_2042 ();
 sg13g2_fill_2 FILLER_51_2049 ();
 sg13g2_fill_1 FILLER_51_2051 ();
 sg13g2_fill_2 FILLER_51_2127 ();
 sg13g2_fill_1 FILLER_51_2143 ();
 sg13g2_fill_1 FILLER_51_2219 ();
 sg13g2_fill_1 FILLER_51_2275 ();
 sg13g2_fill_2 FILLER_51_2283 ();
 sg13g2_fill_1 FILLER_51_2291 ();
 sg13g2_decap_8 FILLER_51_2306 ();
 sg13g2_decap_8 FILLER_51_2313 ();
 sg13g2_decap_4 FILLER_51_2328 ();
 sg13g2_fill_2 FILLER_51_2338 ();
 sg13g2_fill_1 FILLER_51_2340 ();
 sg13g2_decap_4 FILLER_51_2351 ();
 sg13g2_fill_2 FILLER_51_2355 ();
 sg13g2_fill_2 FILLER_51_2361 ();
 sg13g2_fill_1 FILLER_51_2363 ();
 sg13g2_fill_2 FILLER_51_2373 ();
 sg13g2_decap_4 FILLER_51_2406 ();
 sg13g2_fill_1 FILLER_51_2410 ();
 sg13g2_fill_1 FILLER_51_2421 ();
 sg13g2_fill_1 FILLER_51_2428 ();
 sg13g2_fill_1 FILLER_51_2455 ();
 sg13g2_fill_2 FILLER_51_2499 ();
 sg13g2_fill_1 FILLER_51_2527 ();
 sg13g2_decap_8 FILLER_51_2564 ();
 sg13g2_decap_8 FILLER_51_2571 ();
 sg13g2_decap_8 FILLER_51_2578 ();
 sg13g2_decap_8 FILLER_51_2585 ();
 sg13g2_decap_8 FILLER_51_2592 ();
 sg13g2_decap_8 FILLER_51_2599 ();
 sg13g2_decap_8 FILLER_51_2606 ();
 sg13g2_decap_8 FILLER_51_2613 ();
 sg13g2_decap_8 FILLER_51_2620 ();
 sg13g2_decap_8 FILLER_51_2627 ();
 sg13g2_decap_8 FILLER_51_2634 ();
 sg13g2_decap_8 FILLER_51_2641 ();
 sg13g2_decap_8 FILLER_51_2648 ();
 sg13g2_decap_8 FILLER_51_2655 ();
 sg13g2_decap_8 FILLER_51_2662 ();
 sg13g2_fill_1 FILLER_51_2669 ();
 sg13g2_decap_4 FILLER_52_0 ();
 sg13g2_fill_2 FILLER_52_17 ();
 sg13g2_fill_2 FILLER_52_24 ();
 sg13g2_fill_1 FILLER_52_26 ();
 sg13g2_fill_1 FILLER_52_34 ();
 sg13g2_fill_2 FILLER_52_39 ();
 sg13g2_fill_1 FILLER_52_41 ();
 sg13g2_fill_2 FILLER_52_47 ();
 sg13g2_fill_1 FILLER_52_49 ();
 sg13g2_fill_2 FILLER_52_63 ();
 sg13g2_fill_1 FILLER_52_65 ();
 sg13g2_fill_1 FILLER_52_71 ();
 sg13g2_fill_1 FILLER_52_85 ();
 sg13g2_fill_2 FILLER_52_100 ();
 sg13g2_fill_1 FILLER_52_102 ();
 sg13g2_fill_2 FILLER_52_136 ();
 sg13g2_decap_4 FILLER_52_143 ();
 sg13g2_fill_1 FILLER_52_147 ();
 sg13g2_decap_8 FILLER_52_156 ();
 sg13g2_decap_4 FILLER_52_163 ();
 sg13g2_fill_2 FILLER_52_167 ();
 sg13g2_decap_8 FILLER_52_174 ();
 sg13g2_fill_2 FILLER_52_181 ();
 sg13g2_fill_1 FILLER_52_183 ();
 sg13g2_decap_8 FILLER_52_188 ();
 sg13g2_decap_4 FILLER_52_195 ();
 sg13g2_fill_1 FILLER_52_199 ();
 sg13g2_fill_2 FILLER_52_260 ();
 sg13g2_fill_1 FILLER_52_291 ();
 sg13g2_fill_2 FILLER_52_299 ();
 sg13g2_fill_2 FILLER_52_310 ();
 sg13g2_fill_1 FILLER_52_328 ();
 sg13g2_fill_2 FILLER_52_342 ();
 sg13g2_fill_1 FILLER_52_372 ();
 sg13g2_fill_2 FILLER_52_378 ();
 sg13g2_fill_2 FILLER_52_391 ();
 sg13g2_fill_1 FILLER_52_397 ();
 sg13g2_fill_2 FILLER_52_425 ();
 sg13g2_fill_2 FILLER_52_474 ();
 sg13g2_fill_2 FILLER_52_483 ();
 sg13g2_fill_1 FILLER_52_485 ();
 sg13g2_fill_2 FILLER_52_502 ();
 sg13g2_fill_1 FILLER_52_512 ();
 sg13g2_fill_1 FILLER_52_534 ();
 sg13g2_fill_2 FILLER_52_550 ();
 sg13g2_fill_1 FILLER_52_564 ();
 sg13g2_fill_1 FILLER_52_570 ();
 sg13g2_fill_1 FILLER_52_575 ();
 sg13g2_decap_4 FILLER_52_585 ();
 sg13g2_fill_2 FILLER_52_615 ();
 sg13g2_fill_2 FILLER_52_622 ();
 sg13g2_fill_1 FILLER_52_674 ();
 sg13g2_decap_8 FILLER_52_679 ();
 sg13g2_decap_8 FILLER_52_686 ();
 sg13g2_decap_4 FILLER_52_693 ();
 sg13g2_fill_1 FILLER_52_706 ();
 sg13g2_fill_1 FILLER_52_715 ();
 sg13g2_fill_1 FILLER_52_731 ();
 sg13g2_fill_1 FILLER_52_736 ();
 sg13g2_decap_8 FILLER_52_774 ();
 sg13g2_fill_1 FILLER_52_848 ();
 sg13g2_fill_2 FILLER_52_879 ();
 sg13g2_fill_1 FILLER_52_881 ();
 sg13g2_fill_1 FILLER_52_910 ();
 sg13g2_fill_1 FILLER_52_1021 ();
 sg13g2_fill_1 FILLER_52_1095 ();
 sg13g2_fill_1 FILLER_52_1101 ();
 sg13g2_fill_2 FILLER_52_1107 ();
 sg13g2_decap_8 FILLER_52_1190 ();
 sg13g2_fill_2 FILLER_52_1197 ();
 sg13g2_decap_8 FILLER_52_1214 ();
 sg13g2_fill_2 FILLER_52_1221 ();
 sg13g2_fill_2 FILLER_52_1229 ();
 sg13g2_fill_1 FILLER_52_1231 ();
 sg13g2_fill_2 FILLER_52_1246 ();
 sg13g2_fill_1 FILLER_52_1265 ();
 sg13g2_fill_1 FILLER_52_1275 ();
 sg13g2_fill_2 FILLER_52_1280 ();
 sg13g2_decap_8 FILLER_52_1320 ();
 sg13g2_decap_4 FILLER_52_1331 ();
 sg13g2_fill_2 FILLER_52_1335 ();
 sg13g2_fill_2 FILLER_52_1355 ();
 sg13g2_fill_2 FILLER_52_1361 ();
 sg13g2_fill_1 FILLER_52_1368 ();
 sg13g2_fill_1 FILLER_52_1377 ();
 sg13g2_fill_1 FILLER_52_1386 ();
 sg13g2_decap_8 FILLER_52_1391 ();
 sg13g2_decap_4 FILLER_52_1398 ();
 sg13g2_fill_1 FILLER_52_1402 ();
 sg13g2_fill_1 FILLER_52_1417 ();
 sg13g2_fill_1 FILLER_52_1427 ();
 sg13g2_fill_1 FILLER_52_1454 ();
 sg13g2_fill_1 FILLER_52_1459 ();
 sg13g2_fill_1 FILLER_52_1464 ();
 sg13g2_fill_2 FILLER_52_1470 ();
 sg13g2_fill_1 FILLER_52_1472 ();
 sg13g2_decap_4 FILLER_52_1545 ();
 sg13g2_decap_4 FILLER_52_1565 ();
 sg13g2_fill_1 FILLER_52_1569 ();
 sg13g2_fill_2 FILLER_52_1574 ();
 sg13g2_fill_1 FILLER_52_1586 ();
 sg13g2_decap_4 FILLER_52_1596 ();
 sg13g2_decap_8 FILLER_52_1610 ();
 sg13g2_decap_8 FILLER_52_1617 ();
 sg13g2_decap_8 FILLER_52_1624 ();
 sg13g2_decap_4 FILLER_52_1631 ();
 sg13g2_fill_2 FILLER_52_1635 ();
 sg13g2_decap_8 FILLER_52_1641 ();
 sg13g2_fill_2 FILLER_52_1648 ();
 sg13g2_fill_1 FILLER_52_1660 ();
 sg13g2_fill_2 FILLER_52_1665 ();
 sg13g2_fill_1 FILLER_52_1667 ();
 sg13g2_fill_2 FILLER_52_1672 ();
 sg13g2_fill_1 FILLER_52_1674 ();
 sg13g2_decap_8 FILLER_52_1680 ();
 sg13g2_fill_2 FILLER_52_1687 ();
 sg13g2_decap_4 FILLER_52_1693 ();
 sg13g2_fill_1 FILLER_52_1697 ();
 sg13g2_decap_8 FILLER_52_1716 ();
 sg13g2_decap_4 FILLER_52_1723 ();
 sg13g2_fill_1 FILLER_52_1727 ();
 sg13g2_fill_2 FILLER_52_1734 ();
 sg13g2_fill_1 FILLER_52_1736 ();
 sg13g2_fill_2 FILLER_52_1742 ();
 sg13g2_fill_1 FILLER_52_1744 ();
 sg13g2_decap_4 FILLER_52_1770 ();
 sg13g2_decap_8 FILLER_52_1779 ();
 sg13g2_decap_8 FILLER_52_1786 ();
 sg13g2_decap_8 FILLER_52_1793 ();
 sg13g2_decap_8 FILLER_52_1800 ();
 sg13g2_decap_8 FILLER_52_1807 ();
 sg13g2_decap_8 FILLER_52_1814 ();
 sg13g2_fill_2 FILLER_52_1821 ();
 sg13g2_fill_1 FILLER_52_1823 ();
 sg13g2_fill_1 FILLER_52_1864 ();
 sg13g2_fill_1 FILLER_52_1921 ();
 sg13g2_fill_1 FILLER_52_1952 ();
 sg13g2_decap_8 FILLER_52_1979 ();
 sg13g2_fill_2 FILLER_52_2001 ();
 sg13g2_fill_2 FILLER_52_2008 ();
 sg13g2_fill_2 FILLER_52_2014 ();
 sg13g2_decap_8 FILLER_52_2020 ();
 sg13g2_decap_8 FILLER_52_2027 ();
 sg13g2_decap_8 FILLER_52_2034 ();
 sg13g2_fill_1 FILLER_52_2041 ();
 sg13g2_fill_1 FILLER_52_2125 ();
 sg13g2_fill_1 FILLER_52_2152 ();
 sg13g2_fill_1 FILLER_52_2163 ();
 sg13g2_fill_2 FILLER_52_2190 ();
 sg13g2_fill_1 FILLER_52_2211 ();
 sg13g2_decap_4 FILLER_52_2284 ();
 sg13g2_fill_2 FILLER_52_2288 ();
 sg13g2_fill_1 FILLER_52_2326 ();
 sg13g2_fill_2 FILLER_52_2331 ();
 sg13g2_fill_1 FILLER_52_2333 ();
 sg13g2_fill_1 FILLER_52_2360 ();
 sg13g2_fill_2 FILLER_52_2378 ();
 sg13g2_decap_4 FILLER_52_2384 ();
 sg13g2_decap_4 FILLER_52_2394 ();
 sg13g2_fill_2 FILLER_52_2404 ();
 sg13g2_fill_1 FILLER_52_2406 ();
 sg13g2_fill_2 FILLER_52_2443 ();
 sg13g2_fill_1 FILLER_52_2461 ();
 sg13g2_fill_2 FILLER_52_2526 ();
 sg13g2_fill_1 FILLER_52_2541 ();
 sg13g2_decap_8 FILLER_52_2550 ();
 sg13g2_decap_8 FILLER_52_2561 ();
 sg13g2_decap_8 FILLER_52_2568 ();
 sg13g2_decap_8 FILLER_52_2575 ();
 sg13g2_decap_8 FILLER_52_2582 ();
 sg13g2_decap_8 FILLER_52_2589 ();
 sg13g2_decap_8 FILLER_52_2596 ();
 sg13g2_decap_8 FILLER_52_2603 ();
 sg13g2_decap_8 FILLER_52_2610 ();
 sg13g2_decap_8 FILLER_52_2617 ();
 sg13g2_decap_8 FILLER_52_2624 ();
 sg13g2_decap_8 FILLER_52_2631 ();
 sg13g2_decap_8 FILLER_52_2638 ();
 sg13g2_decap_8 FILLER_52_2645 ();
 sg13g2_decap_8 FILLER_52_2652 ();
 sg13g2_decap_8 FILLER_52_2659 ();
 sg13g2_decap_4 FILLER_52_2666 ();
 sg13g2_decap_4 FILLER_53_0 ();
 sg13g2_fill_1 FILLER_53_101 ();
 sg13g2_fill_1 FILLER_53_106 ();
 sg13g2_fill_2 FILLER_53_111 ();
 sg13g2_fill_1 FILLER_53_117 ();
 sg13g2_fill_2 FILLER_53_121 ();
 sg13g2_fill_1 FILLER_53_123 ();
 sg13g2_decap_8 FILLER_53_130 ();
 sg13g2_decap_4 FILLER_53_137 ();
 sg13g2_decap_4 FILLER_53_146 ();
 sg13g2_fill_2 FILLER_53_150 ();
 sg13g2_fill_1 FILLER_53_160 ();
 sg13g2_fill_1 FILLER_53_172 ();
 sg13g2_decap_4 FILLER_53_178 ();
 sg13g2_fill_1 FILLER_53_182 ();
 sg13g2_fill_2 FILLER_53_202 ();
 sg13g2_decap_8 FILLER_53_208 ();
 sg13g2_decap_4 FILLER_53_219 ();
 sg13g2_fill_1 FILLER_53_233 ();
 sg13g2_fill_1 FILLER_53_239 ();
 sg13g2_fill_2 FILLER_53_266 ();
 sg13g2_fill_2 FILLER_53_311 ();
 sg13g2_fill_2 FILLER_53_335 ();
 sg13g2_fill_1 FILLER_53_348 ();
 sg13g2_fill_2 FILLER_53_372 ();
 sg13g2_fill_2 FILLER_53_388 ();
 sg13g2_fill_1 FILLER_53_395 ();
 sg13g2_fill_1 FILLER_53_400 ();
 sg13g2_fill_1 FILLER_53_453 ();
 sg13g2_fill_2 FILLER_53_464 ();
 sg13g2_fill_1 FILLER_53_496 ();
 sg13g2_fill_1 FILLER_53_502 ();
 sg13g2_fill_2 FILLER_53_544 ();
 sg13g2_decap_8 FILLER_53_609 ();
 sg13g2_fill_2 FILLER_53_616 ();
 sg13g2_fill_2 FILLER_53_662 ();
 sg13g2_fill_1 FILLER_53_664 ();
 sg13g2_decap_8 FILLER_53_684 ();
 sg13g2_fill_2 FILLER_53_691 ();
 sg13g2_fill_1 FILLER_53_693 ();
 sg13g2_fill_2 FILLER_53_700 ();
 sg13g2_decap_8 FILLER_53_712 ();
 sg13g2_decap_8 FILLER_53_719 ();
 sg13g2_decap_4 FILLER_53_726 ();
 sg13g2_decap_4 FILLER_53_735 ();
 sg13g2_decap_8 FILLER_53_779 ();
 sg13g2_decap_4 FILLER_53_786 ();
 sg13g2_fill_1 FILLER_53_790 ();
 sg13g2_decap_4 FILLER_53_830 ();
 sg13g2_fill_2 FILLER_53_834 ();
 sg13g2_decap_8 FILLER_53_841 ();
 sg13g2_decap_8 FILLER_53_848 ();
 sg13g2_fill_2 FILLER_53_855 ();
 sg13g2_fill_2 FILLER_53_877 ();
 sg13g2_fill_2 FILLER_53_891 ();
 sg13g2_fill_1 FILLER_53_916 ();
 sg13g2_fill_2 FILLER_53_961 ();
 sg13g2_fill_1 FILLER_53_979 ();
 sg13g2_fill_1 FILLER_53_1002 ();
 sg13g2_fill_2 FILLER_53_1041 ();
 sg13g2_fill_1 FILLER_53_1047 ();
 sg13g2_fill_2 FILLER_53_1065 ();
 sg13g2_fill_1 FILLER_53_1082 ();
 sg13g2_fill_2 FILLER_53_1096 ();
 sg13g2_decap_4 FILLER_53_1149 ();
 sg13g2_fill_1 FILLER_53_1153 ();
 sg13g2_decap_8 FILLER_53_1159 ();
 sg13g2_fill_1 FILLER_53_1166 ();
 sg13g2_fill_2 FILLER_53_1179 ();
 sg13g2_decap_4 FILLER_53_1195 ();
 sg13g2_fill_1 FILLER_53_1203 ();
 sg13g2_fill_1 FILLER_53_1222 ();
 sg13g2_fill_2 FILLER_53_1284 ();
 sg13g2_fill_2 FILLER_53_1298 ();
 sg13g2_fill_1 FILLER_53_1300 ();
 sg13g2_decap_8 FILLER_53_1315 ();
 sg13g2_fill_1 FILLER_53_1322 ();
 sg13g2_fill_1 FILLER_53_1335 ();
 sg13g2_fill_1 FILLER_53_1341 ();
 sg13g2_fill_2 FILLER_53_1355 ();
 sg13g2_fill_1 FILLER_53_1357 ();
 sg13g2_fill_1 FILLER_53_1381 ();
 sg13g2_fill_1 FILLER_53_1386 ();
 sg13g2_fill_1 FILLER_53_1413 ();
 sg13g2_fill_1 FILLER_53_1440 ();
 sg13g2_decap_4 FILLER_53_1445 ();
 sg13g2_fill_2 FILLER_53_1449 ();
 sg13g2_fill_2 FILLER_53_1456 ();
 sg13g2_fill_1 FILLER_53_1500 ();
 sg13g2_fill_1 FILLER_53_1522 ();
 sg13g2_fill_1 FILLER_53_1526 ();
 sg13g2_fill_1 FILLER_53_1532 ();
 sg13g2_fill_1 FILLER_53_1538 ();
 sg13g2_fill_2 FILLER_53_1544 ();
 sg13g2_decap_8 FILLER_53_1577 ();
 sg13g2_fill_1 FILLER_53_1584 ();
 sg13g2_fill_2 FILLER_53_1590 ();
 sg13g2_fill_1 FILLER_53_1592 ();
 sg13g2_decap_8 FILLER_53_1619 ();
 sg13g2_decap_8 FILLER_53_1626 ();
 sg13g2_decap_8 FILLER_53_1633 ();
 sg13g2_decap_4 FILLER_53_1640 ();
 sg13g2_fill_1 FILLER_53_1644 ();
 sg13g2_fill_2 FILLER_53_1653 ();
 sg13g2_fill_1 FILLER_53_1655 ();
 sg13g2_decap_8 FILLER_53_1673 ();
 sg13g2_decap_4 FILLER_53_1680 ();
 sg13g2_fill_1 FILLER_53_1684 ();
 sg13g2_decap_8 FILLER_53_1690 ();
 sg13g2_fill_1 FILLER_53_1706 ();
 sg13g2_decap_4 FILLER_53_1712 ();
 sg13g2_decap_8 FILLER_53_1725 ();
 sg13g2_fill_1 FILLER_53_1737 ();
 sg13g2_fill_2 FILLER_53_1743 ();
 sg13g2_fill_1 FILLER_53_1750 ();
 sg13g2_fill_2 FILLER_53_1756 ();
 sg13g2_fill_1 FILLER_53_1779 ();
 sg13g2_fill_1 FILLER_53_1800 ();
 sg13g2_decap_8 FILLER_53_1862 ();
 sg13g2_fill_1 FILLER_53_1869 ();
 sg13g2_fill_2 FILLER_53_1887 ();
 sg13g2_fill_1 FILLER_53_1889 ();
 sg13g2_fill_1 FILLER_53_1895 ();
 sg13g2_fill_1 FILLER_53_1906 ();
 sg13g2_fill_2 FILLER_53_1933 ();
 sg13g2_fill_1 FILLER_53_1940 ();
 sg13g2_decap_8 FILLER_53_1970 ();
 sg13g2_fill_1 FILLER_53_1977 ();
 sg13g2_fill_1 FILLER_53_1982 ();
 sg13g2_fill_1 FILLER_53_2023 ();
 sg13g2_fill_1 FILLER_53_2054 ();
 sg13g2_fill_2 FILLER_53_2092 ();
 sg13g2_fill_1 FILLER_53_2125 ();
 sg13g2_fill_1 FILLER_53_2136 ();
 sg13g2_fill_1 FILLER_53_2141 ();
 sg13g2_fill_1 FILLER_53_2147 ();
 sg13g2_fill_1 FILLER_53_2158 ();
 sg13g2_fill_1 FILLER_53_2173 ();
 sg13g2_fill_1 FILLER_53_2179 ();
 sg13g2_fill_2 FILLER_53_2247 ();
 sg13g2_fill_1 FILLER_53_2255 ();
 sg13g2_fill_1 FILLER_53_2264 ();
 sg13g2_decap_8 FILLER_53_2286 ();
 sg13g2_fill_2 FILLER_53_2293 ();
 sg13g2_fill_2 FILLER_53_2299 ();
 sg13g2_fill_1 FILLER_53_2301 ();
 sg13g2_fill_1 FILLER_53_2308 ();
 sg13g2_fill_2 FILLER_53_2319 ();
 sg13g2_fill_1 FILLER_53_2321 ();
 sg13g2_decap_8 FILLER_53_2336 ();
 sg13g2_decap_4 FILLER_53_2347 ();
 sg13g2_decap_8 FILLER_53_2381 ();
 sg13g2_decap_4 FILLER_53_2388 ();
 sg13g2_fill_1 FILLER_53_2392 ();
 sg13g2_fill_1 FILLER_53_2435 ();
 sg13g2_fill_1 FILLER_53_2516 ();
 sg13g2_decap_4 FILLER_53_2530 ();
 sg13g2_fill_2 FILLER_53_2534 ();
 sg13g2_decap_8 FILLER_53_2572 ();
 sg13g2_decap_8 FILLER_53_2579 ();
 sg13g2_decap_8 FILLER_53_2586 ();
 sg13g2_decap_8 FILLER_53_2593 ();
 sg13g2_decap_8 FILLER_53_2600 ();
 sg13g2_decap_8 FILLER_53_2607 ();
 sg13g2_decap_8 FILLER_53_2614 ();
 sg13g2_decap_8 FILLER_53_2621 ();
 sg13g2_decap_8 FILLER_53_2628 ();
 sg13g2_decap_8 FILLER_53_2635 ();
 sg13g2_decap_8 FILLER_53_2642 ();
 sg13g2_decap_8 FILLER_53_2649 ();
 sg13g2_decap_8 FILLER_53_2656 ();
 sg13g2_decap_8 FILLER_53_2663 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_7 ();
 sg13g2_fill_1 FILLER_54_9 ();
 sg13g2_decap_4 FILLER_54_14 ();
 sg13g2_fill_1 FILLER_54_27 ();
 sg13g2_fill_1 FILLER_54_33 ();
 sg13g2_fill_1 FILLER_54_38 ();
 sg13g2_fill_1 FILLER_54_44 ();
 sg13g2_fill_2 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_fill_1 FILLER_54_63 ();
 sg13g2_fill_1 FILLER_54_72 ();
 sg13g2_fill_2 FILLER_54_77 ();
 sg13g2_fill_2 FILLER_54_84 ();
 sg13g2_fill_1 FILLER_54_86 ();
 sg13g2_fill_2 FILLER_54_91 ();
 sg13g2_fill_1 FILLER_54_93 ();
 sg13g2_decap_4 FILLER_54_111 ();
 sg13g2_fill_2 FILLER_54_115 ();
 sg13g2_decap_8 FILLER_54_122 ();
 sg13g2_fill_1 FILLER_54_129 ();
 sg13g2_fill_2 FILLER_54_140 ();
 sg13g2_fill_2 FILLER_54_168 ();
 sg13g2_fill_1 FILLER_54_170 ();
 sg13g2_fill_1 FILLER_54_197 ();
 sg13g2_decap_8 FILLER_54_203 ();
 sg13g2_fill_2 FILLER_54_256 ();
 sg13g2_fill_1 FILLER_54_293 ();
 sg13g2_fill_1 FILLER_54_380 ();
 sg13g2_fill_1 FILLER_54_396 ();
 sg13g2_fill_1 FILLER_54_402 ();
 sg13g2_fill_1 FILLER_54_408 ();
 sg13g2_fill_2 FILLER_54_433 ();
 sg13g2_fill_2 FILLER_54_474 ();
 sg13g2_fill_1 FILLER_54_476 ();
 sg13g2_fill_1 FILLER_54_508 ();
 sg13g2_decap_8 FILLER_54_513 ();
 sg13g2_decap_8 FILLER_54_520 ();
 sg13g2_decap_8 FILLER_54_527 ();
 sg13g2_decap_4 FILLER_54_539 ();
 sg13g2_fill_1 FILLER_54_543 ();
 sg13g2_fill_2 FILLER_54_549 ();
 sg13g2_fill_1 FILLER_54_555 ();
 sg13g2_fill_1 FILLER_54_566 ();
 sg13g2_fill_1 FILLER_54_595 ();
 sg13g2_decap_8 FILLER_54_604 ();
 sg13g2_decap_8 FILLER_54_611 ();
 sg13g2_decap_4 FILLER_54_618 ();
 sg13g2_fill_1 FILLER_54_646 ();
 sg13g2_fill_1 FILLER_54_703 ();
 sg13g2_decap_4 FILLER_54_730 ();
 sg13g2_fill_1 FILLER_54_739 ();
 sg13g2_fill_1 FILLER_54_744 ();
 sg13g2_fill_2 FILLER_54_776 ();
 sg13g2_fill_1 FILLER_54_778 ();
 sg13g2_decap_8 FILLER_54_784 ();
 sg13g2_fill_2 FILLER_54_791 ();
 sg13g2_fill_1 FILLER_54_793 ();
 sg13g2_decap_4 FILLER_54_800 ();
 sg13g2_decap_4 FILLER_54_836 ();
 sg13g2_fill_1 FILLER_54_876 ();
 sg13g2_fill_1 FILLER_54_934 ();
 sg13g2_decap_4 FILLER_54_939 ();
 sg13g2_fill_2 FILLER_54_943 ();
 sg13g2_fill_2 FILLER_54_985 ();
 sg13g2_fill_1 FILLER_54_1003 ();
 sg13g2_fill_1 FILLER_54_1010 ();
 sg13g2_fill_1 FILLER_54_1030 ();
 sg13g2_fill_2 FILLER_54_1077 ();
 sg13g2_fill_1 FILLER_54_1083 ();
 sg13g2_fill_2 FILLER_54_1087 ();
 sg13g2_fill_2 FILLER_54_1109 ();
 sg13g2_fill_1 FILLER_54_1116 ();
 sg13g2_fill_1 FILLER_54_1121 ();
 sg13g2_fill_1 FILLER_54_1126 ();
 sg13g2_decap_4 FILLER_54_1144 ();
 sg13g2_decap_8 FILLER_54_1152 ();
 sg13g2_decap_8 FILLER_54_1159 ();
 sg13g2_decap_8 FILLER_54_1166 ();
 sg13g2_fill_2 FILLER_54_1173 ();
 sg13g2_fill_1 FILLER_54_1175 ();
 sg13g2_fill_1 FILLER_54_1181 ();
 sg13g2_fill_1 FILLER_54_1186 ();
 sg13g2_fill_1 FILLER_54_1190 ();
 sg13g2_fill_1 FILLER_54_1211 ();
 sg13g2_fill_1 FILLER_54_1217 ();
 sg13g2_fill_1 FILLER_54_1263 ();
 sg13g2_fill_2 FILLER_54_1273 ();
 sg13g2_decap_8 FILLER_54_1283 ();
 sg13g2_fill_2 FILLER_54_1290 ();
 sg13g2_decap_4 FILLER_54_1304 ();
 sg13g2_fill_2 FILLER_54_1308 ();
 sg13g2_decap_8 FILLER_54_1314 ();
 sg13g2_decap_8 FILLER_54_1321 ();
 sg13g2_decap_8 FILLER_54_1328 ();
 sg13g2_decap_8 FILLER_54_1335 ();
 sg13g2_decap_8 FILLER_54_1342 ();
 sg13g2_decap_8 FILLER_54_1349 ();
 sg13g2_decap_8 FILLER_54_1356 ();
 sg13g2_fill_1 FILLER_54_1363 ();
 sg13g2_fill_2 FILLER_54_1373 ();
 sg13g2_decap_8 FILLER_54_1384 ();
 sg13g2_fill_2 FILLER_54_1391 ();
 sg13g2_fill_1 FILLER_54_1393 ();
 sg13g2_fill_1 FILLER_54_1398 ();
 sg13g2_fill_2 FILLER_54_1445 ();
 sg13g2_decap_4 FILLER_54_1452 ();
 sg13g2_fill_1 FILLER_54_1473 ();
 sg13g2_fill_2 FILLER_54_1484 ();
 sg13g2_fill_1 FILLER_54_1486 ();
 sg13g2_decap_4 FILLER_54_1492 ();
 sg13g2_decap_8 FILLER_54_1539 ();
 sg13g2_fill_1 FILLER_54_1546 ();
 sg13g2_decap_8 FILLER_54_1590 ();
 sg13g2_fill_2 FILLER_54_1597 ();
 sg13g2_fill_2 FILLER_54_1603 ();
 sg13g2_decap_4 FILLER_54_1609 ();
 sg13g2_decap_8 FILLER_54_1623 ();
 sg13g2_decap_4 FILLER_54_1630 ();
 sg13g2_fill_1 FILLER_54_1634 ();
 sg13g2_fill_2 FILLER_54_1655 ();
 sg13g2_decap_4 FILLER_54_1687 ();
 sg13g2_fill_2 FILLER_54_1691 ();
 sg13g2_fill_1 FILLER_54_1722 ();
 sg13g2_fill_1 FILLER_54_1728 ();
 sg13g2_fill_1 FILLER_54_1734 ();
 sg13g2_fill_1 FILLER_54_1740 ();
 sg13g2_fill_1 FILLER_54_1779 ();
 sg13g2_fill_2 FILLER_54_1789 ();
 sg13g2_decap_8 FILLER_54_1834 ();
 sg13g2_decap_4 FILLER_54_1841 ();
 sg13g2_decap_8 FILLER_54_1858 ();
 sg13g2_decap_8 FILLER_54_1865 ();
 sg13g2_decap_4 FILLER_54_1872 ();
 sg13g2_fill_1 FILLER_54_1876 ();
 sg13g2_decap_4 FILLER_54_1882 ();
 sg13g2_decap_4 FILLER_54_1895 ();
 sg13g2_decap_4 FILLER_54_1903 ();
 sg13g2_fill_2 FILLER_54_1913 ();
 sg13g2_fill_2 FILLER_54_1919 ();
 sg13g2_fill_1 FILLER_54_1960 ();
 sg13g2_fill_1 FILLER_54_1991 ();
 sg13g2_fill_2 FILLER_54_2018 ();
 sg13g2_fill_1 FILLER_54_2020 ();
 sg13g2_decap_8 FILLER_54_2051 ();
 sg13g2_fill_2 FILLER_54_2058 ();
 sg13g2_fill_1 FILLER_54_2060 ();
 sg13g2_decap_8 FILLER_54_2073 ();
 sg13g2_fill_1 FILLER_54_2080 ();
 sg13g2_decap_8 FILLER_54_2086 ();
 sg13g2_decap_4 FILLER_54_2093 ();
 sg13g2_fill_2 FILLER_54_2097 ();
 sg13g2_fill_2 FILLER_54_2141 ();
 sg13g2_fill_1 FILLER_54_2162 ();
 sg13g2_fill_2 FILLER_54_2178 ();
 sg13g2_decap_8 FILLER_54_2297 ();
 sg13g2_decap_4 FILLER_54_2304 ();
 sg13g2_fill_1 FILLER_54_2308 ();
 sg13g2_fill_2 FILLER_54_2319 ();
 sg13g2_fill_2 FILLER_54_2372 ();
 sg13g2_fill_1 FILLER_54_2374 ();
 sg13g2_fill_1 FILLER_54_2420 ();
 sg13g2_fill_2 FILLER_54_2425 ();
 sg13g2_fill_2 FILLER_54_2437 ();
 sg13g2_fill_2 FILLER_54_2465 ();
 sg13g2_fill_1 FILLER_54_2467 ();
 sg13g2_fill_2 FILLER_54_2474 ();
 sg13g2_fill_2 FILLER_54_2484 ();
 sg13g2_fill_1 FILLER_54_2499 ();
 sg13g2_fill_1 FILLER_54_2504 ();
 sg13g2_fill_1 FILLER_54_2531 ();
 sg13g2_fill_2 FILLER_54_2571 ();
 sg13g2_fill_1 FILLER_54_2573 ();
 sg13g2_decap_8 FILLER_54_2578 ();
 sg13g2_decap_8 FILLER_54_2585 ();
 sg13g2_decap_8 FILLER_54_2592 ();
 sg13g2_decap_8 FILLER_54_2599 ();
 sg13g2_decap_8 FILLER_54_2606 ();
 sg13g2_decap_8 FILLER_54_2613 ();
 sg13g2_decap_8 FILLER_54_2620 ();
 sg13g2_decap_8 FILLER_54_2627 ();
 sg13g2_decap_8 FILLER_54_2634 ();
 sg13g2_decap_8 FILLER_54_2641 ();
 sg13g2_decap_8 FILLER_54_2648 ();
 sg13g2_decap_8 FILLER_54_2655 ();
 sg13g2_decap_8 FILLER_54_2662 ();
 sg13g2_fill_1 FILLER_54_2669 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_7 ();
 sg13g2_fill_1 FILLER_55_51 ();
 sg13g2_decap_8 FILLER_55_61 ();
 sg13g2_decap_8 FILLER_55_68 ();
 sg13g2_fill_2 FILLER_55_75 ();
 sg13g2_fill_2 FILLER_55_84 ();
 sg13g2_decap_8 FILLER_55_103 ();
 sg13g2_decap_8 FILLER_55_110 ();
 sg13g2_decap_8 FILLER_55_117 ();
 sg13g2_decap_8 FILLER_55_124 ();
 sg13g2_decap_4 FILLER_55_155 ();
 sg13g2_fill_1 FILLER_55_169 ();
 sg13g2_fill_2 FILLER_55_175 ();
 sg13g2_fill_2 FILLER_55_181 ();
 sg13g2_fill_2 FILLER_55_213 ();
 sg13g2_fill_1 FILLER_55_215 ();
 sg13g2_decap_4 FILLER_55_220 ();
 sg13g2_fill_2 FILLER_55_224 ();
 sg13g2_fill_2 FILLER_55_271 ();
 sg13g2_fill_1 FILLER_55_273 ();
 sg13g2_fill_1 FILLER_55_281 ();
 sg13g2_fill_2 FILLER_55_341 ();
 sg13g2_fill_2 FILLER_55_378 ();
 sg13g2_fill_2 FILLER_55_397 ();
 sg13g2_fill_2 FILLER_55_438 ();
 sg13g2_fill_2 FILLER_55_444 ();
 sg13g2_fill_1 FILLER_55_469 ();
 sg13g2_fill_2 FILLER_55_474 ();
 sg13g2_fill_2 FILLER_55_490 ();
 sg13g2_fill_1 FILLER_55_496 ();
 sg13g2_fill_1 FILLER_55_502 ();
 sg13g2_fill_2 FILLER_55_533 ();
 sg13g2_fill_1 FILLER_55_535 ();
 sg13g2_decap_4 FILLER_55_543 ();
 sg13g2_fill_1 FILLER_55_547 ();
 sg13g2_decap_8 FILLER_55_552 ();
 sg13g2_fill_2 FILLER_55_559 ();
 sg13g2_fill_1 FILLER_55_561 ();
 sg13g2_fill_2 FILLER_55_587 ();
 sg13g2_fill_1 FILLER_55_589 ();
 sg13g2_fill_1 FILLER_55_596 ();
 sg13g2_decap_8 FILLER_55_601 ();
 sg13g2_decap_8 FILLER_55_608 ();
 sg13g2_decap_8 FILLER_55_615 ();
 sg13g2_decap_8 FILLER_55_622 ();
 sg13g2_fill_2 FILLER_55_647 ();
 sg13g2_fill_2 FILLER_55_693 ();
 sg13g2_fill_2 FILLER_55_701 ();
 sg13g2_fill_1 FILLER_55_707 ();
 sg13g2_fill_1 FILLER_55_731 ();
 sg13g2_fill_2 FILLER_55_741 ();
 sg13g2_fill_2 FILLER_55_747 ();
 sg13g2_fill_1 FILLER_55_749 ();
 sg13g2_fill_2 FILLER_55_755 ();
 sg13g2_fill_1 FILLER_55_757 ();
 sg13g2_decap_8 FILLER_55_762 ();
 sg13g2_decap_4 FILLER_55_769 ();
 sg13g2_fill_2 FILLER_55_773 ();
 sg13g2_decap_4 FILLER_55_780 ();
 sg13g2_fill_1 FILLER_55_793 ();
 sg13g2_fill_1 FILLER_55_809 ();
 sg13g2_fill_2 FILLER_55_850 ();
 sg13g2_fill_1 FILLER_55_852 ();
 sg13g2_decap_8 FILLER_55_857 ();
 sg13g2_decap_8 FILLER_55_864 ();
 sg13g2_fill_1 FILLER_55_880 ();
 sg13g2_fill_2 FILLER_55_905 ();
 sg13g2_fill_2 FILLER_55_917 ();
 sg13g2_fill_1 FILLER_55_927 ();
 sg13g2_decap_4 FILLER_55_933 ();
 sg13g2_fill_1 FILLER_55_973 ();
 sg13g2_fill_1 FILLER_55_979 ();
 sg13g2_fill_1 FILLER_55_1006 ();
 sg13g2_fill_2 FILLER_55_1016 ();
 sg13g2_fill_1 FILLER_55_1057 ();
 sg13g2_fill_1 FILLER_55_1089 ();
 sg13g2_fill_2 FILLER_55_1126 ();
 sg13g2_fill_2 FILLER_55_1137 ();
 sg13g2_decap_8 FILLER_55_1165 ();
 sg13g2_decap_4 FILLER_55_1172 ();
 sg13g2_fill_1 FILLER_55_1176 ();
 sg13g2_decap_8 FILLER_55_1180 ();
 sg13g2_fill_1 FILLER_55_1187 ();
 sg13g2_decap_4 FILLER_55_1193 ();
 sg13g2_fill_1 FILLER_55_1197 ();
 sg13g2_fill_1 FILLER_55_1211 ();
 sg13g2_fill_1 FILLER_55_1219 ();
 sg13g2_fill_1 FILLER_55_1229 ();
 sg13g2_fill_2 FILLER_55_1240 ();
 sg13g2_decap_8 FILLER_55_1274 ();
 sg13g2_decap_8 FILLER_55_1281 ();
 sg13g2_decap_8 FILLER_55_1288 ();
 sg13g2_fill_2 FILLER_55_1295 ();
 sg13g2_fill_2 FILLER_55_1305 ();
 sg13g2_decap_4 FILLER_55_1311 ();
 sg13g2_fill_2 FILLER_55_1315 ();
 sg13g2_fill_1 FILLER_55_1327 ();
 sg13g2_decap_8 FILLER_55_1332 ();
 sg13g2_decap_8 FILLER_55_1339 ();
 sg13g2_fill_2 FILLER_55_1346 ();
 sg13g2_fill_2 FILLER_55_1352 ();
 sg13g2_fill_1 FILLER_55_1354 ();
 sg13g2_fill_1 FILLER_55_1369 ();
 sg13g2_fill_2 FILLER_55_1378 ();
 sg13g2_fill_1 FILLER_55_1385 ();
 sg13g2_decap_4 FILLER_55_1393 ();
 sg13g2_fill_2 FILLER_55_1397 ();
 sg13g2_fill_1 FILLER_55_1413 ();
 sg13g2_fill_2 FILLER_55_1419 ();
 sg13g2_decap_4 FILLER_55_1426 ();
 sg13g2_fill_1 FILLER_55_1451 ();
 sg13g2_decap_4 FILLER_55_1502 ();
 sg13g2_fill_2 FILLER_55_1519 ();
 sg13g2_decap_8 FILLER_55_1544 ();
 sg13g2_decap_8 FILLER_55_1551 ();
 sg13g2_fill_2 FILLER_55_1558 ();
 sg13g2_fill_2 FILLER_55_1564 ();
 sg13g2_fill_2 FILLER_55_1570 ();
 sg13g2_decap_8 FILLER_55_1576 ();
 sg13g2_decap_8 FILLER_55_1583 ();
 sg13g2_fill_2 FILLER_55_1590 ();
 sg13g2_fill_2 FILLER_55_1596 ();
 sg13g2_fill_1 FILLER_55_1598 ();
 sg13g2_decap_4 FILLER_55_1682 ();
 sg13g2_decap_8 FILLER_55_1691 ();
 sg13g2_fill_2 FILLER_55_1739 ();
 sg13g2_fill_1 FILLER_55_1741 ();
 sg13g2_fill_1 FILLER_55_1775 ();
 sg13g2_fill_1 FILLER_55_1803 ();
 sg13g2_fill_1 FILLER_55_1809 ();
 sg13g2_fill_1 FILLER_55_1815 ();
 sg13g2_fill_1 FILLER_55_1821 ();
 sg13g2_fill_1 FILLER_55_1837 ();
 sg13g2_decap_8 FILLER_55_1842 ();
 sg13g2_decap_8 FILLER_55_1849 ();
 sg13g2_decap_4 FILLER_55_1856 ();
 sg13g2_fill_2 FILLER_55_1891 ();
 sg13g2_decap_4 FILLER_55_1897 ();
 sg13g2_fill_1 FILLER_55_1901 ();
 sg13g2_fill_1 FILLER_55_1912 ();
 sg13g2_fill_1 FILLER_55_1930 ();
 sg13g2_fill_2 FILLER_55_1935 ();
 sg13g2_fill_1 FILLER_55_1949 ();
 sg13g2_decap_4 FILLER_55_1985 ();
 sg13g2_fill_1 FILLER_55_1994 ();
 sg13g2_fill_1 FILLER_55_2004 ();
 sg13g2_fill_2 FILLER_55_2009 ();
 sg13g2_fill_2 FILLER_55_2022 ();
 sg13g2_fill_1 FILLER_55_2029 ();
 sg13g2_fill_2 FILLER_55_2043 ();
 sg13g2_fill_2 FILLER_55_2054 ();
 sg13g2_decap_8 FILLER_55_2095 ();
 sg13g2_fill_2 FILLER_55_2102 ();
 sg13g2_fill_1 FILLER_55_2104 ();
 sg13g2_decap_8 FILLER_55_2109 ();
 sg13g2_decap_4 FILLER_55_2116 ();
 sg13g2_fill_1 FILLER_55_2163 ();
 sg13g2_fill_2 FILLER_55_2232 ();
 sg13g2_fill_2 FILLER_55_2242 ();
 sg13g2_fill_2 FILLER_55_2250 ();
 sg13g2_decap_8 FILLER_55_2295 ();
 sg13g2_decap_4 FILLER_55_2302 ();
 sg13g2_decap_8 FILLER_55_2316 ();
 sg13g2_fill_2 FILLER_55_2323 ();
 sg13g2_fill_1 FILLER_55_2331 ();
 sg13g2_decap_4 FILLER_55_2336 ();
 sg13g2_fill_1 FILLER_55_2340 ();
 sg13g2_decap_4 FILLER_55_2346 ();
 sg13g2_fill_1 FILLER_55_2350 ();
 sg13g2_fill_2 FILLER_55_2393 ();
 sg13g2_fill_2 FILLER_55_2399 ();
 sg13g2_fill_2 FILLER_55_2411 ();
 sg13g2_fill_2 FILLER_55_2423 ();
 sg13g2_fill_1 FILLER_55_2425 ();
 sg13g2_decap_8 FILLER_55_2430 ();
 sg13g2_decap_8 FILLER_55_2437 ();
 sg13g2_decap_8 FILLER_55_2444 ();
 sg13g2_fill_1 FILLER_55_2451 ();
 sg13g2_decap_4 FILLER_55_2457 ();
 sg13g2_fill_2 FILLER_55_2461 ();
 sg13g2_decap_4 FILLER_55_2472 ();
 sg13g2_fill_1 FILLER_55_2526 ();
 sg13g2_decap_8 FILLER_55_2567 ();
 sg13g2_decap_8 FILLER_55_2574 ();
 sg13g2_decap_8 FILLER_55_2581 ();
 sg13g2_decap_8 FILLER_55_2588 ();
 sg13g2_decap_8 FILLER_55_2595 ();
 sg13g2_decap_8 FILLER_55_2602 ();
 sg13g2_decap_8 FILLER_55_2609 ();
 sg13g2_decap_8 FILLER_55_2616 ();
 sg13g2_decap_8 FILLER_55_2623 ();
 sg13g2_decap_8 FILLER_55_2630 ();
 sg13g2_decap_8 FILLER_55_2637 ();
 sg13g2_decap_8 FILLER_55_2644 ();
 sg13g2_decap_8 FILLER_55_2651 ();
 sg13g2_decap_8 FILLER_55_2658 ();
 sg13g2_decap_4 FILLER_55_2665 ();
 sg13g2_fill_1 FILLER_55_2669 ();
 sg13g2_fill_2 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_33 ();
 sg13g2_fill_2 FILLER_56_39 ();
 sg13g2_fill_1 FILLER_56_41 ();
 sg13g2_fill_2 FILLER_56_82 ();
 sg13g2_fill_1 FILLER_56_89 ();
 sg13g2_fill_1 FILLER_56_95 ();
 sg13g2_fill_1 FILLER_56_148 ();
 sg13g2_fill_2 FILLER_56_179 ();
 sg13g2_decap_4 FILLER_56_186 ();
 sg13g2_fill_1 FILLER_56_190 ();
 sg13g2_fill_2 FILLER_56_230 ();
 sg13g2_fill_2 FILLER_56_260 ();
 sg13g2_fill_1 FILLER_56_262 ();
 sg13g2_decap_4 FILLER_56_273 ();
 sg13g2_fill_2 FILLER_56_291 ();
 sg13g2_fill_1 FILLER_56_297 ();
 sg13g2_fill_1 FILLER_56_307 ();
 sg13g2_fill_1 FILLER_56_413 ();
 sg13g2_fill_2 FILLER_56_433 ();
 sg13g2_fill_2 FILLER_56_448 ();
 sg13g2_fill_2 FILLER_56_468 ();
 sg13g2_decap_8 FILLER_56_488 ();
 sg13g2_decap_4 FILLER_56_495 ();
 sg13g2_fill_1 FILLER_56_499 ();
 sg13g2_fill_1 FILLER_56_505 ();
 sg13g2_fill_1 FILLER_56_521 ();
 sg13g2_fill_2 FILLER_56_531 ();
 sg13g2_fill_1 FILLER_56_540 ();
 sg13g2_fill_2 FILLER_56_545 ();
 sg13g2_fill_2 FILLER_56_598 ();
 sg13g2_fill_1 FILLER_56_600 ();
 sg13g2_fill_1 FILLER_56_704 ();
 sg13g2_decap_4 FILLER_56_709 ();
 sg13g2_fill_1 FILLER_56_713 ();
 sg13g2_fill_2 FILLER_56_722 ();
 sg13g2_fill_2 FILLER_56_728 ();
 sg13g2_fill_1 FILLER_56_730 ();
 sg13g2_decap_4 FILLER_56_739 ();
 sg13g2_fill_1 FILLER_56_748 ();
 sg13g2_fill_1 FILLER_56_761 ();
 sg13g2_decap_8 FILLER_56_767 ();
 sg13g2_fill_1 FILLER_56_774 ();
 sg13g2_decap_4 FILLER_56_783 ();
 sg13g2_decap_8 FILLER_56_799 ();
 sg13g2_fill_1 FILLER_56_824 ();
 sg13g2_decap_4 FILLER_56_861 ();
 sg13g2_fill_1 FILLER_56_895 ();
 sg13g2_fill_2 FILLER_56_922 ();
 sg13g2_decap_4 FILLER_56_949 ();
 sg13g2_fill_2 FILLER_56_953 ();
 sg13g2_fill_1 FILLER_56_959 ();
 sg13g2_fill_1 FILLER_56_980 ();
 sg13g2_fill_2 FILLER_56_1007 ();
 sg13g2_fill_2 FILLER_56_1035 ();
 sg13g2_fill_1 FILLER_56_1047 ();
 sg13g2_fill_2 FILLER_56_1067 ();
 sg13g2_fill_1 FILLER_56_1074 ();
 sg13g2_fill_1 FILLER_56_1101 ();
 sg13g2_fill_1 FILLER_56_1107 ();
 sg13g2_fill_1 FILLER_56_1118 ();
 sg13g2_fill_1 FILLER_56_1124 ();
 sg13g2_fill_1 FILLER_56_1130 ();
 sg13g2_decap_8 FILLER_56_1167 ();
 sg13g2_fill_2 FILLER_56_1174 ();
 sg13g2_fill_1 FILLER_56_1176 ();
 sg13g2_fill_1 FILLER_56_1195 ();
 sg13g2_decap_4 FILLER_56_1205 ();
 sg13g2_fill_1 FILLER_56_1209 ();
 sg13g2_fill_2 FILLER_56_1214 ();
 sg13g2_decap_4 FILLER_56_1222 ();
 sg13g2_fill_1 FILLER_56_1272 ();
 sg13g2_decap_8 FILLER_56_1282 ();
 sg13g2_fill_2 FILLER_56_1289 ();
 sg13g2_decap_8 FILLER_56_1295 ();
 sg13g2_fill_1 FILLER_56_1311 ();
 sg13g2_fill_2 FILLER_56_1317 ();
 sg13g2_fill_1 FILLER_56_1319 ();
 sg13g2_fill_1 FILLER_56_1325 ();
 sg13g2_decap_8 FILLER_56_1333 ();
 sg13g2_decap_4 FILLER_56_1340 ();
 sg13g2_fill_2 FILLER_56_1347 ();
 sg13g2_fill_1 FILLER_56_1354 ();
 sg13g2_fill_2 FILLER_56_1360 ();
 sg13g2_fill_1 FILLER_56_1362 ();
 sg13g2_fill_2 FILLER_56_1375 ();
 sg13g2_decap_4 FILLER_56_1407 ();
 sg13g2_fill_2 FILLER_56_1411 ();
 sg13g2_fill_1 FILLER_56_1420 ();
 sg13g2_fill_1 FILLER_56_1436 ();
 sg13g2_fill_1 FILLER_56_1476 ();
 sg13g2_decap_8 FILLER_56_1480 ();
 sg13g2_fill_1 FILLER_56_1487 ();
 sg13g2_decap_8 FILLER_56_1492 ();
 sg13g2_decap_8 FILLER_56_1499 ();
 sg13g2_decap_4 FILLER_56_1506 ();
 sg13g2_fill_2 FILLER_56_1510 ();
 sg13g2_decap_8 FILLER_56_1516 ();
 sg13g2_fill_1 FILLER_56_1523 ();
 sg13g2_fill_2 FILLER_56_1529 ();
 sg13g2_decap_4 FILLER_56_1541 ();
 sg13g2_decap_8 FILLER_56_1555 ();
 sg13g2_decap_8 FILLER_56_1562 ();
 sg13g2_fill_2 FILLER_56_1569 ();
 sg13g2_fill_1 FILLER_56_1610 ();
 sg13g2_fill_2 FILLER_56_1616 ();
 sg13g2_fill_2 FILLER_56_1622 ();
 sg13g2_decap_4 FILLER_56_1658 ();
 sg13g2_decap_4 FILLER_56_1666 ();
 sg13g2_fill_2 FILLER_56_1678 ();
 sg13g2_fill_2 FILLER_56_1686 ();
 sg13g2_fill_1 FILLER_56_1692 ();
 sg13g2_fill_2 FILLER_56_1707 ();
 sg13g2_fill_2 FILLER_56_1714 ();
 sg13g2_fill_2 FILLER_56_1719 ();
 sg13g2_fill_1 FILLER_56_1741 ();
 sg13g2_fill_2 FILLER_56_1747 ();
 sg13g2_decap_4 FILLER_56_1753 ();
 sg13g2_fill_1 FILLER_56_1757 ();
 sg13g2_fill_1 FILLER_56_1793 ();
 sg13g2_decap_4 FILLER_56_1799 ();
 sg13g2_fill_1 FILLER_56_1836 ();
 sg13g2_decap_8 FILLER_56_1851 ();
 sg13g2_decap_8 FILLER_56_1858 ();
 sg13g2_fill_1 FILLER_56_1865 ();
 sg13g2_decap_4 FILLER_56_1870 ();
 sg13g2_fill_1 FILLER_56_1874 ();
 sg13g2_fill_1 FILLER_56_1885 ();
 sg13g2_decap_4 FILLER_56_1922 ();
 sg13g2_fill_1 FILLER_56_1926 ();
 sg13g2_decap_4 FILLER_56_1932 ();
 sg13g2_fill_1 FILLER_56_1936 ();
 sg13g2_fill_2 FILLER_56_1943 ();
 sg13g2_fill_2 FILLER_56_1975 ();
 sg13g2_fill_2 FILLER_56_1983 ();
 sg13g2_fill_1 FILLER_56_1985 ();
 sg13g2_decap_8 FILLER_56_2020 ();
 sg13g2_fill_1 FILLER_56_2027 ();
 sg13g2_decap_8 FILLER_56_2054 ();
 sg13g2_fill_1 FILLER_56_2061 ();
 sg13g2_decap_8 FILLER_56_2088 ();
 sg13g2_decap_8 FILLER_56_2095 ();
 sg13g2_decap_8 FILLER_56_2102 ();
 sg13g2_decap_8 FILLER_56_2109 ();
 sg13g2_fill_2 FILLER_56_2116 ();
 sg13g2_fill_1 FILLER_56_2118 ();
 sg13g2_fill_2 FILLER_56_2124 ();
 sg13g2_fill_2 FILLER_56_2141 ();
 sg13g2_fill_1 FILLER_56_2154 ();
 sg13g2_fill_2 FILLER_56_2165 ();
 sg13g2_fill_1 FILLER_56_2211 ();
 sg13g2_fill_1 FILLER_56_2244 ();
 sg13g2_fill_2 FILLER_56_2265 ();
 sg13g2_fill_1 FILLER_56_2267 ();
 sg13g2_fill_2 FILLER_56_2326 ();
 sg13g2_fill_1 FILLER_56_2354 ();
 sg13g2_fill_1 FILLER_56_2365 ();
 sg13g2_fill_2 FILLER_56_2372 ();
 sg13g2_fill_1 FILLER_56_2374 ();
 sg13g2_decap_8 FILLER_56_2401 ();
 sg13g2_decap_4 FILLER_56_2408 ();
 sg13g2_decap_8 FILLER_56_2416 ();
 sg13g2_decap_8 FILLER_56_2423 ();
 sg13g2_decap_8 FILLER_56_2430 ();
 sg13g2_decap_8 FILLER_56_2437 ();
 sg13g2_decap_8 FILLER_56_2444 ();
 sg13g2_decap_4 FILLER_56_2451 ();
 sg13g2_fill_2 FILLER_56_2455 ();
 sg13g2_decap_8 FILLER_56_2461 ();
 sg13g2_fill_1 FILLER_56_2468 ();
 sg13g2_fill_2 FILLER_56_2474 ();
 sg13g2_fill_1 FILLER_56_2476 ();
 sg13g2_fill_1 FILLER_56_2490 ();
 sg13g2_fill_2 FILLER_56_2509 ();
 sg13g2_decap_8 FILLER_56_2537 ();
 sg13g2_decap_8 FILLER_56_2544 ();
 sg13g2_decap_8 FILLER_56_2551 ();
 sg13g2_decap_8 FILLER_56_2558 ();
 sg13g2_decap_8 FILLER_56_2565 ();
 sg13g2_decap_8 FILLER_56_2572 ();
 sg13g2_decap_8 FILLER_56_2579 ();
 sg13g2_decap_8 FILLER_56_2586 ();
 sg13g2_decap_8 FILLER_56_2593 ();
 sg13g2_decap_8 FILLER_56_2600 ();
 sg13g2_decap_8 FILLER_56_2607 ();
 sg13g2_decap_8 FILLER_56_2614 ();
 sg13g2_decap_8 FILLER_56_2621 ();
 sg13g2_decap_8 FILLER_56_2628 ();
 sg13g2_decap_8 FILLER_56_2635 ();
 sg13g2_decap_8 FILLER_56_2642 ();
 sg13g2_decap_8 FILLER_56_2649 ();
 sg13g2_decap_8 FILLER_56_2656 ();
 sg13g2_decap_8 FILLER_56_2663 ();
 sg13g2_fill_2 FILLER_57_34 ();
 sg13g2_fill_1 FILLER_57_41 ();
 sg13g2_fill_2 FILLER_57_47 ();
 sg13g2_fill_1 FILLER_57_59 ();
 sg13g2_fill_1 FILLER_57_65 ();
 sg13g2_fill_2 FILLER_57_103 ();
 sg13g2_fill_1 FILLER_57_105 ();
 sg13g2_decap_4 FILLER_57_136 ();
 sg13g2_fill_2 FILLER_57_140 ();
 sg13g2_fill_2 FILLER_57_151 ();
 sg13g2_fill_2 FILLER_57_169 ();
 sg13g2_fill_1 FILLER_57_171 ();
 sg13g2_decap_8 FILLER_57_177 ();
 sg13g2_decap_8 FILLER_57_184 ();
 sg13g2_decap_8 FILLER_57_191 ();
 sg13g2_decap_4 FILLER_57_198 ();
 sg13g2_decap_8 FILLER_57_216 ();
 sg13g2_decap_4 FILLER_57_223 ();
 sg13g2_fill_2 FILLER_57_227 ();
 sg13g2_decap_8 FILLER_57_277 ();
 sg13g2_fill_2 FILLER_57_284 ();
 sg13g2_fill_1 FILLER_57_286 ();
 sg13g2_decap_4 FILLER_57_293 ();
 sg13g2_fill_1 FILLER_57_297 ();
 sg13g2_decap_4 FILLER_57_314 ();
 sg13g2_fill_1 FILLER_57_318 ();
 sg13g2_fill_1 FILLER_57_356 ();
 sg13g2_fill_1 FILLER_57_365 ();
 sg13g2_fill_2 FILLER_57_376 ();
 sg13g2_fill_1 FILLER_57_397 ();
 sg13g2_fill_1 FILLER_57_440 ();
 sg13g2_fill_2 FILLER_57_475 ();
 sg13g2_fill_1 FILLER_57_487 ();
 sg13g2_fill_2 FILLER_57_492 ();
 sg13g2_fill_1 FILLER_57_498 ();
 sg13g2_fill_1 FILLER_57_509 ();
 sg13g2_decap_4 FILLER_57_514 ();
 sg13g2_fill_1 FILLER_57_518 ();
 sg13g2_fill_2 FILLER_57_543 ();
 sg13g2_fill_1 FILLER_57_557 ();
 sg13g2_fill_1 FILLER_57_562 ();
 sg13g2_fill_2 FILLER_57_567 ();
 sg13g2_fill_1 FILLER_57_580 ();
 sg13g2_fill_2 FILLER_57_599 ();
 sg13g2_fill_1 FILLER_57_613 ();
 sg13g2_fill_2 FILLER_57_677 ();
 sg13g2_fill_1 FILLER_57_679 ();
 sg13g2_fill_1 FILLER_57_691 ();
 sg13g2_fill_2 FILLER_57_700 ();
 sg13g2_decap_8 FILLER_57_707 ();
 sg13g2_decap_8 FILLER_57_714 ();
 sg13g2_decap_4 FILLER_57_721 ();
 sg13g2_decap_4 FILLER_57_734 ();
 sg13g2_decap_8 FILLER_57_742 ();
 sg13g2_fill_2 FILLER_57_757 ();
 sg13g2_fill_1 FILLER_57_759 ();
 sg13g2_decap_8 FILLER_57_774 ();
 sg13g2_decap_8 FILLER_57_785 ();
 sg13g2_decap_4 FILLER_57_792 ();
 sg13g2_fill_1 FILLER_57_796 ();
 sg13g2_decap_8 FILLER_57_801 ();
 sg13g2_decap_8 FILLER_57_808 ();
 sg13g2_decap_4 FILLER_57_879 ();
 sg13g2_decap_8 FILLER_57_898 ();
 sg13g2_decap_4 FILLER_57_905 ();
 sg13g2_fill_1 FILLER_57_909 ();
 sg13g2_decap_4 FILLER_57_928 ();
 sg13g2_fill_2 FILLER_57_932 ();
 sg13g2_fill_1 FILLER_57_969 ();
 sg13g2_fill_1 FILLER_57_991 ();
 sg13g2_fill_2 FILLER_57_999 ();
 sg13g2_fill_1 FILLER_57_1008 ();
 sg13g2_fill_1 FILLER_57_1014 ();
 sg13g2_fill_1 FILLER_57_1019 ();
 sg13g2_fill_1 FILLER_57_1046 ();
 sg13g2_fill_1 FILLER_57_1055 ();
 sg13g2_fill_2 FILLER_57_1080 ();
 sg13g2_decap_4 FILLER_57_1162 ();
 sg13g2_fill_1 FILLER_57_1166 ();
 sg13g2_fill_1 FILLER_57_1185 ();
 sg13g2_fill_2 FILLER_57_1198 ();
 sg13g2_decap_4 FILLER_57_1204 ();
 sg13g2_decap_4 FILLER_57_1212 ();
 sg13g2_fill_2 FILLER_57_1216 ();
 sg13g2_fill_1 FILLER_57_1233 ();
 sg13g2_fill_1 FILLER_57_1248 ();
 sg13g2_decap_4 FILLER_57_1279 ();
 sg13g2_decap_4 FILLER_57_1290 ();
 sg13g2_fill_2 FILLER_57_1294 ();
 sg13g2_fill_2 FILLER_57_1314 ();
 sg13g2_fill_1 FILLER_57_1335 ();
 sg13g2_decap_4 FILLER_57_1341 ();
 sg13g2_fill_1 FILLER_57_1345 ();
 sg13g2_fill_1 FILLER_57_1355 ();
 sg13g2_fill_1 FILLER_57_1369 ();
 sg13g2_fill_2 FILLER_57_1374 ();
 sg13g2_fill_1 FILLER_57_1376 ();
 sg13g2_fill_1 FILLER_57_1382 ();
 sg13g2_fill_1 FILLER_57_1388 ();
 sg13g2_fill_1 FILLER_57_1399 ();
 sg13g2_fill_2 FILLER_57_1426 ();
 sg13g2_fill_1 FILLER_57_1428 ();
 sg13g2_decap_4 FILLER_57_1493 ();
 sg13g2_fill_1 FILLER_57_1497 ();
 sg13g2_decap_4 FILLER_57_1502 ();
 sg13g2_fill_2 FILLER_57_1526 ();
 sg13g2_fill_1 FILLER_57_1528 ();
 sg13g2_decap_8 FILLER_57_1562 ();
 sg13g2_decap_8 FILLER_57_1569 ();
 sg13g2_decap_8 FILLER_57_1576 ();
 sg13g2_fill_1 FILLER_57_1583 ();
 sg13g2_decap_8 FILLER_57_1597 ();
 sg13g2_decap_4 FILLER_57_1608 ();
 sg13g2_fill_1 FILLER_57_1612 ();
 sg13g2_decap_4 FILLER_57_1622 ();
 sg13g2_fill_1 FILLER_57_1626 ();
 sg13g2_fill_2 FILLER_57_1643 ();
 sg13g2_fill_1 FILLER_57_1645 ();
 sg13g2_decap_8 FILLER_57_1677 ();
 sg13g2_decap_8 FILLER_57_1684 ();
 sg13g2_decap_8 FILLER_57_1691 ();
 sg13g2_decap_8 FILLER_57_1698 ();
 sg13g2_decap_4 FILLER_57_1705 ();
 sg13g2_fill_1 FILLER_57_1709 ();
 sg13g2_decap_8 FILLER_57_1715 ();
 sg13g2_fill_1 FILLER_57_1738 ();
 sg13g2_fill_2 FILLER_57_1761 ();
 sg13g2_fill_2 FILLER_57_1767 ();
 sg13g2_fill_1 FILLER_57_1791 ();
 sg13g2_fill_1 FILLER_57_1806 ();
 sg13g2_decap_4 FILLER_57_1837 ();
 sg13g2_fill_1 FILLER_57_1841 ();
 sg13g2_decap_8 FILLER_57_1847 ();
 sg13g2_fill_1 FILLER_57_1854 ();
 sg13g2_decap_8 FILLER_57_1911 ();
 sg13g2_fill_1 FILLER_57_1918 ();
 sg13g2_decap_8 FILLER_57_1924 ();
 sg13g2_fill_1 FILLER_57_1931 ();
 sg13g2_decap_8 FILLER_57_1973 ();
 sg13g2_fill_2 FILLER_57_1980 ();
 sg13g2_decap_4 FILLER_57_2008 ();
 sg13g2_fill_2 FILLER_57_2021 ();
 sg13g2_decap_4 FILLER_57_2027 ();
 sg13g2_fill_1 FILLER_57_2045 ();
 sg13g2_fill_2 FILLER_57_2056 ();
 sg13g2_decap_8 FILLER_57_2099 ();
 sg13g2_fill_2 FILLER_57_2142 ();
 sg13g2_fill_2 FILLER_57_2191 ();
 sg13g2_fill_2 FILLER_57_2209 ();
 sg13g2_fill_2 FILLER_57_2284 ();
 sg13g2_decap_4 FILLER_57_2290 ();
 sg13g2_fill_2 FILLER_57_2384 ();
 sg13g2_fill_1 FILLER_57_2394 ();
 sg13g2_decap_8 FILLER_57_2400 ();
 sg13g2_fill_1 FILLER_57_2407 ();
 sg13g2_fill_2 FILLER_57_2439 ();
 sg13g2_decap_8 FILLER_57_2578 ();
 sg13g2_decap_8 FILLER_57_2585 ();
 sg13g2_decap_8 FILLER_57_2592 ();
 sg13g2_decap_8 FILLER_57_2599 ();
 sg13g2_decap_8 FILLER_57_2606 ();
 sg13g2_decap_8 FILLER_57_2613 ();
 sg13g2_decap_8 FILLER_57_2620 ();
 sg13g2_decap_8 FILLER_57_2627 ();
 sg13g2_decap_8 FILLER_57_2634 ();
 sg13g2_decap_8 FILLER_57_2641 ();
 sg13g2_decap_8 FILLER_57_2648 ();
 sg13g2_decap_8 FILLER_57_2655 ();
 sg13g2_decap_8 FILLER_57_2662 ();
 sg13g2_fill_1 FILLER_57_2669 ();
 sg13g2_fill_1 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_31 ();
 sg13g2_fill_2 FILLER_58_50 ();
 sg13g2_fill_1 FILLER_58_83 ();
 sg13g2_fill_1 FILLER_58_89 ();
 sg13g2_fill_1 FILLER_58_93 ();
 sg13g2_fill_1 FILLER_58_99 ();
 sg13g2_fill_1 FILLER_58_110 ();
 sg13g2_fill_1 FILLER_58_116 ();
 sg13g2_decap_4 FILLER_58_121 ();
 sg13g2_decap_8 FILLER_58_129 ();
 sg13g2_fill_2 FILLER_58_136 ();
 sg13g2_fill_1 FILLER_58_138 ();
 sg13g2_fill_2 FILLER_58_152 ();
 sg13g2_fill_1 FILLER_58_154 ();
 sg13g2_fill_2 FILLER_58_160 ();
 sg13g2_fill_1 FILLER_58_162 ();
 sg13g2_decap_8 FILLER_58_176 ();
 sg13g2_decap_4 FILLER_58_183 ();
 sg13g2_fill_1 FILLER_58_213 ();
 sg13g2_decap_4 FILLER_58_224 ();
 sg13g2_fill_1 FILLER_58_228 ();
 sg13g2_decap_8 FILLER_58_245 ();
 sg13g2_fill_1 FILLER_58_252 ();
 sg13g2_fill_1 FILLER_58_267 ();
 sg13g2_fill_1 FILLER_58_272 ();
 sg13g2_fill_2 FILLER_58_299 ();
 sg13g2_fill_1 FILLER_58_307 ();
 sg13g2_decap_8 FILLER_58_313 ();
 sg13g2_fill_1 FILLER_58_344 ();
 sg13g2_fill_2 FILLER_58_363 ();
 sg13g2_fill_1 FILLER_58_391 ();
 sg13g2_fill_1 FILLER_58_401 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_fill_1 FILLER_58_415 ();
 sg13g2_fill_1 FILLER_58_423 ();
 sg13g2_fill_1 FILLER_58_429 ();
 sg13g2_fill_2 FILLER_58_437 ();
 sg13g2_fill_1 FILLER_58_465 ();
 sg13g2_fill_1 FILLER_58_471 ();
 sg13g2_fill_2 FILLER_58_477 ();
 sg13g2_fill_2 FILLER_58_505 ();
 sg13g2_fill_1 FILLER_58_507 ();
 sg13g2_fill_2 FILLER_58_513 ();
 sg13g2_fill_1 FILLER_58_548 ();
 sg13g2_fill_2 FILLER_58_569 ();
 sg13g2_fill_1 FILLER_58_571 ();
 sg13g2_decap_4 FILLER_58_595 ();
 sg13g2_decap_8 FILLER_58_606 ();
 sg13g2_fill_1 FILLER_58_642 ();
 sg13g2_decap_4 FILLER_58_647 ();
 sg13g2_decap_4 FILLER_58_668 ();
 sg13g2_fill_1 FILLER_58_714 ();
 sg13g2_decap_8 FILLER_58_719 ();
 sg13g2_fill_2 FILLER_58_762 ();
 sg13g2_fill_1 FILLER_58_764 ();
 sg13g2_fill_1 FILLER_58_805 ();
 sg13g2_fill_2 FILLER_58_810 ();
 sg13g2_fill_1 FILLER_58_812 ();
 sg13g2_fill_2 FILLER_58_839 ();
 sg13g2_fill_2 FILLER_58_874 ();
 sg13g2_fill_1 FILLER_58_876 ();
 sg13g2_fill_2 FILLER_58_882 ();
 sg13g2_decap_4 FILLER_58_889 ();
 sg13g2_fill_1 FILLER_58_893 ();
 sg13g2_decap_8 FILLER_58_898 ();
 sg13g2_decap_4 FILLER_58_905 ();
 sg13g2_fill_1 FILLER_58_909 ();
 sg13g2_fill_2 FILLER_58_930 ();
 sg13g2_fill_1 FILLER_58_937 ();
 sg13g2_fill_2 FILLER_58_943 ();
 sg13g2_fill_1 FILLER_58_950 ();
 sg13g2_fill_2 FILLER_58_956 ();
 sg13g2_fill_1 FILLER_58_962 ();
 sg13g2_fill_2 FILLER_58_975 ();
 sg13g2_fill_2 FILLER_58_990 ();
 sg13g2_fill_1 FILLER_58_1005 ();
 sg13g2_fill_1 FILLER_58_1022 ();
 sg13g2_fill_1 FILLER_58_1028 ();
 sg13g2_fill_1 FILLER_58_1033 ();
 sg13g2_fill_2 FILLER_58_1038 ();
 sg13g2_fill_1 FILLER_58_1044 ();
 sg13g2_fill_1 FILLER_58_1084 ();
 sg13g2_fill_1 FILLER_58_1096 ();
 sg13g2_decap_4 FILLER_58_1153 ();
 sg13g2_decap_8 FILLER_58_1165 ();
 sg13g2_decap_4 FILLER_58_1172 ();
 sg13g2_fill_2 FILLER_58_1180 ();
 sg13g2_fill_1 FILLER_58_1209 ();
 sg13g2_fill_1 FILLER_58_1216 ();
 sg13g2_fill_1 FILLER_58_1221 ();
 sg13g2_fill_1 FILLER_58_1226 ();
 sg13g2_fill_2 FILLER_58_1247 ();
 sg13g2_fill_1 FILLER_58_1249 ();
 sg13g2_decap_4 FILLER_58_1289 ();
 sg13g2_fill_2 FILLER_58_1297 ();
 sg13g2_fill_1 FILLER_58_1299 ();
 sg13g2_fill_2 FILLER_58_1316 ();
 sg13g2_fill_1 FILLER_58_1318 ();
 sg13g2_fill_2 FILLER_58_1326 ();
 sg13g2_fill_2 FILLER_58_1333 ();
 sg13g2_decap_4 FILLER_58_1356 ();
 sg13g2_decap_8 FILLER_58_1370 ();
 sg13g2_fill_2 FILLER_58_1377 ();
 sg13g2_fill_2 FILLER_58_1384 ();
 sg13g2_fill_1 FILLER_58_1386 ();
 sg13g2_fill_1 FILLER_58_1390 ();
 sg13g2_fill_1 FILLER_58_1401 ();
 sg13g2_decap_8 FILLER_58_1406 ();
 sg13g2_fill_2 FILLER_58_1421 ();
 sg13g2_fill_1 FILLER_58_1423 ();
 sg13g2_fill_1 FILLER_58_1479 ();
 sg13g2_fill_1 FILLER_58_1495 ();
 sg13g2_decap_4 FILLER_58_1532 ();
 sg13g2_fill_1 FILLER_58_1541 ();
 sg13g2_decap_8 FILLER_58_1561 ();
 sg13g2_fill_1 FILLER_58_1612 ();
 sg13g2_decap_8 FILLER_58_1631 ();
 sg13g2_decap_8 FILLER_58_1638 ();
 sg13g2_fill_1 FILLER_58_1645 ();
 sg13g2_fill_2 FILLER_58_1650 ();
 sg13g2_decap_4 FILLER_58_1656 ();
 sg13g2_fill_1 FILLER_58_1660 ();
 sg13g2_decap_8 FILLER_58_1680 ();
 sg13g2_fill_2 FILLER_58_1687 ();
 sg13g2_fill_1 FILLER_58_1689 ();
 sg13g2_decap_4 FILLER_58_1695 ();
 sg13g2_fill_1 FILLER_58_1718 ();
 sg13g2_decap_4 FILLER_58_1724 ();
 sg13g2_fill_2 FILLER_58_1728 ();
 sg13g2_fill_2 FILLER_58_1738 ();
 sg13g2_fill_1 FILLER_58_1749 ();
 sg13g2_fill_2 FILLER_58_1758 ();
 sg13g2_fill_1 FILLER_58_1796 ();
 sg13g2_fill_1 FILLER_58_1802 ();
 sg13g2_decap_8 FILLER_58_1816 ();
 sg13g2_fill_1 FILLER_58_1828 ();
 sg13g2_fill_1 FILLER_58_1855 ();
 sg13g2_decap_4 FILLER_58_1887 ();
 sg13g2_fill_1 FILLER_58_1891 ();
 sg13g2_fill_2 FILLER_58_1934 ();
 sg13g2_decap_8 FILLER_58_1969 ();
 sg13g2_decap_8 FILLER_58_1976 ();
 sg13g2_fill_1 FILLER_58_1983 ();
 sg13g2_fill_1 FILLER_58_1993 ();
 sg13g2_decap_8 FILLER_58_1998 ();
 sg13g2_fill_1 FILLER_58_2017 ();
 sg13g2_fill_2 FILLER_58_2082 ();
 sg13g2_fill_2 FILLER_58_2094 ();
 sg13g2_fill_1 FILLER_58_2096 ();
 sg13g2_fill_2 FILLER_58_2131 ();
 sg13g2_fill_1 FILLER_58_2243 ();
 sg13g2_decap_4 FILLER_58_2274 ();
 sg13g2_decap_8 FILLER_58_2294 ();
 sg13g2_fill_2 FILLER_58_2301 ();
 sg13g2_fill_2 FILLER_58_2307 ();
 sg13g2_fill_2 FILLER_58_2315 ();
 sg13g2_fill_1 FILLER_58_2317 ();
 sg13g2_decap_8 FILLER_58_2328 ();
 sg13g2_fill_1 FILLER_58_2335 ();
 sg13g2_fill_1 FILLER_58_2340 ();
 sg13g2_fill_2 FILLER_58_2347 ();
 sg13g2_fill_2 FILLER_58_2355 ();
 sg13g2_fill_2 FILLER_58_2361 ();
 sg13g2_fill_2 FILLER_58_2367 ();
 sg13g2_fill_1 FILLER_58_2369 ();
 sg13g2_fill_1 FILLER_58_2376 ();
 sg13g2_fill_2 FILLER_58_2383 ();
 sg13g2_fill_1 FILLER_58_2420 ();
 sg13g2_fill_2 FILLER_58_2461 ();
 sg13g2_fill_1 FILLER_58_2493 ();
 sg13g2_fill_2 FILLER_58_2504 ();
 sg13g2_fill_2 FILLER_58_2510 ();
 sg13g2_fill_2 FILLER_58_2538 ();
 sg13g2_decap_8 FILLER_58_2576 ();
 sg13g2_decap_8 FILLER_58_2583 ();
 sg13g2_decap_8 FILLER_58_2590 ();
 sg13g2_decap_8 FILLER_58_2597 ();
 sg13g2_decap_8 FILLER_58_2604 ();
 sg13g2_decap_8 FILLER_58_2611 ();
 sg13g2_decap_8 FILLER_58_2618 ();
 sg13g2_decap_8 FILLER_58_2625 ();
 sg13g2_decap_8 FILLER_58_2632 ();
 sg13g2_decap_8 FILLER_58_2639 ();
 sg13g2_decap_8 FILLER_58_2646 ();
 sg13g2_decap_8 FILLER_58_2653 ();
 sg13g2_decap_8 FILLER_58_2660 ();
 sg13g2_fill_2 FILLER_58_2667 ();
 sg13g2_fill_1 FILLER_58_2669 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_fill_1 FILLER_59_36 ();
 sg13g2_decap_4 FILLER_59_51 ();
 sg13g2_fill_2 FILLER_59_55 ();
 sg13g2_decap_4 FILLER_59_61 ();
 sg13g2_fill_1 FILLER_59_69 ();
 sg13g2_fill_2 FILLER_59_88 ();
 sg13g2_fill_2 FILLER_59_102 ();
 sg13g2_decap_4 FILLER_59_112 ();
 sg13g2_fill_2 FILLER_59_116 ();
 sg13g2_fill_1 FILLER_59_123 ();
 sg13g2_fill_1 FILLER_59_129 ();
 sg13g2_fill_1 FILLER_59_135 ();
 sg13g2_fill_1 FILLER_59_140 ();
 sg13g2_fill_1 FILLER_59_146 ();
 sg13g2_fill_1 FILLER_59_173 ();
 sg13g2_decap_4 FILLER_59_195 ();
 sg13g2_decap_8 FILLER_59_214 ();
 sg13g2_decap_4 FILLER_59_221 ();
 sg13g2_decap_8 FILLER_59_230 ();
 sg13g2_decap_4 FILLER_59_237 ();
 sg13g2_fill_1 FILLER_59_241 ();
 sg13g2_fill_2 FILLER_59_277 ();
 sg13g2_fill_1 FILLER_59_279 ();
 sg13g2_decap_4 FILLER_59_284 ();
 sg13g2_fill_2 FILLER_59_288 ();
 sg13g2_fill_1 FILLER_59_295 ();
 sg13g2_fill_1 FILLER_59_301 ();
 sg13g2_fill_1 FILLER_59_306 ();
 sg13g2_fill_1 FILLER_59_315 ();
 sg13g2_decap_4 FILLER_59_325 ();
 sg13g2_fill_1 FILLER_59_329 ();
 sg13g2_fill_1 FILLER_59_356 ();
 sg13g2_fill_2 FILLER_59_365 ();
 sg13g2_fill_1 FILLER_59_417 ();
 sg13g2_fill_2 FILLER_59_529 ();
 sg13g2_fill_1 FILLER_59_583 ();
 sg13g2_fill_1 FILLER_59_588 ();
 sg13g2_decap_8 FILLER_59_603 ();
 sg13g2_decap_8 FILLER_59_610 ();
 sg13g2_fill_2 FILLER_59_617 ();
 sg13g2_decap_4 FILLER_59_634 ();
 sg13g2_fill_1 FILLER_59_638 ();
 sg13g2_decap_8 FILLER_59_644 ();
 sg13g2_fill_2 FILLER_59_651 ();
 sg13g2_fill_1 FILLER_59_653 ();
 sg13g2_decap_4 FILLER_59_659 ();
 sg13g2_fill_1 FILLER_59_663 ();
 sg13g2_decap_4 FILLER_59_672 ();
 sg13g2_fill_2 FILLER_59_676 ();
 sg13g2_fill_2 FILLER_59_723 ();
 sg13g2_fill_2 FILLER_59_729 ();
 sg13g2_fill_1 FILLER_59_731 ();
 sg13g2_fill_1 FILLER_59_768 ();
 sg13g2_fill_1 FILLER_59_795 ();
 sg13g2_fill_1 FILLER_59_834 ();
 sg13g2_fill_2 FILLER_59_871 ();
 sg13g2_decap_8 FILLER_59_899 ();
 sg13g2_decap_4 FILLER_59_906 ();
 sg13g2_fill_1 FILLER_59_910 ();
 sg13g2_fill_1 FILLER_59_920 ();
 sg13g2_fill_1 FILLER_59_932 ();
 sg13g2_fill_1 FILLER_59_938 ();
 sg13g2_fill_1 FILLER_59_943 ();
 sg13g2_fill_2 FILLER_59_951 ();
 sg13g2_fill_1 FILLER_59_953 ();
 sg13g2_fill_2 FILLER_59_963 ();
 sg13g2_fill_1 FILLER_59_965 ();
 sg13g2_fill_1 FILLER_59_971 ();
 sg13g2_fill_1 FILLER_59_982 ();
 sg13g2_fill_2 FILLER_59_1002 ();
 sg13g2_fill_1 FILLER_59_1012 ();
 sg13g2_fill_2 FILLER_59_1016 ();
 sg13g2_fill_2 FILLER_59_1033 ();
 sg13g2_decap_4 FILLER_59_1038 ();
 sg13g2_fill_2 FILLER_59_1042 ();
 sg13g2_fill_1 FILLER_59_1047 ();
 sg13g2_fill_2 FILLER_59_1065 ();
 sg13g2_fill_1 FILLER_59_1112 ();
 sg13g2_fill_2 FILLER_59_1118 ();
 sg13g2_fill_1 FILLER_59_1129 ();
 sg13g2_decap_4 FILLER_59_1136 ();
 sg13g2_decap_4 FILLER_59_1144 ();
 sg13g2_fill_2 FILLER_59_1148 ();
 sg13g2_decap_8 FILLER_59_1154 ();
 sg13g2_fill_2 FILLER_59_1161 ();
 sg13g2_decap_8 FILLER_59_1166 ();
 sg13g2_decap_8 FILLER_59_1173 ();
 sg13g2_fill_1 FILLER_59_1180 ();
 sg13g2_fill_2 FILLER_59_1198 ();
 sg13g2_fill_1 FILLER_59_1200 ();
 sg13g2_decap_4 FILLER_59_1205 ();
 sg13g2_fill_2 FILLER_59_1209 ();
 sg13g2_fill_1 FILLER_59_1226 ();
 sg13g2_fill_2 FILLER_59_1235 ();
 sg13g2_decap_8 FILLER_59_1254 ();
 sg13g2_fill_2 FILLER_59_1261 ();
 sg13g2_fill_1 FILLER_59_1263 ();
 sg13g2_decap_8 FILLER_59_1289 ();
 sg13g2_decap_8 FILLER_59_1296 ();
 sg13g2_fill_1 FILLER_59_1303 ();
 sg13g2_decap_4 FILLER_59_1321 ();
 sg13g2_fill_2 FILLER_59_1325 ();
 sg13g2_decap_8 FILLER_59_1331 ();
 sg13g2_decap_4 FILLER_59_1338 ();
 sg13g2_fill_2 FILLER_59_1342 ();
 sg13g2_decap_8 FILLER_59_1348 ();
 sg13g2_decap_4 FILLER_59_1355 ();
 sg13g2_fill_1 FILLER_59_1364 ();
 sg13g2_fill_2 FILLER_59_1370 ();
 sg13g2_fill_1 FILLER_59_1372 ();
 sg13g2_fill_2 FILLER_59_1378 ();
 sg13g2_fill_1 FILLER_59_1389 ();
 sg13g2_decap_4 FILLER_59_1405 ();
 sg13g2_decap_4 FILLER_59_1419 ();
 sg13g2_fill_1 FILLER_59_1423 ();
 sg13g2_decap_8 FILLER_59_1429 ();
 sg13g2_decap_8 FILLER_59_1436 ();
 sg13g2_decap_4 FILLER_59_1443 ();
 sg13g2_decap_4 FILLER_59_1461 ();
 sg13g2_decap_8 FILLER_59_1477 ();
 sg13g2_decap_8 FILLER_59_1484 ();
 sg13g2_fill_2 FILLER_59_1491 ();
 sg13g2_fill_1 FILLER_59_1493 ();
 sg13g2_fill_1 FILLER_59_1499 ();
 sg13g2_decap_4 FILLER_59_1505 ();
 sg13g2_fill_2 FILLER_59_1509 ();
 sg13g2_fill_2 FILLER_59_1524 ();
 sg13g2_fill_2 FILLER_59_1545 ();
 sg13g2_fill_1 FILLER_59_1547 ();
 sg13g2_fill_2 FILLER_59_1553 ();
 sg13g2_decap_4 FILLER_59_1565 ();
 sg13g2_fill_1 FILLER_59_1569 ();
 sg13g2_fill_2 FILLER_59_1607 ();
 sg13g2_fill_1 FILLER_59_1609 ();
 sg13g2_fill_1 FILLER_59_1614 ();
 sg13g2_fill_1 FILLER_59_1641 ();
 sg13g2_fill_2 FILLER_59_1668 ();
 sg13g2_fill_1 FILLER_59_1696 ();
 sg13g2_fill_1 FILLER_59_1728 ();
 sg13g2_decap_4 FILLER_59_1735 ();
 sg13g2_fill_2 FILLER_59_1739 ();
 sg13g2_fill_1 FILLER_59_1778 ();
 sg13g2_fill_1 FILLER_59_1783 ();
 sg13g2_fill_1 FILLER_59_1789 ();
 sg13g2_fill_1 FILLER_59_1808 ();
 sg13g2_decap_4 FILLER_59_1848 ();
 sg13g2_fill_1 FILLER_59_1872 ();
 sg13g2_fill_1 FILLER_59_1878 ();
 sg13g2_fill_2 FILLER_59_1883 ();
 sg13g2_decap_8 FILLER_59_1893 ();
 sg13g2_decap_4 FILLER_59_1900 ();
 sg13g2_fill_1 FILLER_59_1913 ();
 sg13g2_fill_1 FILLER_59_1918 ();
 sg13g2_fill_2 FILLER_59_1924 ();
 sg13g2_fill_1 FILLER_59_1930 ();
 sg13g2_fill_2 FILLER_59_1945 ();
 sg13g2_fill_2 FILLER_59_1960 ();
 sg13g2_fill_1 FILLER_59_1962 ();
 sg13g2_decap_8 FILLER_59_1969 ();
 sg13g2_decap_4 FILLER_59_1976 ();
 sg13g2_fill_1 FILLER_59_1980 ();
 sg13g2_fill_1 FILLER_59_2011 ();
 sg13g2_fill_1 FILLER_59_2043 ();
 sg13g2_fill_1 FILLER_59_2048 ();
 sg13g2_fill_2 FILLER_59_2101 ();
 sg13g2_fill_2 FILLER_59_2107 ();
 sg13g2_fill_1 FILLER_59_2109 ();
 sg13g2_decap_4 FILLER_59_2137 ();
 sg13g2_fill_1 FILLER_59_2151 ();
 sg13g2_fill_2 FILLER_59_2162 ();
 sg13g2_fill_2 FILLER_59_2168 ();
 sg13g2_fill_2 FILLER_59_2187 ();
 sg13g2_fill_1 FILLER_59_2205 ();
 sg13g2_fill_1 FILLER_59_2209 ();
 sg13g2_fill_1 FILLER_59_2245 ();
 sg13g2_fill_2 FILLER_59_2263 ();
 sg13g2_fill_2 FILLER_59_2282 ();
 sg13g2_decap_8 FILLER_59_2318 ();
 sg13g2_decap_4 FILLER_59_2325 ();
 sg13g2_fill_1 FILLER_59_2329 ();
 sg13g2_decap_8 FILLER_59_2342 ();
 sg13g2_decap_8 FILLER_59_2349 ();
 sg13g2_decap_8 FILLER_59_2356 ();
 sg13g2_fill_1 FILLER_59_2363 ();
 sg13g2_fill_2 FILLER_59_2378 ();
 sg13g2_fill_1 FILLER_59_2380 ();
 sg13g2_fill_2 FILLER_59_2444 ();
 sg13g2_fill_2 FILLER_59_2456 ();
 sg13g2_fill_2 FILLER_59_2468 ();
 sg13g2_fill_2 FILLER_59_2552 ();
 sg13g2_decap_8 FILLER_59_2580 ();
 sg13g2_decap_8 FILLER_59_2587 ();
 sg13g2_decap_8 FILLER_59_2594 ();
 sg13g2_decap_8 FILLER_59_2601 ();
 sg13g2_decap_8 FILLER_59_2608 ();
 sg13g2_decap_8 FILLER_59_2615 ();
 sg13g2_decap_8 FILLER_59_2622 ();
 sg13g2_decap_8 FILLER_59_2629 ();
 sg13g2_decap_8 FILLER_59_2636 ();
 sg13g2_decap_8 FILLER_59_2643 ();
 sg13g2_decap_8 FILLER_59_2650 ();
 sg13g2_decap_8 FILLER_59_2657 ();
 sg13g2_decap_4 FILLER_59_2664 ();
 sg13g2_fill_2 FILLER_59_2668 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_4 FILLER_60_7 ();
 sg13g2_fill_1 FILLER_60_11 ();
 sg13g2_fill_1 FILLER_60_42 ();
 sg13g2_fill_1 FILLER_60_69 ();
 sg13g2_decap_4 FILLER_60_76 ();
 sg13g2_fill_2 FILLER_60_104 ();
 sg13g2_fill_1 FILLER_60_136 ();
 sg13g2_fill_1 FILLER_60_142 ();
 sg13g2_fill_1 FILLER_60_149 ();
 sg13g2_fill_1 FILLER_60_154 ();
 sg13g2_decap_4 FILLER_60_165 ();
 sg13g2_fill_1 FILLER_60_169 ();
 sg13g2_fill_1 FILLER_60_176 ();
 sg13g2_fill_2 FILLER_60_182 ();
 sg13g2_fill_2 FILLER_60_194 ();
 sg13g2_fill_1 FILLER_60_196 ();
 sg13g2_fill_2 FILLER_60_202 ();
 sg13g2_fill_1 FILLER_60_230 ();
 sg13g2_decap_4 FILLER_60_257 ();
 sg13g2_fill_1 FILLER_60_261 ();
 sg13g2_decap_8 FILLER_60_267 ();
 sg13g2_decap_8 FILLER_60_274 ();
 sg13g2_fill_2 FILLER_60_281 ();
 sg13g2_fill_1 FILLER_60_291 ();
 sg13g2_decap_4 FILLER_60_298 ();
 sg13g2_fill_1 FILLER_60_302 ();
 sg13g2_fill_1 FILLER_60_307 ();
 sg13g2_fill_1 FILLER_60_329 ();
 sg13g2_fill_1 FILLER_60_335 ();
 sg13g2_fill_2 FILLER_60_344 ();
 sg13g2_fill_1 FILLER_60_354 ();
 sg13g2_fill_1 FILLER_60_360 ();
 sg13g2_fill_2 FILLER_60_365 ();
 sg13g2_fill_1 FILLER_60_372 ();
 sg13g2_fill_1 FILLER_60_381 ();
 sg13g2_fill_1 FILLER_60_413 ();
 sg13g2_fill_2 FILLER_60_424 ();
 sg13g2_fill_2 FILLER_60_471 ();
 sg13g2_fill_1 FILLER_60_473 ();
 sg13g2_fill_2 FILLER_60_478 ();
 sg13g2_fill_1 FILLER_60_501 ();
 sg13g2_fill_1 FILLER_60_507 ();
 sg13g2_fill_1 FILLER_60_534 ();
 sg13g2_fill_1 FILLER_60_561 ();
 sg13g2_fill_1 FILLER_60_571 ();
 sg13g2_fill_1 FILLER_60_576 ();
 sg13g2_fill_1 FILLER_60_664 ();
 sg13g2_fill_2 FILLER_60_675 ();
 sg13g2_fill_2 FILLER_60_710 ();
 sg13g2_fill_2 FILLER_60_803 ();
 sg13g2_fill_1 FILLER_60_805 ();
 sg13g2_fill_2 FILLER_60_816 ();
 sg13g2_decap_8 FILLER_60_835 ();
 sg13g2_decap_4 FILLER_60_842 ();
 sg13g2_fill_2 FILLER_60_846 ();
 sg13g2_decap_4 FILLER_60_852 ();
 sg13g2_fill_1 FILLER_60_856 ();
 sg13g2_decap_8 FILLER_60_869 ();
 sg13g2_fill_2 FILLER_60_885 ();
 sg13g2_fill_1 FILLER_60_887 ();
 sg13g2_fill_1 FILLER_60_892 ();
 sg13g2_fill_2 FILLER_60_935 ();
 sg13g2_fill_1 FILLER_60_937 ();
 sg13g2_fill_2 FILLER_60_948 ();
 sg13g2_fill_1 FILLER_60_954 ();
 sg13g2_fill_1 FILLER_60_965 ();
 sg13g2_decap_4 FILLER_60_997 ();
 sg13g2_fill_2 FILLER_60_1004 ();
 sg13g2_fill_2 FILLER_60_1017 ();
 sg13g2_decap_8 FILLER_60_1027 ();
 sg13g2_fill_1 FILLER_60_1034 ();
 sg13g2_decap_8 FILLER_60_1040 ();
 sg13g2_decap_4 FILLER_60_1047 ();
 sg13g2_decap_4 FILLER_60_1071 ();
 sg13g2_fill_1 FILLER_60_1088 ();
 sg13g2_fill_2 FILLER_60_1125 ();
 sg13g2_fill_1 FILLER_60_1132 ();
 sg13g2_decap_4 FILLER_60_1138 ();
 sg13g2_fill_1 FILLER_60_1142 ();
 sg13g2_decap_8 FILLER_60_1172 ();
 sg13g2_decap_8 FILLER_60_1179 ();
 sg13g2_fill_2 FILLER_60_1186 ();
 sg13g2_fill_2 FILLER_60_1197 ();
 sg13g2_fill_1 FILLER_60_1204 ();
 sg13g2_fill_1 FILLER_60_1210 ();
 sg13g2_fill_1 FILLER_60_1215 ();
 sg13g2_fill_1 FILLER_60_1226 ();
 sg13g2_decap_8 FILLER_60_1232 ();
 sg13g2_decap_4 FILLER_60_1248 ();
 sg13g2_fill_2 FILLER_60_1252 ();
 sg13g2_fill_1 FILLER_60_1259 ();
 sg13g2_decap_8 FILLER_60_1264 ();
 sg13g2_fill_1 FILLER_60_1271 ();
 sg13g2_fill_1 FILLER_60_1289 ();
 sg13g2_decap_8 FILLER_60_1295 ();
 sg13g2_decap_4 FILLER_60_1302 ();
 sg13g2_fill_1 FILLER_60_1311 ();
 sg13g2_decap_8 FILLER_60_1317 ();
 sg13g2_decap_8 FILLER_60_1324 ();
 sg13g2_decap_4 FILLER_60_1331 ();
 sg13g2_fill_1 FILLER_60_1335 ();
 sg13g2_fill_2 FILLER_60_1340 ();
 sg13g2_fill_1 FILLER_60_1342 ();
 sg13g2_decap_8 FILLER_60_1351 ();
 sg13g2_decap_8 FILLER_60_1363 ();
 sg13g2_decap_4 FILLER_60_1404 ();
 sg13g2_fill_1 FILLER_60_1408 ();
 sg13g2_decap_8 FILLER_60_1414 ();
 sg13g2_decap_8 FILLER_60_1428 ();
 sg13g2_decap_8 FILLER_60_1435 ();
 sg13g2_decap_4 FILLER_60_1442 ();
 sg13g2_fill_1 FILLER_60_1446 ();
 sg13g2_decap_8 FILLER_60_1457 ();
 sg13g2_fill_2 FILLER_60_1464 ();
 sg13g2_fill_1 FILLER_60_1466 ();
 sg13g2_decap_4 FILLER_60_1486 ();
 sg13g2_fill_2 FILLER_60_1490 ();
 sg13g2_decap_8 FILLER_60_1497 ();
 sg13g2_fill_2 FILLER_60_1504 ();
 sg13g2_fill_2 FILLER_60_1510 ();
 sg13g2_fill_1 FILLER_60_1512 ();
 sg13g2_decap_8 FILLER_60_1526 ();
 sg13g2_decap_4 FILLER_60_1533 ();
 sg13g2_fill_1 FILLER_60_1541 ();
 sg13g2_decap_8 FILLER_60_1572 ();
 sg13g2_decap_8 FILLER_60_1579 ();
 sg13g2_fill_1 FILLER_60_1586 ();
 sg13g2_fill_1 FILLER_60_1622 ();
 sg13g2_fill_2 FILLER_60_1633 ();
 sg13g2_fill_2 FILLER_60_1639 ();
 sg13g2_fill_2 FILLER_60_1667 ();
 sg13g2_fill_1 FILLER_60_1669 ();
 sg13g2_fill_1 FILLER_60_1678 ();
 sg13g2_fill_2 FILLER_60_1684 ();
 sg13g2_fill_2 FILLER_60_1708 ();
 sg13g2_fill_1 FILLER_60_1710 ();
 sg13g2_fill_1 FILLER_60_1723 ();
 sg13g2_fill_2 FILLER_60_1737 ();
 sg13g2_fill_1 FILLER_60_1744 ();
 sg13g2_fill_2 FILLER_60_1764 ();
 sg13g2_fill_1 FILLER_60_1771 ();
 sg13g2_fill_1 FILLER_60_1816 ();
 sg13g2_fill_2 FILLER_60_1828 ();
 sg13g2_fill_1 FILLER_60_1835 ();
 sg13g2_fill_1 FILLER_60_1840 ();
 sg13g2_fill_1 FILLER_60_1845 ();
 sg13g2_fill_1 FILLER_60_1850 ();
 sg13g2_fill_2 FILLER_60_1854 ();
 sg13g2_fill_1 FILLER_60_1856 ();
 sg13g2_decap_8 FILLER_60_1895 ();
 sg13g2_decap_4 FILLER_60_1902 ();
 sg13g2_fill_1 FILLER_60_1906 ();
 sg13g2_decap_8 FILLER_60_1974 ();
 sg13g2_fill_2 FILLER_60_1981 ();
 sg13g2_fill_1 FILLER_60_1992 ();
 sg13g2_fill_2 FILLER_60_2022 ();
 sg13g2_decap_4 FILLER_60_2028 ();
 sg13g2_fill_1 FILLER_60_2036 ();
 sg13g2_decap_4 FILLER_60_2045 ();
 sg13g2_decap_8 FILLER_60_2089 ();
 sg13g2_decap_4 FILLER_60_2096 ();
 sg13g2_fill_1 FILLER_60_2100 ();
 sg13g2_decap_8 FILLER_60_2147 ();
 sg13g2_fill_1 FILLER_60_2164 ();
 sg13g2_fill_1 FILLER_60_2169 ();
 sg13g2_fill_2 FILLER_60_2209 ();
 sg13g2_fill_2 FILLER_60_2226 ();
 sg13g2_fill_1 FILLER_60_2260 ();
 sg13g2_fill_1 FILLER_60_2265 ();
 sg13g2_fill_1 FILLER_60_2308 ();
 sg13g2_fill_2 FILLER_60_2314 ();
 sg13g2_fill_1 FILLER_60_2320 ();
 sg13g2_decap_4 FILLER_60_2324 ();
 sg13g2_fill_2 FILLER_60_2328 ();
 sg13g2_fill_1 FILLER_60_2348 ();
 sg13g2_fill_2 FILLER_60_2387 ();
 sg13g2_fill_2 FILLER_60_2395 ();
 sg13g2_fill_2 FILLER_60_2410 ();
 sg13g2_fill_2 FILLER_60_2483 ();
 sg13g2_fill_1 FILLER_60_2485 ();
 sg13g2_decap_4 FILLER_60_2490 ();
 sg13g2_decap_8 FILLER_60_2508 ();
 sg13g2_decap_4 FILLER_60_2515 ();
 sg13g2_decap_4 FILLER_60_2529 ();
 sg13g2_fill_2 FILLER_60_2533 ();
 sg13g2_decap_4 FILLER_60_2539 ();
 sg13g2_decap_4 FILLER_60_2553 ();
 sg13g2_fill_1 FILLER_60_2557 ();
 sg13g2_fill_2 FILLER_60_2562 ();
 sg13g2_fill_1 FILLER_60_2564 ();
 sg13g2_decap_8 FILLER_60_2569 ();
 sg13g2_decap_8 FILLER_60_2576 ();
 sg13g2_decap_8 FILLER_60_2583 ();
 sg13g2_decap_8 FILLER_60_2590 ();
 sg13g2_decap_8 FILLER_60_2597 ();
 sg13g2_decap_8 FILLER_60_2604 ();
 sg13g2_decap_8 FILLER_60_2611 ();
 sg13g2_decap_8 FILLER_60_2618 ();
 sg13g2_decap_8 FILLER_60_2625 ();
 sg13g2_decap_8 FILLER_60_2632 ();
 sg13g2_decap_8 FILLER_60_2639 ();
 sg13g2_decap_8 FILLER_60_2646 ();
 sg13g2_decap_8 FILLER_60_2653 ();
 sg13g2_decap_8 FILLER_60_2660 ();
 sg13g2_fill_2 FILLER_60_2667 ();
 sg13g2_fill_1 FILLER_60_2669 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_fill_2 FILLER_61_17 ();
 sg13g2_decap_4 FILLER_61_29 ();
 sg13g2_fill_2 FILLER_61_94 ();
 sg13g2_decap_4 FILLER_61_147 ();
 sg13g2_fill_1 FILLER_61_151 ();
 sg13g2_decap_4 FILLER_61_162 ();
 sg13g2_fill_1 FILLER_61_183 ();
 sg13g2_fill_1 FILLER_61_198 ();
 sg13g2_fill_2 FILLER_61_213 ();
 sg13g2_decap_8 FILLER_61_219 ();
 sg13g2_fill_2 FILLER_61_266 ();
 sg13g2_fill_1 FILLER_61_317 ();
 sg13g2_decap_8 FILLER_61_327 ();
 sg13g2_fill_1 FILLER_61_334 ();
 sg13g2_fill_2 FILLER_61_355 ();
 sg13g2_decap_8 FILLER_61_370 ();
 sg13g2_decap_8 FILLER_61_377 ();
 sg13g2_fill_1 FILLER_61_384 ();
 sg13g2_fill_1 FILLER_61_398 ();
 sg13g2_decap_4 FILLER_61_428 ();
 sg13g2_fill_1 FILLER_61_432 ();
 sg13g2_decap_4 FILLER_61_436 ();
 sg13g2_fill_1 FILLER_61_440 ();
 sg13g2_fill_1 FILLER_61_453 ();
 sg13g2_decap_8 FILLER_61_457 ();
 sg13g2_decap_4 FILLER_61_464 ();
 sg13g2_decap_4 FILLER_61_475 ();
 sg13g2_fill_1 FILLER_61_479 ();
 sg13g2_decap_4 FILLER_61_485 ();
 sg13g2_fill_2 FILLER_61_520 ();
 sg13g2_decap_8 FILLER_61_572 ();
 sg13g2_fill_2 FILLER_61_579 ();
 sg13g2_fill_1 FILLER_61_591 ();
 sg13g2_fill_2 FILLER_61_623 ();
 sg13g2_fill_1 FILLER_61_625 ();
 sg13g2_fill_1 FILLER_61_662 ();
 sg13g2_fill_1 FILLER_61_673 ();
 sg13g2_fill_1 FILLER_61_682 ();
 sg13g2_fill_1 FILLER_61_686 ();
 sg13g2_fill_1 FILLER_61_691 ();
 sg13g2_fill_1 FILLER_61_696 ();
 sg13g2_fill_2 FILLER_61_775 ();
 sg13g2_fill_2 FILLER_61_787 ();
 sg13g2_fill_2 FILLER_61_803 ();
 sg13g2_fill_2 FILLER_61_810 ();
 sg13g2_decap_4 FILLER_61_820 ();
 sg13g2_fill_1 FILLER_61_835 ();
 sg13g2_decap_8 FILLER_61_858 ();
 sg13g2_decap_4 FILLER_61_865 ();
 sg13g2_fill_2 FILLER_61_869 ();
 sg13g2_decap_8 FILLER_61_889 ();
 sg13g2_decap_8 FILLER_61_896 ();
 sg13g2_fill_1 FILLER_61_903 ();
 sg13g2_fill_1 FILLER_61_980 ();
 sg13g2_decap_4 FILLER_61_987 ();
 sg13g2_fill_2 FILLER_61_991 ();
 sg13g2_decap_8 FILLER_61_997 ();
 sg13g2_decap_4 FILLER_61_1004 ();
 sg13g2_fill_1 FILLER_61_1008 ();
 sg13g2_fill_1 FILLER_61_1012 ();
 sg13g2_decap_4 FILLER_61_1043 ();
 sg13g2_fill_2 FILLER_61_1131 ();
 sg13g2_fill_1 FILLER_61_1133 ();
 sg13g2_decap_8 FILLER_61_1143 ();
 sg13g2_decap_8 FILLER_61_1150 ();
 sg13g2_decap_8 FILLER_61_1157 ();
 sg13g2_decap_8 FILLER_61_1164 ();
 sg13g2_decap_8 FILLER_61_1171 ();
 sg13g2_decap_8 FILLER_61_1178 ();
 sg13g2_fill_1 FILLER_61_1185 ();
 sg13g2_decap_4 FILLER_61_1190 ();
 sg13g2_decap_4 FILLER_61_1203 ();
 sg13g2_fill_1 FILLER_61_1228 ();
 sg13g2_fill_1 FILLER_61_1234 ();
 sg13g2_fill_1 FILLER_61_1244 ();
 sg13g2_decap_8 FILLER_61_1249 ();
 sg13g2_decap_8 FILLER_61_1256 ();
 sg13g2_decap_4 FILLER_61_1263 ();
 sg13g2_fill_2 FILLER_61_1267 ();
 sg13g2_fill_1 FILLER_61_1312 ();
 sg13g2_decap_4 FILLER_61_1317 ();
 sg13g2_decap_8 FILLER_61_1326 ();
 sg13g2_fill_1 FILLER_61_1337 ();
 sg13g2_fill_1 FILLER_61_1350 ();
 sg13g2_fill_2 FILLER_61_1368 ();
 sg13g2_decap_4 FILLER_61_1374 ();
 sg13g2_fill_1 FILLER_61_1385 ();
 sg13g2_decap_8 FILLER_61_1403 ();
 sg13g2_decap_4 FILLER_61_1410 ();
 sg13g2_fill_1 FILLER_61_1414 ();
 sg13g2_decap_8 FILLER_61_1425 ();
 sg13g2_fill_2 FILLER_61_1432 ();
 sg13g2_fill_1 FILLER_61_1434 ();
 sg13g2_decap_4 FILLER_61_1439 ();
 sg13g2_fill_1 FILLER_61_1443 ();
 sg13g2_fill_2 FILLER_61_1449 ();
 sg13g2_decap_8 FILLER_61_1456 ();
 sg13g2_decap_4 FILLER_61_1463 ();
 sg13g2_fill_1 FILLER_61_1472 ();
 sg13g2_decap_8 FILLER_61_1506 ();
 sg13g2_decap_8 FILLER_61_1513 ();
 sg13g2_decap_4 FILLER_61_1520 ();
 sg13g2_fill_1 FILLER_61_1528 ();
 sg13g2_fill_2 FILLER_61_1536 ();
 sg13g2_fill_2 FILLER_61_1559 ();
 sg13g2_fill_1 FILLER_61_1561 ();
 sg13g2_decap_8 FILLER_61_1586 ();
 sg13g2_decap_8 FILLER_61_1593 ();
 sg13g2_fill_2 FILLER_61_1613 ();
 sg13g2_decap_4 FILLER_61_1641 ();
 sg13g2_decap_8 FILLER_61_1654 ();
 sg13g2_fill_1 FILLER_61_1709 ();
 sg13g2_fill_1 FILLER_61_1752 ();
 sg13g2_fill_1 FILLER_61_1769 ();
 sg13g2_fill_1 FILLER_61_1775 ();
 sg13g2_fill_1 FILLER_61_1787 ();
 sg13g2_fill_1 FILLER_61_1798 ();
 sg13g2_fill_2 FILLER_61_1807 ();
 sg13g2_fill_1 FILLER_61_1814 ();
 sg13g2_fill_1 FILLER_61_1820 ();
 sg13g2_fill_1 FILLER_61_1826 ();
 sg13g2_fill_1 FILLER_61_1832 ();
 sg13g2_fill_1 FILLER_61_1846 ();
 sg13g2_fill_1 FILLER_61_1852 ();
 sg13g2_fill_2 FILLER_61_1857 ();
 sg13g2_fill_1 FILLER_61_1864 ();
 sg13g2_decap_8 FILLER_61_1902 ();
 sg13g2_fill_1 FILLER_61_1960 ();
 sg13g2_fill_1 FILLER_61_1965 ();
 sg13g2_decap_8 FILLER_61_1971 ();
 sg13g2_fill_1 FILLER_61_1978 ();
 sg13g2_decap_8 FILLER_61_1984 ();
 sg13g2_fill_2 FILLER_61_1991 ();
 sg13g2_fill_1 FILLER_61_1998 ();
 sg13g2_fill_1 FILLER_61_2003 ();
 sg13g2_fill_1 FILLER_61_2008 ();
 sg13g2_fill_1 FILLER_61_2058 ();
 sg13g2_decap_8 FILLER_61_2063 ();
 sg13g2_fill_1 FILLER_61_2074 ();
 sg13g2_decap_8 FILLER_61_2083 ();
 sg13g2_decap_8 FILLER_61_2090 ();
 sg13g2_decap_8 FILLER_61_2097 ();
 sg13g2_decap_4 FILLER_61_2120 ();
 sg13g2_decap_8 FILLER_61_2128 ();
 sg13g2_fill_2 FILLER_61_2135 ();
 sg13g2_fill_1 FILLER_61_2153 ();
 sg13g2_fill_2 FILLER_61_2195 ();
 sg13g2_fill_1 FILLER_61_2244 ();
 sg13g2_fill_1 FILLER_61_2251 ();
 sg13g2_fill_1 FILLER_61_2257 ();
 sg13g2_fill_1 FILLER_61_2268 ();
 sg13g2_fill_1 FILLER_61_2273 ();
 sg13g2_decap_8 FILLER_61_2283 ();
 sg13g2_decap_8 FILLER_61_2295 ();
 sg13g2_fill_1 FILLER_61_2302 ();
 sg13g2_fill_1 FILLER_61_2310 ();
 sg13g2_fill_1 FILLER_61_2321 ();
 sg13g2_fill_2 FILLER_61_2328 ();
 sg13g2_decap_4 FILLER_61_2362 ();
 sg13g2_fill_2 FILLER_61_2366 ();
 sg13g2_fill_2 FILLER_61_2404 ();
 sg13g2_fill_1 FILLER_61_2406 ();
 sg13g2_fill_1 FILLER_61_2413 ();
 sg13g2_fill_2 FILLER_61_2419 ();
 sg13g2_decap_4 FILLER_61_2427 ();
 sg13g2_fill_2 FILLER_61_2431 ();
 sg13g2_fill_2 FILLER_61_2474 ();
 sg13g2_fill_1 FILLER_61_2476 ();
 sg13g2_fill_1 FILLER_61_2483 ();
 sg13g2_decap_8 FILLER_61_2530 ();
 sg13g2_decap_4 FILLER_61_2537 ();
 sg13g2_fill_1 FILLER_61_2541 ();
 sg13g2_decap_8 FILLER_61_2552 ();
 sg13g2_fill_1 FILLER_61_2559 ();
 sg13g2_decap_8 FILLER_61_2564 ();
 sg13g2_decap_8 FILLER_61_2571 ();
 sg13g2_decap_8 FILLER_61_2578 ();
 sg13g2_decap_8 FILLER_61_2585 ();
 sg13g2_decap_8 FILLER_61_2592 ();
 sg13g2_decap_8 FILLER_61_2599 ();
 sg13g2_decap_8 FILLER_61_2606 ();
 sg13g2_decap_8 FILLER_61_2613 ();
 sg13g2_decap_8 FILLER_61_2620 ();
 sg13g2_decap_8 FILLER_61_2627 ();
 sg13g2_decap_8 FILLER_61_2634 ();
 sg13g2_decap_8 FILLER_61_2641 ();
 sg13g2_decap_8 FILLER_61_2648 ();
 sg13g2_decap_8 FILLER_61_2655 ();
 sg13g2_decap_8 FILLER_61_2662 ();
 sg13g2_fill_1 FILLER_61_2669 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_4 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_37 ();
 sg13g2_fill_1 FILLER_62_58 ();
 sg13g2_fill_1 FILLER_62_121 ();
 sg13g2_fill_1 FILLER_62_127 ();
 sg13g2_decap_8 FILLER_62_163 ();
 sg13g2_decap_8 FILLER_62_170 ();
 sg13g2_decap_8 FILLER_62_177 ();
 sg13g2_decap_4 FILLER_62_184 ();
 sg13g2_decap_8 FILLER_62_214 ();
 sg13g2_fill_1 FILLER_62_221 ();
 sg13g2_fill_1 FILLER_62_226 ();
 sg13g2_fill_2 FILLER_62_238 ();
 sg13g2_fill_2 FILLER_62_244 ();
 sg13g2_fill_1 FILLER_62_251 ();
 sg13g2_fill_2 FILLER_62_257 ();
 sg13g2_fill_2 FILLER_62_277 ();
 sg13g2_fill_1 FILLER_62_279 ();
 sg13g2_decap_8 FILLER_62_322 ();
 sg13g2_fill_1 FILLER_62_329 ();
 sg13g2_decap_8 FILLER_62_335 ();
 sg13g2_fill_2 FILLER_62_342 ();
 sg13g2_fill_1 FILLER_62_344 ();
 sg13g2_decap_8 FILLER_62_355 ();
 sg13g2_decap_8 FILLER_62_362 ();
 sg13g2_fill_1 FILLER_62_369 ();
 sg13g2_fill_1 FILLER_62_413 ();
 sg13g2_fill_1 FILLER_62_417 ();
 sg13g2_fill_1 FILLER_62_422 ();
 sg13g2_fill_1 FILLER_62_428 ();
 sg13g2_fill_2 FILLER_62_434 ();
 sg13g2_fill_1 FILLER_62_436 ();
 sg13g2_fill_1 FILLER_62_442 ();
 sg13g2_fill_2 FILLER_62_481 ();
 sg13g2_fill_1 FILLER_62_497 ();
 sg13g2_decap_8 FILLER_62_512 ();
 sg13g2_decap_8 FILLER_62_519 ();
 sg13g2_decap_8 FILLER_62_526 ();
 sg13g2_decap_8 FILLER_62_533 ();
 sg13g2_decap_8 FILLER_62_540 ();
 sg13g2_fill_1 FILLER_62_551 ();
 sg13g2_fill_2 FILLER_62_569 ();
 sg13g2_fill_2 FILLER_62_575 ();
 sg13g2_fill_1 FILLER_62_577 ();
 sg13g2_fill_1 FILLER_62_588 ();
 sg13g2_fill_2 FILLER_62_615 ();
 sg13g2_fill_2 FILLER_62_643 ();
 sg13g2_fill_2 FILLER_62_671 ();
 sg13g2_fill_1 FILLER_62_673 ();
 sg13g2_decap_8 FILLER_62_700 ();
 sg13g2_decap_8 FILLER_62_707 ();
 sg13g2_decap_8 FILLER_62_714 ();
 sg13g2_fill_1 FILLER_62_726 ();
 sg13g2_fill_1 FILLER_62_731 ();
 sg13g2_decap_4 FILLER_62_771 ();
 sg13g2_fill_2 FILLER_62_775 ();
 sg13g2_fill_2 FILLER_62_786 ();
 sg13g2_fill_1 FILLER_62_788 ();
 sg13g2_fill_2 FILLER_62_796 ();
 sg13g2_fill_1 FILLER_62_825 ();
 sg13g2_fill_1 FILLER_62_832 ();
 sg13g2_fill_1 FILLER_62_839 ();
 sg13g2_fill_2 FILLER_62_844 ();
 sg13g2_fill_2 FILLER_62_851 ();
 sg13g2_fill_1 FILLER_62_853 ();
 sg13g2_fill_1 FILLER_62_862 ();
 sg13g2_fill_2 FILLER_62_867 ();
 sg13g2_fill_1 FILLER_62_877 ();
 sg13g2_fill_2 FILLER_62_884 ();
 sg13g2_fill_2 FILLER_62_891 ();
 sg13g2_fill_1 FILLER_62_893 ();
 sg13g2_fill_1 FILLER_62_902 ();
 sg13g2_decap_4 FILLER_62_913 ();
 sg13g2_fill_1 FILLER_62_921 ();
 sg13g2_fill_1 FILLER_62_934 ();
 sg13g2_fill_2 FILLER_62_940 ();
 sg13g2_decap_4 FILLER_62_947 ();
 sg13g2_fill_1 FILLER_62_951 ();
 sg13g2_fill_2 FILLER_62_962 ();
 sg13g2_fill_1 FILLER_62_964 ();
 sg13g2_fill_1 FILLER_62_970 ();
 sg13g2_fill_2 FILLER_62_987 ();
 sg13g2_fill_1 FILLER_62_989 ();
 sg13g2_fill_1 FILLER_62_1042 ();
 sg13g2_fill_1 FILLER_62_1054 ();
 sg13g2_fill_1 FILLER_62_1066 ();
 sg13g2_fill_1 FILLER_62_1072 ();
 sg13g2_fill_2 FILLER_62_1078 ();
 sg13g2_fill_1 FILLER_62_1092 ();
 sg13g2_fill_2 FILLER_62_1131 ();
 sg13g2_fill_1 FILLER_62_1133 ();
 sg13g2_decap_8 FILLER_62_1169 ();
 sg13g2_decap_4 FILLER_62_1176 ();
 sg13g2_fill_2 FILLER_62_1180 ();
 sg13g2_decap_4 FILLER_62_1195 ();
 sg13g2_fill_1 FILLER_62_1199 ();
 sg13g2_fill_2 FILLER_62_1243 ();
 sg13g2_decap_8 FILLER_62_1249 ();
 sg13g2_decap_8 FILLER_62_1256 ();
 sg13g2_decap_4 FILLER_62_1263 ();
 sg13g2_decap_8 FILLER_62_1273 ();
 sg13g2_decap_4 FILLER_62_1280 ();
 sg13g2_fill_2 FILLER_62_1284 ();
 sg13g2_fill_2 FILLER_62_1290 ();
 sg13g2_fill_1 FILLER_62_1292 ();
 sg13g2_decap_8 FILLER_62_1297 ();
 sg13g2_decap_4 FILLER_62_1304 ();
 sg13g2_fill_2 FILLER_62_1311 ();
 sg13g2_fill_1 FILLER_62_1317 ();
 sg13g2_decap_4 FILLER_62_1364 ();
 sg13g2_fill_2 FILLER_62_1368 ();
 sg13g2_fill_2 FILLER_62_1382 ();
 sg13g2_decap_8 FILLER_62_1400 ();
 sg13g2_decap_8 FILLER_62_1407 ();
 sg13g2_fill_2 FILLER_62_1414 ();
 sg13g2_fill_1 FILLER_62_1416 ();
 sg13g2_fill_2 FILLER_62_1421 ();
 sg13g2_fill_2 FILLER_62_1431 ();
 sg13g2_fill_2 FILLER_62_1443 ();
 sg13g2_decap_8 FILLER_62_1450 ();
 sg13g2_fill_2 FILLER_62_1457 ();
 sg13g2_fill_1 FILLER_62_1491 ();
 sg13g2_fill_1 FILLER_62_1500 ();
 sg13g2_fill_1 FILLER_62_1506 ();
 sg13g2_decap_8 FILLER_62_1515 ();
 sg13g2_fill_2 FILLER_62_1522 ();
 sg13g2_decap_4 FILLER_62_1571 ();
 sg13g2_fill_2 FILLER_62_1575 ();
 sg13g2_decap_4 FILLER_62_1581 ();
 sg13g2_fill_1 FILLER_62_1585 ();
 sg13g2_decap_8 FILLER_62_1612 ();
 sg13g2_fill_2 FILLER_62_1619 ();
 sg13g2_fill_1 FILLER_62_1621 ();
 sg13g2_fill_2 FILLER_62_1629 ();
 sg13g2_fill_2 FILLER_62_1664 ();
 sg13g2_fill_1 FILLER_62_1666 ();
 sg13g2_fill_2 FILLER_62_1691 ();
 sg13g2_fill_2 FILLER_62_1703 ();
 sg13g2_fill_1 FILLER_62_1714 ();
 sg13g2_fill_2 FILLER_62_1729 ();
 sg13g2_fill_2 FILLER_62_1740 ();
 sg13g2_fill_1 FILLER_62_1742 ();
 sg13g2_fill_2 FILLER_62_1748 ();
 sg13g2_fill_2 FILLER_62_1825 ();
 sg13g2_fill_1 FILLER_62_1844 ();
 sg13g2_fill_2 FILLER_62_1852 ();
 sg13g2_fill_1 FILLER_62_1880 ();
 sg13g2_fill_2 FILLER_62_1895 ();
 sg13g2_decap_8 FILLER_62_1901 ();
 sg13g2_decap_4 FILLER_62_1908 ();
 sg13g2_fill_2 FILLER_62_1923 ();
 sg13g2_decap_4 FILLER_62_1951 ();
 sg13g2_decap_4 FILLER_62_1959 ();
 sg13g2_fill_2 FILLER_62_1989 ();
 sg13g2_fill_1 FILLER_62_1991 ();
 sg13g2_decap_8 FILLER_62_1996 ();
 sg13g2_fill_2 FILLER_62_2003 ();
 sg13g2_fill_2 FILLER_62_2028 ();
 sg13g2_decap_4 FILLER_62_2080 ();
 sg13g2_fill_1 FILLER_62_2084 ();
 sg13g2_fill_1 FILLER_62_2111 ();
 sg13g2_fill_2 FILLER_62_2122 ();
 sg13g2_fill_2 FILLER_62_2132 ();
 sg13g2_fill_2 FILLER_62_2139 ();
 sg13g2_fill_1 FILLER_62_2147 ();
 sg13g2_fill_1 FILLER_62_2174 ();
 sg13g2_fill_1 FILLER_62_2220 ();
 sg13g2_fill_2 FILLER_62_2245 ();
 sg13g2_fill_2 FILLER_62_2286 ();
 sg13g2_fill_1 FILLER_62_2288 ();
 sg13g2_fill_1 FILLER_62_2294 ();
 sg13g2_fill_1 FILLER_62_2308 ();
 sg13g2_fill_2 FILLER_62_2331 ();
 sg13g2_decap_4 FILLER_62_2342 ();
 sg13g2_fill_2 FILLER_62_2346 ();
 sg13g2_fill_1 FILLER_62_2384 ();
 sg13g2_decap_8 FILLER_62_2389 ();
 sg13g2_decap_8 FILLER_62_2396 ();
 sg13g2_fill_1 FILLER_62_2403 ();
 sg13g2_fill_2 FILLER_62_2424 ();
 sg13g2_fill_1 FILLER_62_2426 ();
 sg13g2_decap_4 FILLER_62_2461 ();
 sg13g2_fill_2 FILLER_62_2465 ();
 sg13g2_fill_2 FILLER_62_2477 ();
 sg13g2_decap_4 FILLER_62_2528 ();
 sg13g2_decap_4 FILLER_62_2536 ();
 sg13g2_decap_8 FILLER_62_2576 ();
 sg13g2_decap_8 FILLER_62_2583 ();
 sg13g2_decap_8 FILLER_62_2590 ();
 sg13g2_decap_8 FILLER_62_2597 ();
 sg13g2_decap_8 FILLER_62_2604 ();
 sg13g2_decap_8 FILLER_62_2611 ();
 sg13g2_decap_8 FILLER_62_2618 ();
 sg13g2_decap_8 FILLER_62_2625 ();
 sg13g2_decap_8 FILLER_62_2632 ();
 sg13g2_decap_8 FILLER_62_2639 ();
 sg13g2_decap_8 FILLER_62_2646 ();
 sg13g2_decap_8 FILLER_62_2653 ();
 sg13g2_decap_8 FILLER_62_2660 ();
 sg13g2_fill_2 FILLER_62_2667 ();
 sg13g2_fill_1 FILLER_62_2669 ();
 sg13g2_fill_2 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_38 ();
 sg13g2_decap_4 FILLER_63_45 ();
 sg13g2_fill_2 FILLER_63_49 ();
 sg13g2_fill_2 FILLER_63_77 ();
 sg13g2_fill_1 FILLER_63_79 ();
 sg13g2_fill_1 FILLER_63_89 ();
 sg13g2_fill_1 FILLER_63_113 ();
 sg13g2_fill_2 FILLER_63_124 ();
 sg13g2_fill_1 FILLER_63_135 ();
 sg13g2_fill_1 FILLER_63_141 ();
 sg13g2_fill_2 FILLER_63_168 ();
 sg13g2_fill_1 FILLER_63_170 ();
 sg13g2_fill_1 FILLER_63_204 ();
 sg13g2_fill_2 FILLER_63_218 ();
 sg13g2_fill_1 FILLER_63_220 ();
 sg13g2_fill_2 FILLER_63_231 ();
 sg13g2_fill_1 FILLER_63_233 ();
 sg13g2_fill_2 FILLER_63_238 ();
 sg13g2_fill_1 FILLER_63_240 ();
 sg13g2_decap_8 FILLER_63_245 ();
 sg13g2_decap_4 FILLER_63_267 ();
 sg13g2_fill_1 FILLER_63_275 ();
 sg13g2_fill_1 FILLER_63_287 ();
 sg13g2_fill_2 FILLER_63_308 ();
 sg13g2_decap_4 FILLER_63_330 ();
 sg13g2_fill_2 FILLER_63_334 ();
 sg13g2_fill_1 FILLER_63_354 ();
 sg13g2_fill_2 FILLER_63_370 ();
 sg13g2_fill_1 FILLER_63_376 ();
 sg13g2_fill_1 FILLER_63_382 ();
 sg13g2_fill_2 FILLER_63_427 ();
 sg13g2_fill_1 FILLER_63_429 ();
 sg13g2_fill_2 FILLER_63_457 ();
 sg13g2_decap_8 FILLER_63_533 ();
 sg13g2_decap_8 FILLER_63_540 ();
 sg13g2_fill_2 FILLER_63_547 ();
 sg13g2_fill_1 FILLER_63_549 ();
 sg13g2_decap_8 FILLER_63_610 ();
 sg13g2_fill_2 FILLER_63_653 ();
 sg13g2_fill_1 FILLER_63_655 ();
 sg13g2_decap_4 FILLER_63_660 ();
 sg13g2_decap_8 FILLER_63_668 ();
 sg13g2_fill_1 FILLER_63_675 ();
 sg13g2_decap_8 FILLER_63_684 ();
 sg13g2_decap_8 FILLER_63_691 ();
 sg13g2_fill_2 FILLER_63_698 ();
 sg13g2_fill_1 FILLER_63_700 ();
 sg13g2_fill_1 FILLER_63_731 ();
 sg13g2_decap_8 FILLER_63_736 ();
 sg13g2_decap_8 FILLER_63_743 ();
 sg13g2_fill_1 FILLER_63_750 ();
 sg13g2_fill_1 FILLER_63_795 ();
 sg13g2_fill_2 FILLER_63_845 ();
 sg13g2_fill_2 FILLER_63_858 ();
 sg13g2_fill_1 FILLER_63_860 ();
 sg13g2_fill_1 FILLER_63_881 ();
 sg13g2_fill_1 FILLER_63_886 ();
 sg13g2_decap_4 FILLER_63_891 ();
 sg13g2_decap_8 FILLER_63_903 ();
 sg13g2_fill_1 FILLER_63_910 ();
 sg13g2_decap_4 FILLER_63_920 ();
 sg13g2_fill_2 FILLER_63_924 ();
 sg13g2_decap_4 FILLER_63_929 ();
 sg13g2_fill_1 FILLER_63_980 ();
 sg13g2_decap_8 FILLER_63_1040 ();
 sg13g2_decap_8 FILLER_63_1077 ();
 sg13g2_fill_1 FILLER_63_1084 ();
 sg13g2_fill_1 FILLER_63_1099 ();
 sg13g2_fill_1 FILLER_63_1110 ();
 sg13g2_fill_2 FILLER_63_1121 ();
 sg13g2_fill_1 FILLER_63_1123 ();
 sg13g2_decap_4 FILLER_63_1202 ();
 sg13g2_fill_1 FILLER_63_1206 ();
 sg13g2_decap_8 FILLER_63_1250 ();
 sg13g2_decap_8 FILLER_63_1257 ();
 sg13g2_decap_8 FILLER_63_1267 ();
 sg13g2_fill_1 FILLER_63_1274 ();
 sg13g2_fill_2 FILLER_63_1292 ();
 sg13g2_decap_8 FILLER_63_1312 ();
 sg13g2_decap_4 FILLER_63_1319 ();
 sg13g2_decap_8 FILLER_63_1347 ();
 sg13g2_decap_8 FILLER_63_1354 ();
 sg13g2_decap_8 FILLER_63_1361 ();
 sg13g2_fill_2 FILLER_63_1368 ();
 sg13g2_fill_1 FILLER_63_1370 ();
 sg13g2_fill_2 FILLER_63_1379 ();
 sg13g2_fill_1 FILLER_63_1388 ();
 sg13g2_decap_4 FILLER_63_1401 ();
 sg13g2_fill_2 FILLER_63_1405 ();
 sg13g2_fill_2 FILLER_63_1411 ();
 sg13g2_fill_1 FILLER_63_1423 ();
 sg13g2_fill_1 FILLER_63_1432 ();
 sg13g2_fill_1 FILLER_63_1445 ();
 sg13g2_decap_8 FILLER_63_1453 ();
 sg13g2_decap_4 FILLER_63_1460 ();
 sg13g2_fill_2 FILLER_63_1464 ();
 sg13g2_fill_2 FILLER_63_1480 ();
 sg13g2_decap_4 FILLER_63_1496 ();
 sg13g2_fill_1 FILLER_63_1505 ();
 sg13g2_fill_2 FILLER_63_1515 ();
 sg13g2_fill_2 FILLER_63_1525 ();
 sg13g2_fill_1 FILLER_63_1527 ();
 sg13g2_fill_2 FILLER_63_1532 ();
 sg13g2_fill_2 FILLER_63_1538 ();
 sg13g2_fill_1 FILLER_63_1548 ();
 sg13g2_fill_2 FILLER_63_1567 ();
 sg13g2_fill_1 FILLER_63_1569 ();
 sg13g2_decap_4 FILLER_63_1612 ();
 sg13g2_decap_8 FILLER_63_1647 ();
 sg13g2_decap_8 FILLER_63_1654 ();
 sg13g2_decap_8 FILLER_63_1661 ();
 sg13g2_fill_2 FILLER_63_1668 ();
 sg13g2_fill_1 FILLER_63_1670 ();
 sg13g2_fill_1 FILLER_63_1675 ();
 sg13g2_fill_2 FILLER_63_1681 ();
 sg13g2_fill_2 FILLER_63_1687 ();
 sg13g2_fill_1 FILLER_63_1689 ();
 sg13g2_decap_8 FILLER_63_1695 ();
 sg13g2_decap_8 FILLER_63_1702 ();
 sg13g2_fill_2 FILLER_63_1709 ();
 sg13g2_fill_1 FILLER_63_1721 ();
 sg13g2_fill_1 FILLER_63_1726 ();
 sg13g2_fill_2 FILLER_63_1737 ();
 sg13g2_fill_1 FILLER_63_1739 ();
 sg13g2_fill_2 FILLER_63_1745 ();
 sg13g2_fill_2 FILLER_63_1757 ();
 sg13g2_fill_1 FILLER_63_1773 ();
 sg13g2_fill_2 FILLER_63_1787 ();
 sg13g2_fill_1 FILLER_63_1806 ();
 sg13g2_fill_2 FILLER_63_1824 ();
 sg13g2_fill_2 FILLER_63_1846 ();
 sg13g2_fill_1 FILLER_63_1865 ();
 sg13g2_fill_2 FILLER_63_1877 ();
 sg13g2_fill_2 FILLER_63_1912 ();
 sg13g2_fill_1 FILLER_63_1940 ();
 sg13g2_fill_2 FILLER_63_1949 ();
 sg13g2_fill_1 FILLER_63_1967 ();
 sg13g2_fill_2 FILLER_63_1977 ();
 sg13g2_fill_1 FILLER_63_1979 ();
 sg13g2_decap_4 FILLER_63_2000 ();
 sg13g2_fill_1 FILLER_63_2070 ();
 sg13g2_decap_8 FILLER_63_2076 ();
 sg13g2_decap_8 FILLER_63_2083 ();
 sg13g2_fill_2 FILLER_63_2090 ();
 sg13g2_decap_8 FILLER_63_2139 ();
 sg13g2_decap_4 FILLER_63_2146 ();
 sg13g2_fill_2 FILLER_63_2240 ();
 sg13g2_fill_1 FILLER_63_2252 ();
 sg13g2_fill_1 FILLER_63_2279 ();
 sg13g2_fill_2 FILLER_63_2286 ();
 sg13g2_decap_4 FILLER_63_2331 ();
 sg13g2_decap_8 FILLER_63_2339 ();
 sg13g2_decap_8 FILLER_63_2346 ();
 sg13g2_fill_2 FILLER_63_2353 ();
 sg13g2_fill_1 FILLER_63_2355 ();
 sg13g2_decap_8 FILLER_63_2371 ();
 sg13g2_decap_4 FILLER_63_2384 ();
 sg13g2_fill_2 FILLER_63_2388 ();
 sg13g2_fill_1 FILLER_63_2420 ();
 sg13g2_fill_2 FILLER_63_2455 ();
 sg13g2_fill_1 FILLER_63_2462 ();
 sg13g2_decap_4 FILLER_63_2466 ();
 sg13g2_fill_2 FILLER_63_2470 ();
 sg13g2_fill_2 FILLER_63_2478 ();
 sg13g2_fill_1 FILLER_63_2506 ();
 sg13g2_fill_2 FILLER_63_2579 ();
 sg13g2_decap_8 FILLER_63_2585 ();
 sg13g2_decap_8 FILLER_63_2592 ();
 sg13g2_decap_8 FILLER_63_2599 ();
 sg13g2_decap_8 FILLER_63_2606 ();
 sg13g2_decap_8 FILLER_63_2613 ();
 sg13g2_decap_8 FILLER_63_2620 ();
 sg13g2_decap_8 FILLER_63_2627 ();
 sg13g2_decap_8 FILLER_63_2634 ();
 sg13g2_decap_8 FILLER_63_2641 ();
 sg13g2_decap_8 FILLER_63_2648 ();
 sg13g2_decap_8 FILLER_63_2655 ();
 sg13g2_decap_8 FILLER_63_2662 ();
 sg13g2_fill_1 FILLER_63_2669 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_26 ();
 sg13g2_decap_8 FILLER_64_33 ();
 sg13g2_decap_8 FILLER_64_40 ();
 sg13g2_decap_8 FILLER_64_47 ();
 sg13g2_fill_1 FILLER_64_54 ();
 sg13g2_fill_1 FILLER_64_120 ();
 sg13g2_fill_1 FILLER_64_134 ();
 sg13g2_fill_1 FILLER_64_140 ();
 sg13g2_decap_8 FILLER_64_153 ();
 sg13g2_decap_4 FILLER_64_160 ();
 sg13g2_fill_1 FILLER_64_164 ();
 sg13g2_decap_4 FILLER_64_216 ();
 sg13g2_fill_2 FILLER_64_233 ();
 sg13g2_fill_1 FILLER_64_235 ();
 sg13g2_decap_8 FILLER_64_245 ();
 sg13g2_decap_8 FILLER_64_252 ();
 sg13g2_fill_2 FILLER_64_259 ();
 sg13g2_decap_4 FILLER_64_267 ();
 sg13g2_fill_1 FILLER_64_271 ();
 sg13g2_fill_1 FILLER_64_281 ();
 sg13g2_fill_1 FILLER_64_326 ();
 sg13g2_fill_1 FILLER_64_332 ();
 sg13g2_fill_1 FILLER_64_338 ();
 sg13g2_fill_1 FILLER_64_344 ();
 sg13g2_fill_2 FILLER_64_395 ();
 sg13g2_fill_2 FILLER_64_431 ();
 sg13g2_decap_4 FILLER_64_437 ();
 sg13g2_fill_1 FILLER_64_441 ();
 sg13g2_fill_1 FILLER_64_454 ();
 sg13g2_fill_1 FILLER_64_497 ();
 sg13g2_decap_4 FILLER_64_539 ();
 sg13g2_decap_8 FILLER_64_573 ();
 sg13g2_decap_4 FILLER_64_580 ();
 sg13g2_fill_1 FILLER_64_584 ();
 sg13g2_decap_8 FILLER_64_589 ();
 sg13g2_fill_1 FILLER_64_596 ();
 sg13g2_decap_4 FILLER_64_601 ();
 sg13g2_decap_8 FILLER_64_610 ();
 sg13g2_decap_8 FILLER_64_617 ();
 sg13g2_fill_1 FILLER_64_624 ();
 sg13g2_fill_2 FILLER_64_656 ();
 sg13g2_fill_2 FILLER_64_662 ();
 sg13g2_decap_4 FILLER_64_668 ();
 sg13g2_fill_1 FILLER_64_672 ();
 sg13g2_decap_8 FILLER_64_686 ();
 sg13g2_decap_8 FILLER_64_733 ();
 sg13g2_decap_4 FILLER_64_740 ();
 sg13g2_fill_2 FILLER_64_756 ();
 sg13g2_decap_4 FILLER_64_762 ();
 sg13g2_fill_1 FILLER_64_766 ();
 sg13g2_fill_2 FILLER_64_777 ();
 sg13g2_fill_1 FILLER_64_779 ();
 sg13g2_fill_1 FILLER_64_830 ();
 sg13g2_decap_8 FILLER_64_864 ();
 sg13g2_fill_2 FILLER_64_871 ();
 sg13g2_decap_8 FILLER_64_886 ();
 sg13g2_decap_4 FILLER_64_893 ();
 sg13g2_fill_2 FILLER_64_915 ();
 sg13g2_fill_1 FILLER_64_969 ();
 sg13g2_decap_4 FILLER_64_1002 ();
 sg13g2_fill_2 FILLER_64_1006 ();
 sg13g2_decap_8 FILLER_64_1012 ();
 sg13g2_fill_2 FILLER_64_1019 ();
 sg13g2_fill_2 FILLER_64_1029 ();
 sg13g2_fill_1 FILLER_64_1050 ();
 sg13g2_fill_1 FILLER_64_1059 ();
 sg13g2_fill_1 FILLER_64_1082 ();
 sg13g2_fill_2 FILLER_64_1087 ();
 sg13g2_fill_1 FILLER_64_1089 ();
 sg13g2_decap_8 FILLER_64_1095 ();
 sg13g2_decap_4 FILLER_64_1102 ();
 sg13g2_fill_1 FILLER_64_1141 ();
 sg13g2_fill_1 FILLER_64_1178 ();
 sg13g2_fill_1 FILLER_64_1196 ();
 sg13g2_fill_2 FILLER_64_1229 ();
 sg13g2_fill_2 FILLER_64_1237 ();
 sg13g2_decap_8 FILLER_64_1247 ();
 sg13g2_decap_8 FILLER_64_1254 ();
 sg13g2_fill_2 FILLER_64_1261 ();
 sg13g2_fill_2 FILLER_64_1289 ();
 sg13g2_fill_1 FILLER_64_1299 ();
 sg13g2_fill_1 FILLER_64_1308 ();
 sg13g2_decap_4 FILLER_64_1313 ();
 sg13g2_fill_1 FILLER_64_1317 ();
 sg13g2_decap_8 FILLER_64_1323 ();
 sg13g2_fill_1 FILLER_64_1330 ();
 sg13g2_decap_4 FILLER_64_1347 ();
 sg13g2_fill_2 FILLER_64_1351 ();
 sg13g2_fill_1 FILLER_64_1365 ();
 sg13g2_fill_1 FILLER_64_1405 ();
 sg13g2_fill_1 FILLER_64_1415 ();
 sg13g2_decap_8 FILLER_64_1421 ();
 sg13g2_fill_1 FILLER_64_1432 ();
 sg13g2_fill_2 FILLER_64_1438 ();
 sg13g2_fill_1 FILLER_64_1440 ();
 sg13g2_fill_2 FILLER_64_1446 ();
 sg13g2_decap_8 FILLER_64_1452 ();
 sg13g2_decap_4 FILLER_64_1459 ();
 sg13g2_fill_1 FILLER_64_1463 ();
 sg13g2_fill_2 FILLER_64_1481 ();
 sg13g2_fill_1 FILLER_64_1499 ();
 sg13g2_fill_1 FILLER_64_1516 ();
 sg13g2_decap_8 FILLER_64_1568 ();
 sg13g2_decap_8 FILLER_64_1575 ();
 sg13g2_decap_8 FILLER_64_1582 ();
 sg13g2_decap_4 FILLER_64_1589 ();
 sg13g2_fill_1 FILLER_64_1593 ();
 sg13g2_decap_8 FILLER_64_1631 ();
 sg13g2_decap_4 FILLER_64_1651 ();
 sg13g2_decap_8 FILLER_64_1665 ();
 sg13g2_fill_2 FILLER_64_1682 ();
 sg13g2_decap_4 FILLER_64_1689 ();
 sg13g2_fill_1 FILLER_64_1693 ();
 sg13g2_fill_2 FILLER_64_1699 ();
 sg13g2_fill_1 FILLER_64_1701 ();
 sg13g2_fill_1 FILLER_64_1708 ();
 sg13g2_fill_1 FILLER_64_1734 ();
 sg13g2_fill_2 FILLER_64_1740 ();
 sg13g2_fill_1 FILLER_64_1747 ();
 sg13g2_fill_1 FILLER_64_1819 ();
 sg13g2_fill_2 FILLER_64_1857 ();
 sg13g2_fill_1 FILLER_64_1887 ();
 sg13g2_fill_2 FILLER_64_1914 ();
 sg13g2_fill_1 FILLER_64_1920 ();
 sg13g2_fill_2 FILLER_64_1947 ();
 sg13g2_fill_2 FILLER_64_1958 ();
 sg13g2_fill_1 FILLER_64_1964 ();
 sg13g2_fill_1 FILLER_64_1970 ();
 sg13g2_fill_1 FILLER_64_2005 ();
 sg13g2_fill_1 FILLER_64_2020 ();
 sg13g2_fill_2 FILLER_64_2061 ();
 sg13g2_fill_2 FILLER_64_2069 ();
 sg13g2_fill_1 FILLER_64_2071 ();
 sg13g2_decap_8 FILLER_64_2078 ();
 sg13g2_decap_8 FILLER_64_2085 ();
 sg13g2_decap_8 FILLER_64_2092 ();
 sg13g2_fill_2 FILLER_64_2104 ();
 sg13g2_decap_4 FILLER_64_2124 ();
 sg13g2_fill_2 FILLER_64_2128 ();
 sg13g2_decap_8 FILLER_64_2140 ();
 sg13g2_decap_4 FILLER_64_2152 ();
 sg13g2_fill_2 FILLER_64_2170 ();
 sg13g2_fill_1 FILLER_64_2172 ();
 sg13g2_fill_2 FILLER_64_2178 ();
 sg13g2_fill_2 FILLER_64_2209 ();
 sg13g2_fill_1 FILLER_64_2273 ();
 sg13g2_fill_2 FILLER_64_2302 ();
 sg13g2_fill_1 FILLER_64_2304 ();
 sg13g2_fill_1 FILLER_64_2343 ();
 sg13g2_decap_4 FILLER_64_2387 ();
 sg13g2_fill_1 FILLER_64_2391 ();
 sg13g2_fill_2 FILLER_64_2396 ();
 sg13g2_fill_1 FILLER_64_2403 ();
 sg13g2_fill_1 FILLER_64_2414 ();
 sg13g2_fill_1 FILLER_64_2420 ();
 sg13g2_fill_2 FILLER_64_2431 ();
 sg13g2_fill_1 FILLER_64_2443 ();
 sg13g2_fill_2 FILLER_64_2449 ();
 sg13g2_fill_2 FILLER_64_2455 ();
 sg13g2_fill_1 FILLER_64_2457 ();
 sg13g2_fill_1 FILLER_64_2464 ();
 sg13g2_decap_4 FILLER_64_2484 ();
 sg13g2_fill_1 FILLER_64_2488 ();
 sg13g2_decap_8 FILLER_64_2493 ();
 sg13g2_decap_8 FILLER_64_2500 ();
 sg13g2_decap_4 FILLER_64_2507 ();
 sg13g2_fill_2 FILLER_64_2511 ();
 sg13g2_decap_8 FILLER_64_2517 ();
 sg13g2_decap_8 FILLER_64_2524 ();
 sg13g2_fill_2 FILLER_64_2531 ();
 sg13g2_decap_8 FILLER_64_2543 ();
 sg13g2_fill_2 FILLER_64_2550 ();
 sg13g2_fill_1 FILLER_64_2552 ();
 sg13g2_decap_8 FILLER_64_2579 ();
 sg13g2_decap_8 FILLER_64_2586 ();
 sg13g2_decap_8 FILLER_64_2593 ();
 sg13g2_decap_8 FILLER_64_2600 ();
 sg13g2_decap_8 FILLER_64_2607 ();
 sg13g2_decap_8 FILLER_64_2614 ();
 sg13g2_decap_8 FILLER_64_2621 ();
 sg13g2_decap_8 FILLER_64_2628 ();
 sg13g2_decap_8 FILLER_64_2635 ();
 sg13g2_decap_8 FILLER_64_2642 ();
 sg13g2_decap_8 FILLER_64_2649 ();
 sg13g2_decap_8 FILLER_64_2656 ();
 sg13g2_decap_8 FILLER_64_2663 ();
 sg13g2_decap_4 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_4 ();
 sg13g2_decap_4 FILLER_65_15 ();
 sg13g2_fill_1 FILLER_65_45 ();
 sg13g2_fill_2 FILLER_65_82 ();
 sg13g2_fill_1 FILLER_65_84 ();
 sg13g2_fill_1 FILLER_65_89 ();
 sg13g2_fill_1 FILLER_65_116 ();
 sg13g2_fill_2 FILLER_65_123 ();
 sg13g2_fill_1 FILLER_65_156 ();
 sg13g2_fill_1 FILLER_65_163 ();
 sg13g2_decap_4 FILLER_65_172 ();
 sg13g2_fill_2 FILLER_65_227 ();
 sg13g2_fill_1 FILLER_65_229 ();
 sg13g2_fill_1 FILLER_65_240 ();
 sg13g2_fill_1 FILLER_65_277 ();
 sg13g2_fill_1 FILLER_65_339 ();
 sg13g2_decap_4 FILLER_65_345 ();
 sg13g2_fill_2 FILLER_65_349 ();
 sg13g2_fill_2 FILLER_65_357 ();
 sg13g2_decap_4 FILLER_65_374 ();
 sg13g2_fill_1 FILLER_65_382 ();
 sg13g2_fill_1 FILLER_65_392 ();
 sg13g2_decap_8 FILLER_65_405 ();
 sg13g2_decap_8 FILLER_65_412 ();
 sg13g2_decap_8 FILLER_65_419 ();
 sg13g2_fill_1 FILLER_65_426 ();
 sg13g2_fill_2 FILLER_65_435 ();
 sg13g2_decap_8 FILLER_65_446 ();
 sg13g2_fill_1 FILLER_65_453 ();
 sg13g2_fill_2 FILLER_65_471 ();
 sg13g2_fill_1 FILLER_65_473 ();
 sg13g2_decap_8 FILLER_65_482 ();
 sg13g2_decap_4 FILLER_65_489 ();
 sg13g2_fill_2 FILLER_65_508 ();
 sg13g2_fill_2 FILLER_65_514 ();
 sg13g2_decap_4 FILLER_65_526 ();
 sg13g2_fill_2 FILLER_65_530 ();
 sg13g2_fill_2 FILLER_65_536 ();
 sg13g2_fill_2 FILLER_65_542 ();
 sg13g2_fill_1 FILLER_65_544 ();
 sg13g2_decap_4 FILLER_65_548 ();
 sg13g2_fill_2 FILLER_65_552 ();
 sg13g2_decap_8 FILLER_65_561 ();
 sg13g2_decap_8 FILLER_65_568 ();
 sg13g2_fill_1 FILLER_65_582 ();
 sg13g2_decap_8 FILLER_65_587 ();
 sg13g2_decap_8 FILLER_65_594 ();
 sg13g2_fill_2 FILLER_65_601 ();
 sg13g2_decap_8 FILLER_65_608 ();
 sg13g2_decap_4 FILLER_65_615 ();
 sg13g2_fill_1 FILLER_65_619 ();
 sg13g2_decap_8 FILLER_65_624 ();
 sg13g2_decap_4 FILLER_65_631 ();
 sg13g2_fill_2 FILLER_65_641 ();
 sg13g2_fill_1 FILLER_65_643 ();
 sg13g2_fill_1 FILLER_65_649 ();
 sg13g2_fill_2 FILLER_65_654 ();
 sg13g2_fill_1 FILLER_65_656 ();
 sg13g2_fill_1 FILLER_65_662 ();
 sg13g2_fill_2 FILLER_65_668 ();
 sg13g2_fill_2 FILLER_65_713 ();
 sg13g2_fill_2 FILLER_65_727 ();
 sg13g2_fill_2 FILLER_65_737 ();
 sg13g2_fill_1 FILLER_65_739 ();
 sg13g2_fill_2 FILLER_65_753 ();
 sg13g2_fill_1 FILLER_65_759 ();
 sg13g2_decap_8 FILLER_65_765 ();
 sg13g2_decap_8 FILLER_65_772 ();
 sg13g2_decap_8 FILLER_65_779 ();
 sg13g2_decap_4 FILLER_65_786 ();
 sg13g2_decap_4 FILLER_65_794 ();
 sg13g2_fill_1 FILLER_65_798 ();
 sg13g2_fill_1 FILLER_65_803 ();
 sg13g2_fill_1 FILLER_65_834 ();
 sg13g2_fill_1 FILLER_65_843 ();
 sg13g2_fill_1 FILLER_65_870 ();
 sg13g2_fill_2 FILLER_65_876 ();
 sg13g2_fill_1 FILLER_65_883 ();
 sg13g2_fill_2 FILLER_65_888 ();
 sg13g2_fill_1 FILLER_65_905 ();
 sg13g2_decap_8 FILLER_65_1010 ();
 sg13g2_decap_8 FILLER_65_1017 ();
 sg13g2_decap_8 FILLER_65_1024 ();
 sg13g2_fill_2 FILLER_65_1069 ();
 sg13g2_fill_2 FILLER_65_1092 ();
 sg13g2_fill_2 FILLER_65_1100 ();
 sg13g2_fill_2 FILLER_65_1128 ();
 sg13g2_decap_4 FILLER_65_1142 ();
 sg13g2_decap_4 FILLER_65_1152 ();
 sg13g2_fill_1 FILLER_65_1160 ();
 sg13g2_fill_1 FILLER_65_1168 ();
 sg13g2_fill_1 FILLER_65_1173 ();
 sg13g2_fill_1 FILLER_65_1217 ();
 sg13g2_decap_8 FILLER_65_1245 ();
 sg13g2_decap_4 FILLER_65_1252 ();
 sg13g2_fill_1 FILLER_65_1292 ();
 sg13g2_fill_2 FILLER_65_1306 ();
 sg13g2_decap_4 FILLER_65_1313 ();
 sg13g2_decap_8 FILLER_65_1321 ();
 sg13g2_decap_4 FILLER_65_1328 ();
 sg13g2_fill_1 FILLER_65_1332 ();
 sg13g2_decap_8 FILLER_65_1342 ();
 sg13g2_decap_4 FILLER_65_1349 ();
 sg13g2_fill_1 FILLER_65_1364 ();
 sg13g2_fill_2 FILLER_65_1375 ();
 sg13g2_fill_1 FILLER_65_1387 ();
 sg13g2_fill_1 FILLER_65_1405 ();
 sg13g2_decap_4 FILLER_65_1423 ();
 sg13g2_fill_2 FILLER_65_1427 ();
 sg13g2_fill_2 FILLER_65_1438 ();
 sg13g2_decap_8 FILLER_65_1445 ();
 sg13g2_decap_8 FILLER_65_1452 ();
 sg13g2_fill_1 FILLER_65_1459 ();
 sg13g2_decap_4 FILLER_65_1464 ();
 sg13g2_decap_4 FILLER_65_1472 ();
 sg13g2_decap_4 FILLER_65_1493 ();
 sg13g2_fill_1 FILLER_65_1497 ();
 sg13g2_decap_4 FILLER_65_1511 ();
 sg13g2_fill_1 FILLER_65_1515 ();
 sg13g2_decap_4 FILLER_65_1530 ();
 sg13g2_fill_1 FILLER_65_1555 ();
 sg13g2_decap_8 FILLER_65_1560 ();
 sg13g2_decap_8 FILLER_65_1567 ();
 sg13g2_decap_8 FILLER_65_1574 ();
 sg13g2_decap_8 FILLER_65_1581 ();
 sg13g2_decap_4 FILLER_65_1588 ();
 sg13g2_fill_2 FILLER_65_1592 ();
 sg13g2_decap_8 FILLER_65_1598 ();
 sg13g2_decap_8 FILLER_65_1605 ();
 sg13g2_decap_8 FILLER_65_1621 ();
 sg13g2_decap_8 FILLER_65_1661 ();
 sg13g2_fill_1 FILLER_65_1668 ();
 sg13g2_fill_1 FILLER_65_1673 ();
 sg13g2_fill_2 FILLER_65_1697 ();
 sg13g2_fill_1 FILLER_65_1720 ();
 sg13g2_fill_2 FILLER_65_1783 ();
 sg13g2_fill_1 FILLER_65_1821 ();
 sg13g2_fill_2 FILLER_65_1843 ();
 sg13g2_fill_1 FILLER_65_1872 ();
 sg13g2_fill_2 FILLER_65_1880 ();
 sg13g2_fill_2 FILLER_65_1940 ();
 sg13g2_fill_1 FILLER_65_1948 ();
 sg13g2_fill_2 FILLER_65_1993 ();
 sg13g2_fill_1 FILLER_65_2009 ();
 sg13g2_fill_2 FILLER_65_2015 ();
 sg13g2_fill_1 FILLER_65_2063 ();
 sg13g2_decap_8 FILLER_65_2095 ();
 sg13g2_decap_4 FILLER_65_2107 ();
 sg13g2_fill_1 FILLER_65_2111 ();
 sg13g2_decap_4 FILLER_65_2126 ();
 sg13g2_decap_4 FILLER_65_2145 ();
 sg13g2_fill_1 FILLER_65_2149 ();
 sg13g2_fill_2 FILLER_65_2186 ();
 sg13g2_fill_2 FILLER_65_2191 ();
 sg13g2_fill_2 FILLER_65_2237 ();
 sg13g2_fill_1 FILLER_65_2239 ();
 sg13g2_fill_2 FILLER_65_2246 ();
 sg13g2_fill_1 FILLER_65_2248 ();
 sg13g2_fill_2 FILLER_65_2253 ();
 sg13g2_fill_1 FILLER_65_2255 ();
 sg13g2_fill_2 FILLER_65_2260 ();
 sg13g2_fill_2 FILLER_65_2278 ();
 sg13g2_fill_2 FILLER_65_2285 ();
 sg13g2_decap_4 FILLER_65_2292 ();
 sg13g2_fill_2 FILLER_65_2296 ();
 sg13g2_fill_2 FILLER_65_2303 ();
 sg13g2_fill_1 FILLER_65_2311 ();
 sg13g2_fill_2 FILLER_65_2317 ();
 sg13g2_decap_4 FILLER_65_2328 ();
 sg13g2_fill_1 FILLER_65_2332 ();
 sg13g2_decap_8 FILLER_65_2363 ();
 sg13g2_fill_1 FILLER_65_2370 ();
 sg13g2_fill_2 FILLER_65_2409 ();
 sg13g2_decap_4 FILLER_65_2415 ();
 sg13g2_fill_2 FILLER_65_2419 ();
 sg13g2_fill_1 FILLER_65_2426 ();
 sg13g2_decap_8 FILLER_65_2431 ();
 sg13g2_decap_8 FILLER_65_2438 ();
 sg13g2_decap_4 FILLER_65_2445 ();
 sg13g2_fill_2 FILLER_65_2476 ();
 sg13g2_fill_1 FILLER_65_2478 ();
 sg13g2_decap_8 FILLER_65_2489 ();
 sg13g2_decap_4 FILLER_65_2532 ();
 sg13g2_fill_2 FILLER_65_2536 ();
 sg13g2_decap_8 FILLER_65_2552 ();
 sg13g2_decap_8 FILLER_65_2559 ();
 sg13g2_decap_8 FILLER_65_2566 ();
 sg13g2_decap_8 FILLER_65_2573 ();
 sg13g2_decap_8 FILLER_65_2580 ();
 sg13g2_decap_8 FILLER_65_2587 ();
 sg13g2_decap_8 FILLER_65_2594 ();
 sg13g2_decap_8 FILLER_65_2601 ();
 sg13g2_decap_8 FILLER_65_2608 ();
 sg13g2_decap_8 FILLER_65_2615 ();
 sg13g2_decap_8 FILLER_65_2622 ();
 sg13g2_decap_8 FILLER_65_2629 ();
 sg13g2_decap_8 FILLER_65_2636 ();
 sg13g2_decap_8 FILLER_65_2643 ();
 sg13g2_decap_8 FILLER_65_2650 ();
 sg13g2_decap_8 FILLER_65_2657 ();
 sg13g2_decap_4 FILLER_65_2664 ();
 sg13g2_fill_2 FILLER_65_2668 ();
 sg13g2_decap_4 FILLER_66_0 ();
 sg13g2_fill_1 FILLER_66_4 ();
 sg13g2_decap_8 FILLER_66_19 ();
 sg13g2_fill_1 FILLER_66_26 ();
 sg13g2_decap_4 FILLER_66_31 ();
 sg13g2_fill_1 FILLER_66_35 ();
 sg13g2_fill_1 FILLER_66_46 ();
 sg13g2_decap_8 FILLER_66_73 ();
 sg13g2_fill_2 FILLER_66_80 ();
 sg13g2_fill_1 FILLER_66_86 ();
 sg13g2_fill_2 FILLER_66_113 ();
 sg13g2_fill_1 FILLER_66_136 ();
 sg13g2_fill_1 FILLER_66_156 ();
 sg13g2_fill_2 FILLER_66_161 ();
 sg13g2_decap_4 FILLER_66_173 ();
 sg13g2_fill_1 FILLER_66_217 ();
 sg13g2_fill_1 FILLER_66_223 ();
 sg13g2_decap_8 FILLER_66_264 ();
 sg13g2_fill_1 FILLER_66_271 ();
 sg13g2_fill_2 FILLER_66_277 ();
 sg13g2_fill_1 FILLER_66_279 ();
 sg13g2_fill_1 FILLER_66_286 ();
 sg13g2_fill_1 FILLER_66_293 ();
 sg13g2_fill_2 FILLER_66_298 ();
 sg13g2_fill_2 FILLER_66_308 ();
 sg13g2_fill_2 FILLER_66_315 ();
 sg13g2_fill_1 FILLER_66_322 ();
 sg13g2_fill_2 FILLER_66_336 ();
 sg13g2_decap_4 FILLER_66_354 ();
 sg13g2_fill_1 FILLER_66_358 ();
 sg13g2_decap_8 FILLER_66_365 ();
 sg13g2_fill_2 FILLER_66_372 ();
 sg13g2_fill_1 FILLER_66_374 ();
 sg13g2_fill_1 FILLER_66_406 ();
 sg13g2_decap_8 FILLER_66_411 ();
 sg13g2_decap_8 FILLER_66_418 ();
 sg13g2_fill_2 FILLER_66_425 ();
 sg13g2_decap_4 FILLER_66_491 ();
 sg13g2_fill_1 FILLER_66_501 ();
 sg13g2_fill_1 FILLER_66_575 ();
 sg13g2_fill_2 FILLER_66_609 ();
 sg13g2_fill_2 FILLER_66_617 ();
 sg13g2_fill_1 FILLER_66_619 ();
 sg13g2_fill_2 FILLER_66_629 ();
 sg13g2_fill_2 FILLER_66_657 ();
 sg13g2_fill_1 FILLER_66_670 ();
 sg13g2_fill_1 FILLER_66_689 ();
 sg13g2_fill_1 FILLER_66_701 ();
 sg13g2_fill_1 FILLER_66_711 ();
 sg13g2_fill_2 FILLER_66_722 ();
 sg13g2_fill_1 FILLER_66_724 ();
 sg13g2_fill_2 FILLER_66_750 ();
 sg13g2_decap_4 FILLER_66_788 ();
 sg13g2_fill_1 FILLER_66_796 ();
 sg13g2_fill_2 FILLER_66_822 ();
 sg13g2_fill_2 FILLER_66_833 ();
 sg13g2_fill_2 FILLER_66_853 ();
 sg13g2_fill_1 FILLER_66_875 ();
 sg13g2_fill_1 FILLER_66_894 ();
 sg13g2_fill_2 FILLER_66_899 ();
 sg13g2_decap_4 FILLER_66_909 ();
 sg13g2_fill_2 FILLER_66_913 ();
 sg13g2_decap_4 FILLER_66_935 ();
 sg13g2_fill_2 FILLER_66_939 ();
 sg13g2_fill_2 FILLER_66_945 ();
 sg13g2_decap_4 FILLER_66_951 ();
 sg13g2_decap_8 FILLER_66_1003 ();
 sg13g2_fill_2 FILLER_66_1010 ();
 sg13g2_fill_1 FILLER_66_1012 ();
 sg13g2_fill_1 FILLER_66_1038 ();
 sg13g2_fill_2 FILLER_66_1086 ();
 sg13g2_fill_2 FILLER_66_1097 ();
 sg13g2_fill_1 FILLER_66_1099 ();
 sg13g2_decap_8 FILLER_66_1135 ();
 sg13g2_decap_8 FILLER_66_1142 ();
 sg13g2_decap_8 FILLER_66_1149 ();
 sg13g2_fill_2 FILLER_66_1156 ();
 sg13g2_fill_1 FILLER_66_1158 ();
 sg13g2_fill_1 FILLER_66_1192 ();
 sg13g2_fill_1 FILLER_66_1198 ();
 sg13g2_fill_2 FILLER_66_1217 ();
 sg13g2_decap_8 FILLER_66_1232 ();
 sg13g2_decap_8 FILLER_66_1239 ();
 sg13g2_decap_8 FILLER_66_1246 ();
 sg13g2_decap_4 FILLER_66_1274 ();
 sg13g2_fill_1 FILLER_66_1278 ();
 sg13g2_decap_4 FILLER_66_1313 ();
 sg13g2_fill_2 FILLER_66_1317 ();
 sg13g2_fill_1 FILLER_66_1332 ();
 sg13g2_fill_1 FILLER_66_1340 ();
 sg13g2_fill_1 FILLER_66_1354 ();
 sg13g2_fill_1 FILLER_66_1364 ();
 sg13g2_fill_1 FILLER_66_1370 ();
 sg13g2_fill_1 FILLER_66_1375 ();
 sg13g2_fill_1 FILLER_66_1383 ();
 sg13g2_fill_1 FILLER_66_1388 ();
 sg13g2_decap_8 FILLER_66_1394 ();
 sg13g2_fill_2 FILLER_66_1409 ();
 sg13g2_fill_1 FILLER_66_1411 ();
 sg13g2_fill_2 FILLER_66_1422 ();
 sg13g2_decap_8 FILLER_66_1429 ();
 sg13g2_decap_4 FILLER_66_1436 ();
 sg13g2_fill_2 FILLER_66_1440 ();
 sg13g2_decap_4 FILLER_66_1448 ();
 sg13g2_fill_1 FILLER_66_1472 ();
 sg13g2_decap_8 FILLER_66_1485 ();
 sg13g2_decap_8 FILLER_66_1492 ();
 sg13g2_decap_4 FILLER_66_1514 ();
 sg13g2_fill_2 FILLER_66_1531 ();
 sg13g2_fill_1 FILLER_66_1533 ();
 sg13g2_fill_1 FILLER_66_1545 ();
 sg13g2_fill_2 FILLER_66_1561 ();
 sg13g2_fill_1 FILLER_66_1568 ();
 sg13g2_fill_2 FILLER_66_1573 ();
 sg13g2_decap_8 FILLER_66_1580 ();
 sg13g2_decap_8 FILLER_66_1587 ();
 sg13g2_decap_8 FILLER_66_1594 ();
 sg13g2_fill_2 FILLER_66_1601 ();
 sg13g2_fill_1 FILLER_66_1603 ();
 sg13g2_fill_2 FILLER_66_1634 ();
 sg13g2_fill_1 FILLER_66_1636 ();
 sg13g2_fill_2 FILLER_66_1670 ();
 sg13g2_fill_1 FILLER_66_1672 ();
 sg13g2_decap_4 FILLER_66_1698 ();
 sg13g2_fill_2 FILLER_66_1702 ();
 sg13g2_fill_2 FILLER_66_1715 ();
 sg13g2_fill_2 FILLER_66_1741 ();
 sg13g2_fill_1 FILLER_66_1756 ();
 sg13g2_fill_1 FILLER_66_1807 ();
 sg13g2_fill_2 FILLER_66_1820 ();
 sg13g2_fill_2 FILLER_66_1830 ();
 sg13g2_fill_2 FILLER_66_1838 ();
 sg13g2_fill_2 FILLER_66_1858 ();
 sg13g2_fill_2 FILLER_66_1903 ();
 sg13g2_fill_2 FILLER_66_1925 ();
 sg13g2_fill_1 FILLER_66_1931 ();
 sg13g2_decap_8 FILLER_66_1975 ();
 sg13g2_decap_8 FILLER_66_1982 ();
 sg13g2_decap_8 FILLER_66_1989 ();
 sg13g2_fill_1 FILLER_66_2031 ();
 sg13g2_fill_1 FILLER_66_2040 ();
 sg13g2_fill_1 FILLER_66_2045 ();
 sg13g2_fill_1 FILLER_66_2055 ();
 sg13g2_fill_2 FILLER_66_2082 ();
 sg13g2_decap_4 FILLER_66_2140 ();
 sg13g2_fill_1 FILLER_66_2144 ();
 sg13g2_fill_2 FILLER_66_2181 ();
 sg13g2_fill_2 FILLER_66_2217 ();
 sg13g2_fill_1 FILLER_66_2229 ();
 sg13g2_decap_8 FILLER_66_2235 ();
 sg13g2_fill_2 FILLER_66_2242 ();
 sg13g2_decap_8 FILLER_66_2248 ();
 sg13g2_fill_2 FILLER_66_2255 ();
 sg13g2_fill_1 FILLER_66_2257 ();
 sg13g2_fill_2 FILLER_66_2263 ();
 sg13g2_fill_1 FILLER_66_2265 ();
 sg13g2_decap_8 FILLER_66_2289 ();
 sg13g2_decap_8 FILLER_66_2296 ();
 sg13g2_decap_8 FILLER_66_2303 ();
 sg13g2_fill_1 FILLER_66_2310 ();
 sg13g2_decap_8 FILLER_66_2324 ();
 sg13g2_decap_8 FILLER_66_2331 ();
 sg13g2_fill_2 FILLER_66_2338 ();
 sg13g2_decap_4 FILLER_66_2344 ();
 sg13g2_decap_8 FILLER_66_2358 ();
 sg13g2_fill_2 FILLER_66_2382 ();
 sg13g2_fill_1 FILLER_66_2384 ();
 sg13g2_fill_2 FILLER_66_2423 ();
 sg13g2_decap_4 FILLER_66_2438 ();
 sg13g2_fill_1 FILLER_66_2446 ();
 sg13g2_fill_2 FILLER_66_2451 ();
 sg13g2_decap_8 FILLER_66_2494 ();
 sg13g2_fill_2 FILLER_66_2501 ();
 sg13g2_fill_1 FILLER_66_2503 ();
 sg13g2_fill_2 FILLER_66_2508 ();
 sg13g2_fill_1 FILLER_66_2510 ();
 sg13g2_decap_4 FILLER_66_2517 ();
 sg13g2_fill_1 FILLER_66_2521 ();
 sg13g2_decap_8 FILLER_66_2558 ();
 sg13g2_decap_8 FILLER_66_2565 ();
 sg13g2_decap_8 FILLER_66_2572 ();
 sg13g2_decap_8 FILLER_66_2579 ();
 sg13g2_decap_8 FILLER_66_2586 ();
 sg13g2_decap_8 FILLER_66_2593 ();
 sg13g2_decap_8 FILLER_66_2600 ();
 sg13g2_decap_8 FILLER_66_2607 ();
 sg13g2_decap_8 FILLER_66_2614 ();
 sg13g2_decap_8 FILLER_66_2621 ();
 sg13g2_decap_8 FILLER_66_2628 ();
 sg13g2_decap_8 FILLER_66_2635 ();
 sg13g2_decap_8 FILLER_66_2642 ();
 sg13g2_decap_8 FILLER_66_2649 ();
 sg13g2_decap_8 FILLER_66_2656 ();
 sg13g2_decap_8 FILLER_66_2663 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_fill_2 FILLER_67_33 ();
 sg13g2_fill_2 FILLER_67_78 ();
 sg13g2_fill_1 FILLER_67_80 ();
 sg13g2_fill_2 FILLER_67_124 ();
 sg13g2_fill_1 FILLER_67_126 ();
 sg13g2_fill_1 FILLER_67_138 ();
 sg13g2_fill_2 FILLER_67_204 ();
 sg13g2_fill_1 FILLER_67_206 ();
 sg13g2_fill_2 FILLER_67_212 ();
 sg13g2_fill_1 FILLER_67_214 ();
 sg13g2_fill_2 FILLER_67_230 ();
 sg13g2_fill_1 FILLER_67_242 ();
 sg13g2_fill_2 FILLER_67_264 ();
 sg13g2_fill_2 FILLER_67_291 ();
 sg13g2_fill_1 FILLER_67_298 ();
 sg13g2_decap_8 FILLER_67_303 ();
 sg13g2_fill_2 FILLER_67_321 ();
 sg13g2_fill_2 FILLER_67_329 ();
 sg13g2_fill_1 FILLER_67_331 ();
 sg13g2_fill_1 FILLER_67_337 ();
 sg13g2_fill_2 FILLER_67_352 ();
 sg13g2_fill_2 FILLER_67_382 ();
 sg13g2_fill_1 FILLER_67_389 ();
 sg13g2_fill_1 FILLER_67_394 ();
 sg13g2_decap_8 FILLER_67_430 ();
 sg13g2_decap_8 FILLER_67_437 ();
 sg13g2_fill_1 FILLER_67_453 ();
 sg13g2_fill_2 FILLER_67_458 ();
 sg13g2_decap_8 FILLER_67_495 ();
 sg13g2_decap_4 FILLER_67_502 ();
 sg13g2_fill_2 FILLER_67_506 ();
 sg13g2_fill_2 FILLER_67_513 ();
 sg13g2_fill_2 FILLER_67_538 ();
 sg13g2_fill_2 FILLER_67_581 ();
 sg13g2_fill_1 FILLER_67_583 ();
 sg13g2_fill_2 FILLER_67_588 ();
 sg13g2_fill_2 FILLER_67_616 ();
 sg13g2_fill_1 FILLER_67_618 ();
 sg13g2_fill_1 FILLER_67_625 ();
 sg13g2_decap_8 FILLER_67_631 ();
 sg13g2_fill_2 FILLER_67_641 ();
 sg13g2_fill_1 FILLER_67_643 ();
 sg13g2_decap_8 FILLER_67_649 ();
 sg13g2_decap_8 FILLER_67_664 ();
 sg13g2_fill_2 FILLER_67_703 ();
 sg13g2_fill_2 FILLER_67_856 ();
 sg13g2_fill_2 FILLER_67_914 ();
 sg13g2_decap_8 FILLER_67_924 ();
 sg13g2_decap_8 FILLER_67_931 ();
 sg13g2_decap_8 FILLER_67_938 ();
 sg13g2_decap_8 FILLER_67_945 ();
 sg13g2_decap_8 FILLER_67_952 ();
 sg13g2_fill_1 FILLER_67_959 ();
 sg13g2_fill_2 FILLER_67_975 ();
 sg13g2_fill_2 FILLER_67_980 ();
 sg13g2_fill_2 FILLER_67_1016 ();
 sg13g2_fill_2 FILLER_67_1045 ();
 sg13g2_fill_1 FILLER_67_1073 ();
 sg13g2_fill_2 FILLER_67_1093 ();
 sg13g2_fill_1 FILLER_67_1095 ();
 sg13g2_fill_2 FILLER_67_1123 ();
 sg13g2_fill_2 FILLER_67_1130 ();
 sg13g2_decap_8 FILLER_67_1144 ();
 sg13g2_decap_4 FILLER_67_1151 ();
 sg13g2_fill_1 FILLER_67_1155 ();
 sg13g2_decap_8 FILLER_67_1161 ();
 sg13g2_fill_1 FILLER_67_1168 ();
 sg13g2_fill_2 FILLER_67_1183 ();
 sg13g2_fill_1 FILLER_67_1185 ();
 sg13g2_decap_8 FILLER_67_1190 ();
 sg13g2_fill_2 FILLER_67_1203 ();
 sg13g2_fill_1 FILLER_67_1217 ();
 sg13g2_fill_2 FILLER_67_1231 ();
 sg13g2_fill_1 FILLER_67_1249 ();
 sg13g2_fill_2 FILLER_67_1268 ();
 sg13g2_fill_2 FILLER_67_1274 ();
 sg13g2_decap_4 FILLER_67_1304 ();
 sg13g2_decap_8 FILLER_67_1316 ();
 sg13g2_decap_8 FILLER_67_1323 ();
 sg13g2_fill_1 FILLER_67_1348 ();
 sg13g2_decap_8 FILLER_67_1361 ();
 sg13g2_decap_4 FILLER_67_1372 ();
 sg13g2_fill_2 FILLER_67_1376 ();
 sg13g2_fill_1 FILLER_67_1403 ();
 sg13g2_decap_8 FILLER_67_1421 ();
 sg13g2_fill_2 FILLER_67_1428 ();
 sg13g2_fill_1 FILLER_67_1437 ();
 sg13g2_decap_8 FILLER_67_1443 ();
 sg13g2_fill_2 FILLER_67_1450 ();
 sg13g2_fill_1 FILLER_67_1452 ();
 sg13g2_fill_2 FILLER_67_1468 ();
 sg13g2_fill_1 FILLER_67_1470 ();
 sg13g2_decap_8 FILLER_67_1478 ();
 sg13g2_fill_2 FILLER_67_1485 ();
 sg13g2_fill_2 FILLER_67_1492 ();
 sg13g2_decap_4 FILLER_67_1498 ();
 sg13g2_fill_2 FILLER_67_1517 ();
 sg13g2_decap_4 FILLER_67_1524 ();
 sg13g2_fill_2 FILLER_67_1528 ();
 sg13g2_fill_2 FILLER_67_1554 ();
 sg13g2_fill_1 FILLER_67_1556 ();
 sg13g2_fill_2 FILLER_67_1565 ();
 sg13g2_fill_2 FILLER_67_1571 ();
 sg13g2_fill_1 FILLER_67_1573 ();
 sg13g2_fill_2 FILLER_67_1579 ();
 sg13g2_fill_2 FILLER_67_1585 ();
 sg13g2_fill_1 FILLER_67_1587 ();
 sg13g2_fill_2 FILLER_67_1613 ();
 sg13g2_decap_4 FILLER_67_1619 ();
 sg13g2_fill_1 FILLER_67_1623 ();
 sg13g2_fill_1 FILLER_67_1650 ();
 sg13g2_decap_4 FILLER_67_1658 ();
 sg13g2_fill_1 FILLER_67_1662 ();
 sg13g2_fill_1 FILLER_67_1673 ();
 sg13g2_fill_1 FILLER_67_1685 ();
 sg13g2_decap_4 FILLER_67_1691 ();
 sg13g2_fill_1 FILLER_67_1695 ();
 sg13g2_fill_1 FILLER_67_1707 ();
 sg13g2_fill_2 FILLER_67_1728 ();
 sg13g2_fill_1 FILLER_67_1740 ();
 sg13g2_fill_1 FILLER_67_1770 ();
 sg13g2_fill_1 FILLER_67_1789 ();
 sg13g2_fill_1 FILLER_67_1795 ();
 sg13g2_fill_1 FILLER_67_1812 ();
 sg13g2_fill_1 FILLER_67_1816 ();
 sg13g2_fill_2 FILLER_67_1844 ();
 sg13g2_fill_1 FILLER_67_1859 ();
 sg13g2_fill_1 FILLER_67_1888 ();
 sg13g2_fill_1 FILLER_67_1897 ();
 sg13g2_fill_2 FILLER_67_1905 ();
 sg13g2_fill_1 FILLER_67_1987 ();
 sg13g2_fill_1 FILLER_67_1998 ();
 sg13g2_decap_4 FILLER_67_2090 ();
 sg13g2_fill_2 FILLER_67_2094 ();
 sg13g2_fill_2 FILLER_67_2100 ();
 sg13g2_fill_2 FILLER_67_2106 ();
 sg13g2_fill_1 FILLER_67_2108 ();
 sg13g2_decap_4 FILLER_67_2140 ();
 sg13g2_decap_4 FILLER_67_2162 ();
 sg13g2_fill_2 FILLER_67_2172 ();
 sg13g2_fill_1 FILLER_67_2174 ();
 sg13g2_decap_4 FILLER_67_2225 ();
 sg13g2_fill_2 FILLER_67_2265 ();
 sg13g2_fill_1 FILLER_67_2267 ();
 sg13g2_fill_2 FILLER_67_2272 ();
 sg13g2_fill_2 FILLER_67_2297 ();
 sg13g2_fill_2 FILLER_67_2309 ();
 sg13g2_decap_8 FILLER_67_2352 ();
 sg13g2_fill_1 FILLER_67_2359 ();
 sg13g2_fill_2 FILLER_67_2391 ();
 sg13g2_fill_1 FILLER_67_2393 ();
 sg13g2_decap_4 FILLER_67_2479 ();
 sg13g2_decap_8 FILLER_67_2515 ();
 sg13g2_fill_2 FILLER_67_2522 ();
 sg13g2_fill_1 FILLER_67_2524 ();
 sg13g2_decap_8 FILLER_67_2578 ();
 sg13g2_decap_8 FILLER_67_2585 ();
 sg13g2_decap_8 FILLER_67_2592 ();
 sg13g2_decap_8 FILLER_67_2599 ();
 sg13g2_decap_8 FILLER_67_2606 ();
 sg13g2_decap_8 FILLER_67_2613 ();
 sg13g2_decap_8 FILLER_67_2620 ();
 sg13g2_decap_8 FILLER_67_2627 ();
 sg13g2_decap_8 FILLER_67_2634 ();
 sg13g2_decap_8 FILLER_67_2641 ();
 sg13g2_decap_8 FILLER_67_2648 ();
 sg13g2_decap_8 FILLER_67_2655 ();
 sg13g2_decap_8 FILLER_67_2662 ();
 sg13g2_fill_1 FILLER_67_2669 ();
 sg13g2_fill_1 FILLER_68_4 ();
 sg13g2_fill_1 FILLER_68_71 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_fill_2 FILLER_68_84 ();
 sg13g2_fill_1 FILLER_68_86 ();
 sg13g2_decap_4 FILLER_68_91 ();
 sg13g2_fill_2 FILLER_68_99 ();
 sg13g2_fill_1 FILLER_68_105 ();
 sg13g2_fill_1 FILLER_68_111 ();
 sg13g2_decap_4 FILLER_68_164 ();
 sg13g2_decap_8 FILLER_68_194 ();
 sg13g2_decap_4 FILLER_68_201 ();
 sg13g2_fill_2 FILLER_68_205 ();
 sg13g2_decap_8 FILLER_68_212 ();
 sg13g2_fill_1 FILLER_68_219 ();
 sg13g2_decap_4 FILLER_68_228 ();
 sg13g2_fill_1 FILLER_68_237 ();
 sg13g2_fill_1 FILLER_68_244 ();
 sg13g2_fill_1 FILLER_68_250 ();
 sg13g2_fill_1 FILLER_68_256 ();
 sg13g2_fill_1 FILLER_68_262 ();
 sg13g2_decap_8 FILLER_68_299 ();
 sg13g2_decap_8 FILLER_68_306 ();
 sg13g2_fill_2 FILLER_68_313 ();
 sg13g2_fill_1 FILLER_68_315 ();
 sg13g2_fill_2 FILLER_68_326 ();
 sg13g2_fill_1 FILLER_68_328 ();
 sg13g2_fill_1 FILLER_68_345 ();
 sg13g2_fill_1 FILLER_68_371 ();
 sg13g2_fill_2 FILLER_68_376 ();
 sg13g2_fill_1 FILLER_68_378 ();
 sg13g2_fill_1 FILLER_68_405 ();
 sg13g2_fill_1 FILLER_68_410 ();
 sg13g2_fill_2 FILLER_68_415 ();
 sg13g2_fill_2 FILLER_68_421 ();
 sg13g2_fill_2 FILLER_68_449 ();
 sg13g2_decap_4 FILLER_68_455 ();
 sg13g2_fill_2 FILLER_68_459 ();
 sg13g2_fill_1 FILLER_68_466 ();
 sg13g2_fill_1 FILLER_68_471 ();
 sg13g2_fill_2 FILLER_68_485 ();
 sg13g2_fill_1 FILLER_68_487 ();
 sg13g2_decap_4 FILLER_68_497 ();
 sg13g2_fill_1 FILLER_68_501 ();
 sg13g2_fill_2 FILLER_68_571 ();
 sg13g2_fill_1 FILLER_68_573 ();
 sg13g2_fill_2 FILLER_68_589 ();
 sg13g2_fill_1 FILLER_68_591 ();
 sg13g2_fill_1 FILLER_68_602 ();
 sg13g2_decap_8 FILLER_68_652 ();
 sg13g2_decap_4 FILLER_68_659 ();
 sg13g2_fill_2 FILLER_68_698 ();
 sg13g2_fill_1 FILLER_68_788 ();
 sg13g2_fill_1 FILLER_68_815 ();
 sg13g2_decap_4 FILLER_68_899 ();
 sg13g2_fill_1 FILLER_68_903 ();
 sg13g2_decap_8 FILLER_68_912 ();
 sg13g2_fill_1 FILLER_68_919 ();
 sg13g2_decap_4 FILLER_68_933 ();
 sg13g2_decap_8 FILLER_68_941 ();
 sg13g2_fill_1 FILLER_68_948 ();
 sg13g2_fill_2 FILLER_68_972 ();
 sg13g2_fill_1 FILLER_68_974 ();
 sg13g2_fill_1 FILLER_68_1079 ();
 sg13g2_fill_1 FILLER_68_1085 ();
 sg13g2_fill_1 FILLER_68_1090 ();
 sg13g2_fill_2 FILLER_68_1095 ();
 sg13g2_fill_2 FILLER_68_1108 ();
 sg13g2_fill_2 FILLER_68_1163 ();
 sg13g2_decap_4 FILLER_68_1170 ();
 sg13g2_fill_1 FILLER_68_1174 ();
 sg13g2_decap_4 FILLER_68_1204 ();
 sg13g2_fill_1 FILLER_68_1208 ();
 sg13g2_fill_2 FILLER_68_1217 ();
 sg13g2_fill_1 FILLER_68_1219 ();
 sg13g2_fill_2 FILLER_68_1232 ();
 sg13g2_fill_1 FILLER_68_1234 ();
 sg13g2_fill_1 FILLER_68_1239 ();
 sg13g2_fill_2 FILLER_68_1244 ();
 sg13g2_fill_2 FILLER_68_1251 ();
 sg13g2_fill_1 FILLER_68_1253 ();
 sg13g2_fill_1 FILLER_68_1267 ();
 sg13g2_decap_8 FILLER_68_1273 ();
 sg13g2_decap_8 FILLER_68_1280 ();
 sg13g2_fill_1 FILLER_68_1291 ();
 sg13g2_fill_1 FILLER_68_1302 ();
 sg13g2_decap_8 FILLER_68_1307 ();
 sg13g2_fill_2 FILLER_68_1314 ();
 sg13g2_fill_1 FILLER_68_1316 ();
 sg13g2_fill_1 FILLER_68_1341 ();
 sg13g2_decap_8 FILLER_68_1354 ();
 sg13g2_decap_8 FILLER_68_1376 ();
 sg13g2_decap_4 FILLER_68_1433 ();
 sg13g2_fill_2 FILLER_68_1437 ();
 sg13g2_decap_8 FILLER_68_1448 ();
 sg13g2_decap_8 FILLER_68_1455 ();
 sg13g2_decap_4 FILLER_68_1462 ();
 sg13g2_fill_1 FILLER_68_1466 ();
 sg13g2_decap_4 FILLER_68_1483 ();
 sg13g2_fill_2 FILLER_68_1514 ();
 sg13g2_fill_1 FILLER_68_1521 ();
 sg13g2_decap_8 FILLER_68_1526 ();
 sg13g2_fill_2 FILLER_68_1533 ();
 sg13g2_fill_2 FILLER_68_1539 ();
 sg13g2_fill_2 FILLER_68_1566 ();
 sg13g2_fill_2 FILLER_68_1619 ();
 sg13g2_decap_8 FILLER_68_1635 ();
 sg13g2_decap_4 FILLER_68_1642 ();
 sg13g2_decap_8 FILLER_68_1650 ();
 sg13g2_fill_2 FILLER_68_1657 ();
 sg13g2_fill_1 FILLER_68_1659 ();
 sg13g2_fill_1 FILLER_68_1679 ();
 sg13g2_decap_8 FILLER_68_1703 ();
 sg13g2_fill_2 FILLER_68_1710 ();
 sg13g2_decap_8 FILLER_68_1715 ();
 sg13g2_decap_4 FILLER_68_1726 ();
 sg13g2_fill_2 FILLER_68_1730 ();
 sg13g2_fill_2 FILLER_68_1741 ();
 sg13g2_fill_1 FILLER_68_1754 ();
 sg13g2_fill_1 FILLER_68_1772 ();
 sg13g2_fill_1 FILLER_68_1782 ();
 sg13g2_fill_2 FILLER_68_1796 ();
 sg13g2_fill_1 FILLER_68_1812 ();
 sg13g2_fill_2 FILLER_68_1819 ();
 sg13g2_fill_2 FILLER_68_1834 ();
 sg13g2_fill_1 FILLER_68_1894 ();
 sg13g2_fill_1 FILLER_68_1921 ();
 sg13g2_fill_1 FILLER_68_1948 ();
 sg13g2_fill_1 FILLER_68_1970 ();
 sg13g2_fill_2 FILLER_68_1983 ();
 sg13g2_fill_1 FILLER_68_1985 ();
 sg13g2_fill_2 FILLER_68_2021 ();
 sg13g2_fill_2 FILLER_68_2031 ();
 sg13g2_decap_4 FILLER_68_2077 ();
 sg13g2_fill_2 FILLER_68_2081 ();
 sg13g2_decap_8 FILLER_68_2088 ();
 sg13g2_decap_8 FILLER_68_2095 ();
 sg13g2_decap_8 FILLER_68_2102 ();
 sg13g2_fill_2 FILLER_68_2109 ();
 sg13g2_decap_4 FILLER_68_2154 ();
 sg13g2_fill_1 FILLER_68_2158 ();
 sg13g2_fill_1 FILLER_68_2164 ();
 sg13g2_decap_8 FILLER_68_2178 ();
 sg13g2_decap_8 FILLER_68_2185 ();
 sg13g2_fill_1 FILLER_68_2216 ();
 sg13g2_fill_1 FILLER_68_2227 ();
 sg13g2_fill_1 FILLER_68_2264 ();
 sg13g2_fill_2 FILLER_68_2291 ();
 sg13g2_fill_2 FILLER_68_2323 ();
 sg13g2_decap_8 FILLER_68_2334 ();
 sg13g2_decap_8 FILLER_68_2345 ();
 sg13g2_decap_8 FILLER_68_2352 ();
 sg13g2_decap_8 FILLER_68_2359 ();
 sg13g2_decap_4 FILLER_68_2366 ();
 sg13g2_fill_1 FILLER_68_2370 ();
 sg13g2_decap_4 FILLER_68_2375 ();
 sg13g2_fill_1 FILLER_68_2379 ();
 sg13g2_decap_8 FILLER_68_2390 ();
 sg13g2_fill_2 FILLER_68_2397 ();
 sg13g2_decap_8 FILLER_68_2464 ();
 sg13g2_decap_4 FILLER_68_2471 ();
 sg13g2_fill_2 FILLER_68_2507 ();
 sg13g2_decap_8 FILLER_68_2565 ();
 sg13g2_decap_8 FILLER_68_2572 ();
 sg13g2_decap_8 FILLER_68_2579 ();
 sg13g2_decap_8 FILLER_68_2586 ();
 sg13g2_decap_8 FILLER_68_2593 ();
 sg13g2_decap_8 FILLER_68_2600 ();
 sg13g2_decap_8 FILLER_68_2607 ();
 sg13g2_decap_8 FILLER_68_2614 ();
 sg13g2_decap_8 FILLER_68_2621 ();
 sg13g2_decap_8 FILLER_68_2628 ();
 sg13g2_decap_8 FILLER_68_2635 ();
 sg13g2_decap_8 FILLER_68_2642 ();
 sg13g2_decap_8 FILLER_68_2649 ();
 sg13g2_decap_8 FILLER_68_2656 ();
 sg13g2_decap_8 FILLER_68_2663 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_fill_2 FILLER_69_37 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_fill_1 FILLER_69_63 ();
 sg13g2_decap_4 FILLER_69_67 ();
 sg13g2_decap_8 FILLER_69_75 ();
 sg13g2_fill_2 FILLER_69_82 ();
 sg13g2_fill_1 FILLER_69_110 ();
 sg13g2_fill_2 FILLER_69_115 ();
 sg13g2_fill_1 FILLER_69_143 ();
 sg13g2_fill_1 FILLER_69_154 ();
 sg13g2_decap_8 FILLER_69_159 ();
 sg13g2_decap_8 FILLER_69_166 ();
 sg13g2_decap_4 FILLER_69_173 ();
 sg13g2_decap_8 FILLER_69_181 ();
 sg13g2_fill_2 FILLER_69_188 ();
 sg13g2_decap_4 FILLER_69_225 ();
 sg13g2_fill_2 FILLER_69_229 ();
 sg13g2_decap_4 FILLER_69_235 ();
 sg13g2_fill_2 FILLER_69_239 ();
 sg13g2_fill_2 FILLER_69_276 ();
 sg13g2_fill_1 FILLER_69_282 ();
 sg13g2_decap_8 FILLER_69_288 ();
 sg13g2_fill_1 FILLER_69_295 ();
 sg13g2_decap_8 FILLER_69_300 ();
 sg13g2_decap_8 FILLER_69_307 ();
 sg13g2_decap_4 FILLER_69_314 ();
 sg13g2_fill_2 FILLER_69_318 ();
 sg13g2_decap_8 FILLER_69_380 ();
 sg13g2_fill_1 FILLER_69_387 ();
 sg13g2_fill_1 FILLER_69_414 ();
 sg13g2_fill_2 FILLER_69_454 ();
 sg13g2_decap_8 FILLER_69_462 ();
 sg13g2_decap_4 FILLER_69_469 ();
 sg13g2_fill_2 FILLER_69_473 ();
 sg13g2_decap_8 FILLER_69_484 ();
 sg13g2_fill_2 FILLER_69_491 ();
 sg13g2_fill_1 FILLER_69_493 ();
 sg13g2_fill_1 FILLER_69_499 ();
 sg13g2_fill_1 FILLER_69_531 ();
 sg13g2_decap_8 FILLER_69_537 ();
 sg13g2_fill_2 FILLER_69_548 ();
 sg13g2_fill_1 FILLER_69_559 ();
 sg13g2_fill_1 FILLER_69_616 ();
 sg13g2_fill_1 FILLER_69_624 ();
 sg13g2_decap_4 FILLER_69_633 ();
 sg13g2_fill_1 FILLER_69_637 ();
 sg13g2_decap_4 FILLER_69_674 ();
 sg13g2_fill_1 FILLER_69_678 ();
 sg13g2_decap_4 FILLER_69_689 ();
 sg13g2_fill_1 FILLER_69_693 ();
 sg13g2_decap_8 FILLER_69_700 ();
 sg13g2_fill_1 FILLER_69_707 ();
 sg13g2_fill_2 FILLER_69_716 ();
 sg13g2_fill_2 FILLER_69_722 ();
 sg13g2_fill_2 FILLER_69_727 ();
 sg13g2_fill_2 FILLER_69_747 ();
 sg13g2_fill_1 FILLER_69_787 ();
 sg13g2_fill_2 FILLER_69_794 ();
 sg13g2_fill_1 FILLER_69_796 ();
 sg13g2_decap_8 FILLER_69_804 ();
 sg13g2_fill_2 FILLER_69_811 ();
 sg13g2_fill_1 FILLER_69_838 ();
 sg13g2_fill_1 FILLER_69_851 ();
 sg13g2_fill_1 FILLER_69_877 ();
 sg13g2_fill_2 FILLER_69_884 ();
 sg13g2_fill_1 FILLER_69_945 ();
 sg13g2_decap_4 FILLER_69_976 ();
 sg13g2_fill_2 FILLER_69_980 ();
 sg13g2_fill_1 FILLER_69_987 ();
 sg13g2_fill_2 FILLER_69_997 ();
 sg13g2_fill_2 FILLER_69_1003 ();
 sg13g2_fill_2 FILLER_69_1091 ();
 sg13g2_fill_1 FILLER_69_1093 ();
 sg13g2_fill_1 FILLER_69_1103 ();
 sg13g2_decap_8 FILLER_69_1117 ();
 sg13g2_decap_4 FILLER_69_1141 ();
 sg13g2_fill_2 FILLER_69_1149 ();
 sg13g2_decap_4 FILLER_69_1161 ();
 sg13g2_fill_1 FILLER_69_1178 ();
 sg13g2_fill_2 FILLER_69_1188 ();
 sg13g2_decap_4 FILLER_69_1200 ();
 sg13g2_fill_1 FILLER_69_1204 ();
 sg13g2_fill_1 FILLER_69_1233 ();
 sg13g2_fill_1 FILLER_69_1243 ();
 sg13g2_fill_1 FILLER_69_1263 ();
 sg13g2_fill_2 FILLER_69_1269 ();
 sg13g2_fill_1 FILLER_69_1271 ();
 sg13g2_fill_1 FILLER_69_1296 ();
 sg13g2_decap_8 FILLER_69_1315 ();
 sg13g2_decap_8 FILLER_69_1322 ();
 sg13g2_fill_1 FILLER_69_1329 ();
 sg13g2_fill_2 FILLER_69_1339 ();
 sg13g2_fill_1 FILLER_69_1345 ();
 sg13g2_fill_1 FILLER_69_1384 ();
 sg13g2_fill_2 FILLER_69_1390 ();
 sg13g2_fill_2 FILLER_69_1412 ();
 sg13g2_fill_1 FILLER_69_1414 ();
 sg13g2_decap_4 FILLER_69_1430 ();
 sg13g2_fill_2 FILLER_69_1434 ();
 sg13g2_fill_1 FILLER_69_1465 ();
 sg13g2_fill_2 FILLER_69_1470 ();
 sg13g2_fill_1 FILLER_69_1480 ();
 sg13g2_decap_4 FILLER_69_1485 ();
 sg13g2_fill_2 FILLER_69_1489 ();
 sg13g2_decap_4 FILLER_69_1515 ();
 sg13g2_fill_2 FILLER_69_1519 ();
 sg13g2_decap_8 FILLER_69_1525 ();
 sg13g2_fill_2 FILLER_69_1532 ();
 sg13g2_decap_8 FILLER_69_1547 ();
 sg13g2_fill_2 FILLER_69_1554 ();
 sg13g2_fill_1 FILLER_69_1556 ();
 sg13g2_fill_2 FILLER_69_1572 ();
 sg13g2_fill_1 FILLER_69_1585 ();
 sg13g2_fill_1 FILLER_69_1606 ();
 sg13g2_fill_1 FILLER_69_1612 ();
 sg13g2_decap_4 FILLER_69_1623 ();
 sg13g2_fill_1 FILLER_69_1627 ();
 sg13g2_fill_2 FILLER_69_1638 ();
 sg13g2_decap_8 FILLER_69_1650 ();
 sg13g2_decap_8 FILLER_69_1657 ();
 sg13g2_decap_8 FILLER_69_1664 ();
 sg13g2_fill_2 FILLER_69_1671 ();
 sg13g2_fill_1 FILLER_69_1677 ();
 sg13g2_decap_8 FILLER_69_1683 ();
 sg13g2_decap_8 FILLER_69_1716 ();
 sg13g2_fill_2 FILLER_69_1723 ();
 sg13g2_decap_8 FILLER_69_1729 ();
 sg13g2_fill_1 FILLER_69_1736 ();
 sg13g2_decap_8 FILLER_69_1742 ();
 sg13g2_fill_2 FILLER_69_1749 ();
 sg13g2_fill_1 FILLER_69_1755 ();
 sg13g2_fill_1 FILLER_69_1777 ();
 sg13g2_fill_1 FILLER_69_1805 ();
 sg13g2_fill_1 FILLER_69_1809 ();
 sg13g2_fill_2 FILLER_69_1846 ();
 sg13g2_fill_2 FILLER_69_1947 ();
 sg13g2_fill_1 FILLER_69_1949 ();
 sg13g2_fill_2 FILLER_69_1961 ();
 sg13g2_fill_2 FILLER_69_1971 ();
 sg13g2_fill_1 FILLER_69_1973 ();
 sg13g2_decap_4 FILLER_69_1995 ();
 sg13g2_fill_2 FILLER_69_1999 ();
 sg13g2_fill_2 FILLER_69_2050 ();
 sg13g2_decap_8 FILLER_69_2078 ();
 sg13g2_fill_2 FILLER_69_2085 ();
 sg13g2_fill_1 FILLER_69_2087 ();
 sg13g2_decap_8 FILLER_69_2097 ();
 sg13g2_decap_8 FILLER_69_2104 ();
 sg13g2_decap_8 FILLER_69_2111 ();
 sg13g2_fill_2 FILLER_69_2118 ();
 sg13g2_fill_1 FILLER_69_2120 ();
 sg13g2_decap_4 FILLER_69_2131 ();
 sg13g2_decap_8 FILLER_69_2143 ();
 sg13g2_fill_2 FILLER_69_2251 ();
 sg13g2_fill_1 FILLER_69_2253 ();
 sg13g2_decap_4 FILLER_69_2294 ();
 sg13g2_fill_1 FILLER_69_2298 ();
 sg13g2_decap_4 FILLER_69_2319 ();
 sg13g2_fill_1 FILLER_69_2323 ();
 sg13g2_fill_1 FILLER_69_2334 ();
 sg13g2_fill_2 FILLER_69_2371 ();
 sg13g2_fill_2 FILLER_69_2445 ();
 sg13g2_fill_1 FILLER_69_2477 ();
 sg13g2_fill_2 FILLER_69_2492 ();
 sg13g2_fill_1 FILLER_69_2546 ();
 sg13g2_decap_8 FILLER_69_2573 ();
 sg13g2_decap_8 FILLER_69_2580 ();
 sg13g2_decap_8 FILLER_69_2587 ();
 sg13g2_decap_8 FILLER_69_2594 ();
 sg13g2_decap_8 FILLER_69_2601 ();
 sg13g2_decap_8 FILLER_69_2608 ();
 sg13g2_decap_8 FILLER_69_2615 ();
 sg13g2_decap_8 FILLER_69_2622 ();
 sg13g2_decap_8 FILLER_69_2629 ();
 sg13g2_decap_8 FILLER_69_2636 ();
 sg13g2_decap_8 FILLER_69_2643 ();
 sg13g2_decap_8 FILLER_69_2650 ();
 sg13g2_decap_8 FILLER_69_2657 ();
 sg13g2_decap_4 FILLER_69_2664 ();
 sg13g2_fill_2 FILLER_69_2668 ();
 sg13g2_decap_4 FILLER_70_0 ();
 sg13g2_fill_1 FILLER_70_4 ();
 sg13g2_fill_1 FILLER_70_15 ();
 sg13g2_decap_4 FILLER_70_26 ();
 sg13g2_decap_4 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_43 ();
 sg13g2_decap_8 FILLER_70_50 ();
 sg13g2_fill_1 FILLER_70_57 ();
 sg13g2_fill_2 FILLER_70_62 ();
 sg13g2_fill_1 FILLER_70_85 ();
 sg13g2_fill_2 FILLER_70_91 ();
 sg13g2_fill_1 FILLER_70_93 ();
 sg13g2_fill_2 FILLER_70_114 ();
 sg13g2_fill_1 FILLER_70_121 ();
 sg13g2_fill_2 FILLER_70_166 ();
 sg13g2_decap_4 FILLER_70_172 ();
 sg13g2_fill_2 FILLER_70_176 ();
 sg13g2_decap_4 FILLER_70_183 ();
 sg13g2_fill_1 FILLER_70_187 ();
 sg13g2_fill_1 FILLER_70_198 ();
 sg13g2_fill_2 FILLER_70_235 ();
 sg13g2_fill_2 FILLER_70_258 ();
 sg13g2_fill_2 FILLER_70_265 ();
 sg13g2_fill_1 FILLER_70_267 ();
 sg13g2_fill_2 FILLER_70_273 ();
 sg13g2_fill_1 FILLER_70_275 ();
 sg13g2_fill_2 FILLER_70_286 ();
 sg13g2_fill_1 FILLER_70_288 ();
 sg13g2_decap_8 FILLER_70_315 ();
 sg13g2_decap_4 FILLER_70_322 ();
 sg13g2_fill_2 FILLER_70_326 ();
 sg13g2_fill_1 FILLER_70_335 ();
 sg13g2_fill_1 FILLER_70_362 ();
 sg13g2_fill_2 FILLER_70_368 ();
 sg13g2_decap_8 FILLER_70_374 ();
 sg13g2_fill_1 FILLER_70_381 ();
 sg13g2_decap_4 FILLER_70_387 ();
 sg13g2_fill_1 FILLER_70_391 ();
 sg13g2_fill_1 FILLER_70_396 ();
 sg13g2_decap_8 FILLER_70_401 ();
 sg13g2_decap_4 FILLER_70_408 ();
 sg13g2_fill_2 FILLER_70_412 ();
 sg13g2_decap_8 FILLER_70_427 ();
 sg13g2_fill_1 FILLER_70_434 ();
 sg13g2_fill_1 FILLER_70_439 ();
 sg13g2_fill_2 FILLER_70_444 ();
 sg13g2_fill_2 FILLER_70_472 ();
 sg13g2_fill_1 FILLER_70_474 ();
 sg13g2_decap_8 FILLER_70_480 ();
 sg13g2_decap_4 FILLER_70_487 ();
 sg13g2_fill_1 FILLER_70_491 ();
 sg13g2_fill_1 FILLER_70_518 ();
 sg13g2_decap_4 FILLER_70_523 ();
 sg13g2_decap_8 FILLER_70_546 ();
 sg13g2_decap_8 FILLER_70_553 ();
 sg13g2_fill_2 FILLER_70_560 ();
 sg13g2_fill_1 FILLER_70_562 ();
 sg13g2_fill_1 FILLER_70_584 ();
 sg13g2_fill_1 FILLER_70_592 ();
 sg13g2_fill_1 FILLER_70_603 ();
 sg13g2_fill_1 FILLER_70_607 ();
 sg13g2_fill_2 FILLER_70_641 ();
 sg13g2_decap_8 FILLER_70_673 ();
 sg13g2_fill_1 FILLER_70_680 ();
 sg13g2_decap_4 FILLER_70_691 ();
 sg13g2_decap_8 FILLER_70_699 ();
 sg13g2_decap_4 FILLER_70_706 ();
 sg13g2_fill_1 FILLER_70_723 ();
 sg13g2_fill_1 FILLER_70_761 ();
 sg13g2_fill_2 FILLER_70_770 ();
 sg13g2_fill_2 FILLER_70_806 ();
 sg13g2_fill_2 FILLER_70_813 ();
 sg13g2_fill_1 FILLER_70_815 ();
 sg13g2_fill_2 FILLER_70_823 ();
 sg13g2_fill_1 FILLER_70_825 ();
 sg13g2_fill_2 FILLER_70_835 ();
 sg13g2_fill_1 FILLER_70_870 ();
 sg13g2_decap_4 FILLER_70_880 ();
 sg13g2_fill_2 FILLER_70_884 ();
 sg13g2_fill_2 FILLER_70_932 ();
 sg13g2_fill_2 FILLER_70_938 ();
 sg13g2_fill_2 FILLER_70_966 ();
 sg13g2_fill_2 FILLER_70_974 ();
 sg13g2_fill_2 FILLER_70_981 ();
 sg13g2_fill_1 FILLER_70_990 ();
 sg13g2_decap_8 FILLER_70_1001 ();
 sg13g2_decap_4 FILLER_70_1012 ();
 sg13g2_decap_4 FILLER_70_1028 ();
 sg13g2_decap_8 FILLER_70_1036 ();
 sg13g2_fill_2 FILLER_70_1043 ();
 sg13g2_decap_4 FILLER_70_1049 ();
 sg13g2_fill_1 FILLER_70_1053 ();
 sg13g2_fill_2 FILLER_70_1057 ();
 sg13g2_fill_1 FILLER_70_1067 ();
 sg13g2_fill_2 FILLER_70_1088 ();
 sg13g2_decap_8 FILLER_70_1130 ();
 sg13g2_fill_1 FILLER_70_1137 ();
 sg13g2_decap_8 FILLER_70_1143 ();
 sg13g2_fill_2 FILLER_70_1150 ();
 sg13g2_fill_1 FILLER_70_1152 ();
 sg13g2_fill_1 FILLER_70_1166 ();
 sg13g2_fill_1 FILLER_70_1171 ();
 sg13g2_fill_2 FILLER_70_1188 ();
 sg13g2_fill_1 FILLER_70_1190 ();
 sg13g2_fill_1 FILLER_70_1209 ();
 sg13g2_fill_1 FILLER_70_1216 ();
 sg13g2_fill_1 FILLER_70_1245 ();
 sg13g2_fill_1 FILLER_70_1271 ();
 sg13g2_decap_8 FILLER_70_1277 ();
 sg13g2_decap_8 FILLER_70_1284 ();
 sg13g2_decap_8 FILLER_70_1291 ();
 sg13g2_decap_4 FILLER_70_1298 ();
 sg13g2_decap_4 FILLER_70_1312 ();
 sg13g2_fill_2 FILLER_70_1316 ();
 sg13g2_fill_2 FILLER_70_1326 ();
 sg13g2_fill_1 FILLER_70_1341 ();
 sg13g2_fill_1 FILLER_70_1349 ();
 sg13g2_fill_2 FILLER_70_1364 ();
 sg13g2_fill_1 FILLER_70_1366 ();
 sg13g2_fill_1 FILLER_70_1396 ();
 sg13g2_fill_1 FILLER_70_1402 ();
 sg13g2_fill_1 FILLER_70_1416 ();
 sg13g2_fill_2 FILLER_70_1422 ();
 sg13g2_fill_1 FILLER_70_1424 ();
 sg13g2_fill_2 FILLER_70_1431 ();
 sg13g2_fill_1 FILLER_70_1433 ();
 sg13g2_fill_2 FILLER_70_1438 ();
 sg13g2_fill_2 FILLER_70_1445 ();
 sg13g2_fill_1 FILLER_70_1447 ();
 sg13g2_fill_1 FILLER_70_1453 ();
 sg13g2_fill_1 FILLER_70_1492 ();
 sg13g2_fill_2 FILLER_70_1497 ();
 sg13g2_fill_1 FILLER_70_1499 ();
 sg13g2_fill_2 FILLER_70_1513 ();
 sg13g2_fill_2 FILLER_70_1520 ();
 sg13g2_fill_2 FILLER_70_1527 ();
 sg13g2_decap_4 FILLER_70_1567 ();
 sg13g2_fill_2 FILLER_70_1571 ();
 sg13g2_fill_1 FILLER_70_1582 ();
 sg13g2_fill_2 FILLER_70_1590 ();
 sg13g2_fill_2 FILLER_70_1596 ();
 sg13g2_fill_1 FILLER_70_1598 ();
 sg13g2_fill_2 FILLER_70_1603 ();
 sg13g2_decap_4 FILLER_70_1609 ();
 sg13g2_fill_2 FILLER_70_1617 ();
 sg13g2_decap_4 FILLER_70_1650 ();
 sg13g2_fill_1 FILLER_70_1654 ();
 sg13g2_decap_4 FILLER_70_1662 ();
 sg13g2_fill_1 FILLER_70_1666 ();
 sg13g2_decap_4 FILLER_70_1679 ();
 sg13g2_fill_1 FILLER_70_1683 ();
 sg13g2_fill_1 FILLER_70_1692 ();
 sg13g2_decap_8 FILLER_70_1697 ();
 sg13g2_decap_8 FILLER_70_1704 ();
 sg13g2_decap_8 FILLER_70_1711 ();
 sg13g2_decap_8 FILLER_70_1726 ();
 sg13g2_fill_2 FILLER_70_1804 ();
 sg13g2_decap_4 FILLER_70_1819 ();
 sg13g2_fill_1 FILLER_70_1831 ();
 sg13g2_fill_2 FILLER_70_1847 ();
 sg13g2_fill_1 FILLER_70_1894 ();
 sg13g2_fill_2 FILLER_70_1900 ();
 sg13g2_fill_1 FILLER_70_1931 ();
 sg13g2_decap_8 FILLER_70_1939 ();
 sg13g2_fill_2 FILLER_70_1946 ();
 sg13g2_fill_1 FILLER_70_1948 ();
 sg13g2_fill_2 FILLER_70_1963 ();
 sg13g2_fill_2 FILLER_70_2012 ();
 sg13g2_fill_1 FILLER_70_2014 ();
 sg13g2_fill_1 FILLER_70_2020 ();
 sg13g2_fill_2 FILLER_70_2026 ();
 sg13g2_fill_2 FILLER_70_2071 ();
 sg13g2_decap_8 FILLER_70_2164 ();
 sg13g2_decap_8 FILLER_70_2171 ();
 sg13g2_fill_1 FILLER_70_2178 ();
 sg13g2_decap_4 FILLER_70_2183 ();
 sg13g2_fill_2 FILLER_70_2187 ();
 sg13g2_fill_2 FILLER_70_2249 ();
 sg13g2_decap_4 FILLER_70_2267 ();
 sg13g2_fill_2 FILLER_70_2275 ();
 sg13g2_decap_8 FILLER_70_2294 ();
 sg13g2_decap_4 FILLER_70_2313 ();
 sg13g2_fill_2 FILLER_70_2317 ();
 sg13g2_fill_1 FILLER_70_2365 ();
 sg13g2_fill_2 FILLER_70_2370 ();
 sg13g2_fill_1 FILLER_70_2372 ();
 sg13g2_decap_8 FILLER_70_2385 ();
 sg13g2_decap_4 FILLER_70_2392 ();
 sg13g2_fill_1 FILLER_70_2396 ();
 sg13g2_decap_4 FILLER_70_2403 ();
 sg13g2_fill_2 FILLER_70_2407 ();
 sg13g2_fill_1 FILLER_70_2434 ();
 sg13g2_fill_1 FILLER_70_2438 ();
 sg13g2_decap_4 FILLER_70_2449 ();
 sg13g2_fill_1 FILLER_70_2453 ();
 sg13g2_decap_8 FILLER_70_2458 ();
 sg13g2_decap_8 FILLER_70_2465 ();
 sg13g2_decap_8 FILLER_70_2472 ();
 sg13g2_fill_2 FILLER_70_2479 ();
 sg13g2_decap_4 FILLER_70_2485 ();
 sg13g2_fill_1 FILLER_70_2499 ();
 sg13g2_decap_4 FILLER_70_2504 ();
 sg13g2_fill_2 FILLER_70_2508 ();
 sg13g2_decap_4 FILLER_70_2516 ();
 sg13g2_fill_2 FILLER_70_2520 ();
 sg13g2_fill_2 FILLER_70_2526 ();
 sg13g2_fill_1 FILLER_70_2528 ();
 sg13g2_decap_8 FILLER_70_2533 ();
 sg13g2_decap_8 FILLER_70_2540 ();
 sg13g2_decap_4 FILLER_70_2547 ();
 sg13g2_fill_1 FILLER_70_2551 ();
 sg13g2_decap_8 FILLER_70_2556 ();
 sg13g2_decap_8 FILLER_70_2563 ();
 sg13g2_decap_8 FILLER_70_2570 ();
 sg13g2_decap_8 FILLER_70_2577 ();
 sg13g2_decap_8 FILLER_70_2584 ();
 sg13g2_decap_8 FILLER_70_2591 ();
 sg13g2_decap_8 FILLER_70_2598 ();
 sg13g2_decap_8 FILLER_70_2605 ();
 sg13g2_decap_8 FILLER_70_2612 ();
 sg13g2_decap_8 FILLER_70_2619 ();
 sg13g2_decap_8 FILLER_70_2626 ();
 sg13g2_decap_8 FILLER_70_2633 ();
 sg13g2_decap_8 FILLER_70_2640 ();
 sg13g2_decap_8 FILLER_70_2647 ();
 sg13g2_decap_8 FILLER_70_2654 ();
 sg13g2_decap_8 FILLER_70_2661 ();
 sg13g2_fill_2 FILLER_70_2668 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_fill_2 FILLER_71_14 ();
 sg13g2_fill_2 FILLER_71_44 ();
 sg13g2_fill_2 FILLER_71_54 ();
 sg13g2_fill_1 FILLER_71_56 ();
 sg13g2_fill_1 FILLER_71_96 ();
 sg13g2_fill_1 FILLER_71_102 ();
 sg13g2_fill_1 FILLER_71_108 ();
 sg13g2_fill_1 FILLER_71_121 ();
 sg13g2_decap_8 FILLER_71_148 ();
 sg13g2_fill_2 FILLER_71_155 ();
 sg13g2_fill_1 FILLER_71_188 ();
 sg13g2_decap_4 FILLER_71_215 ();
 sg13g2_decap_8 FILLER_71_246 ();
 sg13g2_decap_4 FILLER_71_253 ();
 sg13g2_fill_1 FILLER_71_257 ();
 sg13g2_fill_2 FILLER_71_299 ();
 sg13g2_decap_8 FILLER_71_390 ();
 sg13g2_decap_8 FILLER_71_397 ();
 sg13g2_decap_8 FILLER_71_404 ();
 sg13g2_decap_4 FILLER_71_411 ();
 sg13g2_decap_8 FILLER_71_423 ();
 sg13g2_fill_2 FILLER_71_434 ();
 sg13g2_fill_1 FILLER_71_444 ();
 sg13g2_fill_2 FILLER_71_450 ();
 sg13g2_decap_4 FILLER_71_495 ();
 sg13g2_fill_2 FILLER_71_499 ();
 sg13g2_decap_4 FILLER_71_505 ();
 sg13g2_fill_2 FILLER_71_509 ();
 sg13g2_decap_8 FILLER_71_515 ();
 sg13g2_fill_2 FILLER_71_522 ();
 sg13g2_decap_4 FILLER_71_529 ();
 sg13g2_fill_2 FILLER_71_537 ();
 sg13g2_fill_1 FILLER_71_539 ();
 sg13g2_decap_4 FILLER_71_553 ();
 sg13g2_fill_1 FILLER_71_557 ();
 sg13g2_fill_2 FILLER_71_611 ();
 sg13g2_fill_2 FILLER_71_622 ();
 sg13g2_fill_2 FILLER_71_634 ();
 sg13g2_decap_4 FILLER_71_641 ();
 sg13g2_fill_1 FILLER_71_649 ();
 sg13g2_fill_2 FILLER_71_658 ();
 sg13g2_fill_1 FILLER_71_686 ();
 sg13g2_fill_2 FILLER_71_697 ();
 sg13g2_fill_2 FILLER_71_728 ();
 sg13g2_fill_2 FILLER_71_779 ();
 sg13g2_fill_2 FILLER_71_785 ();
 sg13g2_fill_1 FILLER_71_787 ();
 sg13g2_fill_2 FILLER_71_792 ();
 sg13g2_fill_1 FILLER_71_798 ();
 sg13g2_fill_2 FILLER_71_809 ();
 sg13g2_fill_1 FILLER_71_816 ();
 sg13g2_fill_2 FILLER_71_827 ();
 sg13g2_fill_1 FILLER_71_829 ();
 sg13g2_fill_2 FILLER_71_897 ();
 sg13g2_fill_1 FILLER_71_910 ();
 sg13g2_fill_2 FILLER_71_915 ();
 sg13g2_fill_1 FILLER_71_917 ();
 sg13g2_fill_2 FILLER_71_922 ();
 sg13g2_fill_2 FILLER_71_950 ();
 sg13g2_fill_1 FILLER_71_952 ();
 sg13g2_fill_2 FILLER_71_957 ();
 sg13g2_fill_1 FILLER_71_959 ();
 sg13g2_fill_2 FILLER_71_970 ();
 sg13g2_fill_1 FILLER_71_972 ();
 sg13g2_decap_4 FILLER_71_977 ();
 sg13g2_fill_2 FILLER_71_981 ();
 sg13g2_decap_4 FILLER_71_1027 ();
 sg13g2_fill_1 FILLER_71_1031 ();
 sg13g2_decap_8 FILLER_71_1037 ();
 sg13g2_decap_8 FILLER_71_1044 ();
 sg13g2_decap_8 FILLER_71_1051 ();
 sg13g2_fill_2 FILLER_71_1058 ();
 sg13g2_fill_1 FILLER_71_1060 ();
 sg13g2_fill_1 FILLER_71_1090 ();
 sg13g2_fill_1 FILLER_71_1124 ();
 sg13g2_decap_4 FILLER_71_1129 ();
 sg13g2_fill_2 FILLER_71_1133 ();
 sg13g2_fill_1 FILLER_71_1170 ();
 sg13g2_decap_4 FILLER_71_1188 ();
 sg13g2_fill_1 FILLER_71_1192 ();
 sg13g2_fill_1 FILLER_71_1217 ();
 sg13g2_fill_1 FILLER_71_1228 ();
 sg13g2_decap_4 FILLER_71_1240 ();
 sg13g2_fill_1 FILLER_71_1244 ();
 sg13g2_fill_1 FILLER_71_1272 ();
 sg13g2_decap_8 FILLER_71_1284 ();
 sg13g2_fill_1 FILLER_71_1291 ();
 sg13g2_decap_8 FILLER_71_1296 ();
 sg13g2_decap_8 FILLER_71_1303 ();
 sg13g2_fill_1 FILLER_71_1310 ();
 sg13g2_fill_1 FILLER_71_1332 ();
 sg13g2_fill_2 FILLER_71_1345 ();
 sg13g2_fill_2 FILLER_71_1351 ();
 sg13g2_fill_1 FILLER_71_1353 ();
 sg13g2_fill_1 FILLER_71_1370 ();
 sg13g2_fill_1 FILLER_71_1375 ();
 sg13g2_fill_1 FILLER_71_1380 ();
 sg13g2_fill_2 FILLER_71_1404 ();
 sg13g2_fill_1 FILLER_71_1406 ();
 sg13g2_fill_2 FILLER_71_1412 ();
 sg13g2_decap_4 FILLER_71_1432 ();
 sg13g2_fill_2 FILLER_71_1458 ();
 sg13g2_fill_1 FILLER_71_1464 ();
 sg13g2_fill_2 FILLER_71_1470 ();
 sg13g2_fill_1 FILLER_71_1476 ();
 sg13g2_fill_1 FILLER_71_1488 ();
 sg13g2_decap_4 FILLER_71_1520 ();
 sg13g2_fill_1 FILLER_71_1524 ();
 sg13g2_fill_2 FILLER_71_1547 ();
 sg13g2_fill_1 FILLER_71_1549 ();
 sg13g2_fill_2 FILLER_71_1567 ();
 sg13g2_fill_1 FILLER_71_1583 ();
 sg13g2_decap_4 FILLER_71_1588 ();
 sg13g2_fill_1 FILLER_71_1596 ();
 sg13g2_fill_1 FILLER_71_1601 ();
 sg13g2_decap_4 FILLER_71_1606 ();
 sg13g2_decap_8 FILLER_71_1615 ();
 sg13g2_decap_8 FILLER_71_1622 ();
 sg13g2_decap_4 FILLER_71_1629 ();
 sg13g2_fill_1 FILLER_71_1637 ();
 sg13g2_fill_1 FILLER_71_1669 ();
 sg13g2_decap_8 FILLER_71_1696 ();
 sg13g2_decap_8 FILLER_71_1708 ();
 sg13g2_fill_1 FILLER_71_1741 ();
 sg13g2_fill_1 FILLER_71_1752 ();
 sg13g2_fill_1 FILLER_71_1757 ();
 sg13g2_decap_8 FILLER_71_1790 ();
 sg13g2_fill_2 FILLER_71_1797 ();
 sg13g2_decap_8 FILLER_71_1808 ();
 sg13g2_decap_8 FILLER_71_1829 ();
 sg13g2_fill_2 FILLER_71_1836 ();
 sg13g2_fill_1 FILLER_71_1838 ();
 sg13g2_fill_1 FILLER_71_1849 ();
 sg13g2_fill_1 FILLER_71_1882 ();
 sg13g2_fill_1 FILLER_71_1888 ();
 sg13g2_fill_1 FILLER_71_1916 ();
 sg13g2_decap_4 FILLER_71_1933 ();
 sg13g2_fill_1 FILLER_71_1937 ();
 sg13g2_fill_2 FILLER_71_1942 ();
 sg13g2_fill_1 FILLER_71_1944 ();
 sg13g2_fill_1 FILLER_71_1950 ();
 sg13g2_decap_4 FILLER_71_1964 ();
 sg13g2_fill_1 FILLER_71_1968 ();
 sg13g2_fill_1 FILLER_71_2013 ();
 sg13g2_fill_1 FILLER_71_2020 ();
 sg13g2_fill_2 FILLER_71_2026 ();
 sg13g2_fill_1 FILLER_71_2028 ();
 sg13g2_fill_1 FILLER_71_2041 ();
 sg13g2_fill_1 FILLER_71_2061 ();
 sg13g2_fill_2 FILLER_71_2114 ();
 sg13g2_fill_1 FILLER_71_2116 ();
 sg13g2_decap_8 FILLER_71_2121 ();
 sg13g2_decap_8 FILLER_71_2128 ();
 sg13g2_fill_2 FILLER_71_2135 ();
 sg13g2_decap_8 FILLER_71_2160 ();
 sg13g2_decap_8 FILLER_71_2167 ();
 sg13g2_decap_4 FILLER_71_2174 ();
 sg13g2_fill_1 FILLER_71_2178 ();
 sg13g2_fill_2 FILLER_71_2183 ();
 sg13g2_decap_4 FILLER_71_2195 ();
 sg13g2_fill_1 FILLER_71_2199 ();
 sg13g2_fill_2 FILLER_71_2213 ();
 sg13g2_fill_1 FILLER_71_2215 ();
 sg13g2_decap_8 FILLER_71_2243 ();
 sg13g2_decap_8 FILLER_71_2250 ();
 sg13g2_fill_1 FILLER_71_2257 ();
 sg13g2_decap_8 FILLER_71_2270 ();
 sg13g2_decap_8 FILLER_71_2277 ();
 sg13g2_fill_2 FILLER_71_2284 ();
 sg13g2_fill_1 FILLER_71_2286 ();
 sg13g2_decap_8 FILLER_71_2292 ();
 sg13g2_decap_8 FILLER_71_2303 ();
 sg13g2_fill_2 FILLER_71_2310 ();
 sg13g2_decap_4 FILLER_71_2318 ();
 sg13g2_fill_1 FILLER_71_2342 ();
 sg13g2_fill_1 FILLER_71_2353 ();
 sg13g2_fill_2 FILLER_71_2360 ();
 sg13g2_fill_1 FILLER_71_2388 ();
 sg13g2_decap_4 FILLER_71_2395 ();
 sg13g2_decap_4 FILLER_71_2405 ();
 sg13g2_fill_1 FILLER_71_2409 ();
 sg13g2_decap_4 FILLER_71_2433 ();
 sg13g2_fill_2 FILLER_71_2437 ();
 sg13g2_decap_8 FILLER_71_2454 ();
 sg13g2_decap_4 FILLER_71_2461 ();
 sg13g2_fill_2 FILLER_71_2465 ();
 sg13g2_decap_4 FILLER_71_2499 ();
 sg13g2_fill_2 FILLER_71_2503 ();
 sg13g2_decap_8 FILLER_71_2515 ();
 sg13g2_fill_1 FILLER_71_2522 ();
 sg13g2_decap_8 FILLER_71_2559 ();
 sg13g2_decap_8 FILLER_71_2566 ();
 sg13g2_decap_8 FILLER_71_2573 ();
 sg13g2_decap_8 FILLER_71_2580 ();
 sg13g2_decap_8 FILLER_71_2587 ();
 sg13g2_decap_8 FILLER_71_2594 ();
 sg13g2_decap_8 FILLER_71_2601 ();
 sg13g2_decap_8 FILLER_71_2608 ();
 sg13g2_decap_8 FILLER_71_2615 ();
 sg13g2_decap_8 FILLER_71_2622 ();
 sg13g2_decap_8 FILLER_71_2629 ();
 sg13g2_decap_8 FILLER_71_2636 ();
 sg13g2_decap_8 FILLER_71_2643 ();
 sg13g2_decap_8 FILLER_71_2650 ();
 sg13g2_decap_8 FILLER_71_2657 ();
 sg13g2_decap_4 FILLER_71_2664 ();
 sg13g2_fill_2 FILLER_71_2668 ();
 sg13g2_fill_2 FILLER_72_0 ();
 sg13g2_fill_2 FILLER_72_40 ();
 sg13g2_fill_1 FILLER_72_42 ();
 sg13g2_decap_4 FILLER_72_57 ();
 sg13g2_fill_2 FILLER_72_61 ();
 sg13g2_fill_2 FILLER_72_67 ();
 sg13g2_fill_1 FILLER_72_69 ();
 sg13g2_fill_2 FILLER_72_106 ();
 sg13g2_fill_1 FILLER_72_108 ();
 sg13g2_fill_2 FILLER_72_114 ();
 sg13g2_fill_2 FILLER_72_120 ();
 sg13g2_fill_2 FILLER_72_148 ();
 sg13g2_fill_1 FILLER_72_150 ();
 sg13g2_decap_4 FILLER_72_161 ();
 sg13g2_fill_2 FILLER_72_165 ();
 sg13g2_decap_8 FILLER_72_193 ();
 sg13g2_fill_2 FILLER_72_200 ();
 sg13g2_fill_1 FILLER_72_202 ();
 sg13g2_decap_8 FILLER_72_207 ();
 sg13g2_decap_4 FILLER_72_214 ();
 sg13g2_decap_8 FILLER_72_244 ();
 sg13g2_decap_8 FILLER_72_251 ();
 sg13g2_fill_2 FILLER_72_258 ();
 sg13g2_fill_1 FILLER_72_275 ();
 sg13g2_decap_8 FILLER_72_291 ();
 sg13g2_fill_2 FILLER_72_348 ();
 sg13g2_fill_2 FILLER_72_364 ();
 sg13g2_decap_8 FILLER_72_392 ();
 sg13g2_decap_8 FILLER_72_399 ();
 sg13g2_decap_4 FILLER_72_406 ();
 sg13g2_fill_2 FILLER_72_449 ();
 sg13g2_decap_8 FILLER_72_494 ();
 sg13g2_fill_2 FILLER_72_501 ();
 sg13g2_fill_1 FILLER_72_503 ();
 sg13g2_fill_2 FILLER_72_534 ();
 sg13g2_fill_1 FILLER_72_545 ();
 sg13g2_fill_2 FILLER_72_550 ();
 sg13g2_fill_2 FILLER_72_576 ();
 sg13g2_fill_2 FILLER_72_594 ();
 sg13g2_fill_1 FILLER_72_599 ();
 sg13g2_fill_1 FILLER_72_620 ();
 sg13g2_decap_8 FILLER_72_651 ();
 sg13g2_fill_1 FILLER_72_734 ();
 sg13g2_decap_4 FILLER_72_779 ();
 sg13g2_fill_2 FILLER_72_783 ();
 sg13g2_fill_2 FILLER_72_798 ();
 sg13g2_fill_1 FILLER_72_800 ();
 sg13g2_fill_2 FILLER_72_807 ();
 sg13g2_fill_1 FILLER_72_809 ();
 sg13g2_fill_1 FILLER_72_836 ();
 sg13g2_fill_2 FILLER_72_841 ();
 sg13g2_fill_1 FILLER_72_843 ();
 sg13g2_decap_4 FILLER_72_864 ();
 sg13g2_fill_2 FILLER_72_868 ();
 sg13g2_fill_2 FILLER_72_875 ();
 sg13g2_fill_2 FILLER_72_893 ();
 sg13g2_decap_4 FILLER_72_905 ();
 sg13g2_fill_2 FILLER_72_909 ();
 sg13g2_fill_1 FILLER_72_915 ();
 sg13g2_fill_2 FILLER_72_922 ();
 sg13g2_fill_2 FILLER_72_934 ();
 sg13g2_fill_2 FILLER_72_940 ();
 sg13g2_fill_1 FILLER_72_942 ();
 sg13g2_decap_8 FILLER_72_947 ();
 sg13g2_fill_2 FILLER_72_954 ();
 sg13g2_decap_4 FILLER_72_1003 ();
 sg13g2_fill_1 FILLER_72_1007 ();
 sg13g2_decap_8 FILLER_72_1044 ();
 sg13g2_decap_8 FILLER_72_1051 ();
 sg13g2_fill_2 FILLER_72_1058 ();
 sg13g2_fill_1 FILLER_72_1060 ();
 sg13g2_decap_4 FILLER_72_1066 ();
 sg13g2_fill_2 FILLER_72_1070 ();
 sg13g2_decap_8 FILLER_72_1076 ();
 sg13g2_decap_8 FILLER_72_1114 ();
 sg13g2_decap_8 FILLER_72_1121 ();
 sg13g2_decap_4 FILLER_72_1136 ();
 sg13g2_fill_1 FILLER_72_1140 ();
 sg13g2_decap_8 FILLER_72_1150 ();
 sg13g2_decap_8 FILLER_72_1157 ();
 sg13g2_fill_2 FILLER_72_1164 ();
 sg13g2_fill_1 FILLER_72_1166 ();
 sg13g2_fill_1 FILLER_72_1172 ();
 sg13g2_decap_4 FILLER_72_1192 ();
 sg13g2_fill_1 FILLER_72_1204 ();
 sg13g2_fill_2 FILLER_72_1214 ();
 sg13g2_fill_1 FILLER_72_1228 ();
 sg13g2_decap_8 FILLER_72_1240 ();
 sg13g2_decap_8 FILLER_72_1247 ();
 sg13g2_fill_2 FILLER_72_1254 ();
 sg13g2_fill_1 FILLER_72_1256 ();
 sg13g2_fill_2 FILLER_72_1265 ();
 sg13g2_decap_8 FILLER_72_1272 ();
 sg13g2_decap_8 FILLER_72_1279 ();
 sg13g2_decap_8 FILLER_72_1286 ();
 sg13g2_decap_8 FILLER_72_1293 ();
 sg13g2_decap_8 FILLER_72_1300 ();
 sg13g2_decap_8 FILLER_72_1307 ();
 sg13g2_fill_2 FILLER_72_1314 ();
 sg13g2_fill_1 FILLER_72_1316 ();
 sg13g2_fill_1 FILLER_72_1351 ();
 sg13g2_fill_1 FILLER_72_1356 ();
 sg13g2_decap_8 FILLER_72_1362 ();
 sg13g2_decap_4 FILLER_72_1382 ();
 sg13g2_fill_1 FILLER_72_1390 ();
 sg13g2_decap_8 FILLER_72_1408 ();
 sg13g2_decap_4 FILLER_72_1415 ();
 sg13g2_decap_4 FILLER_72_1423 ();
 sg13g2_fill_2 FILLER_72_1427 ();
 sg13g2_fill_1 FILLER_72_1437 ();
 sg13g2_decap_4 FILLER_72_1443 ();
 sg13g2_fill_1 FILLER_72_1447 ();
 sg13g2_fill_2 FILLER_72_1459 ();
 sg13g2_fill_2 FILLER_72_1482 ();
 sg13g2_decap_4 FILLER_72_1489 ();
 sg13g2_fill_2 FILLER_72_1502 ();
 sg13g2_fill_1 FILLER_72_1504 ();
 sg13g2_fill_2 FILLER_72_1517 ();
 sg13g2_fill_1 FILLER_72_1519 ();
 sg13g2_decap_4 FILLER_72_1534 ();
 sg13g2_fill_1 FILLER_72_1586 ();
 sg13g2_decap_4 FILLER_72_1601 ();
 sg13g2_fill_1 FILLER_72_1605 ();
 sg13g2_decap_4 FILLER_72_1618 ();
 sg13g2_decap_4 FILLER_72_1626 ();
 sg13g2_fill_2 FILLER_72_1630 ();
 sg13g2_fill_2 FILLER_72_1658 ();
 sg13g2_decap_8 FILLER_72_1691 ();
 sg13g2_fill_1 FILLER_72_1698 ();
 sg13g2_decap_8 FILLER_72_1729 ();
 sg13g2_decap_4 FILLER_72_1736 ();
 sg13g2_fill_1 FILLER_72_1740 ();
 sg13g2_fill_1 FILLER_72_1747 ();
 sg13g2_decap_4 FILLER_72_1758 ();
 sg13g2_fill_2 FILLER_72_1788 ();
 sg13g2_decap_4 FILLER_72_1800 ();
 sg13g2_fill_1 FILLER_72_1835 ();
 sg13g2_decap_8 FILLER_72_1842 ();
 sg13g2_decap_8 FILLER_72_1849 ();
 sg13g2_fill_1 FILLER_72_1856 ();
 sg13g2_fill_1 FILLER_72_1872 ();
 sg13g2_fill_2 FILLER_72_1885 ();
 sg13g2_fill_2 FILLER_72_1895 ();
 sg13g2_fill_1 FILLER_72_1897 ();
 sg13g2_fill_1 FILLER_72_1924 ();
 sg13g2_fill_2 FILLER_72_1929 ();
 sg13g2_fill_1 FILLER_72_1931 ();
 sg13g2_decap_8 FILLER_72_1962 ();
 sg13g2_decap_4 FILLER_72_1969 ();
 sg13g2_fill_1 FILLER_72_1973 ();
 sg13g2_decap_4 FILLER_72_1978 ();
 sg13g2_fill_1 FILLER_72_1982 ();
 sg13g2_fill_2 FILLER_72_1988 ();
 sg13g2_fill_1 FILLER_72_1990 ();
 sg13g2_decap_4 FILLER_72_1995 ();
 sg13g2_fill_1 FILLER_72_1999 ();
 sg13g2_fill_2 FILLER_72_2010 ();
 sg13g2_fill_1 FILLER_72_2046 ();
 sg13g2_fill_1 FILLER_72_2073 ();
 sg13g2_fill_1 FILLER_72_2079 ();
 sg13g2_fill_1 FILLER_72_2096 ();
 sg13g2_fill_1 FILLER_72_2106 ();
 sg13g2_fill_2 FILLER_72_2125 ();
 sg13g2_decap_8 FILLER_72_2132 ();
 sg13g2_decap_4 FILLER_72_2139 ();
 sg13g2_fill_2 FILLER_72_2143 ();
 sg13g2_fill_2 FILLER_72_2149 ();
 sg13g2_fill_2 FILLER_72_2159 ();
 sg13g2_fill_1 FILLER_72_2161 ();
 sg13g2_fill_2 FILLER_72_2172 ();
 sg13g2_fill_2 FILLER_72_2200 ();
 sg13g2_fill_2 FILLER_72_2218 ();
 sg13g2_fill_1 FILLER_72_2220 ();
 sg13g2_decap_4 FILLER_72_2227 ();
 sg13g2_fill_2 FILLER_72_2241 ();
 sg13g2_decap_8 FILLER_72_2247 ();
 sg13g2_fill_1 FILLER_72_2254 ();
 sg13g2_fill_2 FILLER_72_2281 ();
 sg13g2_decap_8 FILLER_72_2289 ();
 sg13g2_decap_8 FILLER_72_2296 ();
 sg13g2_decap_4 FILLER_72_2303 ();
 sg13g2_fill_1 FILLER_72_2307 ();
 sg13g2_fill_1 FILLER_72_2334 ();
 sg13g2_fill_1 FILLER_72_2339 ();
 sg13g2_fill_2 FILLER_72_2348 ();
 sg13g2_decap_4 FILLER_72_2360 ();
 sg13g2_fill_2 FILLER_72_2373 ();
 sg13g2_fill_1 FILLER_72_2375 ();
 sg13g2_decap_4 FILLER_72_2380 ();
 sg13g2_fill_1 FILLER_72_2384 ();
 sg13g2_fill_1 FILLER_72_2395 ();
 sg13g2_fill_1 FILLER_72_2406 ();
 sg13g2_fill_1 FILLER_72_2417 ();
 sg13g2_decap_4 FILLER_72_2454 ();
 sg13g2_fill_2 FILLER_72_2458 ();
 sg13g2_fill_2 FILLER_72_2496 ();
 sg13g2_decap_8 FILLER_72_2564 ();
 sg13g2_decap_8 FILLER_72_2571 ();
 sg13g2_decap_8 FILLER_72_2578 ();
 sg13g2_decap_8 FILLER_72_2585 ();
 sg13g2_decap_8 FILLER_72_2592 ();
 sg13g2_decap_8 FILLER_72_2599 ();
 sg13g2_decap_8 FILLER_72_2606 ();
 sg13g2_decap_8 FILLER_72_2613 ();
 sg13g2_decap_8 FILLER_72_2620 ();
 sg13g2_decap_8 FILLER_72_2627 ();
 sg13g2_decap_8 FILLER_72_2634 ();
 sg13g2_decap_8 FILLER_72_2641 ();
 sg13g2_decap_8 FILLER_72_2648 ();
 sg13g2_decap_8 FILLER_72_2655 ();
 sg13g2_decap_8 FILLER_72_2662 ();
 sg13g2_fill_1 FILLER_72_2669 ();
 sg13g2_fill_2 FILLER_73_0 ();
 sg13g2_fill_1 FILLER_73_62 ();
 sg13g2_decap_8 FILLER_73_68 ();
 sg13g2_decap_4 FILLER_73_75 ();
 sg13g2_fill_2 FILLER_73_83 ();
 sg13g2_fill_2 FILLER_73_114 ();
 sg13g2_fill_1 FILLER_73_116 ();
 sg13g2_decap_4 FILLER_73_126 ();
 sg13g2_fill_1 FILLER_73_130 ();
 sg13g2_decap_8 FILLER_73_135 ();
 sg13g2_decap_8 FILLER_73_207 ();
 sg13g2_fill_1 FILLER_73_214 ();
 sg13g2_fill_1 FILLER_73_272 ();
 sg13g2_decap_8 FILLER_73_277 ();
 sg13g2_fill_2 FILLER_73_284 ();
 sg13g2_fill_1 FILLER_73_286 ();
 sg13g2_decap_4 FILLER_73_313 ();
 sg13g2_fill_2 FILLER_73_317 ();
 sg13g2_fill_1 FILLER_73_371 ();
 sg13g2_fill_1 FILLER_73_398 ();
 sg13g2_fill_2 FILLER_73_455 ();
 sg13g2_fill_1 FILLER_73_468 ();
 sg13g2_fill_2 FILLER_73_481 ();
 sg13g2_fill_1 FILLER_73_483 ();
 sg13g2_decap_4 FILLER_73_492 ();
 sg13g2_fill_2 FILLER_73_496 ();
 sg13g2_fill_2 FILLER_73_508 ();
 sg13g2_fill_1 FILLER_73_510 ();
 sg13g2_decap_4 FILLER_73_514 ();
 sg13g2_fill_1 FILLER_73_518 ();
 sg13g2_fill_2 FILLER_73_524 ();
 sg13g2_fill_1 FILLER_73_526 ();
 sg13g2_fill_2 FILLER_73_536 ();
 sg13g2_fill_1 FILLER_73_547 ();
 sg13g2_fill_1 FILLER_73_566 ();
 sg13g2_fill_1 FILLER_73_577 ();
 sg13g2_fill_1 FILLER_73_583 ();
 sg13g2_fill_1 FILLER_73_592 ();
 sg13g2_fill_2 FILLER_73_627 ();
 sg13g2_fill_1 FILLER_73_629 ();
 sg13g2_decap_8 FILLER_73_634 ();
 sg13g2_decap_8 FILLER_73_641 ();
 sg13g2_decap_8 FILLER_73_648 ();
 sg13g2_decap_8 FILLER_73_655 ();
 sg13g2_fill_1 FILLER_73_662 ();
 sg13g2_fill_1 FILLER_73_730 ();
 sg13g2_fill_1 FILLER_73_761 ();
 sg13g2_fill_1 FILLER_73_931 ();
 sg13g2_decap_4 FILLER_73_946 ();
 sg13g2_decap_4 FILLER_73_978 ();
 sg13g2_fill_1 FILLER_73_982 ();
 sg13g2_decap_8 FILLER_73_991 ();
 sg13g2_fill_1 FILLER_73_1003 ();
 sg13g2_fill_2 FILLER_73_1029 ();
 sg13g2_fill_1 FILLER_73_1031 ();
 sg13g2_decap_8 FILLER_73_1040 ();
 sg13g2_decap_8 FILLER_73_1051 ();
 sg13g2_decap_4 FILLER_73_1058 ();
 sg13g2_fill_2 FILLER_73_1088 ();
 sg13g2_fill_2 FILLER_73_1094 ();
 sg13g2_fill_1 FILLER_73_1096 ();
 sg13g2_fill_2 FILLER_73_1101 ();
 sg13g2_fill_1 FILLER_73_1103 ();
 sg13g2_fill_2 FILLER_73_1123 ();
 sg13g2_fill_1 FILLER_73_1125 ();
 sg13g2_fill_2 FILLER_73_1156 ();
 sg13g2_fill_1 FILLER_73_1158 ();
 sg13g2_decap_4 FILLER_73_1168 ();
 sg13g2_fill_2 FILLER_73_1172 ();
 sg13g2_decap_4 FILLER_73_1203 ();
 sg13g2_fill_1 FILLER_73_1207 ();
 sg13g2_fill_2 FILLER_73_1235 ();
 sg13g2_fill_1 FILLER_73_1237 ();
 sg13g2_decap_4 FILLER_73_1242 ();
 sg13g2_fill_2 FILLER_73_1246 ();
 sg13g2_decap_8 FILLER_73_1265 ();
 sg13g2_decap_4 FILLER_73_1272 ();
 sg13g2_fill_2 FILLER_73_1276 ();
 sg13g2_decap_8 FILLER_73_1283 ();
 sg13g2_decap_4 FILLER_73_1298 ();
 sg13g2_decap_4 FILLER_73_1306 ();
 sg13g2_decap_8 FILLER_73_1324 ();
 sg13g2_fill_2 FILLER_73_1331 ();
 sg13g2_fill_1 FILLER_73_1365 ();
 sg13g2_decap_4 FILLER_73_1371 ();
 sg13g2_fill_1 FILLER_73_1375 ();
 sg13g2_fill_2 FILLER_73_1397 ();
 sg13g2_decap_4 FILLER_73_1413 ();
 sg13g2_fill_2 FILLER_73_1417 ();
 sg13g2_fill_1 FILLER_73_1432 ();
 sg13g2_fill_1 FILLER_73_1438 ();
 sg13g2_fill_1 FILLER_73_1443 ();
 sg13g2_fill_1 FILLER_73_1454 ();
 sg13g2_decap_4 FILLER_73_1463 ();
 sg13g2_fill_1 FILLER_73_1471 ();
 sg13g2_fill_1 FILLER_73_1477 ();
 sg13g2_fill_2 FILLER_73_1503 ();
 sg13g2_decap_4 FILLER_73_1510 ();
 sg13g2_fill_2 FILLER_73_1514 ();
 sg13g2_fill_2 FILLER_73_1521 ();
 sg13g2_fill_1 FILLER_73_1523 ();
 sg13g2_decap_4 FILLER_73_1533 ();
 sg13g2_fill_1 FILLER_73_1541 ();
 sg13g2_fill_2 FILLER_73_1547 ();
 sg13g2_decap_4 FILLER_73_1559 ();
 sg13g2_fill_2 FILLER_73_1584 ();
 sg13g2_decap_4 FILLER_73_1590 ();
 sg13g2_fill_2 FILLER_73_1594 ();
 sg13g2_fill_2 FILLER_73_1601 ();
 sg13g2_fill_1 FILLER_73_1603 ();
 sg13g2_decap_4 FILLER_73_1628 ();
 sg13g2_fill_1 FILLER_73_1632 ();
 sg13g2_fill_2 FILLER_73_1637 ();
 sg13g2_fill_1 FILLER_73_1639 ();
 sg13g2_fill_1 FILLER_73_1644 ();
 sg13g2_decap_8 FILLER_73_1649 ();
 sg13g2_decap_8 FILLER_73_1656 ();
 sg13g2_decap_4 FILLER_73_1663 ();
 sg13g2_fill_2 FILLER_73_1667 ();
 sg13g2_decap_8 FILLER_73_1690 ();
 sg13g2_fill_2 FILLER_73_1697 ();
 sg13g2_fill_1 FILLER_73_1699 ();
 sg13g2_fill_2 FILLER_73_1710 ();
 sg13g2_fill_1 FILLER_73_1712 ();
 sg13g2_decap_8 FILLER_73_1854 ();
 sg13g2_fill_2 FILLER_73_1861 ();
 sg13g2_decap_4 FILLER_73_1868 ();
 sg13g2_fill_2 FILLER_73_1872 ();
 sg13g2_fill_2 FILLER_73_1879 ();
 sg13g2_fill_1 FILLER_73_1881 ();
 sg13g2_fill_1 FILLER_73_1886 ();
 sg13g2_fill_1 FILLER_73_1913 ();
 sg13g2_fill_2 FILLER_73_1924 ();
 sg13g2_fill_1 FILLER_73_1926 ();
 sg13g2_decap_8 FILLER_73_1957 ();
 sg13g2_decap_8 FILLER_73_1964 ();
 sg13g2_fill_1 FILLER_73_1971 ();
 sg13g2_fill_1 FILLER_73_2011 ();
 sg13g2_decap_4 FILLER_73_2018 ();
 sg13g2_fill_2 FILLER_73_2022 ();
 sg13g2_fill_1 FILLER_73_2030 ();
 sg13g2_fill_2 FILLER_73_2041 ();
 sg13g2_fill_1 FILLER_73_2043 ();
 sg13g2_fill_2 FILLER_73_2078 ();
 sg13g2_fill_2 FILLER_73_2101 ();
 sg13g2_fill_1 FILLER_73_2103 ();
 sg13g2_decap_8 FILLER_73_2118 ();
 sg13g2_decap_8 FILLER_73_2125 ();
 sg13g2_fill_2 FILLER_73_2136 ();
 sg13g2_fill_1 FILLER_73_2138 ();
 sg13g2_fill_1 FILLER_73_2169 ();
 sg13g2_fill_2 FILLER_73_2338 ();
 sg13g2_fill_1 FILLER_73_2366 ();
 sg13g2_fill_1 FILLER_73_2373 ();
 sg13g2_decap_4 FILLER_73_2506 ();
 sg13g2_fill_2 FILLER_73_2510 ();
 sg13g2_fill_2 FILLER_73_2516 ();
 sg13g2_fill_1 FILLER_73_2518 ();
 sg13g2_fill_2 FILLER_73_2524 ();
 sg13g2_fill_1 FILLER_73_2526 ();
 sg13g2_fill_2 FILLER_73_2541 ();
 sg13g2_fill_1 FILLER_73_2543 ();
 sg13g2_decap_8 FILLER_73_2548 ();
 sg13g2_decap_8 FILLER_73_2555 ();
 sg13g2_decap_8 FILLER_73_2562 ();
 sg13g2_decap_8 FILLER_73_2569 ();
 sg13g2_decap_8 FILLER_73_2576 ();
 sg13g2_decap_8 FILLER_73_2583 ();
 sg13g2_decap_8 FILLER_73_2590 ();
 sg13g2_decap_8 FILLER_73_2597 ();
 sg13g2_decap_8 FILLER_73_2604 ();
 sg13g2_decap_8 FILLER_73_2611 ();
 sg13g2_decap_8 FILLER_73_2618 ();
 sg13g2_decap_8 FILLER_73_2625 ();
 sg13g2_decap_8 FILLER_73_2632 ();
 sg13g2_decap_8 FILLER_73_2639 ();
 sg13g2_decap_8 FILLER_73_2646 ();
 sg13g2_decap_8 FILLER_73_2653 ();
 sg13g2_decap_8 FILLER_73_2660 ();
 sg13g2_fill_2 FILLER_73_2667 ();
 sg13g2_fill_1 FILLER_73_2669 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_4 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_61 ();
 sg13g2_decap_8 FILLER_74_68 ();
 sg13g2_fill_2 FILLER_74_75 ();
 sg13g2_fill_1 FILLER_74_107 ();
 sg13g2_decap_8 FILLER_74_121 ();
 sg13g2_decap_8 FILLER_74_128 ();
 sg13g2_decap_8 FILLER_74_135 ();
 sg13g2_decap_4 FILLER_74_142 ();
 sg13g2_decap_4 FILLER_74_162 ();
 sg13g2_fill_1 FILLER_74_166 ();
 sg13g2_decap_4 FILLER_74_198 ();
 sg13g2_fill_1 FILLER_74_202 ();
 sg13g2_decap_4 FILLER_74_208 ();
 sg13g2_decap_8 FILLER_74_241 ();
 sg13g2_decap_4 FILLER_74_248 ();
 sg13g2_fill_2 FILLER_74_252 ();
 sg13g2_decap_4 FILLER_74_264 ();
 sg13g2_fill_2 FILLER_74_268 ();
 sg13g2_decap_8 FILLER_74_274 ();
 sg13g2_decap_8 FILLER_74_281 ();
 sg13g2_decap_4 FILLER_74_288 ();
 sg13g2_fill_2 FILLER_74_292 ();
 sg13g2_fill_2 FILLER_74_298 ();
 sg13g2_fill_2 FILLER_74_379 ();
 sg13g2_decap_8 FILLER_74_390 ();
 sg13g2_decap_8 FILLER_74_397 ();
 sg13g2_fill_2 FILLER_74_404 ();
 sg13g2_fill_1 FILLER_74_437 ();
 sg13g2_fill_2 FILLER_74_442 ();
 sg13g2_decap_8 FILLER_74_484 ();
 sg13g2_decap_8 FILLER_74_491 ();
 sg13g2_decap_8 FILLER_74_498 ();
 sg13g2_fill_1 FILLER_74_505 ();
 sg13g2_fill_2 FILLER_74_535 ();
 sg13g2_fill_2 FILLER_74_546 ();
 sg13g2_fill_1 FILLER_74_548 ();
 sg13g2_fill_2 FILLER_74_560 ();
 sg13g2_fill_1 FILLER_74_562 ();
 sg13g2_fill_1 FILLER_74_623 ();
 sg13g2_decap_8 FILLER_74_654 ();
 sg13g2_decap_8 FILLER_74_661 ();
 sg13g2_decap_4 FILLER_74_668 ();
 sg13g2_fill_2 FILLER_74_696 ();
 sg13g2_fill_2 FILLER_74_703 ();
 sg13g2_fill_1 FILLER_74_705 ();
 sg13g2_fill_2 FILLER_74_732 ();
 sg13g2_fill_2 FILLER_74_744 ();
 sg13g2_fill_1 FILLER_74_746 ();
 sg13g2_fill_1 FILLER_74_773 ();
 sg13g2_fill_1 FILLER_74_778 ();
 sg13g2_fill_1 FILLER_74_783 ();
 sg13g2_fill_1 FILLER_74_810 ();
 sg13g2_fill_2 FILLER_74_817 ();
 sg13g2_fill_1 FILLER_74_819 ();
 sg13g2_fill_1 FILLER_74_847 ();
 sg13g2_fill_2 FILLER_74_887 ();
 sg13g2_fill_1 FILLER_74_889 ();
 sg13g2_fill_2 FILLER_74_920 ();
 sg13g2_fill_1 FILLER_74_927 ();
 sg13g2_decap_8 FILLER_74_972 ();
 sg13g2_fill_1 FILLER_74_979 ();
 sg13g2_fill_2 FILLER_74_996 ();
 sg13g2_fill_2 FILLER_74_1047 ();
 sg13g2_fill_1 FILLER_74_1049 ();
 sg13g2_fill_1 FILLER_74_1063 ();
 sg13g2_fill_2 FILLER_74_1073 ();
 sg13g2_decap_8 FILLER_74_1079 ();
 sg13g2_decap_8 FILLER_74_1086 ();
 sg13g2_decap_8 FILLER_74_1093 ();
 sg13g2_decap_8 FILLER_74_1100 ();
 sg13g2_decap_8 FILLER_74_1107 ();
 sg13g2_fill_1 FILLER_74_1114 ();
 sg13g2_decap_4 FILLER_74_1123 ();
 sg13g2_fill_2 FILLER_74_1153 ();
 sg13g2_fill_1 FILLER_74_1155 ();
 sg13g2_fill_1 FILLER_74_1184 ();
 sg13g2_fill_1 FILLER_74_1190 ();
 sg13g2_decap_4 FILLER_74_1232 ();
 sg13g2_fill_1 FILLER_74_1249 ();
 sg13g2_decap_8 FILLER_74_1269 ();
 sg13g2_decap_8 FILLER_74_1276 ();
 sg13g2_fill_2 FILLER_74_1283 ();
 sg13g2_fill_2 FILLER_74_1290 ();
 sg13g2_fill_2 FILLER_74_1304 ();
 sg13g2_decap_8 FILLER_74_1322 ();
 sg13g2_decap_8 FILLER_74_1329 ();
 sg13g2_decap_8 FILLER_74_1336 ();
 sg13g2_fill_2 FILLER_74_1343 ();
 sg13g2_fill_1 FILLER_74_1345 ();
 sg13g2_decap_4 FILLER_74_1371 ();
 sg13g2_fill_2 FILLER_74_1375 ();
 sg13g2_decap_8 FILLER_74_1383 ();
 sg13g2_decap_8 FILLER_74_1390 ();
 sg13g2_decap_4 FILLER_74_1397 ();
 sg13g2_fill_2 FILLER_74_1412 ();
 sg13g2_fill_1 FILLER_74_1414 ();
 sg13g2_fill_1 FILLER_74_1419 ();
 sg13g2_decap_8 FILLER_74_1425 ();
 sg13g2_fill_1 FILLER_74_1432 ();
 sg13g2_fill_1 FILLER_74_1437 ();
 sg13g2_fill_2 FILLER_74_1443 ();
 sg13g2_fill_1 FILLER_74_1445 ();
 sg13g2_decap_4 FILLER_74_1456 ();
 sg13g2_fill_1 FILLER_74_1460 ();
 sg13g2_fill_2 FILLER_74_1478 ();
 sg13g2_fill_1 FILLER_74_1480 ();
 sg13g2_fill_2 FILLER_74_1518 ();
 sg13g2_fill_2 FILLER_74_1531 ();
 sg13g2_fill_1 FILLER_74_1537 ();
 sg13g2_fill_1 FILLER_74_1550 ();
 sg13g2_decap_8 FILLER_74_1555 ();
 sg13g2_decap_4 FILLER_74_1562 ();
 sg13g2_fill_1 FILLER_74_1581 ();
 sg13g2_decap_4 FILLER_74_1607 ();
 sg13g2_fill_2 FILLER_74_1617 ();
 sg13g2_fill_1 FILLER_74_1619 ();
 sg13g2_fill_1 FILLER_74_1651 ();
 sg13g2_fill_2 FILLER_74_1656 ();
 sg13g2_fill_1 FILLER_74_1658 ();
 sg13g2_decap_4 FILLER_74_1695 ();
 sg13g2_fill_1 FILLER_74_1699 ();
 sg13g2_decap_4 FILLER_74_1705 ();
 sg13g2_fill_2 FILLER_74_1719 ();
 sg13g2_decap_8 FILLER_74_1735 ();
 sg13g2_fill_1 FILLER_74_1742 ();
 sg13g2_fill_2 FILLER_74_1747 ();
 sg13g2_fill_1 FILLER_74_1749 ();
 sg13g2_fill_2 FILLER_74_1755 ();
 sg13g2_fill_2 FILLER_74_1763 ();
 sg13g2_fill_1 FILLER_74_1765 ();
 sg13g2_fill_2 FILLER_74_1776 ();
 sg13g2_fill_1 FILLER_74_1825 ();
 sg13g2_fill_1 FILLER_74_1830 ();
 sg13g2_fill_2 FILLER_74_1887 ();
 sg13g2_fill_1 FILLER_74_1900 ();
 sg13g2_fill_1 FILLER_74_1911 ();
 sg13g2_fill_2 FILLER_74_1930 ();
 sg13g2_fill_1 FILLER_74_1932 ();
 sg13g2_fill_2 FILLER_74_1966 ();
 sg13g2_fill_2 FILLER_74_1973 ();
 sg13g2_fill_1 FILLER_74_1979 ();
 sg13g2_fill_2 FILLER_74_2006 ();
 sg13g2_decap_4 FILLER_74_2034 ();
 sg13g2_fill_2 FILLER_74_2038 ();
 sg13g2_decap_4 FILLER_74_2046 ();
 sg13g2_decap_8 FILLER_74_2060 ();
 sg13g2_fill_2 FILLER_74_2092 ();
 sg13g2_fill_1 FILLER_74_2094 ();
 sg13g2_fill_2 FILLER_74_2121 ();
 sg13g2_decap_8 FILLER_74_2195 ();
 sg13g2_fill_2 FILLER_74_2202 ();
 sg13g2_fill_1 FILLER_74_2204 ();
 sg13g2_fill_2 FILLER_74_2209 ();
 sg13g2_fill_1 FILLER_74_2211 ();
 sg13g2_fill_1 FILLER_74_2218 ();
 sg13g2_fill_1 FILLER_74_2269 ();
 sg13g2_fill_2 FILLER_74_2320 ();
 sg13g2_fill_2 FILLER_74_2458 ();
 sg13g2_fill_1 FILLER_74_2460 ();
 sg13g2_decap_8 FILLER_74_2503 ();
 sg13g2_decap_4 FILLER_74_2510 ();
 sg13g2_fill_2 FILLER_74_2514 ();
 sg13g2_decap_8 FILLER_74_2533 ();
 sg13g2_decap_8 FILLER_74_2540 ();
 sg13g2_decap_8 FILLER_74_2547 ();
 sg13g2_decap_8 FILLER_74_2554 ();
 sg13g2_decap_8 FILLER_74_2561 ();
 sg13g2_decap_8 FILLER_74_2568 ();
 sg13g2_decap_8 FILLER_74_2575 ();
 sg13g2_decap_8 FILLER_74_2582 ();
 sg13g2_decap_8 FILLER_74_2589 ();
 sg13g2_decap_8 FILLER_74_2596 ();
 sg13g2_decap_8 FILLER_74_2603 ();
 sg13g2_decap_8 FILLER_74_2610 ();
 sg13g2_decap_8 FILLER_74_2617 ();
 sg13g2_decap_8 FILLER_74_2624 ();
 sg13g2_decap_8 FILLER_74_2631 ();
 sg13g2_decap_8 FILLER_74_2638 ();
 sg13g2_decap_8 FILLER_74_2645 ();
 sg13g2_decap_8 FILLER_74_2652 ();
 sg13g2_decap_8 FILLER_74_2659 ();
 sg13g2_decap_4 FILLER_74_2666 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_fill_1 FILLER_75_14 ();
 sg13g2_fill_1 FILLER_75_38 ();
 sg13g2_fill_1 FILLER_75_55 ();
 sg13g2_decap_8 FILLER_75_61 ();
 sg13g2_fill_2 FILLER_75_68 ();
 sg13g2_fill_1 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_114 ();
 sg13g2_decap_4 FILLER_75_121 ();
 sg13g2_decap_4 FILLER_75_135 ();
 sg13g2_fill_2 FILLER_75_169 ();
 sg13g2_fill_1 FILLER_75_191 ();
 sg13g2_fill_2 FILLER_75_203 ();
 sg13g2_decap_4 FILLER_75_209 ();
 sg13g2_fill_2 FILLER_75_213 ();
 sg13g2_fill_1 FILLER_75_241 ();
 sg13g2_decap_8 FILLER_75_293 ();
 sg13g2_fill_2 FILLER_75_300 ();
 sg13g2_decap_4 FILLER_75_305 ();
 sg13g2_fill_1 FILLER_75_309 ();
 sg13g2_decap_8 FILLER_75_320 ();
 sg13g2_decap_4 FILLER_75_331 ();
 sg13g2_decap_8 FILLER_75_365 ();
 sg13g2_decap_8 FILLER_75_372 ();
 sg13g2_decap_8 FILLER_75_379 ();
 sg13g2_decap_8 FILLER_75_386 ();
 sg13g2_decap_8 FILLER_75_393 ();
 sg13g2_decap_8 FILLER_75_400 ();
 sg13g2_fill_1 FILLER_75_407 ();
 sg13g2_decap_4 FILLER_75_413 ();
 sg13g2_fill_1 FILLER_75_417 ();
 sg13g2_decap_8 FILLER_75_422 ();
 sg13g2_fill_1 FILLER_75_429 ();
 sg13g2_decap_8 FILLER_75_434 ();
 sg13g2_fill_2 FILLER_75_441 ();
 sg13g2_fill_2 FILLER_75_455 ();
 sg13g2_fill_1 FILLER_75_466 ();
 sg13g2_fill_1 FILLER_75_475 ();
 sg13g2_fill_1 FILLER_75_480 ();
 sg13g2_fill_2 FILLER_75_496 ();
 sg13g2_fill_1 FILLER_75_498 ();
 sg13g2_fill_1 FILLER_75_517 ();
 sg13g2_fill_2 FILLER_75_533 ();
 sg13g2_decap_4 FILLER_75_539 ();
 sg13g2_fill_2 FILLER_75_543 ();
 sg13g2_decap_8 FILLER_75_553 ();
 sg13g2_decap_4 FILLER_75_560 ();
 sg13g2_fill_1 FILLER_75_605 ();
 sg13g2_fill_1 FILLER_75_620 ();
 sg13g2_fill_2 FILLER_75_624 ();
 sg13g2_fill_1 FILLER_75_631 ();
 sg13g2_decap_8 FILLER_75_649 ();
 sg13g2_decap_4 FILLER_75_656 ();
 sg13g2_fill_2 FILLER_75_660 ();
 sg13g2_fill_2 FILLER_75_696 ();
 sg13g2_fill_2 FILLER_75_710 ();
 sg13g2_decap_8 FILLER_75_729 ();
 sg13g2_decap_8 FILLER_75_736 ();
 sg13g2_decap_8 FILLER_75_766 ();
 sg13g2_decap_8 FILLER_75_773 ();
 sg13g2_decap_8 FILLER_75_780 ();
 sg13g2_fill_2 FILLER_75_787 ();
 sg13g2_decap_4 FILLER_75_793 ();
 sg13g2_fill_1 FILLER_75_797 ();
 sg13g2_decap_8 FILLER_75_824 ();
 sg13g2_fill_2 FILLER_75_831 ();
 sg13g2_fill_1 FILLER_75_833 ();
 sg13g2_decap_4 FILLER_75_874 ();
 sg13g2_fill_2 FILLER_75_878 ();
 sg13g2_fill_1 FILLER_75_892 ();
 sg13g2_fill_2 FILLER_75_897 ();
 sg13g2_fill_1 FILLER_75_899 ();
 sg13g2_fill_1 FILLER_75_910 ();
 sg13g2_fill_2 FILLER_75_945 ();
 sg13g2_decap_8 FILLER_75_1018 ();
 sg13g2_decap_4 FILLER_75_1099 ();
 sg13g2_decap_8 FILLER_75_1147 ();
 sg13g2_decap_4 FILLER_75_1154 ();
 sg13g2_fill_2 FILLER_75_1169 ();
 sg13g2_fill_1 FILLER_75_1175 ();
 sg13g2_fill_1 FILLER_75_1199 ();
 sg13g2_fill_2 FILLER_75_1205 ();
 sg13g2_fill_2 FILLER_75_1216 ();
 sg13g2_fill_1 FILLER_75_1218 ();
 sg13g2_fill_1 FILLER_75_1229 ();
 sg13g2_decap_8 FILLER_75_1244 ();
 sg13g2_decap_4 FILLER_75_1251 ();
 sg13g2_fill_1 FILLER_75_1285 ();
 sg13g2_decap_4 FILLER_75_1291 ();
 sg13g2_fill_1 FILLER_75_1295 ();
 sg13g2_fill_1 FILLER_75_1302 ();
 sg13g2_fill_1 FILLER_75_1311 ();
 sg13g2_fill_2 FILLER_75_1316 ();
 sg13g2_decap_8 FILLER_75_1331 ();
 sg13g2_decap_8 FILLER_75_1338 ();
 sg13g2_fill_1 FILLER_75_1345 ();
 sg13g2_fill_1 FILLER_75_1373 ();
 sg13g2_decap_8 FILLER_75_1380 ();
 sg13g2_fill_2 FILLER_75_1387 ();
 sg13g2_fill_1 FILLER_75_1389 ();
 sg13g2_decap_4 FILLER_75_1400 ();
 sg13g2_fill_1 FILLER_75_1413 ();
 sg13g2_fill_2 FILLER_75_1451 ();
 sg13g2_fill_2 FILLER_75_1457 ();
 sg13g2_fill_1 FILLER_75_1459 ();
 sg13g2_fill_2 FILLER_75_1470 ();
 sg13g2_fill_1 FILLER_75_1472 ();
 sg13g2_fill_2 FILLER_75_1479 ();
 sg13g2_decap_4 FILLER_75_1495 ();
 sg13g2_fill_2 FILLER_75_1504 ();
 sg13g2_fill_2 FILLER_75_1553 ();
 sg13g2_fill_2 FILLER_75_1571 ();
 sg13g2_fill_1 FILLER_75_1573 ();
 sg13g2_fill_1 FILLER_75_1616 ();
 sg13g2_fill_2 FILLER_75_1621 ();
 sg13g2_fill_1 FILLER_75_1623 ();
 sg13g2_decap_4 FILLER_75_1650 ();
 sg13g2_decap_8 FILLER_75_1658 ();
 sg13g2_fill_1 FILLER_75_1665 ();
 sg13g2_decap_8 FILLER_75_1676 ();
 sg13g2_fill_2 FILLER_75_1683 ();
 sg13g2_decap_8 FILLER_75_1695 ();
 sg13g2_decap_8 FILLER_75_1732 ();
 sg13g2_decap_4 FILLER_75_1739 ();
 sg13g2_fill_1 FILLER_75_1743 ();
 sg13g2_fill_2 FILLER_75_1761 ();
 sg13g2_fill_2 FILLER_75_1773 ();
 sg13g2_fill_1 FILLER_75_1775 ();
 sg13g2_fill_2 FILLER_75_1780 ();
 sg13g2_decap_8 FILLER_75_1788 ();
 sg13g2_decap_8 FILLER_75_1809 ();
 sg13g2_decap_4 FILLER_75_1832 ();
 sg13g2_fill_2 FILLER_75_1836 ();
 sg13g2_decap_4 FILLER_75_1842 ();
 sg13g2_fill_1 FILLER_75_1846 ();
 sg13g2_decap_8 FILLER_75_1853 ();
 sg13g2_decap_4 FILLER_75_1860 ();
 sg13g2_decap_8 FILLER_75_1868 ();
 sg13g2_decap_4 FILLER_75_1875 ();
 sg13g2_fill_2 FILLER_75_1884 ();
 sg13g2_fill_2 FILLER_75_1913 ();
 sg13g2_fill_1 FILLER_75_1915 ();
 sg13g2_fill_2 FILLER_75_1962 ();
 sg13g2_fill_2 FILLER_75_1968 ();
 sg13g2_fill_2 FILLER_75_2000 ();
 sg13g2_fill_1 FILLER_75_2002 ();
 sg13g2_decap_8 FILLER_75_2032 ();
 sg13g2_decap_8 FILLER_75_2039 ();
 sg13g2_decap_8 FILLER_75_2046 ();
 sg13g2_decap_4 FILLER_75_2053 ();
 sg13g2_fill_1 FILLER_75_2057 ();
 sg13g2_fill_2 FILLER_75_2062 ();
 sg13g2_fill_1 FILLER_75_2064 ();
 sg13g2_fill_1 FILLER_75_2069 ();
 sg13g2_fill_2 FILLER_75_2075 ();
 sg13g2_fill_1 FILLER_75_2122 ();
 sg13g2_fill_2 FILLER_75_2132 ();
 sg13g2_decap_8 FILLER_75_2163 ();
 sg13g2_fill_1 FILLER_75_2174 ();
 sg13g2_decap_8 FILLER_75_2189 ();
 sg13g2_decap_8 FILLER_75_2196 ();
 sg13g2_decap_4 FILLER_75_2203 ();
 sg13g2_fill_2 FILLER_75_2207 ();
 sg13g2_decap_4 FILLER_75_2219 ();
 sg13g2_fill_2 FILLER_75_2223 ();
 sg13g2_fill_2 FILLER_75_2233 ();
 sg13g2_fill_1 FILLER_75_2255 ();
 sg13g2_fill_2 FILLER_75_2260 ();
 sg13g2_fill_2 FILLER_75_2266 ();
 sg13g2_fill_1 FILLER_75_2274 ();
 sg13g2_fill_2 FILLER_75_2318 ();
 sg13g2_decap_4 FILLER_75_2361 ();
 sg13g2_decap_4 FILLER_75_2369 ();
 sg13g2_decap_4 FILLER_75_2378 ();
 sg13g2_fill_2 FILLER_75_2382 ();
 sg13g2_fill_1 FILLER_75_2390 ();
 sg13g2_decap_8 FILLER_75_2399 ();
 sg13g2_decap_4 FILLER_75_2406 ();
 sg13g2_fill_1 FILLER_75_2410 ();
 sg13g2_fill_2 FILLER_75_2416 ();
 sg13g2_fill_2 FILLER_75_2424 ();
 sg13g2_decap_8 FILLER_75_2434 ();
 sg13g2_fill_1 FILLER_75_2441 ();
 sg13g2_decap_8 FILLER_75_2446 ();
 sg13g2_fill_1 FILLER_75_2453 ();
 sg13g2_decap_4 FILLER_75_2466 ();
 sg13g2_fill_2 FILLER_75_2470 ();
 sg13g2_fill_1 FILLER_75_2494 ();
 sg13g2_fill_1 FILLER_75_2505 ();
 sg13g2_fill_1 FILLER_75_2512 ();
 sg13g2_decap_8 FILLER_75_2539 ();
 sg13g2_decap_8 FILLER_75_2546 ();
 sg13g2_decap_8 FILLER_75_2553 ();
 sg13g2_decap_8 FILLER_75_2560 ();
 sg13g2_decap_8 FILLER_75_2567 ();
 sg13g2_decap_8 FILLER_75_2574 ();
 sg13g2_decap_8 FILLER_75_2581 ();
 sg13g2_decap_8 FILLER_75_2588 ();
 sg13g2_decap_8 FILLER_75_2595 ();
 sg13g2_decap_8 FILLER_75_2602 ();
 sg13g2_decap_8 FILLER_75_2609 ();
 sg13g2_decap_8 FILLER_75_2616 ();
 sg13g2_decap_8 FILLER_75_2623 ();
 sg13g2_decap_8 FILLER_75_2630 ();
 sg13g2_decap_8 FILLER_75_2637 ();
 sg13g2_decap_8 FILLER_75_2644 ();
 sg13g2_decap_8 FILLER_75_2651 ();
 sg13g2_decap_8 FILLER_75_2658 ();
 sg13g2_decap_4 FILLER_75_2665 ();
 sg13g2_fill_1 FILLER_75_2669 ();
 sg13g2_fill_2 FILLER_76_0 ();
 sg13g2_fill_1 FILLER_76_42 ();
 sg13g2_fill_2 FILLER_76_69 ();
 sg13g2_fill_2 FILLER_76_108 ();
 sg13g2_fill_1 FILLER_76_110 ();
 sg13g2_fill_2 FILLER_76_115 ();
 sg13g2_fill_1 FILLER_76_150 ();
 sg13g2_fill_2 FILLER_76_170 ();
 sg13g2_fill_1 FILLER_76_207 ();
 sg13g2_fill_2 FILLER_76_212 ();
 sg13g2_fill_1 FILLER_76_214 ();
 sg13g2_decap_4 FILLER_76_248 ();
 sg13g2_fill_1 FILLER_76_252 ();
 sg13g2_fill_1 FILLER_76_281 ();
 sg13g2_decap_8 FILLER_76_308 ();
 sg13g2_decap_8 FILLER_76_315 ();
 sg13g2_decap_8 FILLER_76_322 ();
 sg13g2_decap_4 FILLER_76_334 ();
 sg13g2_fill_1 FILLER_76_363 ();
 sg13g2_fill_2 FILLER_76_367 ();
 sg13g2_fill_2 FILLER_76_379 ();
 sg13g2_decap_8 FILLER_76_385 ();
 sg13g2_decap_8 FILLER_76_392 ();
 sg13g2_decap_4 FILLER_76_399 ();
 sg13g2_fill_1 FILLER_76_403 ();
 sg13g2_decap_4 FILLER_76_435 ();
 sg13g2_decap_8 FILLER_76_443 ();
 sg13g2_fill_1 FILLER_76_450 ();
 sg13g2_fill_1 FILLER_76_456 ();
 sg13g2_fill_1 FILLER_76_465 ();
 sg13g2_fill_2 FILLER_76_476 ();
 sg13g2_decap_8 FILLER_76_486 ();
 sg13g2_fill_1 FILLER_76_493 ();
 sg13g2_fill_1 FILLER_76_532 ();
 sg13g2_fill_2 FILLER_76_543 ();
 sg13g2_fill_1 FILLER_76_545 ();
 sg13g2_fill_2 FILLER_76_549 ();
 sg13g2_fill_1 FILLER_76_551 ();
 sg13g2_fill_2 FILLER_76_560 ();
 sg13g2_fill_2 FILLER_76_588 ();
 sg13g2_fill_1 FILLER_76_594 ();
 sg13g2_fill_2 FILLER_76_612 ();
 sg13g2_decap_8 FILLER_76_641 ();
 sg13g2_decap_8 FILLER_76_648 ();
 sg13g2_decap_4 FILLER_76_655 ();
 sg13g2_fill_2 FILLER_76_695 ();
 sg13g2_decap_8 FILLER_76_707 ();
 sg13g2_decap_4 FILLER_76_714 ();
 sg13g2_fill_1 FILLER_76_718 ();
 sg13g2_fill_2 FILLER_76_729 ();
 sg13g2_decap_8 FILLER_76_762 ();
 sg13g2_decap_8 FILLER_76_769 ();
 sg13g2_decap_8 FILLER_76_776 ();
 sg13g2_fill_1 FILLER_76_783 ();
 sg13g2_decap_8 FILLER_76_794 ();
 sg13g2_decap_4 FILLER_76_801 ();
 sg13g2_fill_1 FILLER_76_805 ();
 sg13g2_fill_2 FILLER_76_810 ();
 sg13g2_decap_4 FILLER_76_828 ();
 sg13g2_decap_4 FILLER_76_840 ();
 sg13g2_decap_8 FILLER_76_848 ();
 sg13g2_decap_8 FILLER_76_855 ();
 sg13g2_decap_4 FILLER_76_862 ();
 sg13g2_fill_1 FILLER_76_866 ();
 sg13g2_decap_4 FILLER_76_877 ();
 sg13g2_decap_8 FILLER_76_891 ();
 sg13g2_decap_8 FILLER_76_908 ();
 sg13g2_decap_8 FILLER_76_915 ();
 sg13g2_fill_1 FILLER_76_922 ();
 sg13g2_decap_8 FILLER_76_939 ();
 sg13g2_decap_4 FILLER_76_946 ();
 sg13g2_fill_2 FILLER_76_973 ();
 sg13g2_fill_2 FILLER_76_989 ();
 sg13g2_fill_1 FILLER_76_1014 ();
 sg13g2_decap_8 FILLER_76_1051 ();
 sg13g2_decap_8 FILLER_76_1058 ();
 sg13g2_fill_2 FILLER_76_1065 ();
 sg13g2_fill_1 FILLER_76_1067 ();
 sg13g2_fill_2 FILLER_76_1109 ();
 sg13g2_fill_2 FILLER_76_1136 ();
 sg13g2_decap_8 FILLER_76_1142 ();
 sg13g2_decap_8 FILLER_76_1149 ();
 sg13g2_decap_4 FILLER_76_1156 ();
 sg13g2_decap_8 FILLER_76_1166 ();
 sg13g2_fill_2 FILLER_76_1173 ();
 sg13g2_fill_1 FILLER_76_1175 ();
 sg13g2_fill_1 FILLER_76_1185 ();
 sg13g2_fill_1 FILLER_76_1190 ();
 sg13g2_fill_1 FILLER_76_1195 ();
 sg13g2_fill_2 FILLER_76_1205 ();
 sg13g2_fill_1 FILLER_76_1207 ();
 sg13g2_fill_2 FILLER_76_1215 ();
 sg13g2_fill_1 FILLER_76_1226 ();
 sg13g2_fill_1 FILLER_76_1236 ();
 sg13g2_decap_4 FILLER_76_1250 ();
 sg13g2_fill_1 FILLER_76_1254 ();
 sg13g2_decap_8 FILLER_76_1264 ();
 sg13g2_fill_2 FILLER_76_1271 ();
 sg13g2_fill_2 FILLER_76_1282 ();
 sg13g2_fill_1 FILLER_76_1284 ();
 sg13g2_fill_1 FILLER_76_1297 ();
 sg13g2_fill_1 FILLER_76_1328 ();
 sg13g2_fill_1 FILLER_76_1333 ();
 sg13g2_fill_2 FILLER_76_1344 ();
 sg13g2_fill_1 FILLER_76_1358 ();
 sg13g2_fill_1 FILLER_76_1384 ();
 sg13g2_fill_2 FILLER_76_1423 ();
 sg13g2_fill_1 FILLER_76_1425 ();
 sg13g2_fill_1 FILLER_76_1434 ();
 sg13g2_fill_2 FILLER_76_1440 ();
 sg13g2_fill_1 FILLER_76_1446 ();
 sg13g2_fill_1 FILLER_76_1491 ();
 sg13g2_fill_1 FILLER_76_1548 ();
 sg13g2_fill_2 FILLER_76_1598 ();
 sg13g2_fill_2 FILLER_76_1604 ();
 sg13g2_fill_1 FILLER_76_1606 ();
 sg13g2_decap_4 FILLER_76_1623 ();
 sg13g2_decap_4 FILLER_76_1635 ();
 sg13g2_fill_1 FILLER_76_1639 ();
 sg13g2_decap_4 FILLER_76_1671 ();
 sg13g2_fill_1 FILLER_76_1675 ();
 sg13g2_decap_8 FILLER_76_1686 ();
 sg13g2_fill_2 FILLER_76_1693 ();
 sg13g2_decap_4 FILLER_76_1705 ();
 sg13g2_decap_8 FILLER_76_1749 ();
 sg13g2_decap_8 FILLER_76_1762 ();
 sg13g2_decap_4 FILLER_76_1779 ();
 sg13g2_fill_1 FILLER_76_1809 ();
 sg13g2_fill_2 FILLER_76_1820 ();
 sg13g2_fill_2 FILLER_76_1832 ();
 sg13g2_fill_2 FILLER_76_1840 ();
 sg13g2_fill_1 FILLER_76_1842 ();
 sg13g2_decap_8 FILLER_76_1863 ();
 sg13g2_decap_4 FILLER_76_1870 ();
 sg13g2_fill_1 FILLER_76_1874 ();
 sg13g2_decap_4 FILLER_76_1881 ();
 sg13g2_fill_2 FILLER_76_1890 ();
 sg13g2_decap_4 FILLER_76_1938 ();
 sg13g2_decap_4 FILLER_76_1978 ();
 sg13g2_fill_1 FILLER_76_1982 ();
 sg13g2_fill_1 FILLER_76_2000 ();
 sg13g2_fill_2 FILLER_76_2006 ();
 sg13g2_fill_1 FILLER_76_2008 ();
 sg13g2_fill_1 FILLER_76_2017 ();
 sg13g2_fill_2 FILLER_76_2024 ();
 sg13g2_fill_1 FILLER_76_2026 ();
 sg13g2_fill_1 FILLER_76_2039 ();
 sg13g2_fill_1 FILLER_76_2066 ();
 sg13g2_decap_4 FILLER_76_2096 ();
 sg13g2_fill_1 FILLER_76_2110 ();
 sg13g2_decap_8 FILLER_76_2115 ();
 sg13g2_fill_1 FILLER_76_2122 ();
 sg13g2_fill_1 FILLER_76_2131 ();
 sg13g2_fill_2 FILLER_76_2136 ();
 sg13g2_fill_1 FILLER_76_2142 ();
 sg13g2_decap_8 FILLER_76_2161 ();
 sg13g2_fill_2 FILLER_76_2168 ();
 sg13g2_fill_1 FILLER_76_2170 ();
 sg13g2_decap_8 FILLER_76_2187 ();
 sg13g2_decap_8 FILLER_76_2194 ();
 sg13g2_decap_8 FILLER_76_2201 ();
 sg13g2_decap_8 FILLER_76_2208 ();
 sg13g2_fill_2 FILLER_76_2215 ();
 sg13g2_fill_1 FILLER_76_2217 ();
 sg13g2_fill_2 FILLER_76_2250 ();
 sg13g2_fill_1 FILLER_76_2293 ();
 sg13g2_fill_2 FILLER_76_2303 ();
 sg13g2_fill_2 FILLER_76_2311 ();
 sg13g2_fill_1 FILLER_76_2313 ();
 sg13g2_fill_2 FILLER_76_2320 ();
 sg13g2_fill_1 FILLER_76_2322 ();
 sg13g2_fill_2 FILLER_76_2333 ();
 sg13g2_fill_1 FILLER_76_2335 ();
 sg13g2_decap_8 FILLER_76_2341 ();
 sg13g2_fill_1 FILLER_76_2348 ();
 sg13g2_fill_1 FILLER_76_2354 ();
 sg13g2_decap_8 FILLER_76_2365 ();
 sg13g2_fill_1 FILLER_76_2372 ();
 sg13g2_fill_1 FILLER_76_2377 ();
 sg13g2_decap_8 FILLER_76_2404 ();
 sg13g2_fill_2 FILLER_76_2411 ();
 sg13g2_decap_4 FILLER_76_2423 ();
 sg13g2_decap_4 FILLER_76_2433 ();
 sg13g2_fill_2 FILLER_76_2437 ();
 sg13g2_decap_8 FILLER_76_2449 ();
 sg13g2_decap_8 FILLER_76_2456 ();
 sg13g2_decap_8 FILLER_76_2463 ();
 sg13g2_decap_8 FILLER_76_2470 ();
 sg13g2_fill_2 FILLER_76_2477 ();
 sg13g2_fill_1 FILLER_76_2479 ();
 sg13g2_decap_4 FILLER_76_2490 ();
 sg13g2_decap_8 FILLER_76_2530 ();
 sg13g2_decap_8 FILLER_76_2537 ();
 sg13g2_decap_8 FILLER_76_2544 ();
 sg13g2_decap_8 FILLER_76_2551 ();
 sg13g2_decap_8 FILLER_76_2558 ();
 sg13g2_decap_8 FILLER_76_2565 ();
 sg13g2_decap_8 FILLER_76_2572 ();
 sg13g2_decap_8 FILLER_76_2579 ();
 sg13g2_decap_8 FILLER_76_2586 ();
 sg13g2_decap_8 FILLER_76_2593 ();
 sg13g2_decap_8 FILLER_76_2600 ();
 sg13g2_decap_8 FILLER_76_2607 ();
 sg13g2_decap_8 FILLER_76_2614 ();
 sg13g2_decap_8 FILLER_76_2621 ();
 sg13g2_decap_8 FILLER_76_2628 ();
 sg13g2_decap_8 FILLER_76_2635 ();
 sg13g2_decap_8 FILLER_76_2642 ();
 sg13g2_decap_8 FILLER_76_2649 ();
 sg13g2_decap_8 FILLER_76_2656 ();
 sg13g2_decap_8 FILLER_76_2663 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_fill_2 FILLER_77_7 ();
 sg13g2_decap_4 FILLER_77_13 ();
 sg13g2_fill_2 FILLER_77_42 ();
 sg13g2_fill_2 FILLER_77_61 ();
 sg13g2_fill_1 FILLER_77_63 ();
 sg13g2_fill_1 FILLER_77_90 ();
 sg13g2_fill_1 FILLER_77_99 ();
 sg13g2_fill_1 FILLER_77_105 ();
 sg13g2_fill_2 FILLER_77_114 ();
 sg13g2_fill_2 FILLER_77_152 ();
 sg13g2_fill_2 FILLER_77_203 ();
 sg13g2_decap_8 FILLER_77_218 ();
 sg13g2_decap_4 FILLER_77_251 ();
 sg13g2_fill_2 FILLER_77_255 ();
 sg13g2_fill_1 FILLER_77_281 ();
 sg13g2_fill_2 FILLER_77_300 ();
 sg13g2_fill_1 FILLER_77_318 ();
 sg13g2_decap_8 FILLER_77_323 ();
 sg13g2_fill_1 FILLER_77_335 ();
 sg13g2_fill_2 FILLER_77_371 ();
 sg13g2_fill_1 FILLER_77_373 ();
 sg13g2_fill_2 FILLER_77_417 ();
 sg13g2_fill_1 FILLER_77_445 ();
 sg13g2_fill_1 FILLER_77_476 ();
 sg13g2_fill_2 FILLER_77_606 ();
 sg13g2_decap_8 FILLER_77_639 ();
 sg13g2_decap_8 FILLER_77_646 ();
 sg13g2_decap_8 FILLER_77_653 ();
 sg13g2_fill_1 FILLER_77_660 ();
 sg13g2_decap_8 FILLER_77_669 ();
 sg13g2_decap_8 FILLER_77_676 ();
 sg13g2_decap_8 FILLER_77_683 ();
 sg13g2_decap_4 FILLER_77_716 ();
 sg13g2_fill_1 FILLER_77_750 ();
 sg13g2_decap_8 FILLER_77_777 ();
 sg13g2_fill_2 FILLER_77_784 ();
 sg13g2_decap_4 FILLER_77_812 ();
 sg13g2_fill_1 FILLER_77_816 ();
 sg13g2_decap_4 FILLER_77_827 ();
 sg13g2_decap_8 FILLER_77_857 ();
 sg13g2_fill_2 FILLER_77_894 ();
 sg13g2_fill_1 FILLER_77_896 ();
 sg13g2_fill_2 FILLER_77_928 ();
 sg13g2_decap_4 FILLER_77_966 ();
 sg13g2_fill_1 FILLER_77_970 ();
 sg13g2_fill_2 FILLER_77_1015 ();
 sg13g2_fill_2 FILLER_77_1027 ();
 sg13g2_fill_2 FILLER_77_1037 ();
 sg13g2_decap_8 FILLER_77_1043 ();
 sg13g2_fill_2 FILLER_77_1050 ();
 sg13g2_decap_8 FILLER_77_1056 ();
 sg13g2_decap_8 FILLER_77_1063 ();
 sg13g2_fill_2 FILLER_77_1070 ();
 sg13g2_fill_1 FILLER_77_1072 ();
 sg13g2_fill_1 FILLER_77_1078 ();
 sg13g2_decap_8 FILLER_77_1109 ();
 sg13g2_fill_2 FILLER_77_1116 ();
 sg13g2_fill_2 FILLER_77_1122 ();
 sg13g2_fill_1 FILLER_77_1150 ();
 sg13g2_fill_2 FILLER_77_1156 ();
 sg13g2_fill_1 FILLER_77_1217 ();
 sg13g2_fill_1 FILLER_77_1232 ();
 sg13g2_decap_8 FILLER_77_1249 ();
 sg13g2_decap_8 FILLER_77_1256 ();
 sg13g2_decap_4 FILLER_77_1263 ();
 sg13g2_fill_2 FILLER_77_1307 ();
 sg13g2_fill_1 FILLER_77_1322 ();
 sg13g2_fill_2 FILLER_77_1371 ();
 sg13g2_fill_1 FILLER_77_1379 ();
 sg13g2_fill_1 FILLER_77_1389 ();
 sg13g2_fill_1 FILLER_77_1428 ();
 sg13g2_fill_2 FILLER_77_1448 ();
 sg13g2_fill_1 FILLER_77_1507 ();
 sg13g2_fill_1 FILLER_77_1516 ();
 sg13g2_fill_1 FILLER_77_1548 ();
 sg13g2_fill_1 FILLER_77_1555 ();
 sg13g2_fill_1 FILLER_77_1564 ();
 sg13g2_fill_1 FILLER_77_1571 ();
 sg13g2_fill_1 FILLER_77_1580 ();
 sg13g2_fill_2 FILLER_77_1598 ();
 sg13g2_fill_2 FILLER_77_1612 ();
 sg13g2_fill_1 FILLER_77_1614 ();
 sg13g2_fill_1 FILLER_77_1668 ();
 sg13g2_fill_1 FILLER_77_1673 ();
 sg13g2_fill_2 FILLER_77_1700 ();
 sg13g2_fill_1 FILLER_77_1712 ();
 sg13g2_fill_1 FILLER_77_1740 ();
 sg13g2_decap_4 FILLER_77_1767 ();
 sg13g2_fill_1 FILLER_77_1771 ();
 sg13g2_decap_4 FILLER_77_1896 ();
 sg13g2_decap_4 FILLER_77_1930 ();
 sg13g2_fill_1 FILLER_77_1964 ();
 sg13g2_fill_2 FILLER_77_1969 ();
 sg13g2_fill_2 FILLER_77_2023 ();
 sg13g2_fill_2 FILLER_77_2065 ();
 sg13g2_fill_1 FILLER_77_2067 ();
 sg13g2_fill_2 FILLER_77_2082 ();
 sg13g2_fill_1 FILLER_77_2084 ();
 sg13g2_decap_4 FILLER_77_2122 ();
 sg13g2_fill_1 FILLER_77_2126 ();
 sg13g2_fill_2 FILLER_77_2153 ();
 sg13g2_fill_1 FILLER_77_2155 ();
 sg13g2_fill_1 FILLER_77_2166 ();
 sg13g2_decap_8 FILLER_77_2193 ();
 sg13g2_decap_8 FILLER_77_2200 ();
 sg13g2_fill_2 FILLER_77_2207 ();
 sg13g2_fill_1 FILLER_77_2209 ();
 sg13g2_decap_4 FILLER_77_2220 ();
 sg13g2_decap_8 FILLER_77_2228 ();
 sg13g2_fill_2 FILLER_77_2235 ();
 sg13g2_fill_1 FILLER_77_2237 ();
 sg13g2_decap_8 FILLER_77_2278 ();
 sg13g2_fill_1 FILLER_77_2285 ();
 sg13g2_fill_2 FILLER_77_2312 ();
 sg13g2_fill_1 FILLER_77_2314 ();
 sg13g2_decap_4 FILLER_77_2356 ();
 sg13g2_fill_2 FILLER_77_2386 ();
 sg13g2_fill_1 FILLER_77_2388 ();
 sg13g2_fill_2 FILLER_77_2438 ();
 sg13g2_decap_8 FILLER_77_2480 ();
 sg13g2_fill_1 FILLER_77_2487 ();
 sg13g2_fill_1 FILLER_77_2514 ();
 sg13g2_decap_8 FILLER_77_2519 ();
 sg13g2_decap_8 FILLER_77_2526 ();
 sg13g2_decap_8 FILLER_77_2533 ();
 sg13g2_decap_8 FILLER_77_2540 ();
 sg13g2_decap_8 FILLER_77_2547 ();
 sg13g2_decap_8 FILLER_77_2554 ();
 sg13g2_decap_8 FILLER_77_2561 ();
 sg13g2_decap_8 FILLER_77_2568 ();
 sg13g2_decap_8 FILLER_77_2575 ();
 sg13g2_decap_8 FILLER_77_2582 ();
 sg13g2_decap_8 FILLER_77_2589 ();
 sg13g2_decap_8 FILLER_77_2596 ();
 sg13g2_decap_8 FILLER_77_2603 ();
 sg13g2_decap_8 FILLER_77_2610 ();
 sg13g2_decap_8 FILLER_77_2617 ();
 sg13g2_decap_8 FILLER_77_2624 ();
 sg13g2_decap_8 FILLER_77_2631 ();
 sg13g2_decap_8 FILLER_77_2638 ();
 sg13g2_decap_8 FILLER_77_2645 ();
 sg13g2_decap_8 FILLER_77_2652 ();
 sg13g2_decap_8 FILLER_77_2659 ();
 sg13g2_decap_4 FILLER_77_2666 ();
 sg13g2_fill_1 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_27 ();
 sg13g2_fill_1 FILLER_78_33 ();
 sg13g2_fill_2 FILLER_78_39 ();
 sg13g2_fill_2 FILLER_78_46 ();
 sg13g2_fill_1 FILLER_78_48 ();
 sg13g2_fill_2 FILLER_78_155 ();
 sg13g2_fill_1 FILLER_78_205 ();
 sg13g2_decap_4 FILLER_78_247 ();
 sg13g2_fill_1 FILLER_78_296 ();
 sg13g2_fill_1 FILLER_78_301 ();
 sg13g2_fill_1 FILLER_78_338 ();
 sg13g2_fill_1 FILLER_78_344 ();
 sg13g2_fill_1 FILLER_78_376 ();
 sg13g2_fill_2 FILLER_78_403 ();
 sg13g2_fill_1 FILLER_78_409 ();
 sg13g2_fill_1 FILLER_78_423 ();
 sg13g2_fill_2 FILLER_78_469 ();
 sg13g2_decap_8 FILLER_78_476 ();
 sg13g2_decap_4 FILLER_78_483 ();
 sg13g2_fill_2 FILLER_78_487 ();
 sg13g2_decap_4 FILLER_78_493 ();
 sg13g2_fill_1 FILLER_78_497 ();
 sg13g2_fill_2 FILLER_78_532 ();
 sg13g2_fill_1 FILLER_78_534 ();
 sg13g2_fill_2 FILLER_78_543 ();
 sg13g2_fill_1 FILLER_78_545 ();
 sg13g2_fill_1 FILLER_78_550 ();
 sg13g2_fill_2 FILLER_78_561 ();
 sg13g2_fill_1 FILLER_78_563 ();
 sg13g2_fill_1 FILLER_78_574 ();
 sg13g2_fill_1 FILLER_78_580 ();
 sg13g2_fill_1 FILLER_78_585 ();
 sg13g2_fill_1 FILLER_78_612 ();
 sg13g2_fill_1 FILLER_78_623 ();
 sg13g2_decap_8 FILLER_78_650 ();
 sg13g2_fill_2 FILLER_78_693 ();
 sg13g2_decap_4 FILLER_78_777 ();
 sg13g2_fill_2 FILLER_78_827 ();
 sg13g2_fill_1 FILLER_78_895 ();
 sg13g2_decap_8 FILLER_78_922 ();
 sg13g2_fill_1 FILLER_78_929 ();
 sg13g2_fill_1 FILLER_78_992 ();
 sg13g2_fill_1 FILLER_78_1019 ();
 sg13g2_fill_1 FILLER_78_1024 ();
 sg13g2_decap_4 FILLER_78_1064 ();
 sg13g2_fill_1 FILLER_78_1068 ();
 sg13g2_fill_1 FILLER_78_1157 ();
 sg13g2_fill_1 FILLER_78_1170 ();
 sg13g2_fill_1 FILLER_78_1198 ();
 sg13g2_fill_2 FILLER_78_1204 ();
 sg13g2_fill_1 FILLER_78_1217 ();
 sg13g2_fill_1 FILLER_78_1229 ();
 sg13g2_decap_8 FILLER_78_1254 ();
 sg13g2_decap_4 FILLER_78_1261 ();
 sg13g2_fill_1 FILLER_78_1265 ();
 sg13g2_fill_2 FILLER_78_1270 ();
 sg13g2_fill_1 FILLER_78_1309 ();
 sg13g2_fill_1 FILLER_78_1315 ();
 sg13g2_fill_1 FILLER_78_1324 ();
 sg13g2_decap_4 FILLER_78_1344 ();
 sg13g2_fill_2 FILLER_78_1353 ();
 sg13g2_fill_1 FILLER_78_1355 ();
 sg13g2_fill_1 FILLER_78_1368 ();
 sg13g2_fill_1 FILLER_78_1374 ();
 sg13g2_fill_1 FILLER_78_1384 ();
 sg13g2_decap_4 FILLER_78_1397 ();
 sg13g2_fill_1 FILLER_78_1401 ();
 sg13g2_fill_1 FILLER_78_1431 ();
 sg13g2_fill_1 FILLER_78_1441 ();
 sg13g2_fill_1 FILLER_78_1457 ();
 sg13g2_fill_2 FILLER_78_1463 ();
 sg13g2_fill_1 FILLER_78_1465 ();
 sg13g2_fill_1 FILLER_78_1519 ();
 sg13g2_fill_1 FILLER_78_1534 ();
 sg13g2_fill_1 FILLER_78_1550 ();
 sg13g2_fill_1 FILLER_78_1590 ();
 sg13g2_fill_1 FILLER_78_1601 ();
 sg13g2_decap_8 FILLER_78_1606 ();
 sg13g2_decap_8 FILLER_78_1613 ();
 sg13g2_fill_2 FILLER_78_1620 ();
 sg13g2_fill_1 FILLER_78_1622 ();
 sg13g2_decap_4 FILLER_78_1628 ();
 sg13g2_fill_2 FILLER_78_1636 ();
 sg13g2_fill_1 FILLER_78_1638 ();
 sg13g2_fill_1 FILLER_78_1643 ();
 sg13g2_fill_2 FILLER_78_1703 ();
 sg13g2_fill_2 FILLER_78_1709 ();
 sg13g2_fill_2 FILLER_78_1793 ();
 sg13g2_fill_1 FILLER_78_1795 ();
 sg13g2_fill_1 FILLER_78_1862 ();
 sg13g2_fill_1 FILLER_78_1867 ();
 sg13g2_fill_1 FILLER_78_1899 ();
 sg13g2_fill_1 FILLER_78_1941 ();
 sg13g2_decap_4 FILLER_78_1973 ();
 sg13g2_fill_2 FILLER_78_1982 ();
 sg13g2_fill_1 FILLER_78_1988 ();
 sg13g2_decap_8 FILLER_78_1992 ();
 sg13g2_fill_1 FILLER_78_2051 ();
 sg13g2_fill_2 FILLER_78_2135 ();
 sg13g2_fill_1 FILLER_78_2173 ();
 sg13g2_fill_2 FILLER_78_2178 ();
 sg13g2_fill_1 FILLER_78_2190 ();
 sg13g2_decap_4 FILLER_78_2227 ();
 sg13g2_fill_2 FILLER_78_2231 ();
 sg13g2_decap_8 FILLER_78_2341 ();
 sg13g2_fill_2 FILLER_78_2348 ();
 sg13g2_fill_2 FILLER_78_2376 ();
 sg13g2_fill_1 FILLER_78_2378 ();
 sg13g2_decap_4 FILLER_78_2467 ();
 sg13g2_decap_8 FILLER_78_2475 ();
 sg13g2_fill_2 FILLER_78_2482 ();
 sg13g2_decap_8 FILLER_78_2514 ();
 sg13g2_decap_8 FILLER_78_2521 ();
 sg13g2_decap_8 FILLER_78_2528 ();
 sg13g2_decap_8 FILLER_78_2535 ();
 sg13g2_decap_8 FILLER_78_2542 ();
 sg13g2_decap_8 FILLER_78_2549 ();
 sg13g2_decap_8 FILLER_78_2556 ();
 sg13g2_decap_8 FILLER_78_2563 ();
 sg13g2_decap_8 FILLER_78_2570 ();
 sg13g2_decap_8 FILLER_78_2577 ();
 sg13g2_decap_8 FILLER_78_2584 ();
 sg13g2_decap_8 FILLER_78_2591 ();
 sg13g2_decap_8 FILLER_78_2598 ();
 sg13g2_decap_8 FILLER_78_2605 ();
 sg13g2_decap_8 FILLER_78_2612 ();
 sg13g2_decap_8 FILLER_78_2619 ();
 sg13g2_decap_8 FILLER_78_2626 ();
 sg13g2_decap_8 FILLER_78_2633 ();
 sg13g2_decap_8 FILLER_78_2640 ();
 sg13g2_decap_8 FILLER_78_2647 ();
 sg13g2_decap_8 FILLER_78_2654 ();
 sg13g2_decap_8 FILLER_78_2661 ();
 sg13g2_fill_2 FILLER_78_2668 ();
 sg13g2_decap_4 FILLER_79_0 ();
 sg13g2_fill_2 FILLER_79_34 ();
 sg13g2_fill_1 FILLER_79_36 ();
 sg13g2_decap_8 FILLER_79_71 ();
 sg13g2_fill_1 FILLER_79_78 ();
 sg13g2_fill_1 FILLER_79_87 ();
 sg13g2_fill_1 FILLER_79_119 ();
 sg13g2_fill_1 FILLER_79_130 ();
 sg13g2_fill_2 FILLER_79_135 ();
 sg13g2_fill_2 FILLER_79_194 ();
 sg13g2_fill_1 FILLER_79_202 ();
 sg13g2_decap_4 FILLER_79_246 ();
 sg13g2_fill_1 FILLER_79_250 ();
 sg13g2_fill_1 FILLER_79_300 ();
 sg13g2_decap_4 FILLER_79_327 ();
 sg13g2_fill_1 FILLER_79_331 ();
 sg13g2_decap_8 FILLER_79_337 ();
 sg13g2_decap_8 FILLER_79_344 ();
 sg13g2_decap_8 FILLER_79_364 ();
 sg13g2_decap_8 FILLER_79_371 ();
 sg13g2_decap_8 FILLER_79_378 ();
 sg13g2_fill_1 FILLER_79_385 ();
 sg13g2_decap_8 FILLER_79_390 ();
 sg13g2_fill_1 FILLER_79_397 ();
 sg13g2_decap_8 FILLER_79_429 ();
 sg13g2_fill_1 FILLER_79_436 ();
 sg13g2_fill_2 FILLER_79_441 ();
 sg13g2_fill_1 FILLER_79_469 ();
 sg13g2_fill_1 FILLER_79_475 ();
 sg13g2_fill_2 FILLER_79_502 ();
 sg13g2_fill_2 FILLER_79_508 ();
 sg13g2_fill_2 FILLER_79_620 ();
 sg13g2_fill_2 FILLER_79_655 ();
 sg13g2_decap_4 FILLER_79_693 ();
 sg13g2_fill_2 FILLER_79_697 ();
 sg13g2_fill_2 FILLER_79_725 ();
 sg13g2_fill_1 FILLER_79_727 ();
 sg13g2_fill_2 FILLER_79_754 ();
 sg13g2_fill_1 FILLER_79_797 ();
 sg13g2_fill_1 FILLER_79_802 ();
 sg13g2_fill_2 FILLER_79_813 ();
 sg13g2_fill_2 FILLER_79_841 ();
 sg13g2_decap_4 FILLER_79_853 ();
 sg13g2_fill_2 FILLER_79_857 ();
 sg13g2_decap_8 FILLER_79_956 ();
 sg13g2_decap_8 FILLER_79_963 ();
 sg13g2_fill_2 FILLER_79_970 ();
 sg13g2_decap_8 FILLER_79_980 ();
 sg13g2_fill_1 FILLER_79_987 ();
 sg13g2_fill_1 FILLER_79_1002 ();
 sg13g2_fill_2 FILLER_79_1039 ();
 sg13g2_decap_4 FILLER_79_1067 ();
 sg13g2_fill_2 FILLER_79_1071 ();
 sg13g2_fill_1 FILLER_79_1103 ();
 sg13g2_fill_2 FILLER_79_1108 ();
 sg13g2_fill_2 FILLER_79_1136 ();
 sg13g2_decap_4 FILLER_79_1142 ();
 sg13g2_fill_1 FILLER_79_1146 ();
 sg13g2_fill_2 FILLER_79_1157 ();
 sg13g2_decap_4 FILLER_79_1195 ();
 sg13g2_fill_1 FILLER_79_1203 ();
 sg13g2_fill_1 FILLER_79_1209 ();
 sg13g2_fill_1 FILLER_79_1215 ();
 sg13g2_fill_1 FILLER_79_1239 ();
 sg13g2_decap_8 FILLER_79_1249 ();
 sg13g2_decap_8 FILLER_79_1261 ();
 sg13g2_decap_8 FILLER_79_1268 ();
 sg13g2_decap_4 FILLER_79_1275 ();
 sg13g2_fill_1 FILLER_79_1279 ();
 sg13g2_fill_1 FILLER_79_1305 ();
 sg13g2_fill_2 FILLER_79_1311 ();
 sg13g2_fill_2 FILLER_79_1321 ();
 sg13g2_decap_8 FILLER_79_1332 ();
 sg13g2_decap_8 FILLER_79_1339 ();
 sg13g2_decap_8 FILLER_79_1346 ();
 sg13g2_decap_4 FILLER_79_1353 ();
 sg13g2_fill_2 FILLER_79_1357 ();
 sg13g2_decap_8 FILLER_79_1374 ();
 sg13g2_fill_1 FILLER_79_1381 ();
 sg13g2_decap_8 FILLER_79_1386 ();
 sg13g2_decap_8 FILLER_79_1393 ();
 sg13g2_decap_4 FILLER_79_1400 ();
 sg13g2_fill_2 FILLER_79_1408 ();
 sg13g2_fill_1 FILLER_79_1424 ();
 sg13g2_decap_4 FILLER_79_1438 ();
 sg13g2_fill_1 FILLER_79_1457 ();
 sg13g2_fill_1 FILLER_79_1477 ();
 sg13g2_fill_1 FILLER_79_1514 ();
 sg13g2_fill_1 FILLER_79_1545 ();
 sg13g2_decap_4 FILLER_79_1586 ();
 sg13g2_decap_4 FILLER_79_1595 ();
 sg13g2_fill_2 FILLER_79_1599 ();
 sg13g2_decap_8 FILLER_79_1631 ();
 sg13g2_decap_8 FILLER_79_1638 ();
 sg13g2_decap_8 FILLER_79_1645 ();
 sg13g2_decap_4 FILLER_79_1652 ();
 sg13g2_fill_1 FILLER_79_1656 ();
 sg13g2_decap_8 FILLER_79_1661 ();
 sg13g2_fill_2 FILLER_79_1678 ();
 sg13g2_decap_4 FILLER_79_1690 ();
 sg13g2_fill_1 FILLER_79_1730 ();
 sg13g2_fill_1 FILLER_79_1741 ();
 sg13g2_fill_2 FILLER_79_1746 ();
 sg13g2_fill_1 FILLER_79_1752 ();
 sg13g2_fill_2 FILLER_79_1773 ();
 sg13g2_fill_2 FILLER_79_1785 ();
 sg13g2_fill_2 FILLER_79_1812 ();
 sg13g2_fill_1 FILLER_79_1814 ();
 sg13g2_decap_4 FILLER_79_1833 ();
 sg13g2_fill_2 FILLER_79_1837 ();
 sg13g2_decap_8 FILLER_79_1843 ();
 sg13g2_decap_8 FILLER_79_1850 ();
 sg13g2_decap_4 FILLER_79_1857 ();
 sg13g2_fill_1 FILLER_79_1861 ();
 sg13g2_fill_2 FILLER_79_1866 ();
 sg13g2_fill_2 FILLER_79_1882 ();
 sg13g2_fill_2 FILLER_79_1897 ();
 sg13g2_fill_2 FILLER_79_1939 ();
 sg13g2_decap_8 FILLER_79_1945 ();
 sg13g2_decap_4 FILLER_79_1952 ();
 sg13g2_fill_2 FILLER_79_1956 ();
 sg13g2_fill_2 FILLER_79_1984 ();
 sg13g2_fill_2 FILLER_79_2038 ();
 sg13g2_fill_1 FILLER_79_2040 ();
 sg13g2_fill_2 FILLER_79_2080 ();
 sg13g2_fill_1 FILLER_79_2082 ();
 sg13g2_fill_2 FILLER_79_2087 ();
 sg13g2_fill_2 FILLER_79_2098 ();
 sg13g2_fill_1 FILLER_79_2126 ();
 sg13g2_decap_4 FILLER_79_2131 ();
 sg13g2_fill_2 FILLER_79_2135 ();
 sg13g2_decap_4 FILLER_79_2163 ();
 sg13g2_fill_1 FILLER_79_2227 ();
 sg13g2_fill_2 FILLER_79_2238 ();
 sg13g2_fill_1 FILLER_79_2240 ();
 sg13g2_decap_4 FILLER_79_2268 ();
 sg13g2_fill_2 FILLER_79_2272 ();
 sg13g2_fill_1 FILLER_79_2278 ();
 sg13g2_fill_1 FILLER_79_2289 ();
 sg13g2_fill_2 FILLER_79_2300 ();
 sg13g2_fill_1 FILLER_79_2302 ();
 sg13g2_fill_1 FILLER_79_2322 ();
 sg13g2_fill_1 FILLER_79_2327 ();
 sg13g2_fill_2 FILLER_79_2364 ();
 sg13g2_fill_1 FILLER_79_2366 ();
 sg13g2_decap_8 FILLER_79_2371 ();
 sg13g2_decap_8 FILLER_79_2378 ();
 sg13g2_fill_2 FILLER_79_2385 ();
 sg13g2_fill_2 FILLER_79_2419 ();
 sg13g2_fill_2 FILLER_79_2460 ();
 sg13g2_fill_1 FILLER_79_2462 ();
 sg13g2_fill_1 FILLER_79_2489 ();
 sg13g2_fill_2 FILLER_79_2500 ();
 sg13g2_fill_1 FILLER_79_2502 ();
 sg13g2_decap_8 FILLER_79_2507 ();
 sg13g2_decap_8 FILLER_79_2514 ();
 sg13g2_decap_8 FILLER_79_2521 ();
 sg13g2_decap_8 FILLER_79_2528 ();
 sg13g2_decap_8 FILLER_79_2535 ();
 sg13g2_decap_8 FILLER_79_2542 ();
 sg13g2_decap_8 FILLER_79_2549 ();
 sg13g2_decap_8 FILLER_79_2556 ();
 sg13g2_decap_8 FILLER_79_2563 ();
 sg13g2_decap_8 FILLER_79_2570 ();
 sg13g2_decap_8 FILLER_79_2577 ();
 sg13g2_decap_8 FILLER_79_2584 ();
 sg13g2_decap_8 FILLER_79_2591 ();
 sg13g2_decap_8 FILLER_79_2598 ();
 sg13g2_decap_8 FILLER_79_2605 ();
 sg13g2_decap_8 FILLER_79_2612 ();
 sg13g2_decap_8 FILLER_79_2619 ();
 sg13g2_decap_8 FILLER_79_2626 ();
 sg13g2_decap_8 FILLER_79_2633 ();
 sg13g2_decap_8 FILLER_79_2640 ();
 sg13g2_decap_8 FILLER_79_2647 ();
 sg13g2_decap_8 FILLER_79_2654 ();
 sg13g2_decap_8 FILLER_79_2661 ();
 sg13g2_fill_2 FILLER_79_2668 ();
 sg13g2_fill_2 FILLER_80_0 ();
 sg13g2_fill_1 FILLER_80_2 ();
 sg13g2_decap_4 FILLER_80_6 ();
 sg13g2_fill_1 FILLER_80_10 ();
 sg13g2_fill_2 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_46 ();
 sg13g2_fill_1 FILLER_80_53 ();
 sg13g2_decap_8 FILLER_80_62 ();
 sg13g2_decap_8 FILLER_80_69 ();
 sg13g2_fill_2 FILLER_80_76 ();
 sg13g2_fill_2 FILLER_80_157 ();
 sg13g2_fill_2 FILLER_80_183 ();
 sg13g2_fill_1 FILLER_80_195 ();
 sg13g2_fill_1 FILLER_80_207 ();
 sg13g2_fill_1 FILLER_80_212 ();
 sg13g2_fill_1 FILLER_80_217 ();
 sg13g2_fill_1 FILLER_80_222 ();
 sg13g2_fill_1 FILLER_80_231 ();
 sg13g2_fill_2 FILLER_80_245 ();
 sg13g2_fill_2 FILLER_80_268 ();
 sg13g2_decap_4 FILLER_80_287 ();
 sg13g2_decap_4 FILLER_80_299 ();
 sg13g2_fill_1 FILLER_80_303 ();
 sg13g2_decap_8 FILLER_80_313 ();
 sg13g2_decap_4 FILLER_80_324 ();
 sg13g2_decap_8 FILLER_80_332 ();
 sg13g2_decap_8 FILLER_80_339 ();
 sg13g2_fill_1 FILLER_80_346 ();
 sg13g2_fill_1 FILLER_80_352 ();
 sg13g2_fill_2 FILLER_80_370 ();
 sg13g2_decap_4 FILLER_80_390 ();
 sg13g2_fill_1 FILLER_80_394 ();
 sg13g2_decap_8 FILLER_80_402 ();
 sg13g2_decap_8 FILLER_80_409 ();
 sg13g2_decap_8 FILLER_80_420 ();
 sg13g2_decap_8 FILLER_80_427 ();
 sg13g2_decap_8 FILLER_80_434 ();
 sg13g2_decap_8 FILLER_80_441 ();
 sg13g2_fill_2 FILLER_80_448 ();
 sg13g2_fill_1 FILLER_80_454 ();
 sg13g2_decap_8 FILLER_80_459 ();
 sg13g2_decap_4 FILLER_80_466 ();
 sg13g2_decap_4 FILLER_80_474 ();
 sg13g2_decap_8 FILLER_80_499 ();
 sg13g2_decap_8 FILLER_80_506 ();
 sg13g2_decap_4 FILLER_80_513 ();
 sg13g2_fill_1 FILLER_80_517 ();
 sg13g2_decap_4 FILLER_80_526 ();
 sg13g2_decap_8 FILLER_80_534 ();
 sg13g2_decap_4 FILLER_80_541 ();
 sg13g2_decap_8 FILLER_80_549 ();
 sg13g2_decap_8 FILLER_80_556 ();
 sg13g2_decap_4 FILLER_80_563 ();
 sg13g2_fill_2 FILLER_80_567 ();
 sg13g2_decap_8 FILLER_80_573 ();
 sg13g2_decap_4 FILLER_80_580 ();
 sg13g2_fill_2 FILLER_80_584 ();
 sg13g2_fill_2 FILLER_80_590 ();
 sg13g2_decap_4 FILLER_80_596 ();
 sg13g2_decap_4 FILLER_80_604 ();
 sg13g2_decap_8 FILLER_80_648 ();
 sg13g2_decap_8 FILLER_80_655 ();
 sg13g2_decap_4 FILLER_80_662 ();
 sg13g2_decap_8 FILLER_80_670 ();
 sg13g2_decap_4 FILLER_80_677 ();
 sg13g2_decap_8 FILLER_80_691 ();
 sg13g2_decap_4 FILLER_80_698 ();
 sg13g2_fill_1 FILLER_80_702 ();
 sg13g2_decap_4 FILLER_80_711 ();
 sg13g2_decap_8 FILLER_80_725 ();
 sg13g2_decap_8 FILLER_80_732 ();
 sg13g2_decap_8 FILLER_80_739 ();
 sg13g2_decap_4 FILLER_80_746 ();
 sg13g2_fill_1 FILLER_80_750 ();
 sg13g2_decap_8 FILLER_80_795 ();
 sg13g2_decap_8 FILLER_80_802 ();
 sg13g2_decap_8 FILLER_80_809 ();
 sg13g2_decap_8 FILLER_80_816 ();
 sg13g2_fill_1 FILLER_80_823 ();
 sg13g2_decap_8 FILLER_80_828 ();
 sg13g2_fill_1 FILLER_80_835 ();
 sg13g2_decap_8 FILLER_80_844 ();
 sg13g2_fill_2 FILLER_80_851 ();
 sg13g2_fill_1 FILLER_80_853 ();
 sg13g2_decap_4 FILLER_80_864 ();
 sg13g2_decap_8 FILLER_80_872 ();
 sg13g2_decap_8 FILLER_80_879 ();
 sg13g2_fill_2 FILLER_80_886 ();
 sg13g2_fill_2 FILLER_80_902 ();
 sg13g2_fill_1 FILLER_80_904 ();
 sg13g2_fill_1 FILLER_80_914 ();
 sg13g2_decap_4 FILLER_80_919 ();
 sg13g2_fill_1 FILLER_80_923 ();
 sg13g2_decap_8 FILLER_80_950 ();
 sg13g2_decap_8 FILLER_80_957 ();
 sg13g2_decap_8 FILLER_80_964 ();
 sg13g2_decap_8 FILLER_80_971 ();
 sg13g2_decap_8 FILLER_80_978 ();
 sg13g2_decap_8 FILLER_80_985 ();
 sg13g2_decap_8 FILLER_80_992 ();
 sg13g2_decap_8 FILLER_80_999 ();
 sg13g2_fill_1 FILLER_80_1006 ();
 sg13g2_decap_8 FILLER_80_1012 ();
 sg13g2_fill_1 FILLER_80_1019 ();
 sg13g2_decap_8 FILLER_80_1056 ();
 sg13g2_decap_8 FILLER_80_1063 ();
 sg13g2_decap_8 FILLER_80_1070 ();
 sg13g2_decap_8 FILLER_80_1077 ();
 sg13g2_decap_8 FILLER_80_1088 ();
 sg13g2_decap_8 FILLER_80_1095 ();
 sg13g2_decap_8 FILLER_80_1102 ();
 sg13g2_fill_2 FILLER_80_1109 ();
 sg13g2_fill_1 FILLER_80_1111 ();
 sg13g2_decap_8 FILLER_80_1120 ();
 sg13g2_decap_4 FILLER_80_1127 ();
 sg13g2_decap_8 FILLER_80_1135 ();
 sg13g2_decap_8 FILLER_80_1142 ();
 sg13g2_decap_8 FILLER_80_1149 ();
 sg13g2_decap_8 FILLER_80_1156 ();
 sg13g2_decap_8 FILLER_80_1163 ();
 sg13g2_decap_8 FILLER_80_1170 ();
 sg13g2_decap_8 FILLER_80_1177 ();
 sg13g2_decap_8 FILLER_80_1184 ();
 sg13g2_decap_8 FILLER_80_1191 ();
 sg13g2_fill_2 FILLER_80_1198 ();
 sg13g2_fill_1 FILLER_80_1200 ();
 sg13g2_fill_2 FILLER_80_1206 ();
 sg13g2_fill_1 FILLER_80_1219 ();
 sg13g2_fill_1 FILLER_80_1231 ();
 sg13g2_decap_8 FILLER_80_1236 ();
 sg13g2_decap_8 FILLER_80_1243 ();
 sg13g2_decap_8 FILLER_80_1250 ();
 sg13g2_decap_8 FILLER_80_1257 ();
 sg13g2_decap_8 FILLER_80_1264 ();
 sg13g2_decap_8 FILLER_80_1271 ();
 sg13g2_decap_8 FILLER_80_1278 ();
 sg13g2_decap_8 FILLER_80_1285 ();
 sg13g2_decap_4 FILLER_80_1292 ();
 sg13g2_fill_1 FILLER_80_1296 ();
 sg13g2_fill_2 FILLER_80_1310 ();
 sg13g2_decap_8 FILLER_80_1316 ();
 sg13g2_fill_2 FILLER_80_1323 ();
 sg13g2_fill_1 FILLER_80_1325 ();
 sg13g2_decap_8 FILLER_80_1330 ();
 sg13g2_decap_8 FILLER_80_1337 ();
 sg13g2_decap_8 FILLER_80_1344 ();
 sg13g2_decap_8 FILLER_80_1351 ();
 sg13g2_decap_8 FILLER_80_1358 ();
 sg13g2_decap_8 FILLER_80_1365 ();
 sg13g2_decap_8 FILLER_80_1372 ();
 sg13g2_decap_8 FILLER_80_1379 ();
 sg13g2_decap_8 FILLER_80_1386 ();
 sg13g2_decap_8 FILLER_80_1393 ();
 sg13g2_decap_8 FILLER_80_1400 ();
 sg13g2_decap_8 FILLER_80_1407 ();
 sg13g2_decap_8 FILLER_80_1414 ();
 sg13g2_decap_8 FILLER_80_1421 ();
 sg13g2_decap_8 FILLER_80_1428 ();
 sg13g2_fill_2 FILLER_80_1435 ();
 sg13g2_fill_1 FILLER_80_1437 ();
 sg13g2_decap_8 FILLER_80_1443 ();
 sg13g2_decap_8 FILLER_80_1450 ();
 sg13g2_decap_8 FILLER_80_1457 ();
 sg13g2_decap_8 FILLER_80_1464 ();
 sg13g2_decap_8 FILLER_80_1471 ();
 sg13g2_decap_8 FILLER_80_1478 ();
 sg13g2_fill_2 FILLER_80_1485 ();
 sg13g2_decap_8 FILLER_80_1492 ();
 sg13g2_fill_2 FILLER_80_1499 ();
 sg13g2_fill_1 FILLER_80_1501 ();
 sg13g2_decap_8 FILLER_80_1506 ();
 sg13g2_decap_8 FILLER_80_1513 ();
 sg13g2_decap_8 FILLER_80_1520 ();
 sg13g2_decap_8 FILLER_80_1527 ();
 sg13g2_decap_8 FILLER_80_1534 ();
 sg13g2_decap_8 FILLER_80_1541 ();
 sg13g2_decap_8 FILLER_80_1548 ();
 sg13g2_decap_4 FILLER_80_1555 ();
 sg13g2_fill_2 FILLER_80_1559 ();
 sg13g2_decap_8 FILLER_80_1565 ();
 sg13g2_decap_8 FILLER_80_1572 ();
 sg13g2_decap_8 FILLER_80_1579 ();
 sg13g2_decap_8 FILLER_80_1586 ();
 sg13g2_decap_8 FILLER_80_1593 ();
 sg13g2_decap_8 FILLER_80_1600 ();
 sg13g2_decap_4 FILLER_80_1607 ();
 sg13g2_fill_1 FILLER_80_1611 ();
 sg13g2_decap_8 FILLER_80_1642 ();
 sg13g2_fill_1 FILLER_80_1649 ();
 sg13g2_fill_2 FILLER_80_1654 ();
 sg13g2_fill_1 FILLER_80_1656 ();
 sg13g2_decap_8 FILLER_80_1687 ();
 sg13g2_decap_8 FILLER_80_1694 ();
 sg13g2_decap_8 FILLER_80_1701 ();
 sg13g2_decap_8 FILLER_80_1708 ();
 sg13g2_decap_8 FILLER_80_1729 ();
 sg13g2_decap_8 FILLER_80_1736 ();
 sg13g2_decap_8 FILLER_80_1769 ();
 sg13g2_decap_4 FILLER_80_1776 ();
 sg13g2_fill_1 FILLER_80_1780 ();
 sg13g2_decap_8 FILLER_80_1785 ();
 sg13g2_decap_8 FILLER_80_1796 ();
 sg13g2_decap_8 FILLER_80_1803 ();
 sg13g2_decap_8 FILLER_80_1810 ();
 sg13g2_decap_8 FILLER_80_1843 ();
 sg13g2_fill_2 FILLER_80_1850 ();
 sg13g2_fill_1 FILLER_80_1852 ();
 sg13g2_decap_8 FILLER_80_1879 ();
 sg13g2_decap_8 FILLER_80_1886 ();
 sg13g2_decap_8 FILLER_80_1893 ();
 sg13g2_decap_8 FILLER_80_1900 ();
 sg13g2_decap_8 FILLER_80_1911 ();
 sg13g2_fill_2 FILLER_80_1918 ();
 sg13g2_decap_8 FILLER_80_1928 ();
 sg13g2_decap_8 FILLER_80_1935 ();
 sg13g2_decap_8 FILLER_80_1942 ();
 sg13g2_decap_8 FILLER_80_1949 ();
 sg13g2_decap_8 FILLER_80_1956 ();
 sg13g2_decap_4 FILLER_80_1963 ();
 sg13g2_decap_8 FILLER_80_1971 ();
 sg13g2_fill_1 FILLER_80_1982 ();
 sg13g2_fill_2 FILLER_80_2004 ();
 sg13g2_decap_4 FILLER_80_2010 ();
 sg13g2_fill_2 FILLER_80_2014 ();
 sg13g2_fill_2 FILLER_80_2028 ();
 sg13g2_fill_1 FILLER_80_2030 ();
 sg13g2_fill_2 FILLER_80_2035 ();
 sg13g2_fill_1 FILLER_80_2037 ();
 sg13g2_fill_2 FILLER_80_2042 ();
 sg13g2_fill_1 FILLER_80_2048 ();
 sg13g2_decap_4 FILLER_80_2053 ();
 sg13g2_fill_2 FILLER_80_2057 ();
 sg13g2_fill_1 FILLER_80_2063 ();
 sg13g2_decap_8 FILLER_80_2068 ();
 sg13g2_decap_8 FILLER_80_2075 ();
 sg13g2_fill_2 FILLER_80_2082 ();
 sg13g2_fill_2 FILLER_80_2088 ();
 sg13g2_fill_1 FILLER_80_2090 ();
 sg13g2_decap_8 FILLER_80_2125 ();
 sg13g2_decap_8 FILLER_80_2132 ();
 sg13g2_fill_2 FILLER_80_2139 ();
 sg13g2_decap_8 FILLER_80_2149 ();
 sg13g2_decap_8 FILLER_80_2156 ();
 sg13g2_decap_8 FILLER_80_2163 ();
 sg13g2_fill_2 FILLER_80_2170 ();
 sg13g2_fill_1 FILLER_80_2172 ();
 sg13g2_decap_8 FILLER_80_2177 ();
 sg13g2_decap_8 FILLER_80_2184 ();
 sg13g2_decap_8 FILLER_80_2191 ();
 sg13g2_decap_4 FILLER_80_2198 ();
 sg13g2_fill_1 FILLER_80_2202 ();
 sg13g2_decap_8 FILLER_80_2233 ();
 sg13g2_fill_1 FILLER_80_2240 ();
 sg13g2_fill_2 FILLER_80_2251 ();
 sg13g2_decap_8 FILLER_80_2279 ();
 sg13g2_decap_8 FILLER_80_2286 ();
 sg13g2_decap_8 FILLER_80_2297 ();
 sg13g2_decap_8 FILLER_80_2304 ();
 sg13g2_decap_8 FILLER_80_2311 ();
 sg13g2_decap_8 FILLER_80_2318 ();
 sg13g2_decap_4 FILLER_80_2325 ();
 sg13g2_fill_2 FILLER_80_2329 ();
 sg13g2_fill_1 FILLER_80_2335 ();
 sg13g2_decap_8 FILLER_80_2340 ();
 sg13g2_decap_8 FILLER_80_2347 ();
 sg13g2_fill_2 FILLER_80_2354 ();
 sg13g2_fill_1 FILLER_80_2356 ();
 sg13g2_decap_8 FILLER_80_2397 ();
 sg13g2_decap_4 FILLER_80_2404 ();
 sg13g2_fill_2 FILLER_80_2408 ();
 sg13g2_decap_8 FILLER_80_2418 ();
 sg13g2_fill_2 FILLER_80_2425 ();
 sg13g2_fill_1 FILLER_80_2427 ();
 sg13g2_fill_2 FILLER_80_2432 ();
 sg13g2_fill_1 FILLER_80_2434 ();
 sg13g2_decap_8 FILLER_80_2469 ();
 sg13g2_decap_8 FILLER_80_2476 ();
 sg13g2_decap_8 FILLER_80_2483 ();
 sg13g2_decap_8 FILLER_80_2490 ();
 sg13g2_decap_8 FILLER_80_2497 ();
 sg13g2_decap_8 FILLER_80_2504 ();
 sg13g2_decap_8 FILLER_80_2511 ();
 sg13g2_decap_8 FILLER_80_2518 ();
 sg13g2_decap_8 FILLER_80_2525 ();
 sg13g2_decap_8 FILLER_80_2532 ();
 sg13g2_decap_8 FILLER_80_2539 ();
 sg13g2_decap_8 FILLER_80_2546 ();
 sg13g2_decap_8 FILLER_80_2553 ();
 sg13g2_decap_8 FILLER_80_2560 ();
 sg13g2_decap_8 FILLER_80_2567 ();
 sg13g2_decap_8 FILLER_80_2574 ();
 sg13g2_decap_8 FILLER_80_2581 ();
 sg13g2_decap_8 FILLER_80_2588 ();
 sg13g2_decap_8 FILLER_80_2595 ();
 sg13g2_decap_8 FILLER_80_2602 ();
 sg13g2_decap_8 FILLER_80_2609 ();
 sg13g2_decap_8 FILLER_80_2616 ();
 sg13g2_decap_8 FILLER_80_2623 ();
 sg13g2_decap_8 FILLER_80_2630 ();
 sg13g2_decap_8 FILLER_80_2637 ();
 sg13g2_decap_8 FILLER_80_2644 ();
 sg13g2_decap_8 FILLER_80_2651 ();
 sg13g2_decap_8 FILLER_80_2658 ();
 sg13g2_decap_4 FILLER_80_2665 ();
 sg13g2_fill_1 FILLER_80_2669 ();
endmodule
