module tt_um_tomkeddie_a (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire clknet_0_clk;
 wire net58;
 wire b0;
 wire g0;
 wire hs;
 wire \vga.blank_h ;
 wire \vga.blank_v ;
 wire \vga.car_pos_h[0] ;
 wire \vga.car_pos_h[1] ;
 wire \vga.car_pos_h[2] ;
 wire \vga.car_pos_h[3] ;
 wire \vga.car_pos_h[4] ;
 wire \vga.car_pos_h[5] ;
 wire \vga.car_pos_h[6] ;
 wire \vga.car_pos_h[7] ;
 wire \vga.car_pos_h[8] ;
 wire \vga.car_pos_h[9] ;
 wire \vga.count_h[0] ;
 wire \vga.count_h[1] ;
 wire \vga.count_h[2] ;
 wire \vga.count_h[3] ;
 wire \vga.count_h[4] ;
 wire \vga.count_h[5] ;
 wire \vga.count_h[6] ;
 wire \vga.count_h[7] ;
 wire \vga.count_h[8] ;
 wire \vga.count_h[9] ;
 wire \vga.count_v[0] ;
 wire \vga.count_v[1] ;
 wire \vga.count_v[2] ;
 wire \vga.count_v[3] ;
 wire \vga.count_v[4] ;
 wire \vga.count_v[5] ;
 wire \vga.count_v[6] ;
 wire \vga.count_v[7] ;
 wire \vga.count_v[8] ;
 wire \vga.count_v[9] ;
 wire \vga.hs_out ;
 wire \vga.interval_counter[0] ;
 wire \vga.interval_counter[10] ;
 wire \vga.interval_counter[11] ;
 wire \vga.interval_counter[12] ;
 wire \vga.interval_counter[13] ;
 wire \vga.interval_counter[14] ;
 wire \vga.interval_counter[15] ;
 wire \vga.interval_counter[16] ;
 wire \vga.interval_counter[17] ;
 wire \vga.interval_counter[18] ;
 wire \vga.interval_counter[19] ;
 wire \vga.interval_counter[1] ;
 wire \vga.interval_counter[20] ;
 wire \vga.interval_counter[21] ;
 wire \vga.interval_counter[22] ;
 wire \vga.interval_counter[23] ;
 wire \vga.interval_counter[24] ;
 wire \vga.interval_counter[2] ;
 wire \vga.interval_counter[3] ;
 wire \vga.interval_counter[4] ;
 wire \vga.interval_counter[5] ;
 wire \vga.interval_counter[6] ;
 wire \vga.interval_counter[7] ;
 wire \vga.interval_counter[8] ;
 wire \vga.interval_counter[9] ;
 wire \vga.left_1d ;
 wire \vga.left_pressed ;
 wire \vga.right_1d ;
 wire \vga.right_pressed ;
 wire \vga.score[0] ;
 wire \vga.score_ten_enable ;
 wire \vga.score_unit_pixels[1] ;
 wire \vga.score_unit_pixels[2] ;
 wire \vga.speed_lsb_1d ;
 wire \vga.speed_msb_1d ;
 wire \vga.vs ;
 wire \vga.vs_out ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sg13g2_inv_1 _0624_ (.Y(_0093_),
    .A(\vga.score[0] ));
 sg13g2_buf_2 _0625_ (.A(rst_n),
    .X(_0094_));
 sg13g2_o21ai_1 _0626_ (.B1(_0094_),
    .Y(_0000_),
    .A1(_0093_),
    .A2(net3));
 sg13g2_inv_1 _0627_ (.Y(_0001_),
    .A(_0000_));
 sg13g2_buf_1 _0628_ (.A(\vga.count_v[3] ),
    .X(_0095_));
 sg13g2_buf_1 _0629_ (.A(\vga.count_v[1] ),
    .X(_0096_));
 sg13g2_nand2b_1 _0630_ (.Y(_0097_),
    .B(net54),
    .A_N(net55));
 sg13g2_buf_1 _0631_ (.A(\vga.count_v[5] ),
    .X(_0098_));
 sg13g2_buf_1 _0632_ (.A(\vga.count_v[2] ),
    .X(_0099_));
 sg13g2_buf_1 _0633_ (.A(\vga.count_v[4] ),
    .X(_0100_));
 sg13g2_inv_1 _0634_ (.Y(_0101_),
    .A(_0100_));
 sg13g2_nand3_1 _0635_ (.B(net52),
    .C(_0101_),
    .A(net53),
    .Y(_0102_));
 sg13g2_nor2_1 _0636_ (.A(_0097_),
    .B(_0102_),
    .Y(_0103_));
 sg13g2_inv_1 _0637_ (.Y(_0104_),
    .A(net52));
 sg13g2_nor2_1 _0638_ (.A(_0104_),
    .B(net54),
    .Y(_0105_));
 sg13g2_nand2_1 _0639_ (.Y(_0106_),
    .A(net55),
    .B(_0105_));
 sg13g2_nand3b_1 _0640_ (.B(_0104_),
    .C(net54),
    .Y(_0107_),
    .A_N(net55));
 sg13g2_nand2b_1 _0641_ (.Y(_0108_),
    .B(_0100_),
    .A_N(net53));
 sg13g2_a21oi_1 _0642_ (.A1(_0106_),
    .A2(_0107_),
    .Y(_0109_),
    .B1(_0108_));
 sg13g2_buf_2 _0643_ (.A(\vga.count_v[6] ),
    .X(_0110_));
 sg13g2_buf_2 _0644_ (.A(\vga.count_v[0] ),
    .X(_0111_));
 sg13g2_or3_1 _0645_ (.A(\vga.count_v[9] ),
    .B(\vga.count_v[8] ),
    .C(\vga.count_v[7] ),
    .X(_0112_));
 sg13g2_nor3_1 _0646_ (.A(_0110_),
    .B(_0111_),
    .C(_0112_),
    .Y(_0113_));
 sg13g2_o21ai_1 _0647_ (.B1(_0113_),
    .Y(_0114_),
    .A1(_0103_),
    .A2(_0109_));
 sg13g2_xor2_1 _0648_ (.B(_0096_),
    .A(net55),
    .X(_0115_));
 sg13g2_nor3_1 _0649_ (.A(net52),
    .B(_0101_),
    .C(_0115_),
    .Y(_0116_));
 sg13g2_and3_1 _0650_ (.X(_0117_),
    .A(net53),
    .B(_0113_),
    .C(_0116_));
 sg13g2_nor2_1 _0651_ (.A(\vga.score_unit_pixels[1] ),
    .B(_0117_),
    .Y(_0118_));
 sg13g2_inv_1 _0652_ (.Y(_0119_),
    .A(_0102_));
 sg13g2_nor2_1 _0653_ (.A(net52),
    .B(_0108_),
    .Y(_0120_));
 sg13g2_a21oi_1 _0654_ (.A1(_0002_),
    .A2(_0119_),
    .Y(_0121_),
    .B1(_0120_));
 sg13g2_o21ai_1 _0655_ (.B1(_0113_),
    .Y(_0122_),
    .A1(_0097_),
    .A2(_0121_));
 sg13g2_inv_1 _0656_ (.Y(_0123_),
    .A(net54));
 sg13g2_o21ai_1 _0657_ (.B1(net55),
    .Y(_0124_),
    .A1(_0123_),
    .A2(_0004_));
 sg13g2_and2_1 _0658_ (.A(_0097_),
    .B(_0124_),
    .X(_0125_));
 sg13g2_nor4_1 _0659_ (.A(net53),
    .B(net55),
    .C(_0123_),
    .D(_0004_),
    .Y(_0126_));
 sg13g2_a21oi_1 _0660_ (.A1(net53),
    .A2(_0125_),
    .Y(_0127_),
    .B1(_0126_));
 sg13g2_nand3b_1 _0661_ (.B(net55),
    .C(_0105_),
    .Y(_0128_),
    .A_N(net53));
 sg13g2_o21ai_1 _0662_ (.B1(_0128_),
    .Y(_0129_),
    .A1(net52),
    .A2(_0127_));
 sg13g2_a21oi_1 _0663_ (.A1(_0100_),
    .A2(_0129_),
    .Y(_0130_),
    .B1(_0103_));
 sg13g2_nor2_1 _0664_ (.A(_0122_),
    .B(_0130_),
    .Y(_0131_));
 sg13g2_a21oi_1 _0665_ (.A1(_0114_),
    .A2(_0118_),
    .Y(_0088_),
    .B1(_0131_));
 sg13g2_nand2b_1 _0666_ (.Y(_0132_),
    .B(\vga.score_unit_pixels[2] ),
    .A_N(_0117_));
 sg13g2_nand2_1 _0667_ (.Y(_0133_),
    .A(_0003_),
    .B(_0117_));
 sg13g2_nand3_1 _0668_ (.B(_0132_),
    .C(_0133_),
    .A(_0114_),
    .Y(_0089_));
 sg13g2_nor4_1 _0669_ (.A(\vga.interval_counter[20] ),
    .B(\vga.interval_counter[23] ),
    .C(\vga.interval_counter[22] ),
    .D(\vga.interval_counter[24] ),
    .Y(_0134_));
 sg13g2_nor2b_1 _0670_ (.A(\vga.interval_counter[21] ),
    .B_N(_0134_),
    .Y(_0135_));
 sg13g2_nor3_1 _0671_ (.A(\vga.interval_counter[17] ),
    .B(\vga.interval_counter[19] ),
    .C(\vga.interval_counter[18] ),
    .Y(_0136_));
 sg13g2_buf_2 _0672_ (.A(\vga.interval_counter[16] ),
    .X(_0137_));
 sg13g2_nor4_1 _0673_ (.A(\vga.interval_counter[8] ),
    .B(\vga.interval_counter[10] ),
    .C(\vga.interval_counter[14] ),
    .D(_0137_),
    .Y(_0138_));
 sg13g2_nand2_1 _0674_ (.Y(_0139_),
    .A(_0136_),
    .B(_0138_));
 sg13g2_nor2_1 _0675_ (.A(\vga.interval_counter[2] ),
    .B(\vga.interval_counter[6] ),
    .Y(_0140_));
 sg13g2_buf_8 _0676_ (.A(\vga.interval_counter[1] ),
    .X(_0141_));
 sg13g2_buf_8 _0677_ (.A(\vga.interval_counter[0] ),
    .X(_0142_));
 sg13g2_nor4_1 _0678_ (.A(_0141_),
    .B(_0142_),
    .C(\vga.interval_counter[3] ),
    .D(\vga.interval_counter[9] ),
    .Y(_0143_));
 sg13g2_nand2_1 _0679_ (.Y(_0144_),
    .A(_0140_),
    .B(_0143_));
 sg13g2_inv_1 _0680_ (.Y(_0145_),
    .A(\vga.interval_counter[5] ));
 sg13g2_buf_2 _0681_ (.A(\vga.interval_counter[13] ),
    .X(_0146_));
 sg13g2_buf_2 _0682_ (.A(\vga.interval_counter[12] ),
    .X(_0147_));
 sg13g2_buf_2 _0683_ (.A(\vga.interval_counter[15] ),
    .X(_0148_));
 sg13g2_nor4_1 _0684_ (.A(\vga.interval_counter[11] ),
    .B(_0146_),
    .C(_0147_),
    .D(_0148_),
    .Y(_0149_));
 sg13g2_nand3b_1 _0685_ (.B(_0145_),
    .C(_0149_),
    .Y(_0150_),
    .A_N(\vga.interval_counter[4] ));
 sg13g2_nor4_1 _0686_ (.A(\vga.interval_counter[7] ),
    .B(_0139_),
    .C(_0144_),
    .D(_0150_),
    .Y(_0151_));
 sg13g2_and2_1 _0687_ (.A(_0135_),
    .B(_0151_),
    .X(_0152_));
 sg13g2_buf_1 _0688_ (.A(_0152_),
    .X(_0153_));
 sg13g2_mux2_1 _0689_ (.A0(\vga.left_1d ),
    .A1(net1),
    .S(_0153_),
    .X(_0081_));
 sg13g2_mux2_1 _0690_ (.A0(\vga.right_1d ),
    .A1(net2),
    .S(_0153_),
    .X(_0084_));
 sg13g2_inv_1 _0691_ (.Y(_0021_),
    .A(_0000_));
 sg13g2_nor2b_1 _0692_ (.A(\vga.count_h[8] ),
    .B_N(\vga.count_h[9] ),
    .Y(_0154_));
 sg13g2_buf_1 _0693_ (.A(\vga.count_h[7] ),
    .X(_0155_));
 sg13g2_buf_1 _0694_ (.A(\vga.count_h[6] ),
    .X(_0156_));
 sg13g2_buf_1 _0695_ (.A(\vga.count_h[5] ),
    .X(_0157_));
 sg13g2_buf_1 _0696_ (.A(\vga.count_h[4] ),
    .X(_0158_));
 sg13g2_inv_1 _0697_ (.Y(_0159_),
    .A(net48));
 sg13g2_buf_2 _0698_ (.A(\vga.count_h[0] ),
    .X(_0160_));
 sg13g2_buf_1 _0699_ (.A(\vga.count_h[2] ),
    .X(_0161_));
 sg13g2_buf_1 _0700_ (.A(\vga.count_h[1] ),
    .X(_0162_));
 sg13g2_buf_1 _0701_ (.A(\vga.count_h[3] ),
    .X(_0163_));
 sg13g2_and4_1 _0702_ (.A(_0160_),
    .B(net47),
    .C(net46),
    .D(_0163_),
    .X(_0164_));
 sg13g2_buf_2 _0703_ (.A(_0164_),
    .X(_0165_));
 sg13g2_nand3_1 _0704_ (.B(_0165_),
    .C(_0154_),
    .A(_0159_),
    .Y(_0166_));
 sg13g2_o21ai_1 _0705_ (.B1(_0166_),
    .Y(_0167_),
    .A1(_0159_),
    .A2(_0007_));
 sg13g2_nand4_1 _0706_ (.B(net50),
    .C(net49),
    .A(net51),
    .Y(_0168_),
    .D(_0167_));
 sg13g2_o21ai_1 _0707_ (.B1(_0168_),
    .Y(_0169_),
    .A1(_0007_),
    .A2(_0154_));
 sg13g2_nor4_1 _0708_ (.A(net50),
    .B(net49),
    .C(net48),
    .D(_0165_),
    .Y(_0170_));
 sg13g2_nand2b_1 _0709_ (.Y(_0171_),
    .B(net51),
    .A_N(_0170_));
 sg13g2_a21oi_1 _0710_ (.A1(_0154_),
    .A2(_0171_),
    .Y(_0172_),
    .B1(_0007_));
 sg13g2_nand2_1 _0711_ (.Y(_0173_),
    .A(_0094_),
    .B(_0172_));
 sg13g2_nor2_1 _0712_ (.A(_0169_),
    .B(_0173_),
    .Y(_0055_));
 sg13g2_inv_1 _0713_ (.Y(_0174_),
    .A(_0020_));
 sg13g2_nand4_1 _0714_ (.B(\vga.interval_counter[9] ),
    .C(\vga.interval_counter[11] ),
    .A(\vga.interval_counter[8] ),
    .Y(_0175_),
    .D(\vga.interval_counter[10] ));
 sg13g2_nor2_1 _0715_ (.A(_0147_),
    .B(_0137_),
    .Y(_0176_));
 sg13g2_nand3_1 _0716_ (.B(_0140_),
    .C(_0176_),
    .A(_0142_),
    .Y(_0177_));
 sg13g2_inv_1 _0717_ (.Y(_0178_),
    .A(\vga.interval_counter[14] ));
 sg13g2_nand4_1 _0718_ (.B(_0145_),
    .C(_0178_),
    .A(\vga.interval_counter[4] ),
    .Y(_0179_),
    .D(_0148_));
 sg13g2_inv_1 _0719_ (.Y(_0180_),
    .A(_0141_));
 sg13g2_nand4_1 _0720_ (.B(_0180_),
    .C(\vga.interval_counter[3] ),
    .A(net4),
    .Y(_0181_),
    .D(\vga.interval_counter[7] ));
 sg13g2_nor4_1 _0721_ (.A(_0175_),
    .B(_0177_),
    .C(_0179_),
    .D(_0181_),
    .Y(_0182_));
 sg13g2_or3_1 _0722_ (.A(net4),
    .B(\vga.interval_counter[7] ),
    .C(\vga.interval_counter[11] ),
    .X(_0183_));
 sg13g2_inv_1 _0723_ (.Y(_0184_),
    .A(\vga.interval_counter[10] ));
 sg13g2_nand2_1 _0724_ (.Y(_0185_),
    .A(\vga.interval_counter[8] ),
    .B(\vga.interval_counter[9] ));
 sg13g2_nand2_1 _0725_ (.Y(_0186_),
    .A(\vga.interval_counter[6] ),
    .B(\vga.interval_counter[14] ));
 sg13g2_nand2b_1 _0726_ (.Y(_0187_),
    .B(\vga.interval_counter[2] ),
    .A_N(_0142_));
 sg13g2_or4_1 _0727_ (.A(_0184_),
    .B(_0185_),
    .C(_0186_),
    .D(_0187_),
    .X(_0188_));
 sg13g2_nand4_1 _0728_ (.B(_0147_),
    .C(_0148_),
    .A(\vga.interval_counter[5] ),
    .Y(_0189_),
    .D(_0137_));
 sg13g2_or3_1 _0729_ (.A(_0180_),
    .B(\vga.interval_counter[3] ),
    .C(\vga.interval_counter[4] ),
    .X(_0190_));
 sg13g2_nor4_1 _0730_ (.A(_0183_),
    .B(_0188_),
    .C(_0189_),
    .D(_0190_),
    .Y(_0191_));
 sg13g2_inv_1 _0731_ (.Y(_0192_),
    .A(\vga.interval_counter[17] ));
 sg13g2_nor4_1 _0732_ (.A(_0146_),
    .B(_0192_),
    .C(\vga.interval_counter[19] ),
    .D(\vga.interval_counter[18] ),
    .Y(_0193_));
 sg13g2_o21ai_1 _0733_ (.B1(_0193_),
    .Y(_0194_),
    .A1(_0182_),
    .A2(_0191_));
 sg13g2_nand4_1 _0734_ (.B(\vga.interval_counter[10] ),
    .C(_0146_),
    .A(\vga.interval_counter[8] ),
    .Y(_0195_),
    .D(_0147_));
 sg13g2_nor4_1 _0735_ (.A(_0144_),
    .B(_0179_),
    .C(_0183_),
    .D(_0195_),
    .Y(_0196_));
 sg13g2_nor3_1 _0736_ (.A(_0150_),
    .B(_0181_),
    .C(_0188_),
    .Y(_0197_));
 sg13g2_or2_1 _0737_ (.X(_0198_),
    .B(_0197_),
    .A(_0196_));
 sg13g2_nand4_1 _0738_ (.B(_0137_),
    .C(_0136_),
    .A(net5),
    .Y(_0199_),
    .D(_0198_));
 sg13g2_o21ai_1 _0739_ (.B1(_0199_),
    .Y(_0200_),
    .A1(net5),
    .A2(_0194_));
 sg13g2_xnor2_1 _0740_ (.Y(_0201_),
    .A(\vga.speed_msb_1d ),
    .B(net5));
 sg13g2_xnor2_1 _0741_ (.Y(_0202_),
    .A(\vga.speed_lsb_1d ),
    .B(net4));
 sg13g2_nand3_1 _0742_ (.B(_0201_),
    .C(_0202_),
    .A(_0094_),
    .Y(_0203_));
 sg13g2_a21o_1 _0743_ (.A2(_0200_),
    .A1(_0135_),
    .B1(_0203_),
    .X(_0204_));
 sg13g2_buf_2 _0744_ (.A(_0204_),
    .X(_0205_));
 sg13g2_buf_1 _0745_ (.A(_0205_),
    .X(_0206_));
 sg13g2_nor2_1 _0746_ (.A(_0174_),
    .B(net29),
    .Y(_0056_));
 sg13g2_and4_1 _0747_ (.A(_0141_),
    .B(_0142_),
    .C(\vga.interval_counter[3] ),
    .D(\vga.interval_counter[2] ),
    .X(_0207_));
 sg13g2_and3_1 _0748_ (.X(_0208_),
    .A(\vga.interval_counter[4] ),
    .B(\vga.interval_counter[5] ),
    .C(_0207_));
 sg13g2_nand3_1 _0749_ (.B(\vga.interval_counter[6] ),
    .C(_0208_),
    .A(\vga.interval_counter[7] ),
    .Y(_0209_));
 sg13g2_buf_2 _0750_ (.A(_0209_),
    .X(_0210_));
 sg13g2_nor2_1 _0751_ (.A(_0185_),
    .B(_0210_),
    .Y(_0211_));
 sg13g2_xnor2_1 _0752_ (.Y(_0212_),
    .A(\vga.interval_counter[10] ),
    .B(_0211_));
 sg13g2_nor2_1 _0753_ (.A(net29),
    .B(_0212_),
    .Y(_0057_));
 sg13g2_nor3_1 _0754_ (.A(_0184_),
    .B(_0185_),
    .C(_0210_),
    .Y(_0213_));
 sg13g2_xnor2_1 _0755_ (.Y(_0214_),
    .A(\vga.interval_counter[11] ),
    .B(_0213_));
 sg13g2_nor2_1 _0756_ (.A(net29),
    .B(_0214_),
    .Y(_0058_));
 sg13g2_nor2_1 _0757_ (.A(_0175_),
    .B(_0210_),
    .Y(_0215_));
 sg13g2_xnor2_1 _0758_ (.Y(_0216_),
    .A(_0147_),
    .B(_0215_));
 sg13g2_nor2_1 _0759_ (.A(_0206_),
    .B(_0216_),
    .Y(_0059_));
 sg13g2_nand2_1 _0760_ (.Y(_0217_),
    .A(_0147_),
    .B(_0215_));
 sg13g2_xor2_1 _0761_ (.B(_0217_),
    .A(_0146_),
    .X(_0218_));
 sg13g2_nor2_1 _0762_ (.A(_0206_),
    .B(_0218_),
    .Y(_0060_));
 sg13g2_nand3_1 _0763_ (.B(_0147_),
    .C(_0215_),
    .A(_0146_),
    .Y(_0219_));
 sg13g2_xnor2_1 _0764_ (.Y(_0220_),
    .A(_0178_),
    .B(_0219_));
 sg13g2_nor2_1 _0765_ (.A(net29),
    .B(_0220_),
    .Y(_0061_));
 sg13g2_nand3_1 _0766_ (.B(_0147_),
    .C(\vga.interval_counter[14] ),
    .A(_0146_),
    .Y(_0221_));
 sg13g2_nor3_1 _0767_ (.A(_0175_),
    .B(_0210_),
    .C(_0221_),
    .Y(_0222_));
 sg13g2_xnor2_1 _0768_ (.Y(_0223_),
    .A(_0148_),
    .B(_0222_));
 sg13g2_nor2_1 _0769_ (.A(net29),
    .B(_0223_),
    .Y(_0062_));
 sg13g2_nand2_1 _0770_ (.Y(_0224_),
    .A(_0148_),
    .B(_0222_));
 sg13g2_xor2_1 _0771_ (.B(_0224_),
    .A(_0137_),
    .X(_0225_));
 sg13g2_nor2_1 _0772_ (.A(net29),
    .B(_0225_),
    .Y(_0063_));
 sg13g2_nand2_1 _0773_ (.Y(_0226_),
    .A(_0148_),
    .B(_0137_));
 sg13g2_nor4_2 _0774_ (.A(_0175_),
    .B(_0226_),
    .C(_0210_),
    .Y(_0227_),
    .D(_0221_));
 sg13g2_xnor2_1 _0775_ (.Y(_0228_),
    .A(\vga.interval_counter[17] ),
    .B(_0227_));
 sg13g2_nor2_1 _0776_ (.A(net29),
    .B(_0228_),
    .Y(_0064_));
 sg13g2_nand2_1 _0777_ (.Y(_0229_),
    .A(\vga.interval_counter[17] ),
    .B(_0227_));
 sg13g2_xor2_1 _0778_ (.B(_0229_),
    .A(\vga.interval_counter[18] ),
    .X(_0230_));
 sg13g2_nor2_1 _0779_ (.A(net29),
    .B(_0230_),
    .Y(_0065_));
 sg13g2_buf_1 _0780_ (.A(_0205_),
    .X(_0231_));
 sg13g2_and2_1 _0781_ (.A(\vga.interval_counter[17] ),
    .B(\vga.interval_counter[18] ),
    .X(_0232_));
 sg13g2_nand2_1 _0782_ (.Y(_0233_),
    .A(_0227_),
    .B(_0232_));
 sg13g2_xor2_1 _0783_ (.B(_0233_),
    .A(\vga.interval_counter[19] ),
    .X(_0234_));
 sg13g2_nor2_1 _0784_ (.A(_0231_),
    .B(_0234_),
    .Y(_0066_));
 sg13g2_xnor2_1 _0785_ (.Y(_0235_),
    .A(_0141_),
    .B(_0142_));
 sg13g2_nor2_1 _0786_ (.A(net28),
    .B(_0235_),
    .Y(_0067_));
 sg13g2_nand3_1 _0787_ (.B(_0227_),
    .C(_0232_),
    .A(\vga.interval_counter[19] ),
    .Y(_0236_));
 sg13g2_xor2_1 _0788_ (.B(_0236_),
    .A(\vga.interval_counter[20] ),
    .X(_0237_));
 sg13g2_nor2_1 _0789_ (.A(net28),
    .B(_0237_),
    .Y(_0068_));
 sg13g2_and4_1 _0790_ (.A(\vga.interval_counter[19] ),
    .B(\vga.interval_counter[20] ),
    .C(_0227_),
    .D(_0232_),
    .X(_0238_));
 sg13g2_buf_8 _0791_ (.A(_0238_),
    .X(_0239_));
 sg13g2_xnor2_1 _0792_ (.Y(_0240_),
    .A(\vga.interval_counter[21] ),
    .B(_0239_));
 sg13g2_nor2_1 _0793_ (.A(net28),
    .B(_0240_),
    .Y(_0069_));
 sg13g2_nand2_1 _0794_ (.Y(_0241_),
    .A(\vga.interval_counter[21] ),
    .B(_0239_));
 sg13g2_xor2_1 _0795_ (.B(_0241_),
    .A(\vga.interval_counter[22] ),
    .X(_0242_));
 sg13g2_nor2_1 _0796_ (.A(_0231_),
    .B(_0242_),
    .Y(_0070_));
 sg13g2_nand3_1 _0797_ (.B(\vga.interval_counter[22] ),
    .C(_0239_),
    .A(\vga.interval_counter[21] ),
    .Y(_0243_));
 sg13g2_xor2_1 _0798_ (.B(_0243_),
    .A(\vga.interval_counter[23] ),
    .X(_0244_));
 sg13g2_nor2_1 _0799_ (.A(net28),
    .B(_0244_),
    .Y(_0071_));
 sg13g2_nand4_1 _0800_ (.B(\vga.interval_counter[23] ),
    .C(\vga.interval_counter[22] ),
    .A(\vga.interval_counter[21] ),
    .Y(_0245_),
    .D(_0239_));
 sg13g2_xor2_1 _0801_ (.B(_0245_),
    .A(\vga.interval_counter[24] ),
    .X(_0246_));
 sg13g2_nor2_1 _0802_ (.A(net28),
    .B(_0246_),
    .Y(_0072_));
 sg13g2_nand2_1 _0803_ (.Y(_0247_),
    .A(_0141_),
    .B(_0142_));
 sg13g2_xor2_1 _0804_ (.B(_0247_),
    .A(\vga.interval_counter[2] ),
    .X(_0248_));
 sg13g2_nor2_1 _0805_ (.A(net28),
    .B(_0248_),
    .Y(_0073_));
 sg13g2_nand3_1 _0806_ (.B(_0142_),
    .C(\vga.interval_counter[2] ),
    .A(_0141_),
    .Y(_0249_));
 sg13g2_xor2_1 _0807_ (.B(_0249_),
    .A(\vga.interval_counter[3] ),
    .X(_0250_));
 sg13g2_nor2_1 _0808_ (.A(net28),
    .B(_0250_),
    .Y(_0074_));
 sg13g2_xnor2_1 _0809_ (.Y(_0251_),
    .A(\vga.interval_counter[4] ),
    .B(_0207_));
 sg13g2_nor2_1 _0810_ (.A(net28),
    .B(_0251_),
    .Y(_0075_));
 sg13g2_nand2_1 _0811_ (.Y(_0252_),
    .A(\vga.interval_counter[4] ),
    .B(_0207_));
 sg13g2_xnor2_1 _0812_ (.Y(_0253_),
    .A(_0145_),
    .B(_0252_));
 sg13g2_nor2_1 _0813_ (.A(_0205_),
    .B(_0253_),
    .Y(_0076_));
 sg13g2_xnor2_1 _0814_ (.Y(_0254_),
    .A(\vga.interval_counter[6] ),
    .B(_0208_));
 sg13g2_nor2_1 _0815_ (.A(_0205_),
    .B(_0254_),
    .Y(_0077_));
 sg13g2_nand2_1 _0816_ (.Y(_0255_),
    .A(\vga.interval_counter[6] ),
    .B(_0208_));
 sg13g2_xor2_1 _0817_ (.B(_0255_),
    .A(\vga.interval_counter[7] ),
    .X(_0256_));
 sg13g2_nor2_1 _0818_ (.A(_0205_),
    .B(_0256_),
    .Y(_0078_));
 sg13g2_inv_1 _0819_ (.Y(_0257_),
    .A(\vga.interval_counter[8] ));
 sg13g2_xnor2_1 _0820_ (.Y(_0258_),
    .A(_0257_),
    .B(_0210_));
 sg13g2_nor2_1 _0821_ (.A(_0205_),
    .B(_0258_),
    .Y(_0079_));
 sg13g2_nor2_1 _0822_ (.A(_0257_),
    .B(_0210_),
    .Y(_0259_));
 sg13g2_xnor2_1 _0823_ (.Y(_0260_),
    .A(\vga.interval_counter[9] ),
    .B(_0259_));
 sg13g2_nor2_1 _0824_ (.A(_0205_),
    .B(_0260_),
    .Y(_0080_));
 sg13g2_and3_1 _0825_ (.X(_0082_),
    .A(\vga.left_1d ),
    .B(net1),
    .C(_0153_));
 sg13g2_nand2_1 _0826_ (.Y(_0261_),
    .A(_0123_),
    .B(_0111_));
 sg13g2_a21oi_1 _0827_ (.A1(_0008_),
    .A2(_0261_),
    .Y(_0262_),
    .B1(_0104_));
 sg13g2_nor3_1 _0828_ (.A(\vga.count_v[5] ),
    .B(\vga.count_v[3] ),
    .C(_0100_),
    .Y(_0263_));
 sg13g2_nor2b_1 _0829_ (.A(_0262_),
    .B_N(_0263_),
    .Y(_0264_));
 sg13g2_nor2b_1 _0830_ (.A(_0264_),
    .B_N(_0110_),
    .Y(_0265_));
 sg13g2_nand2_1 _0831_ (.Y(_0266_),
    .A(net54),
    .B(_0111_));
 sg13g2_nor2_1 _0832_ (.A(_0095_),
    .B(_0099_),
    .Y(_0267_));
 sg13g2_a21oi_1 _0833_ (.A1(_0266_),
    .A2(_0267_),
    .Y(_0268_),
    .B1(_0101_));
 sg13g2_nor3_1 _0834_ (.A(_0110_),
    .B(net53),
    .C(_0268_),
    .Y(_0269_));
 sg13g2_nor3_1 _0835_ (.A(_0112_),
    .B(_0265_),
    .C(_0269_),
    .Y(_0270_));
 sg13g2_nor2_1 _0836_ (.A(_0160_),
    .B(net46),
    .Y(_0271_));
 sg13g2_and2_1 _0837_ (.A(net47),
    .B(net45),
    .X(_0272_));
 sg13g2_nand2b_1 _0838_ (.Y(_0273_),
    .B(_0272_),
    .A_N(_0271_));
 sg13g2_buf_1 _0839_ (.A(\vga.count_h[8] ),
    .X(_0274_));
 sg13g2_nand2_1 _0840_ (.Y(_0275_),
    .A(net50),
    .B(\vga.count_h[5] ));
 sg13g2_nand2b_1 _0841_ (.Y(_0276_),
    .B(_0275_),
    .A_N(\vga.count_h[7] ));
 sg13g2_buf_1 _0842_ (.A(\vga.count_h[9] ),
    .X(_0277_));
 sg13g2_a21oi_1 _0843_ (.A1(net44),
    .A2(_0276_),
    .Y(_0278_),
    .B1(_0277_));
 sg13g2_nand2b_1 _0844_ (.Y(_0279_),
    .B(net44),
    .A_N(\vga.count_h[7] ));
 sg13g2_nor4_1 _0845_ (.A(\vga.count_h[9] ),
    .B(net48),
    .C(_0275_),
    .D(_0279_),
    .Y(_0280_));
 sg13g2_nand3_1 _0846_ (.B(_0271_),
    .C(_0280_),
    .A(_0272_),
    .Y(_0281_));
 sg13g2_o21ai_1 _0847_ (.B1(_0281_),
    .Y(_0282_),
    .A1(_0273_),
    .A2(_0278_));
 sg13g2_a21oi_1 _0848_ (.A1(_0155_),
    .A2(net44),
    .Y(_0283_),
    .B1(\vga.count_h[9] ));
 sg13g2_nand4_1 _0849_ (.B(net50),
    .C(\vga.count_h[5] ),
    .A(_0274_),
    .Y(_0284_),
    .D(net48));
 sg13g2_and2_1 _0850_ (.A(_0283_),
    .B(_0284_),
    .X(_0285_));
 sg13g2_inv_1 _0851_ (.Y(_0286_),
    .A(net50));
 sg13g2_or3_1 _0852_ (.A(_0286_),
    .B(_0277_),
    .C(_0279_),
    .X(_0287_));
 sg13g2_nor2_1 _0853_ (.A(_0287_),
    .B(_0285_),
    .Y(_0288_));
 sg13g2_nand3b_1 _0854_ (.B(_0158_),
    .C(_0157_),
    .Y(_0289_),
    .A_N(net46));
 sg13g2_a21oi_1 _0855_ (.A1(net47),
    .A2(_0289_),
    .Y(_0290_),
    .B1(net45));
 sg13g2_a22oi_1 _0856_ (.Y(_0291_),
    .B1(_0288_),
    .B2(_0290_),
    .A2(_0285_),
    .A1(_0282_));
 sg13g2_inv_1 _0857_ (.Y(_0292_),
    .A(\vga.score_ten_enable ));
 sg13g2_nand2_1 _0858_ (.Y(_0293_),
    .A(_0160_),
    .B(net46));
 sg13g2_nand2b_1 _0859_ (.Y(_0294_),
    .B(_0293_),
    .A_N(net47));
 sg13g2_o21ai_1 _0860_ (.B1(_0273_),
    .Y(_0295_),
    .A1(net45),
    .A2(_0294_));
 sg13g2_nor4_1 _0861_ (.A(net49),
    .B(_0159_),
    .C(_0295_),
    .D(_0287_),
    .Y(_0296_));
 sg13g2_nor2b_1 _0862_ (.A(_0282_),
    .B_N(_0285_),
    .Y(_0297_));
 sg13g2_inv_1 _0863_ (.Y(_0298_),
    .A(\vga.score_unit_pixels[2] ));
 sg13g2_nor3_1 _0864_ (.A(net47),
    .B(net46),
    .C(net45),
    .Y(_0299_));
 sg13g2_a21oi_1 _0865_ (.A1(_0280_),
    .A2(_0299_),
    .Y(_0300_),
    .B1(_0278_));
 sg13g2_and2_1 _0866_ (.A(_0298_),
    .B(_0300_),
    .X(_0301_));
 sg13g2_a22oi_1 _0867_ (.Y(_0302_),
    .B1(_0297_),
    .B2(_0301_),
    .A2(_0296_),
    .A1(_0292_));
 sg13g2_o21ai_1 _0868_ (.B1(_0302_),
    .Y(_0303_),
    .A1(\vga.score_unit_pixels[1] ),
    .A2(_0291_));
 sg13g2_and2_1 _0869_ (.A(\vga.car_pos_h[5] ),
    .B(\vga.car_pos_h[4] ),
    .X(_0304_));
 sg13g2_buf_2 _0870_ (.A(_0304_),
    .X(_0305_));
 sg13g2_buf_1 _0871_ (.A(\vga.car_pos_h[5] ),
    .X(_0306_));
 sg13g2_nor2_2 _0872_ (.A(net42),
    .B(\vga.car_pos_h[4] ),
    .Y(_0307_));
 sg13g2_inv_1 _0873_ (.Y(_0308_),
    .A(_0014_));
 sg13g2_mux2_1 _0874_ (.A0(_0305_),
    .A1(_0307_),
    .S(_0308_),
    .X(_0309_));
 sg13g2_buf_1 _0875_ (.A(\vga.car_pos_h[4] ),
    .X(_0310_));
 sg13g2_xnor2_1 _0876_ (.Y(_0311_),
    .A(_0306_),
    .B(net41));
 sg13g2_nor3_1 _0877_ (.A(_0005_),
    .B(_0014_),
    .C(_0311_),
    .Y(_0312_));
 sg13g2_a221oi_1 _0878_ (.B2(_0005_),
    .C1(_0312_),
    .B1(_0309_),
    .A1(net50),
    .Y(_0313_),
    .A2(_0305_));
 sg13g2_nor2b_1 _0879_ (.A(_0017_),
    .B_N(_0313_),
    .Y(_0314_));
 sg13g2_mux2_1 _0880_ (.A0(_0305_),
    .A1(_0307_),
    .S(_0014_),
    .X(_0315_));
 sg13g2_nor2_1 _0881_ (.A(_0005_),
    .B(_0308_),
    .Y(_0316_));
 sg13g2_xor2_1 _0882_ (.B(net41),
    .A(net42),
    .X(_0317_));
 sg13g2_o21ai_1 _0883_ (.B1(_0017_),
    .Y(_0318_),
    .A1(_0286_),
    .A2(_0305_));
 sg13g2_a221oi_1 _0884_ (.B2(_0317_),
    .C1(_0318_),
    .B1(_0316_),
    .A1(_0005_),
    .Y(_0319_),
    .A2(_0315_));
 sg13g2_xor2_1 _0885_ (.B(_0017_),
    .A(_0014_),
    .X(_0320_));
 sg13g2_nor3_1 _0886_ (.A(_0005_),
    .B(net42),
    .C(_0320_),
    .Y(_0321_));
 sg13g2_a21o_1 _0887_ (.A2(_0320_),
    .A1(_0305_),
    .B1(_0321_),
    .X(_0322_));
 sg13g2_nand2_1 _0888_ (.Y(_0323_),
    .A(net49),
    .B(_0322_));
 sg13g2_o21ai_1 _0889_ (.B1(_0323_),
    .Y(_0324_),
    .A1(_0314_),
    .A2(_0319_));
 sg13g2_xor2_1 _0890_ (.B(_0305_),
    .A(_0017_),
    .X(_0325_));
 sg13g2_a22oi_1 _0891_ (.Y(_0326_),
    .B1(_0325_),
    .B2(net50),
    .A2(_0311_),
    .A1(net49));
 sg13g2_inv_1 _0892_ (.Y(_0327_),
    .A(_0310_));
 sg13g2_buf_1 _0893_ (.A(\vga.car_pos_h[3] ),
    .X(_0328_));
 sg13g2_xor2_1 _0894_ (.B(net40),
    .A(net45),
    .X(_0329_));
 sg13g2_buf_1 _0895_ (.A(\vga.car_pos_h[1] ),
    .X(_0330_));
 sg13g2_nor2b_1 _0896_ (.A(net46),
    .B_N(_0330_),
    .Y(_0331_));
 sg13g2_nor2_1 _0897_ (.A(_0329_),
    .B(_0331_),
    .Y(_0332_));
 sg13g2_nand2b_1 _0898_ (.Y(_0333_),
    .B(net46),
    .A_N(_0330_));
 sg13g2_nor2b_1 _0899_ (.A(_0160_),
    .B_N(\vga.car_pos_h[0] ),
    .Y(_0334_));
 sg13g2_xor2_1 _0900_ (.B(\vga.car_pos_h[2] ),
    .A(net47),
    .X(_0335_));
 sg13g2_a21oi_1 _0901_ (.A1(_0333_),
    .A2(_0334_),
    .Y(_0336_),
    .B1(_0335_));
 sg13g2_nor2b_1 _0902_ (.A(net45),
    .B_N(net40),
    .Y(_0337_));
 sg13g2_nand2b_1 _0903_ (.Y(_0338_),
    .B(net47),
    .A_N(\vga.car_pos_h[2] ));
 sg13g2_nand2b_1 _0904_ (.Y(_0339_),
    .B(net45),
    .A_N(_0328_));
 sg13g2_o21ai_1 _0905_ (.B1(_0339_),
    .Y(_0340_),
    .A1(_0337_),
    .A2(_0338_));
 sg13g2_a21oi_1 _0906_ (.A1(_0332_),
    .A2(_0336_),
    .Y(_0341_),
    .B1(_0340_));
 sg13g2_nor3_1 _0907_ (.A(_0327_),
    .B(_0329_),
    .C(_0331_),
    .Y(_0342_));
 sg13g2_a221oi_1 _0908_ (.B2(_0336_),
    .C1(net48),
    .B1(_0342_),
    .A1(net41),
    .Y(_0343_),
    .A2(_0340_));
 sg13g2_a21o_1 _0909_ (.A2(_0341_),
    .A1(_0327_),
    .B1(_0343_),
    .X(_0344_));
 sg13g2_nand2_1 _0910_ (.Y(_0345_),
    .A(_0326_),
    .B(_0344_));
 sg13g2_buf_1 _0911_ (.A(\vga.car_pos_h[6] ),
    .X(_0346_));
 sg13g2_and3_1 _0912_ (.X(_0347_),
    .A(net38),
    .B(net42),
    .C(\vga.car_pos_h[4] ));
 sg13g2_xor2_1 _0913_ (.B(_0347_),
    .A(_0016_),
    .X(_0348_));
 sg13g2_buf_2 _0914_ (.A(_0011_),
    .X(_0349_));
 sg13g2_buf_1 _0915_ (.A(\vga.car_pos_h[8] ),
    .X(_0350_));
 sg13g2_buf_1 _0916_ (.A(\vga.car_pos_h[7] ),
    .X(_0351_));
 sg13g2_nand3_1 _0917_ (.B(net36),
    .C(_0347_),
    .A(net37),
    .Y(_0352_));
 sg13g2_xnor2_1 _0918_ (.Y(_0353_),
    .A(_0349_),
    .B(_0352_));
 sg13g2_nand4_1 _0919_ (.B(net38),
    .C(_0306_),
    .A(net36),
    .Y(_0354_),
    .D(net41));
 sg13g2_xor2_1 _0920_ (.B(_0354_),
    .A(_0015_),
    .X(_0355_));
 sg13g2_nor2_1 _0921_ (.A(_0013_),
    .B(_0355_),
    .Y(_0356_));
 sg13g2_a21o_1 _0922_ (.A2(_0353_),
    .A1(net43),
    .B1(_0356_),
    .X(_0357_));
 sg13g2_a221oi_1 _0923_ (.B2(_0155_),
    .C1(_0357_),
    .B1(_0348_),
    .A1(_0324_),
    .Y(_0358_),
    .A2(_0345_));
 sg13g2_nand2_1 _0924_ (.Y(_0359_),
    .A(_0013_),
    .B(_0355_));
 sg13g2_a21o_1 _0925_ (.A2(_0359_),
    .A1(_0007_),
    .B1(net43),
    .X(_0360_));
 sg13g2_inv_1 _0926_ (.Y(_0361_),
    .A(\vga.car_pos_h[9] ));
 sg13g2_nand2b_1 _0927_ (.Y(_0362_),
    .B(_0361_),
    .A_N(_0352_));
 sg13g2_nand2_1 _0928_ (.Y(_0363_),
    .A(_0349_),
    .B(_0352_));
 sg13g2_o21ai_1 _0929_ (.B1(_0363_),
    .Y(_0364_),
    .A1(_0349_),
    .A2(_0362_));
 sg13g2_nor2_1 _0930_ (.A(_0349_),
    .B(_0352_),
    .Y(_0365_));
 sg13g2_a21oi_1 _0931_ (.A1(_0349_),
    .A2(_0362_),
    .Y(_0366_),
    .B1(_0365_));
 sg13g2_a21oi_1 _0932_ (.A1(_0013_),
    .A2(_0355_),
    .Y(_0367_),
    .B1(_0007_));
 sg13g2_a22oi_1 _0933_ (.Y(_0368_),
    .B1(_0366_),
    .B2(_0367_),
    .A2(_0364_),
    .A1(_0360_));
 sg13g2_nor3_1 _0934_ (.A(net51),
    .B(_0357_),
    .C(_0348_),
    .Y(_0369_));
 sg13g2_or2_1 _0935_ (.X(_0370_),
    .B(_0369_),
    .A(_0368_));
 sg13g2_or4_1 _0936_ (.A(net36),
    .B(\vga.car_pos_h[6] ),
    .C(\vga.car_pos_h[5] ),
    .D(\vga.car_pos_h[4] ),
    .X(_0371_));
 sg13g2_buf_1 _0937_ (.A(_0371_),
    .X(_0372_));
 sg13g2_nor2_1 _0938_ (.A(net37),
    .B(_0372_),
    .Y(_0373_));
 sg13g2_mux2_1 _0939_ (.A0(_0373_),
    .A1(_0372_),
    .S(_0349_),
    .X(_0374_));
 sg13g2_nor2_1 _0940_ (.A(net37),
    .B(_0013_),
    .Y(_0375_));
 sg13g2_nand2_1 _0941_ (.Y(_0376_),
    .A(\vga.count_h[9] ),
    .B(_0349_));
 sg13g2_o21ai_1 _0942_ (.B1(_0376_),
    .Y(_0377_),
    .A1(_0013_),
    .A2(_0372_));
 sg13g2_and2_1 _0943_ (.A(net37),
    .B(_0377_),
    .X(_0378_));
 sg13g2_a221oi_1 _0944_ (.B2(_0372_),
    .C1(_0378_),
    .B1(_0375_),
    .A1(net43),
    .Y(_0379_),
    .A2(_0374_));
 sg13g2_inv_1 _0945_ (.Y(_0380_),
    .A(_0012_));
 sg13g2_xnor2_1 _0946_ (.Y(_0381_),
    .A(net44),
    .B(net37));
 sg13g2_nand2_1 _0947_ (.Y(_0382_),
    .A(_0351_),
    .B(_0381_));
 sg13g2_o21ai_1 _0948_ (.B1(_0382_),
    .Y(_0383_),
    .A1(_0372_),
    .A2(_0381_));
 sg13g2_or2_1 _0949_ (.X(_0384_),
    .B(net41),
    .A(net42));
 sg13g2_o21ai_1 _0950_ (.B1(net36),
    .Y(_0385_),
    .A1(net38),
    .A2(_0384_));
 sg13g2_and2_1 _0951_ (.A(_0372_),
    .B(_0385_),
    .X(_0386_));
 sg13g2_a22oi_1 _0952_ (.Y(_0387_),
    .B1(_0386_),
    .B2(_0381_),
    .A2(_0383_),
    .A1(_0380_));
 sg13g2_nor3_1 _0953_ (.A(_0329_),
    .B(_0331_),
    .C(_0335_),
    .Y(_0388_));
 sg13g2_o21ai_1 _0954_ (.B1(_0333_),
    .Y(_0389_),
    .A1(net48),
    .A2(_0310_));
 sg13g2_buf_1 _0955_ (.A(\vga.car_pos_h[0] ),
    .X(_0390_));
 sg13g2_nor2b_1 _0956_ (.A(net35),
    .B_N(_0160_),
    .Y(_0391_));
 sg13g2_nor3_1 _0957_ (.A(_0334_),
    .B(_0389_),
    .C(_0391_),
    .Y(_0392_));
 sg13g2_a22oi_1 _0958_ (.Y(_0393_),
    .B1(_0388_),
    .B2(_0392_),
    .A2(_0317_),
    .A1(net49));
 sg13g2_xor2_1 _0959_ (.B(_0346_),
    .A(net50),
    .X(_0394_));
 sg13g2_nand2_1 _0960_ (.Y(_0395_),
    .A(_0307_),
    .B(_0394_));
 sg13g2_o21ai_1 _0961_ (.B1(_0395_),
    .Y(_0396_),
    .A1(_0327_),
    .A2(_0394_));
 sg13g2_nor2_1 _0962_ (.A(_0311_),
    .B(_0394_),
    .Y(_0397_));
 sg13g2_a21oi_1 _0963_ (.A1(net49),
    .A2(_0396_),
    .Y(_0398_),
    .B1(_0397_));
 sg13g2_a21o_1 _0964_ (.A2(_0393_),
    .A1(_0344_),
    .B1(_0398_),
    .X(_0399_));
 sg13g2_xnor2_1 _0965_ (.Y(_0400_),
    .A(net38),
    .B(_0307_));
 sg13g2_a22oi_1 _0966_ (.Y(_0401_),
    .B1(_0400_),
    .B2(_0308_),
    .A2(_0386_),
    .A1(_0380_));
 sg13g2_and2_1 _0967_ (.A(_0379_),
    .B(_0401_),
    .X(_0402_));
 sg13g2_xor2_1 _0968_ (.B(_0373_),
    .A(_0349_),
    .X(_0403_));
 sg13g2_nand3_1 _0969_ (.B(net54),
    .C(_0111_),
    .A(net52),
    .Y(_0404_));
 sg13g2_nand3_1 _0970_ (.B(\vga.count_v[7] ),
    .C(_0110_),
    .A(\vga.count_v[8] ),
    .Y(_0405_));
 sg13g2_a21o_1 _0971_ (.A2(_0404_),
    .A1(_0263_),
    .B1(_0405_),
    .X(_0406_));
 sg13g2_inv_1 _0972_ (.Y(_0407_),
    .A(\vga.count_v[9] ));
 sg13g2_a22oi_1 _0973_ (.Y(_0408_),
    .B1(_0406_),
    .B2(_0407_),
    .A2(_0373_),
    .A1(_0361_));
 sg13g2_o21ai_1 _0974_ (.B1(_0408_),
    .Y(_0409_),
    .A1(net43),
    .A2(_0403_));
 sg13g2_a221oi_1 _0975_ (.B2(_0402_),
    .C1(_0409_),
    .B1(_0399_),
    .A1(_0379_),
    .Y(_0410_),
    .A2(_0387_));
 sg13g2_o21ai_1 _0976_ (.B1(_0410_),
    .Y(_0411_),
    .A1(_0358_),
    .A2(_0370_));
 sg13g2_nand2_1 _0977_ (.Y(_0412_),
    .A(\vga.score_unit_pixels[2] ),
    .B(_0300_));
 sg13g2_a221oi_1 _0978_ (.B2(_0412_),
    .C1(net43),
    .B1(_0297_),
    .A1(net51),
    .Y(_0413_),
    .A2(_0274_));
 sg13g2_o21ai_1 _0979_ (.B1(_0270_),
    .Y(_0414_),
    .A1(_0296_),
    .A2(_0413_));
 sg13g2_inv_2 _0980_ (.Y(_0415_),
    .A(_0094_));
 sg13g2_or3_1 _0981_ (.A(_0415_),
    .B(\vga.blank_h ),
    .C(\vga.blank_v ),
    .X(_0416_));
 sg13g2_a221oi_1 _0982_ (.B2(_0414_),
    .C1(_0416_),
    .B1(_0411_),
    .A1(_0270_),
    .Y(_0083_),
    .A2(_0303_));
 sg13g2_and3_1 _0983_ (.X(_0085_),
    .A(\vga.right_1d ),
    .B(net2),
    .C(_0153_));
 sg13g2_nand2_1 _0984_ (.Y(_0417_),
    .A(net48),
    .B(_0165_));
 sg13g2_nor2_2 _0985_ (.A(_0275_),
    .B(_0417_),
    .Y(_0418_));
 sg13g2_nor2b_1 _0986_ (.A(_0007_),
    .B_N(_0170_),
    .Y(_0419_));
 sg13g2_mux2_1 _0987_ (.A0(_0418_),
    .A1(_0419_),
    .S(net51),
    .X(_0420_));
 sg13g2_a21o_1 _0988_ (.A2(_0420_),
    .A1(_0154_),
    .B1(_0415_),
    .X(_0421_));
 sg13g2_inv_1 _0989_ (.Y(_0422_),
    .A(_0005_));
 sg13g2_nor3_1 _0990_ (.A(\vga.count_h[7] ),
    .B(_0156_),
    .C(_0422_),
    .Y(_0423_));
 sg13g2_o21ai_1 _0991_ (.B1(_0423_),
    .Y(_0424_),
    .A1(\vga.count_h[5] ),
    .A2(_0417_));
 sg13g2_and3_1 _0992_ (.X(_0425_),
    .A(net44),
    .B(net43),
    .C(_0424_));
 sg13g2_buf_2 _0993_ (.A(_0425_),
    .X(_0426_));
 sg13g2_and2_1 _0994_ (.A(_0169_),
    .B(_0426_),
    .X(_0427_));
 sg13g2_buf_1 _0995_ (.A(_0427_),
    .X(_0428_));
 sg13g2_nand2b_1 _0996_ (.Y(_0429_),
    .B(\vga.blank_h ),
    .A_N(net30));
 sg13g2_nand2b_1 _0997_ (.Y(_0022_),
    .B(_0429_),
    .A_N(_0421_));
 sg13g2_buf_1 _0998_ (.A(_0094_),
    .X(_0430_));
 sg13g2_nand4_1 _0999_ (.B(net52),
    .C(net54),
    .A(\vga.count_v[3] ),
    .Y(_0431_),
    .D(_0111_));
 sg13g2_nor4_1 _1000_ (.A(\vga.count_v[8] ),
    .B(\vga.count_v[7] ),
    .C(\vga.count_v[5] ),
    .D(_0100_),
    .Y(_0432_));
 sg13g2_nand3b_1 _1001_ (.B(_0432_),
    .C(\vga.count_v[9] ),
    .Y(_0433_),
    .A_N(_0110_));
 sg13g2_mux2_1 _1002_ (.A0(_0431_),
    .A1(_0006_),
    .S(_0433_),
    .X(_0434_));
 sg13g2_nor2_1 _1003_ (.A(_0101_),
    .B(_0431_),
    .Y(_0435_));
 sg13g2_nor2_1 _1004_ (.A(_0098_),
    .B(_0435_),
    .Y(_0436_));
 sg13g2_o21ai_1 _1005_ (.B1(_0407_),
    .Y(_0437_),
    .A1(_0405_),
    .A2(_0436_));
 sg13g2_nand3_1 _1006_ (.B(_0434_),
    .C(_0437_),
    .A(_0426_),
    .Y(_0438_));
 sg13g2_nand2_1 _1007_ (.Y(_0439_),
    .A(_0426_),
    .B(_0437_));
 sg13g2_nand2_1 _1008_ (.Y(_0440_),
    .A(\vga.blank_v ),
    .B(_0439_));
 sg13g2_nand3_1 _1009_ (.B(_0438_),
    .C(_0440_),
    .A(net34),
    .Y(_0023_));
 sg13g2_inv_1 _1010_ (.Y(_0024_),
    .A(_0416_));
 sg13g2_nor4_1 _1011_ (.A(\vga.car_pos_h[9] ),
    .B(_0350_),
    .C(net36),
    .D(net38),
    .Y(_0441_));
 sg13g2_nor2b_1 _1012_ (.A(net42),
    .B_N(_0441_),
    .Y(_0442_));
 sg13g2_nor4_1 _1013_ (.A(net39),
    .B(net35),
    .C(_0328_),
    .D(\vga.car_pos_h[2] ),
    .Y(_0443_));
 sg13g2_nand2b_1 _1014_ (.Y(_0444_),
    .B(net41),
    .A_N(_0443_));
 sg13g2_inv_1 _1015_ (.Y(_0445_),
    .A(\vga.left_pressed ));
 sg13g2_a21oi_2 _1016_ (.B1(_0445_),
    .Y(_0446_),
    .A2(_0444_),
    .A1(_0442_));
 sg13g2_and2_1 _1017_ (.A(net39),
    .B(\vga.car_pos_h[0] ),
    .X(_0447_));
 sg13g2_and4_1 _1018_ (.A(net38),
    .B(\vga.car_pos_h[5] ),
    .C(\vga.car_pos_h[3] ),
    .D(\vga.car_pos_h[2] ),
    .X(_0448_));
 sg13g2_or2_1 _1019_ (.X(_0449_),
    .B(_0351_),
    .A(net37));
 sg13g2_a221oi_1 _1020_ (.B2(_0448_),
    .C1(_0449_),
    .B1(_0447_),
    .A1(_0346_),
    .Y(_0450_),
    .A2(_0305_));
 sg13g2_o21ai_1 _1021_ (.B1(\vga.right_pressed ),
    .Y(_0451_),
    .A1(_0361_),
    .A2(_0450_));
 sg13g2_inv_1 _1022_ (.Y(_0452_),
    .A(_0451_));
 sg13g2_nor2_1 _1023_ (.A(_0446_),
    .B(_0452_),
    .Y(_0453_));
 sg13g2_nand2_1 _1024_ (.Y(_0454_),
    .A(net35),
    .B(_0453_));
 sg13g2_o21ai_1 _1025_ (.B1(_0019_),
    .Y(_0455_),
    .A1(_0446_),
    .A2(_0452_));
 sg13g2_nand3_1 _1026_ (.B(_0454_),
    .C(_0455_),
    .A(net34),
    .Y(_0025_));
 sg13g2_buf_1 _1027_ (.A(_0094_),
    .X(_0456_));
 sg13g2_buf_1 _1028_ (.A(_0451_),
    .X(_0457_));
 sg13g2_nand3_1 _1029_ (.B(_0446_),
    .C(net31),
    .A(_0019_),
    .Y(_0458_));
 sg13g2_o21ai_1 _1030_ (.B1(_0458_),
    .Y(_0459_),
    .A1(_0019_),
    .A2(net31));
 sg13g2_xnor2_1 _1031_ (.Y(_0460_),
    .A(net39),
    .B(_0459_));
 sg13g2_nand2_1 _1032_ (.Y(_0026_),
    .A(net33),
    .B(_0460_));
 sg13g2_buf_1 _1033_ (.A(_0018_),
    .X(_0461_));
 sg13g2_nor2_1 _1034_ (.A(net39),
    .B(_0461_),
    .Y(_0462_));
 sg13g2_a21o_1 _1035_ (.A2(_0446_),
    .A1(net35),
    .B1(_0452_),
    .X(_0463_));
 sg13g2_a22oi_1 _1036_ (.Y(_0464_),
    .B1(_0462_),
    .B2(_0463_),
    .A2(_0453_),
    .A1(\vga.car_pos_h[2] ));
 sg13g2_nand2_1 _1037_ (.Y(_0465_),
    .A(_0446_),
    .B(net31));
 sg13g2_nand3_1 _1038_ (.B(_0461_),
    .C(_0452_),
    .A(_0390_),
    .Y(_0466_));
 sg13g2_o21ai_1 _1039_ (.B1(_0466_),
    .Y(_0467_),
    .A1(_0461_),
    .A2(_0465_));
 sg13g2_and2_1 _1040_ (.A(_0446_),
    .B(net31),
    .X(_0468_));
 sg13g2_nor2b_1 _1041_ (.A(net39),
    .B_N(_0461_),
    .Y(_0469_));
 sg13g2_nor2_1 _1042_ (.A(_0461_),
    .B(_0457_),
    .Y(_0470_));
 sg13g2_a21oi_1 _1043_ (.A1(_0468_),
    .A2(_0469_),
    .Y(_0471_),
    .B1(_0470_));
 sg13g2_nor2_1 _1044_ (.A(_0390_),
    .B(_0471_),
    .Y(_0472_));
 sg13g2_a21oi_1 _1045_ (.A1(net39),
    .A2(_0467_),
    .Y(_0473_),
    .B1(_0472_));
 sg13g2_nand3_1 _1046_ (.B(_0464_),
    .C(_0473_),
    .A(net34),
    .Y(_0027_));
 sg13g2_nor2b_1 _1047_ (.A(net35),
    .B_N(_0469_),
    .Y(_0474_));
 sg13g2_a22oi_1 _1048_ (.Y(_0475_),
    .B1(_0474_),
    .B2(_0468_),
    .A2(_0470_),
    .A1(_0447_));
 sg13g2_xor2_1 _1049_ (.B(_0475_),
    .A(net40),
    .X(_0476_));
 sg13g2_nand2_1 _1050_ (.Y(_0028_),
    .A(net33),
    .B(_0476_));
 sg13g2_inv_1 _1051_ (.Y(_0477_),
    .A(_0461_));
 sg13g2_nor3_1 _1052_ (.A(net35),
    .B(net40),
    .C(_0477_),
    .Y(_0478_));
 sg13g2_nor2b_1 _1053_ (.A(_0461_),
    .B_N(net40),
    .Y(_0479_));
 sg13g2_and2_1 _1054_ (.A(net35),
    .B(_0479_),
    .X(_0480_));
 sg13g2_o21ai_1 _1055_ (.B1(net39),
    .Y(_0481_),
    .A1(_0451_),
    .A2(_0480_));
 sg13g2_o21ai_1 _1056_ (.B1(_0481_),
    .Y(_0482_),
    .A1(_0452_),
    .A2(_0478_));
 sg13g2_mux2_1 _1057_ (.A0(_0465_),
    .A1(net31),
    .S(_0482_),
    .X(_0483_));
 sg13g2_xnor2_1 _1058_ (.Y(_0484_),
    .A(_0327_),
    .B(_0483_));
 sg13g2_nand2_1 _1059_ (.Y(_0029_),
    .A(net33),
    .B(_0484_));
 sg13g2_nor2_1 _1060_ (.A(_0327_),
    .B(_0019_),
    .Y(_0485_));
 sg13g2_nand4_1 _1061_ (.B(net40),
    .C(_0470_),
    .A(net39),
    .Y(_0486_),
    .D(_0485_));
 sg13g2_nor2_1 _1062_ (.A(net41),
    .B(net40),
    .Y(_0487_));
 sg13g2_nand4_1 _1063_ (.B(_0457_),
    .C(_0469_),
    .A(_0019_),
    .Y(_0488_),
    .D(_0487_));
 sg13g2_a21oi_1 _1064_ (.A1(_0486_),
    .A2(_0488_),
    .Y(_0489_),
    .B1(_0453_));
 sg13g2_xnor2_1 _1065_ (.Y(_0490_),
    .A(net42),
    .B(_0489_));
 sg13g2_nand2_1 _1066_ (.Y(_0030_),
    .A(net33),
    .B(_0490_));
 sg13g2_nor2_1 _1067_ (.A(_0384_),
    .B(_0465_),
    .Y(_0491_));
 sg13g2_and2_1 _1068_ (.A(_0305_),
    .B(_0452_),
    .X(_0492_));
 sg13g2_mux2_1 _1069_ (.A0(_0491_),
    .A1(_0492_),
    .S(_0482_),
    .X(_0493_));
 sg13g2_xnor2_1 _1070_ (.Y(_0494_),
    .A(net38),
    .B(_0493_));
 sg13g2_nor2_1 _1071_ (.A(_0415_),
    .B(_0494_),
    .Y(_0031_));
 sg13g2_nand3_1 _1072_ (.B(_0447_),
    .C(_0479_),
    .A(_0347_),
    .Y(_0495_));
 sg13g2_nor4_1 _1073_ (.A(net42),
    .B(net41),
    .C(net35),
    .D(net40),
    .Y(_0496_));
 sg13g2_a21oi_1 _1074_ (.A1(_0469_),
    .A2(_0496_),
    .Y(_0497_),
    .B1(net38));
 sg13g2_nor2b_1 _1075_ (.A(_0497_),
    .B_N(_0017_),
    .Y(_0498_));
 sg13g2_nand3_1 _1076_ (.B(net31),
    .C(_0498_),
    .A(_0446_),
    .Y(_0499_));
 sg13g2_o21ai_1 _1077_ (.B1(_0499_),
    .Y(_0500_),
    .A1(net31),
    .A2(_0495_));
 sg13g2_xnor2_1 _1078_ (.Y(_0501_),
    .A(net36),
    .B(_0500_));
 sg13g2_nor2_1 _1079_ (.A(_0415_),
    .B(_0501_),
    .Y(_0032_));
 sg13g2_o21ai_1 _1080_ (.B1(_0016_),
    .Y(_0502_),
    .A1(net36),
    .A2(_0498_));
 sg13g2_nor2_1 _1081_ (.A(_0465_),
    .B(_0502_),
    .Y(_0503_));
 sg13g2_inv_1 _1082_ (.Y(_0504_),
    .A(net36));
 sg13g2_nor3_1 _1083_ (.A(_0504_),
    .B(net31),
    .C(_0495_),
    .Y(_0505_));
 sg13g2_nor2_1 _1084_ (.A(_0503_),
    .B(_0505_),
    .Y(_0506_));
 sg13g2_xor2_1 _1085_ (.B(_0506_),
    .A(net37),
    .X(_0507_));
 sg13g2_nand2_1 _1086_ (.Y(_0033_),
    .A(net33),
    .B(_0507_));
 sg13g2_a21o_1 _1087_ (.A2(_0468_),
    .A1(_0015_),
    .B1(_0505_),
    .X(_0508_));
 sg13g2_a22oi_1 _1088_ (.Y(_0509_),
    .B1(_0508_),
    .B2(net37),
    .A2(_0503_),
    .A1(_0015_));
 sg13g2_xnor2_1 _1089_ (.Y(_0510_),
    .A(_0361_),
    .B(_0509_));
 sg13g2_nor2_1 _1090_ (.A(_0415_),
    .B(_0510_),
    .Y(_0034_));
 sg13g2_nand2_1 _1091_ (.Y(_0511_),
    .A(_0169_),
    .B(_0172_));
 sg13g2_nand2_1 _1092_ (.Y(_0512_),
    .A(_0009_),
    .B(_0511_));
 sg13g2_or3_1 _1093_ (.A(_0160_),
    .B(_0426_),
    .C(_0511_),
    .X(_0513_));
 sg13g2_nand3_1 _1094_ (.B(_0512_),
    .C(_0513_),
    .A(net34),
    .Y(_0035_));
 sg13g2_xnor2_1 _1095_ (.Y(_0514_),
    .A(_0160_),
    .B(net46));
 sg13g2_o21ai_1 _1096_ (.B1(net33),
    .Y(_0036_),
    .A1(net30),
    .A2(_0514_));
 sg13g2_xor2_1 _1097_ (.B(_0293_),
    .A(_0161_),
    .X(_0515_));
 sg13g2_o21ai_1 _1098_ (.B1(_0456_),
    .Y(_0037_),
    .A1(net30),
    .A2(_0515_));
 sg13g2_nand3_1 _1099_ (.B(net47),
    .C(_0162_),
    .A(_0160_),
    .Y(_0516_));
 sg13g2_xor2_1 _1100_ (.B(_0516_),
    .A(net45),
    .X(_0517_));
 sg13g2_o21ai_1 _1101_ (.B1(net33),
    .Y(_0038_),
    .A1(_0428_),
    .A2(_0517_));
 sg13g2_xnor2_1 _1102_ (.Y(_0518_),
    .A(_0158_),
    .B(_0165_));
 sg13g2_o21ai_1 _1103_ (.B1(_0456_),
    .Y(_0039_),
    .A1(_0428_),
    .A2(_0518_));
 sg13g2_xor2_1 _1104_ (.B(_0417_),
    .A(net49),
    .X(_0519_));
 sg13g2_o21ai_1 _1105_ (.B1(net33),
    .Y(_0040_),
    .A1(net30),
    .A2(_0519_));
 sg13g2_nand3_1 _1106_ (.B(net48),
    .C(_0165_),
    .A(_0157_),
    .Y(_0520_));
 sg13g2_xnor2_1 _1107_ (.Y(_0521_),
    .A(_0286_),
    .B(_0520_));
 sg13g2_buf_1 _1108_ (.A(_0094_),
    .X(_0522_));
 sg13g2_o21ai_1 _1109_ (.B1(net32),
    .Y(_0041_),
    .A1(net30),
    .A2(_0521_));
 sg13g2_xnor2_1 _1110_ (.Y(_0523_),
    .A(net51),
    .B(_0418_));
 sg13g2_o21ai_1 _1111_ (.B1(net32),
    .Y(_0042_),
    .A1(net30),
    .A2(_0523_));
 sg13g2_inv_1 _1112_ (.Y(_0524_),
    .A(net44));
 sg13g2_nand2_1 _1113_ (.Y(_0525_),
    .A(net51),
    .B(_0418_));
 sg13g2_xnor2_1 _1114_ (.Y(_0526_),
    .A(_0524_),
    .B(_0525_));
 sg13g2_o21ai_1 _1115_ (.B1(_0522_),
    .Y(_0043_),
    .A1(net30),
    .A2(_0526_));
 sg13g2_nand3_1 _1116_ (.B(net44),
    .C(_0418_),
    .A(net51),
    .Y(_0527_));
 sg13g2_xor2_1 _1117_ (.B(_0527_),
    .A(net43),
    .X(_0528_));
 sg13g2_o21ai_1 _1118_ (.B1(_0522_),
    .Y(_0044_),
    .A1(net30),
    .A2(_0528_));
 sg13g2_nor2b_1 _1119_ (.A(_0111_),
    .B_N(_0434_),
    .Y(_0529_));
 sg13g2_mux2_1 _1120_ (.A0(_0010_),
    .A1(_0529_),
    .S(_0437_),
    .X(_0530_));
 sg13g2_nand2_1 _1121_ (.Y(_0531_),
    .A(_0426_),
    .B(_0530_));
 sg13g2_nand3_1 _1122_ (.B(net43),
    .C(_0424_),
    .A(net44),
    .Y(_0532_));
 sg13g2_buf_2 _1123_ (.A(_0532_),
    .X(_0533_));
 sg13g2_nand2_1 _1124_ (.Y(_0534_),
    .A(_0111_),
    .B(_0533_));
 sg13g2_nand3_1 _1125_ (.B(_0531_),
    .C(_0534_),
    .A(net34),
    .Y(_0045_));
 sg13g2_nor2b_1 _1126_ (.A(_0434_),
    .B_N(_0437_),
    .Y(_0535_));
 sg13g2_or3_1 _1127_ (.A(_0261_),
    .B(_0533_),
    .C(_0535_),
    .X(_0536_));
 sg13g2_o21ai_1 _1128_ (.B1(_0426_),
    .Y(_0537_),
    .A1(_0111_),
    .A2(_0535_));
 sg13g2_nand2_1 _1129_ (.Y(_0538_),
    .A(net54),
    .B(_0537_));
 sg13g2_nand3_1 _1130_ (.B(_0536_),
    .C(_0538_),
    .A(net34),
    .Y(_0046_));
 sg13g2_nor2_2 _1131_ (.A(_0434_),
    .B(_0439_),
    .Y(_0539_));
 sg13g2_nor2_1 _1132_ (.A(_0266_),
    .B(_0533_),
    .Y(_0540_));
 sg13g2_xnor2_1 _1133_ (.Y(_0541_),
    .A(net52),
    .B(_0540_));
 sg13g2_o21ai_1 _1134_ (.B1(net32),
    .Y(_0047_),
    .A1(_0539_),
    .A2(_0541_));
 sg13g2_nor2_1 _1135_ (.A(_0404_),
    .B(_0533_),
    .Y(_0542_));
 sg13g2_xnor2_1 _1136_ (.Y(_0543_),
    .A(net55),
    .B(_0542_));
 sg13g2_o21ai_1 _1137_ (.B1(net32),
    .Y(_0048_),
    .A1(_0539_),
    .A2(_0543_));
 sg13g2_nor2_1 _1138_ (.A(_0533_),
    .B(_0431_),
    .Y(_0544_));
 sg13g2_xnor2_1 _1139_ (.Y(_0545_),
    .A(_0100_),
    .B(_0544_));
 sg13g2_o21ai_1 _1140_ (.B1(net32),
    .Y(_0049_),
    .A1(_0539_),
    .A2(_0545_));
 sg13g2_and2_1 _1141_ (.A(_0426_),
    .B(_0435_),
    .X(_0546_));
 sg13g2_xnor2_1 _1142_ (.Y(_0547_),
    .A(net53),
    .B(_0546_));
 sg13g2_o21ai_1 _1143_ (.B1(net32),
    .Y(_0050_),
    .A1(_0539_),
    .A2(_0547_));
 sg13g2_nand2_1 _1144_ (.Y(_0548_),
    .A(_0098_),
    .B(_0435_));
 sg13g2_nor2_1 _1145_ (.A(_0533_),
    .B(_0548_),
    .Y(_0549_));
 sg13g2_xnor2_1 _1146_ (.Y(_0550_),
    .A(_0110_),
    .B(_0549_));
 sg13g2_o21ai_1 _1147_ (.B1(net32),
    .Y(_0051_),
    .A1(_0539_),
    .A2(_0550_));
 sg13g2_nand2_1 _1148_ (.Y(_0551_),
    .A(_0110_),
    .B(_0549_));
 sg13g2_xor2_1 _1149_ (.B(_0551_),
    .A(\vga.count_v[7] ),
    .X(_0552_));
 sg13g2_o21ai_1 _1150_ (.B1(net32),
    .Y(_0052_),
    .A1(_0539_),
    .A2(_0552_));
 sg13g2_nand3_1 _1151_ (.B(_0110_),
    .C(_0549_),
    .A(\vga.count_v[7] ),
    .Y(_0553_));
 sg13g2_xor2_1 _1152_ (.B(_0553_),
    .A(\vga.count_v[8] ),
    .X(_0554_));
 sg13g2_o21ai_1 _1153_ (.B1(net34),
    .Y(_0053_),
    .A1(_0539_),
    .A2(_0554_));
 sg13g2_nor2_1 _1154_ (.A(_0405_),
    .B(_0548_),
    .Y(_0555_));
 sg13g2_xor2_1 _1155_ (.B(_0555_),
    .A(_0006_),
    .X(_0556_));
 sg13g2_nor3_1 _1156_ (.A(_0533_),
    .B(_0535_),
    .C(_0556_),
    .Y(_0557_));
 sg13g2_a21oi_1 _1157_ (.A1(\vga.count_v[9] ),
    .A2(_0533_),
    .Y(_0558_),
    .B1(_0557_));
 sg13g2_nor2_1 _1158_ (.A(_0415_),
    .B(_0558_),
    .Y(_0054_));
 sg13g2_o21ai_1 _1159_ (.B1(net34),
    .Y(_0086_),
    .A1(_0093_),
    .A2(net3));
 sg13g2_nor2_1 _1160_ (.A(_0415_),
    .B(_0093_),
    .Y(_0087_));
 sg13g2_and2_1 _1161_ (.A(_0430_),
    .B(net4),
    .X(_0090_));
 sg13g2_and2_1 _1162_ (.A(_0430_),
    .B(net5),
    .X(_0091_));
 sg13g2_nand2_1 _1163_ (.Y(_0559_),
    .A(_0407_),
    .B(_0095_));
 sg13g2_nor4_1 _1164_ (.A(_0008_),
    .B(_0102_),
    .C(_0405_),
    .D(_0559_),
    .Y(_0560_));
 sg13g2_nand2b_1 _1165_ (.Y(_0561_),
    .B(_0560_),
    .A_N(_0438_));
 sg13g2_nand2_1 _1166_ (.Y(_0562_),
    .A(\vga.vs_out ),
    .B(_0438_));
 sg13g2_a21oi_1 _1167_ (.A1(_0561_),
    .A2(_0562_),
    .Y(_0092_),
    .B1(_0415_));
 sg13g2_buf_1 _1168_ (.A(ui_in[7]),
    .X(_0563_));
 sg13g2_inv_1 _1169_ (.Y(net13),
    .A(_0563_));
 sg13g2_nor2b_1 _1170_ (.A(_0563_),
    .B_N(g0),
    .Y(_0564_));
 sg13g2_a21o_1 _1171_ (.A2(b0),
    .A1(_0563_),
    .B1(_0564_),
    .X(net22));
 sg13g2_a21o_1 _1172_ (.A2(\vga.vs ),
    .A1(_0563_),
    .B1(_0564_),
    .X(net23));
 sg13g2_nor2b_1 _1173_ (.A(_0563_),
    .B_N(b0),
    .Y(_0565_));
 sg13g2_a21o_1 _1174_ (.A2(g0),
    .A1(_0563_),
    .B1(_0565_),
    .X(net25));
 sg13g2_a21o_1 _1175_ (.A2(hs),
    .A1(_0563_),
    .B1(_0565_),
    .X(net27));
 sg13g2_dfrbp_1 _1176_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net58),
    .D(_0001_),
    .Q_N(_0621_),
    .Q(_0003_));
 sg13g2_dfrbp_1 _1177_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net59),
    .D(_0000_),
    .Q_N(_0620_),
    .Q(_0002_));
 sg13g2_dfrbp_1 _1178_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net60),
    .D(_0021_),
    .Q_N(_0619_),
    .Q(_0004_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _1176__58 (.L_HI(net58));
 sg13g2_buf_1 _1181_ (.A(net13),
    .X(net6));
 sg13g2_buf_1 _1182_ (.A(net13),
    .X(net7));
 sg13g2_buf_1 _1183_ (.A(net13),
    .X(net8));
 sg13g2_buf_1 _1184_ (.A(net13),
    .X(net9));
 sg13g2_buf_1 _1185_ (.A(net13),
    .X(net10));
 sg13g2_buf_1 _1186_ (.A(net13),
    .X(net11));
 sg13g2_buf_1 _1187_ (.A(net13),
    .X(net12));
 sg13g2_buf_1 _1188_ (.A(g0),
    .X(net14));
 sg13g2_buf_1 _1189_ (.A(g0),
    .X(net15));
 sg13g2_buf_1 _1190_ (.A(g0),
    .X(net16));
 sg13g2_buf_1 _1191_ (.A(g0),
    .X(net17));
 sg13g2_buf_1 _1192_ (.A(hs),
    .X(net18));
 sg13g2_buf_1 _1193_ (.A(\vga.vs ),
    .X(net19));
 sg13g2_buf_1 _1194_ (.A(net56),
    .X(uio_out[6]));
 sg13g2_buf_1 _1195_ (.A(net57),
    .X(uio_out[7]));
 sg13g2_buf_1 _1196_ (.A(g0),
    .X(net20));
 sg13g2_buf_1 _1197_ (.A(g0),
    .X(net21));
 sg13g2_buf_1 _1198_ (.A(net25),
    .X(net24));
 sg13g2_buf_1 _1199_ (.A(b0),
    .X(net26));
 sg13g2_dfrbp_1 \vga.blank_h$_SDFFE_PN1P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net61),
    .D(_0022_),
    .Q_N(_0618_),
    .Q(\vga.blank_h ));
 sg13g2_dfrbp_1 \vga.blank_v$_SDFFE_PN1P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net62),
    .D(_0023_),
    .Q_N(_0617_),
    .Q(\vga.blank_v ));
 sg13g2_dfrbp_1 \vga.blu$_SDFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net63),
    .D(_0024_),
    .Q_N(_0616_),
    .Q(b0));
 sg13g2_dfrbp_1 \vga.car_pos_h[0]$_SDFFE_PN1P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net64),
    .D(_0025_),
    .Q_N(_0019_),
    .Q(\vga.car_pos_h[0] ));
 sg13g2_dfrbp_1 \vga.car_pos_h[1]$_SDFFE_PN1P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net65),
    .D(_0026_),
    .Q_N(_0615_),
    .Q(\vga.car_pos_h[1] ));
 sg13g2_dfrbp_1 \vga.car_pos_h[2]$_SDFFE_PN1P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net66),
    .D(_0027_),
    .Q_N(_0018_),
    .Q(\vga.car_pos_h[2] ));
 sg13g2_dfrbp_1 \vga.car_pos_h[3]$_SDFFE_PN1P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net67),
    .D(_0028_),
    .Q_N(_0614_),
    .Q(\vga.car_pos_h[3] ));
 sg13g2_dfrbp_1 \vga.car_pos_h[4]$_SDFFE_PN1P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net68),
    .D(_0029_),
    .Q_N(_0613_),
    .Q(\vga.car_pos_h[4] ));
 sg13g2_dfrbp_1 \vga.car_pos_h[5]$_SDFFE_PN1P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net69),
    .D(_0030_),
    .Q_N(_0612_),
    .Q(\vga.car_pos_h[5] ));
 sg13g2_dfrbp_1 \vga.car_pos_h[6]$_SDFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net70),
    .D(_0031_),
    .Q_N(_0017_),
    .Q(\vga.car_pos_h[6] ));
 sg13g2_dfrbp_1 \vga.car_pos_h[7]$_SDFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net71),
    .D(_0032_),
    .Q_N(_0016_),
    .Q(\vga.car_pos_h[7] ));
 sg13g2_dfrbp_1 \vga.car_pos_h[8]$_SDFFE_PN1P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net72),
    .D(_0033_),
    .Q_N(_0015_),
    .Q(\vga.car_pos_h[8] ));
 sg13g2_dfrbp_1 \vga.car_pos_h[9]$_SDFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net73),
    .D(_0034_),
    .Q_N(_0011_),
    .Q(\vga.car_pos_h[9] ));
 sg13g2_dfrbp_1 \vga.count_h[0]$_SDFF_PN1_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net74),
    .D(_0035_),
    .Q_N(_0009_),
    .Q(\vga.count_h[0] ));
 sg13g2_dfrbp_1 \vga.count_h[1]$_SDFF_PN1_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net75),
    .D(_0036_),
    .Q_N(_0611_),
    .Q(\vga.count_h[1] ));
 sg13g2_dfrbp_1 \vga.count_h[2]$_SDFF_PN1_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net76),
    .D(_0037_),
    .Q_N(_0610_),
    .Q(\vga.count_h[2] ));
 sg13g2_dfrbp_1 \vga.count_h[3]$_SDFF_PN1_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net77),
    .D(_0038_),
    .Q_N(_0609_),
    .Q(\vga.count_h[3] ));
 sg13g2_dfrbp_1 \vga.count_h[4]$_SDFF_PN1_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net78),
    .D(_0039_),
    .Q_N(_0608_),
    .Q(\vga.count_h[4] ));
 sg13g2_dfrbp_1 \vga.count_h[5]$_SDFF_PN1_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net79),
    .D(_0040_),
    .Q_N(_0005_),
    .Q(\vga.count_h[5] ));
 sg13g2_dfrbp_1 \vga.count_h[6]$_SDFF_PN1_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net80),
    .D(_0041_),
    .Q_N(_0014_),
    .Q(\vga.count_h[6] ));
 sg13g2_dfrbp_1 \vga.count_h[7]$_SDFF_PN1_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net81),
    .D(_0042_),
    .Q_N(_0012_),
    .Q(\vga.count_h[7] ));
 sg13g2_dfrbp_1 \vga.count_h[8]$_SDFF_PN1_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net82),
    .D(_0043_),
    .Q_N(_0013_),
    .Q(\vga.count_h[8] ));
 sg13g2_dfrbp_1 \vga.count_h[9]$_SDFF_PN1_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net83),
    .D(_0044_),
    .Q_N(_0007_),
    .Q(\vga.count_h[9] ));
 sg13g2_dfrbp_1 \vga.count_v[0]$_SDFFE_PN1N_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net84),
    .D(_0045_),
    .Q_N(_0010_),
    .Q(\vga.count_v[0] ));
 sg13g2_dfrbp_1 \vga.count_v[1]$_SDFFE_PN1N_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net85),
    .D(_0046_),
    .Q_N(_0008_),
    .Q(\vga.count_v[1] ));
 sg13g2_dfrbp_1 \vga.count_v[2]$_SDFFE_PN1N_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net86),
    .D(_0047_),
    .Q_N(_0607_),
    .Q(\vga.count_v[2] ));
 sg13g2_dfrbp_1 \vga.count_v[3]$_SDFFE_PN1N_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net87),
    .D(_0048_),
    .Q_N(_0606_),
    .Q(\vga.count_v[3] ));
 sg13g2_dfrbp_1 \vga.count_v[4]$_SDFFE_PN1N_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net88),
    .D(_0049_),
    .Q_N(_0605_),
    .Q(\vga.count_v[4] ));
 sg13g2_dfrbp_1 \vga.count_v[5]$_SDFFE_PN1N_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net89),
    .D(_0050_),
    .Q_N(_0604_),
    .Q(\vga.count_v[5] ));
 sg13g2_dfrbp_1 \vga.count_v[6]$_SDFFE_PN1N_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net90),
    .D(_0051_),
    .Q_N(_0603_),
    .Q(\vga.count_v[6] ));
 sg13g2_dfrbp_1 \vga.count_v[7]$_SDFFE_PN1N_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net91),
    .D(_0052_),
    .Q_N(_0602_),
    .Q(\vga.count_v[7] ));
 sg13g2_dfrbp_1 \vga.count_v[8]$_SDFFE_PN1N_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net92),
    .D(_0053_),
    .Q_N(_0601_),
    .Q(\vga.count_v[8] ));
 sg13g2_dfrbp_1 \vga.count_v[9]$_SDFFE_PN0N_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net93),
    .D(_0054_),
    .Q_N(_0006_),
    .Q(\vga.count_v[9] ));
 sg13g2_dfrbp_1 \vga.hs_out$_SDFF_PP0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net94),
    .D(_0055_),
    .Q_N(hs),
    .Q(\vga.hs_out ));
 sg13g2_dfrbp_1 \vga.interval_counter[0]$_SDFF_PP0_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net95),
    .D(_0056_),
    .Q_N(_0020_),
    .Q(\vga.interval_counter[0] ));
 sg13g2_dfrbp_1 \vga.interval_counter[10]$_SDFF_PP0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net96),
    .D(_0057_),
    .Q_N(_0600_),
    .Q(\vga.interval_counter[10] ));
 sg13g2_dfrbp_1 \vga.interval_counter[11]$_SDFF_PP0_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net97),
    .D(_0058_),
    .Q_N(_0599_),
    .Q(\vga.interval_counter[11] ));
 sg13g2_dfrbp_1 \vga.interval_counter[12]$_SDFF_PP0_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net98),
    .D(_0059_),
    .Q_N(_0598_),
    .Q(\vga.interval_counter[12] ));
 sg13g2_dfrbp_1 \vga.interval_counter[13]$_SDFF_PP0_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net99),
    .D(_0060_),
    .Q_N(_0597_),
    .Q(\vga.interval_counter[13] ));
 sg13g2_dfrbp_1 \vga.interval_counter[14]$_SDFF_PP0_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net100),
    .D(_0061_),
    .Q_N(_0596_),
    .Q(\vga.interval_counter[14] ));
 sg13g2_dfrbp_1 \vga.interval_counter[15]$_SDFF_PP0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net101),
    .D(_0062_),
    .Q_N(_0595_),
    .Q(\vga.interval_counter[15] ));
 sg13g2_dfrbp_1 \vga.interval_counter[16]$_SDFF_PP0_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net102),
    .D(_0063_),
    .Q_N(_0594_),
    .Q(\vga.interval_counter[16] ));
 sg13g2_dfrbp_1 \vga.interval_counter[17]$_SDFF_PP0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net103),
    .D(_0064_),
    .Q_N(_0593_),
    .Q(\vga.interval_counter[17] ));
 sg13g2_dfrbp_1 \vga.interval_counter[18]$_SDFF_PP0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net104),
    .D(_0065_),
    .Q_N(_0592_),
    .Q(\vga.interval_counter[18] ));
 sg13g2_dfrbp_1 \vga.interval_counter[19]$_SDFF_PP0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net105),
    .D(_0066_),
    .Q_N(_0591_),
    .Q(\vga.interval_counter[19] ));
 sg13g2_dfrbp_1 \vga.interval_counter[1]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net106),
    .D(_0067_),
    .Q_N(_0590_),
    .Q(\vga.interval_counter[1] ));
 sg13g2_dfrbp_1 \vga.interval_counter[20]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net107),
    .D(_0068_),
    .Q_N(_0589_),
    .Q(\vga.interval_counter[20] ));
 sg13g2_dfrbp_1 \vga.interval_counter[21]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net108),
    .D(_0069_),
    .Q_N(_0588_),
    .Q(\vga.interval_counter[21] ));
 sg13g2_dfrbp_1 \vga.interval_counter[22]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net109),
    .D(_0070_),
    .Q_N(_0587_),
    .Q(\vga.interval_counter[22] ));
 sg13g2_dfrbp_1 \vga.interval_counter[23]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net110),
    .D(_0071_),
    .Q_N(_0586_),
    .Q(\vga.interval_counter[23] ));
 sg13g2_dfrbp_1 \vga.interval_counter[24]$_SDFF_PP0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net111),
    .D(_0072_),
    .Q_N(_0585_),
    .Q(\vga.interval_counter[24] ));
 sg13g2_dfrbp_1 \vga.interval_counter[2]$_SDFF_PP0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net112),
    .D(_0073_),
    .Q_N(_0584_),
    .Q(\vga.interval_counter[2] ));
 sg13g2_dfrbp_1 \vga.interval_counter[3]$_SDFF_PP0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net113),
    .D(_0074_),
    .Q_N(_0583_),
    .Q(\vga.interval_counter[3] ));
 sg13g2_dfrbp_1 \vga.interval_counter[4]$_SDFF_PP0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net114),
    .D(_0075_),
    .Q_N(_0582_),
    .Q(\vga.interval_counter[4] ));
 sg13g2_dfrbp_1 \vga.interval_counter[5]$_SDFF_PP0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net115),
    .D(_0076_),
    .Q_N(_0581_),
    .Q(\vga.interval_counter[5] ));
 sg13g2_dfrbp_1 \vga.interval_counter[6]$_SDFF_PP0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net116),
    .D(_0077_),
    .Q_N(_0580_),
    .Q(\vga.interval_counter[6] ));
 sg13g2_dfrbp_1 \vga.interval_counter[7]$_SDFF_PP0_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net117),
    .D(_0078_),
    .Q_N(_0579_),
    .Q(\vga.interval_counter[7] ));
 sg13g2_dfrbp_1 \vga.interval_counter[8]$_SDFF_PP0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net118),
    .D(_0079_),
    .Q_N(_0578_),
    .Q(\vga.interval_counter[8] ));
 sg13g2_dfrbp_1 \vga.interval_counter[9]$_SDFF_PP0_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net119),
    .D(_0080_),
    .Q_N(_0577_),
    .Q(\vga.interval_counter[9] ));
 sg13g2_dfrbp_1 \vga.left_1d$_DFFE_PN_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net120),
    .D(_0081_),
    .Q_N(_0576_),
    .Q(\vga.left_1d ));
 sg13g2_dfrbp_1 \vga.left_pressed$_SDFF_PP0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net121),
    .D(_0082_),
    .Q_N(_0575_),
    .Q(\vga.left_pressed ));
 sg13g2_dfrbp_1 \vga.red$_SDFF_PP0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net122),
    .D(_0083_),
    .Q_N(_0574_),
    .Q(g0));
 sg13g2_dfrbp_1 \vga.right_1d$_DFFE_PN_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net123),
    .D(_0084_),
    .Q_N(_0573_),
    .Q(\vga.right_1d ));
 sg13g2_dfrbp_1 \vga.right_pressed$_SDFF_PP0_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net124),
    .D(_0085_),
    .Q_N(_0572_),
    .Q(\vga.right_pressed ));
 sg13g2_dfrbp_1 \vga.score[1]$_SDFFE_PN1P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net125),
    .D(_0086_),
    .Q_N(_0571_),
    .Q(\vga.score[0] ));
 sg13g2_dfrbp_1 \vga.score_ten_enable$_SDFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net126),
    .D(_0087_),
    .Q_N(_0570_),
    .Q(\vga.score_ten_enable ));
 sg13g2_dfrbp_1 \vga.score_unit_pixels[1]$_SDFFCE_PP1P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net127),
    .D(_0088_),
    .Q_N(_0569_),
    .Q(\vga.score_unit_pixels[1] ));
 sg13g2_dfrbp_1 \vga.score_unit_pixels[2]$_SDFFCE_PP1P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net128),
    .D(_0089_),
    .Q_N(_0568_),
    .Q(\vga.score_unit_pixels[2] ));
 sg13g2_dfrbp_1 \vga.speed_lsb_1d$_SDFF_PN0_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net129),
    .D(_0090_),
    .Q_N(_0567_),
    .Q(\vga.speed_lsb_1d ));
 sg13g2_dfrbp_1 \vga.speed_msb_1d$_SDFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net130),
    .D(_0091_),
    .Q_N(_0566_),
    .Q(\vga.speed_msb_1d ));
 sg13g2_dfrbp_1 \vga.vs_out$_SDFFE_PN0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net131),
    .D(_0092_),
    .Q_N(\vga.vs ),
    .Q(\vga.vs_out ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[5]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[6]),
    .X(net5));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_oe[0]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_oe[1]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_oe[2]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_oe[3]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_oe[4]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_oe[5]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_oe[6]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_oe[7]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[0]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_out[1]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_out[2]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_out[3]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_out[4]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uio_out[5]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[0]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[1]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[2]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[3]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[4]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[5]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uo_out[6]));
 sg13g2_buf_1 output27 (.A(net27),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout28 (.A(_0231_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0206_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0428_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0457_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0522_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0456_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0430_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0390_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0351_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0350_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0346_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0330_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0328_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0310_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0306_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0277_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0274_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0163_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0162_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_0161_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_0158_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_0157_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0156_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0155_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0099_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0098_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_0096_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0095_),
    .X(net55));
 sg13g2_tielo _1194__56 (.L_LO(net56));
 sg13g2_tielo _1195__57 (.L_LO(net57));
 sg13g2_tiehi _1177__59 (.L_HI(net59));
 sg13g2_tiehi _1178__60 (.L_HI(net60));
 sg13g2_tiehi \vga.blank_h$_SDFFE_PN1P__61  (.L_HI(net61));
 sg13g2_tiehi \vga.blank_v$_SDFFE_PN1P__62  (.L_HI(net62));
 sg13g2_tiehi \vga.blu$_SDFF_PN0__63  (.L_HI(net63));
 sg13g2_tiehi \vga.car_pos_h[0]$_SDFFE_PN1P__64  (.L_HI(net64));
 sg13g2_tiehi \vga.car_pos_h[1]$_SDFFE_PN1P__65  (.L_HI(net65));
 sg13g2_tiehi \vga.car_pos_h[2]$_SDFFE_PN1P__66  (.L_HI(net66));
 sg13g2_tiehi \vga.car_pos_h[3]$_SDFFE_PN1P__67  (.L_HI(net67));
 sg13g2_tiehi \vga.car_pos_h[4]$_SDFFE_PN1P__68  (.L_HI(net68));
 sg13g2_tiehi \vga.car_pos_h[5]$_SDFFE_PN1P__69  (.L_HI(net69));
 sg13g2_tiehi \vga.car_pos_h[6]$_SDFFE_PN0P__70  (.L_HI(net70));
 sg13g2_tiehi \vga.car_pos_h[7]$_SDFFE_PN0P__71  (.L_HI(net71));
 sg13g2_tiehi \vga.car_pos_h[8]$_SDFFE_PN1P__72  (.L_HI(net72));
 sg13g2_tiehi \vga.car_pos_h[9]$_SDFFE_PN0P__73  (.L_HI(net73));
 sg13g2_tiehi \vga.count_h[0]$_SDFF_PN1__74  (.L_HI(net74));
 sg13g2_tiehi \vga.count_h[1]$_SDFF_PN1__75  (.L_HI(net75));
 sg13g2_tiehi \vga.count_h[2]$_SDFF_PN1__76  (.L_HI(net76));
 sg13g2_tiehi \vga.count_h[3]$_SDFF_PN1__77  (.L_HI(net77));
 sg13g2_tiehi \vga.count_h[4]$_SDFF_PN1__78  (.L_HI(net78));
 sg13g2_tiehi \vga.count_h[5]$_SDFF_PN1__79  (.L_HI(net79));
 sg13g2_tiehi \vga.count_h[6]$_SDFF_PN1__80  (.L_HI(net80));
 sg13g2_tiehi \vga.count_h[7]$_SDFF_PN1__81  (.L_HI(net81));
 sg13g2_tiehi \vga.count_h[8]$_SDFF_PN1__82  (.L_HI(net82));
 sg13g2_tiehi \vga.count_h[9]$_SDFF_PN1__83  (.L_HI(net83));
 sg13g2_tiehi \vga.count_v[0]$_SDFFE_PN1N__84  (.L_HI(net84));
 sg13g2_tiehi \vga.count_v[1]$_SDFFE_PN1N__85  (.L_HI(net85));
 sg13g2_tiehi \vga.count_v[2]$_SDFFE_PN1N__86  (.L_HI(net86));
 sg13g2_tiehi \vga.count_v[3]$_SDFFE_PN1N__87  (.L_HI(net87));
 sg13g2_tiehi \vga.count_v[4]$_SDFFE_PN1N__88  (.L_HI(net88));
 sg13g2_tiehi \vga.count_v[5]$_SDFFE_PN1N__89  (.L_HI(net89));
 sg13g2_tiehi \vga.count_v[6]$_SDFFE_PN1N__90  (.L_HI(net90));
 sg13g2_tiehi \vga.count_v[7]$_SDFFE_PN1N__91  (.L_HI(net91));
 sg13g2_tiehi \vga.count_v[8]$_SDFFE_PN1N__92  (.L_HI(net92));
 sg13g2_tiehi \vga.count_v[9]$_SDFFE_PN0N__93  (.L_HI(net93));
 sg13g2_tiehi \vga.hs_out$_SDFF_PP0__94  (.L_HI(net94));
 sg13g2_tiehi \vga.interval_counter[0]$_SDFF_PP0__95  (.L_HI(net95));
 sg13g2_tiehi \vga.interval_counter[10]$_SDFF_PP0__96  (.L_HI(net96));
 sg13g2_tiehi \vga.interval_counter[11]$_SDFF_PP0__97  (.L_HI(net97));
 sg13g2_tiehi \vga.interval_counter[12]$_SDFF_PP0__98  (.L_HI(net98));
 sg13g2_tiehi \vga.interval_counter[13]$_SDFF_PP0__99  (.L_HI(net99));
 sg13g2_tiehi \vga.interval_counter[14]$_SDFF_PP0__100  (.L_HI(net100));
 sg13g2_tiehi \vga.interval_counter[15]$_SDFF_PP0__101  (.L_HI(net101));
 sg13g2_tiehi \vga.interval_counter[16]$_SDFF_PP0__102  (.L_HI(net102));
 sg13g2_tiehi \vga.interval_counter[17]$_SDFF_PP0__103  (.L_HI(net103));
 sg13g2_tiehi \vga.interval_counter[18]$_SDFF_PP0__104  (.L_HI(net104));
 sg13g2_tiehi \vga.interval_counter[19]$_SDFF_PP0__105  (.L_HI(net105));
 sg13g2_tiehi \vga.interval_counter[1]$_SDFF_PP0__106  (.L_HI(net106));
 sg13g2_tiehi \vga.interval_counter[20]$_SDFF_PP0__107  (.L_HI(net107));
 sg13g2_tiehi \vga.interval_counter[21]$_SDFF_PP0__108  (.L_HI(net108));
 sg13g2_tiehi \vga.interval_counter[22]$_SDFF_PP0__109  (.L_HI(net109));
 sg13g2_tiehi \vga.interval_counter[23]$_SDFF_PP0__110  (.L_HI(net110));
 sg13g2_tiehi \vga.interval_counter[24]$_SDFF_PP0__111  (.L_HI(net111));
 sg13g2_tiehi \vga.interval_counter[2]$_SDFF_PP0__112  (.L_HI(net112));
 sg13g2_tiehi \vga.interval_counter[3]$_SDFF_PP0__113  (.L_HI(net113));
 sg13g2_tiehi \vga.interval_counter[4]$_SDFF_PP0__114  (.L_HI(net114));
 sg13g2_tiehi \vga.interval_counter[5]$_SDFF_PP0__115  (.L_HI(net115));
 sg13g2_tiehi \vga.interval_counter[6]$_SDFF_PP0__116  (.L_HI(net116));
 sg13g2_tiehi \vga.interval_counter[7]$_SDFF_PP0__117  (.L_HI(net117));
 sg13g2_tiehi \vga.interval_counter[8]$_SDFF_PP0__118  (.L_HI(net118));
 sg13g2_tiehi \vga.interval_counter[9]$_SDFF_PP0__119  (.L_HI(net119));
 sg13g2_tiehi \vga.left_1d$_DFFE_PN__120  (.L_HI(net120));
 sg13g2_tiehi \vga.left_pressed$_SDFF_PP0__121  (.L_HI(net121));
 sg13g2_tiehi \vga.red$_SDFF_PP0__122  (.L_HI(net122));
 sg13g2_tiehi \vga.right_1d$_DFFE_PN__123  (.L_HI(net123));
 sg13g2_tiehi \vga.right_pressed$_SDFF_PP0__124  (.L_HI(net124));
 sg13g2_tiehi \vga.score[1]$_SDFFE_PN1P__125  (.L_HI(net125));
 sg13g2_tiehi \vga.score_ten_enable$_SDFF_PN0__126  (.L_HI(net126));
 sg13g2_tiehi \vga.score_unit_pixels[1]$_SDFFCE_PP1P__127  (.L_HI(net127));
 sg13g2_tiehi \vga.score_unit_pixels[2]$_SDFFCE_PP1P__128  (.L_HI(net128));
 sg13g2_tiehi \vga.speed_lsb_1d$_SDFF_PN0__129  (.L_HI(net129));
 sg13g2_tiehi \vga.speed_msb_1d$_SDFF_PN0__130  (.L_HI(net130));
 sg13g2_tiehi \vga.vs_out$_SDFFE_PN0P__131  (.L_HI(net131));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_15_0_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_2 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_fill_2 FILLER_4_427 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_fill_2 FILLER_5_427 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_fill_2 FILLER_7_427 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_fill_2 FILLER_8_427 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_fill_2 FILLER_9_427 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_fill_2 FILLER_10_427 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_fill_2 FILLER_11_427 ();
 sg13g2_fill_1 FILLER_11_429 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_fill_2 FILLER_12_427 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_fill_2 FILLER_13_427 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_fill_2 FILLER_14_427 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_fill_2 FILLER_15_427 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_4 FILLER_16_259 ();
 sg13g2_fill_1 FILLER_16_263 ();
 sg13g2_decap_8 FILLER_16_268 ();
 sg13g2_decap_8 FILLER_16_275 ();
 sg13g2_decap_8 FILLER_16_282 ();
 sg13g2_decap_8 FILLER_16_289 ();
 sg13g2_decap_8 FILLER_16_296 ();
 sg13g2_decap_8 FILLER_16_303 ();
 sg13g2_decap_8 FILLER_16_310 ();
 sg13g2_decap_8 FILLER_16_317 ();
 sg13g2_decap_8 FILLER_16_324 ();
 sg13g2_decap_8 FILLER_16_331 ();
 sg13g2_decap_8 FILLER_16_338 ();
 sg13g2_decap_8 FILLER_16_345 ();
 sg13g2_decap_8 FILLER_16_352 ();
 sg13g2_decap_8 FILLER_16_359 ();
 sg13g2_decap_8 FILLER_16_366 ();
 sg13g2_decap_8 FILLER_16_373 ();
 sg13g2_decap_8 FILLER_16_380 ();
 sg13g2_decap_8 FILLER_16_387 ();
 sg13g2_decap_8 FILLER_16_394 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_decap_8 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_16_415 ();
 sg13g2_decap_8 FILLER_16_422 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_4 FILLER_17_161 ();
 sg13g2_fill_2 FILLER_17_165 ();
 sg13g2_decap_8 FILLER_17_171 ();
 sg13g2_decap_4 FILLER_17_178 ();
 sg13g2_fill_2 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_188 ();
 sg13g2_fill_1 FILLER_17_195 ();
 sg13g2_decap_8 FILLER_17_200 ();
 sg13g2_decap_8 FILLER_17_211 ();
 sg13g2_decap_4 FILLER_17_218 ();
 sg13g2_fill_1 FILLER_17_222 ();
 sg13g2_decap_4 FILLER_17_249 ();
 sg13g2_decap_8 FILLER_17_283 ();
 sg13g2_decap_8 FILLER_17_290 ();
 sg13g2_decap_8 FILLER_17_297 ();
 sg13g2_decap_8 FILLER_17_304 ();
 sg13g2_fill_2 FILLER_17_311 ();
 sg13g2_decap_8 FILLER_17_317 ();
 sg13g2_decap_8 FILLER_17_324 ();
 sg13g2_decap_8 FILLER_17_331 ();
 sg13g2_decap_8 FILLER_17_338 ();
 sg13g2_decap_8 FILLER_17_345 ();
 sg13g2_decap_8 FILLER_17_352 ();
 sg13g2_decap_8 FILLER_17_359 ();
 sg13g2_fill_2 FILLER_17_366 ();
 sg13g2_decap_8 FILLER_17_372 ();
 sg13g2_decap_8 FILLER_17_379 ();
 sg13g2_decap_8 FILLER_17_386 ();
 sg13g2_decap_8 FILLER_17_393 ();
 sg13g2_decap_8 FILLER_17_400 ();
 sg13g2_decap_8 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_17_414 ();
 sg13g2_decap_8 FILLER_17_421 ();
 sg13g2_fill_2 FILLER_17_428 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_fill_1 FILLER_18_147 ();
 sg13g2_fill_2 FILLER_18_186 ();
 sg13g2_fill_1 FILLER_18_218 ();
 sg13g2_fill_2 FILLER_18_228 ();
 sg13g2_fill_1 FILLER_18_230 ();
 sg13g2_fill_2 FILLER_18_235 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_fill_1 FILLER_18_252 ();
 sg13g2_decap_4 FILLER_18_270 ();
 sg13g2_decap_8 FILLER_18_278 ();
 sg13g2_decap_8 FILLER_18_285 ();
 sg13g2_fill_2 FILLER_18_304 ();
 sg13g2_decap_8 FILLER_18_332 ();
 sg13g2_decap_8 FILLER_18_339 ();
 sg13g2_decap_8 FILLER_18_346 ();
 sg13g2_decap_8 FILLER_18_353 ();
 sg13g2_fill_1 FILLER_18_360 ();
 sg13g2_decap_8 FILLER_18_387 ();
 sg13g2_decap_8 FILLER_18_394 ();
 sg13g2_decap_8 FILLER_18_401 ();
 sg13g2_fill_2 FILLER_18_408 ();
 sg13g2_fill_1 FILLER_18_410 ();
 sg13g2_decap_8 FILLER_18_415 ();
 sg13g2_decap_8 FILLER_18_422 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_137 ();
 sg13g2_decap_8 FILLER_19_144 ();
 sg13g2_decap_8 FILLER_19_151 ();
 sg13g2_decap_8 FILLER_19_158 ();
 sg13g2_decap_4 FILLER_19_165 ();
 sg13g2_fill_2 FILLER_19_169 ();
 sg13g2_fill_1 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_188 ();
 sg13g2_decap_4 FILLER_19_195 ();
 sg13g2_fill_1 FILLER_19_199 ();
 sg13g2_fill_2 FILLER_19_217 ();
 sg13g2_fill_1 FILLER_19_242 ();
 sg13g2_fill_1 FILLER_19_248 ();
 sg13g2_fill_1 FILLER_19_255 ();
 sg13g2_fill_1 FILLER_19_276 ();
 sg13g2_fill_1 FILLER_19_287 ();
 sg13g2_fill_2 FILLER_19_303 ();
 sg13g2_decap_4 FILLER_19_310 ();
 sg13g2_fill_2 FILLER_19_314 ();
 sg13g2_fill_1 FILLER_19_320 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_fill_2 FILLER_19_350 ();
 sg13g2_fill_1 FILLER_19_352 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_fill_1 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_fill_1 FILLER_20_156 ();
 sg13g2_fill_2 FILLER_20_218 ();
 sg13g2_fill_2 FILLER_20_225 ();
 sg13g2_fill_1 FILLER_20_227 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_fill_2 FILLER_20_245 ();
 sg13g2_fill_1 FILLER_20_247 ();
 sg13g2_decap_4 FILLER_20_253 ();
 sg13g2_fill_2 FILLER_20_261 ();
 sg13g2_fill_1 FILLER_20_268 ();
 sg13g2_fill_1 FILLER_20_288 ();
 sg13g2_fill_2 FILLER_20_307 ();
 sg13g2_fill_1 FILLER_20_309 ();
 sg13g2_decap_4 FILLER_20_336 ();
 sg13g2_fill_2 FILLER_20_340 ();
 sg13g2_fill_1 FILLER_20_372 ();
 sg13g2_fill_1 FILLER_20_381 ();
 sg13g2_fill_1 FILLER_20_388 ();
 sg13g2_fill_2 FILLER_20_395 ();
 sg13g2_fill_1 FILLER_20_397 ();
 sg13g2_decap_4 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_410 ();
 sg13g2_decap_8 FILLER_20_415 ();
 sg13g2_decap_8 FILLER_20_422 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_67 ();
 sg13g2_fill_2 FILLER_21_74 ();
 sg13g2_decap_8 FILLER_21_81 ();
 sg13g2_decap_8 FILLER_21_88 ();
 sg13g2_decap_8 FILLER_21_95 ();
 sg13g2_decap_8 FILLER_21_102 ();
 sg13g2_decap_8 FILLER_21_109 ();
 sg13g2_decap_8 FILLER_21_116 ();
 sg13g2_fill_2 FILLER_21_123 ();
 sg13g2_fill_1 FILLER_21_125 ();
 sg13g2_fill_1 FILLER_21_130 ();
 sg13g2_fill_2 FILLER_21_143 ();
 sg13g2_fill_1 FILLER_21_145 ();
 sg13g2_decap_4 FILLER_21_151 ();
 sg13g2_fill_2 FILLER_21_160 ();
 sg13g2_fill_1 FILLER_21_162 ();
 sg13g2_fill_1 FILLER_21_171 ();
 sg13g2_decap_4 FILLER_21_181 ();
 sg13g2_fill_2 FILLER_21_185 ();
 sg13g2_decap_4 FILLER_21_191 ();
 sg13g2_fill_2 FILLER_21_221 ();
 sg13g2_decap_4 FILLER_21_237 ();
 sg13g2_fill_2 FILLER_21_241 ();
 sg13g2_decap_4 FILLER_21_251 ();
 sg13g2_fill_1 FILLER_21_255 ();
 sg13g2_decap_4 FILLER_21_274 ();
 sg13g2_fill_2 FILLER_21_278 ();
 sg13g2_fill_1 FILLER_21_288 ();
 sg13g2_fill_1 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_312 ();
 sg13g2_decap_4 FILLER_21_319 ();
 sg13g2_decap_8 FILLER_21_353 ();
 sg13g2_decap_8 FILLER_21_368 ();
 sg13g2_fill_1 FILLER_21_375 ();
 sg13g2_fill_2 FILLER_21_389 ();
 sg13g2_fill_1 FILLER_21_391 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_32 ();
 sg13g2_decap_8 FILLER_22_39 ();
 sg13g2_decap_8 FILLER_22_46 ();
 sg13g2_fill_2 FILLER_22_53 ();
 sg13g2_fill_1 FILLER_22_55 ();
 sg13g2_fill_2 FILLER_22_82 ();
 sg13g2_fill_2 FILLER_22_89 ();
 sg13g2_decap_8 FILLER_22_95 ();
 sg13g2_decap_8 FILLER_22_102 ();
 sg13g2_fill_1 FILLER_22_109 ();
 sg13g2_fill_2 FILLER_22_136 ();
 sg13g2_fill_1 FILLER_22_138 ();
 sg13g2_fill_1 FILLER_22_146 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_4 FILLER_22_168 ();
 sg13g2_fill_1 FILLER_22_172 ();
 sg13g2_fill_1 FILLER_22_181 ();
 sg13g2_fill_1 FILLER_22_187 ();
 sg13g2_fill_1 FILLER_22_198 ();
 sg13g2_fill_1 FILLER_22_204 ();
 sg13g2_decap_4 FILLER_22_211 ();
 sg13g2_fill_1 FILLER_22_215 ();
 sg13g2_decap_8 FILLER_22_221 ();
 sg13g2_decap_8 FILLER_22_228 ();
 sg13g2_fill_2 FILLER_22_248 ();
 sg13g2_fill_1 FILLER_22_250 ();
 sg13g2_decap_4 FILLER_22_256 ();
 sg13g2_fill_1 FILLER_22_260 ();
 sg13g2_fill_2 FILLER_22_267 ();
 sg13g2_decap_4 FILLER_22_274 ();
 sg13g2_fill_1 FILLER_22_278 ();
 sg13g2_decap_4 FILLER_22_289 ();
 sg13g2_fill_2 FILLER_22_293 ();
 sg13g2_decap_4 FILLER_22_300 ();
 sg13g2_fill_1 FILLER_22_304 ();
 sg13g2_decap_8 FILLER_22_310 ();
 sg13g2_decap_8 FILLER_22_317 ();
 sg13g2_decap_4 FILLER_22_324 ();
 sg13g2_fill_2 FILLER_22_328 ();
 sg13g2_decap_8 FILLER_22_334 ();
 sg13g2_fill_2 FILLER_22_341 ();
 sg13g2_fill_1 FILLER_22_343 ();
 sg13g2_decap_4 FILLER_22_383 ();
 sg13g2_fill_2 FILLER_22_387 ();
 sg13g2_decap_8 FILLER_22_406 ();
 sg13g2_decap_8 FILLER_22_413 ();
 sg13g2_decap_8 FILLER_22_420 ();
 sg13g2_fill_2 FILLER_22_427 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_fill_2 FILLER_23_14 ();
 sg13g2_fill_1 FILLER_23_51 ();
 sg13g2_decap_4 FILLER_23_65 ();
 sg13g2_fill_1 FILLER_23_74 ();
 sg13g2_fill_2 FILLER_23_83 ();
 sg13g2_decap_4 FILLER_23_111 ();
 sg13g2_fill_1 FILLER_23_115 ();
 sg13g2_decap_8 FILLER_23_120 ();
 sg13g2_fill_2 FILLER_23_127 ();
 sg13g2_fill_2 FILLER_23_134 ();
 sg13g2_fill_1 FILLER_23_136 ();
 sg13g2_fill_2 FILLER_23_153 ();
 sg13g2_decap_8 FILLER_23_171 ();
 sg13g2_decap_8 FILLER_23_178 ();
 sg13g2_decap_4 FILLER_23_185 ();
 sg13g2_fill_1 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_195 ();
 sg13g2_fill_1 FILLER_23_202 ();
 sg13g2_decap_4 FILLER_23_211 ();
 sg13g2_fill_1 FILLER_23_215 ();
 sg13g2_decap_8 FILLER_23_234 ();
 sg13g2_fill_2 FILLER_23_241 ();
 sg13g2_fill_1 FILLER_23_243 ();
 sg13g2_decap_8 FILLER_23_249 ();
 sg13g2_decap_8 FILLER_23_256 ();
 sg13g2_decap_4 FILLER_23_276 ();
 sg13g2_fill_2 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_317 ();
 sg13g2_fill_2 FILLER_23_324 ();
 sg13g2_fill_1 FILLER_23_326 ();
 sg13g2_fill_2 FILLER_23_339 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_4 FILLER_23_378 ();
 sg13g2_fill_1 FILLER_23_395 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_4 ();
 sg13g2_decap_8 FILLER_24_37 ();
 sg13g2_decap_4 FILLER_24_44 ();
 sg13g2_fill_2 FILLER_24_48 ();
 sg13g2_decap_4 FILLER_24_68 ();
 sg13g2_fill_1 FILLER_24_72 ();
 sg13g2_decap_8 FILLER_24_80 ();
 sg13g2_decap_8 FILLER_24_87 ();
 sg13g2_decap_4 FILLER_24_94 ();
 sg13g2_decap_8 FILLER_24_102 ();
 sg13g2_decap_8 FILLER_24_109 ();
 sg13g2_decap_8 FILLER_24_116 ();
 sg13g2_decap_4 FILLER_24_123 ();
 sg13g2_fill_2 FILLER_24_135 ();
 sg13g2_fill_1 FILLER_24_137 ();
 sg13g2_fill_1 FILLER_24_151 ();
 sg13g2_fill_1 FILLER_24_159 ();
 sg13g2_fill_2 FILLER_24_170 ();
 sg13g2_fill_1 FILLER_24_172 ();
 sg13g2_decap_4 FILLER_24_178 ();
 sg13g2_fill_1 FILLER_24_182 ();
 sg13g2_decap_4 FILLER_24_192 ();
 sg13g2_fill_1 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_4 FILLER_24_210 ();
 sg13g2_decap_4 FILLER_24_224 ();
 sg13g2_fill_1 FILLER_24_228 ();
 sg13g2_decap_8 FILLER_24_255 ();
 sg13g2_decap_8 FILLER_24_262 ();
 sg13g2_decap_4 FILLER_24_269 ();
 sg13g2_decap_4 FILLER_24_283 ();
 sg13g2_fill_2 FILLER_24_287 ();
 sg13g2_decap_4 FILLER_24_293 ();
 sg13g2_decap_4 FILLER_24_301 ();
 sg13g2_decap_4 FILLER_24_369 ();
 sg13g2_fill_1 FILLER_24_385 ();
 sg13g2_fill_2 FILLER_24_391 ();
 sg13g2_fill_2 FILLER_24_397 ();
 sg13g2_fill_1 FILLER_24_399 ();
 sg13g2_fill_2 FILLER_24_408 ();
 sg13g2_fill_1 FILLER_24_410 ();
 sg13g2_decap_8 FILLER_24_415 ();
 sg13g2_decap_8 FILLER_24_422 ();
 sg13g2_fill_1 FILLER_24_429 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_fill_2 FILLER_25_28 ();
 sg13g2_decap_4 FILLER_25_60 ();
 sg13g2_fill_1 FILLER_25_80 ();
 sg13g2_decap_4 FILLER_25_119 ();
 sg13g2_fill_2 FILLER_25_134 ();
 sg13g2_fill_2 FILLER_25_153 ();
 sg13g2_fill_2 FILLER_25_160 ();
 sg13g2_fill_1 FILLER_25_162 ();
 sg13g2_fill_2 FILLER_25_170 ();
 sg13g2_fill_1 FILLER_25_172 ();
 sg13g2_fill_2 FILLER_25_181 ();
 sg13g2_decap_8 FILLER_25_197 ();
 sg13g2_decap_4 FILLER_25_204 ();
 sg13g2_fill_1 FILLER_25_208 ();
 sg13g2_fill_2 FILLER_25_235 ();
 sg13g2_fill_1 FILLER_25_237 ();
 sg13g2_decap_8 FILLER_25_254 ();
 sg13g2_decap_8 FILLER_25_261 ();
 sg13g2_fill_2 FILLER_25_268 ();
 sg13g2_decap_8 FILLER_25_290 ();
 sg13g2_decap_8 FILLER_25_297 ();
 sg13g2_decap_8 FILLER_25_308 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_decap_8 FILLER_25_322 ();
 sg13g2_decap_4 FILLER_25_329 ();
 sg13g2_decap_4 FILLER_25_346 ();
 sg13g2_decap_8 FILLER_25_354 ();
 sg13g2_fill_1 FILLER_25_366 ();
 sg13g2_fill_2 FILLER_25_401 ();
 sg13g2_fill_1 FILLER_25_403 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_fill_1 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_19 ();
 sg13g2_decap_8 FILLER_26_26 ();
 sg13g2_fill_1 FILLER_26_33 ();
 sg13g2_fill_2 FILLER_26_46 ();
 sg13g2_decap_4 FILLER_26_52 ();
 sg13g2_fill_1 FILLER_26_56 ();
 sg13g2_fill_1 FILLER_26_71 ();
 sg13g2_fill_2 FILLER_26_76 ();
 sg13g2_fill_2 FILLER_26_88 ();
 sg13g2_decap_8 FILLER_26_103 ();
 sg13g2_decap_8 FILLER_26_110 ();
 sg13g2_decap_8 FILLER_26_117 ();
 sg13g2_decap_8 FILLER_26_124 ();
 sg13g2_decap_4 FILLER_26_131 ();
 sg13g2_fill_1 FILLER_26_135 ();
 sg13g2_decap_4 FILLER_26_140 ();
 sg13g2_fill_1 FILLER_26_144 ();
 sg13g2_fill_1 FILLER_26_168 ();
 sg13g2_decap_4 FILLER_26_177 ();
 sg13g2_decap_8 FILLER_26_185 ();
 sg13g2_decap_8 FILLER_26_192 ();
 sg13g2_decap_8 FILLER_26_199 ();
 sg13g2_fill_2 FILLER_26_206 ();
 sg13g2_fill_1 FILLER_26_208 ();
 sg13g2_fill_2 FILLER_26_244 ();
 sg13g2_decap_4 FILLER_26_259 ();
 sg13g2_fill_2 FILLER_26_263 ();
 sg13g2_fill_2 FILLER_26_282 ();
 sg13g2_fill_1 FILLER_26_284 ();
 sg13g2_decap_8 FILLER_26_290 ();
 sg13g2_fill_2 FILLER_26_336 ();
 sg13g2_fill_1 FILLER_26_338 ();
 sg13g2_fill_2 FILLER_26_377 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_4 FILLER_26_399 ();
 sg13g2_decap_4 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_26_415 ();
 sg13g2_decap_8 FILLER_26_422 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_fill_2 FILLER_27_42 ();
 sg13g2_fill_2 FILLER_27_49 ();
 sg13g2_fill_1 FILLER_27_51 ();
 sg13g2_decap_4 FILLER_27_60 ();
 sg13g2_fill_1 FILLER_27_77 ();
 sg13g2_fill_1 FILLER_27_83 ();
 sg13g2_decap_8 FILLER_27_89 ();
 sg13g2_decap_4 FILLER_27_96 ();
 sg13g2_decap_4 FILLER_27_105 ();
 sg13g2_fill_2 FILLER_27_109 ();
 sg13g2_fill_1 FILLER_27_116 ();
 sg13g2_fill_2 FILLER_27_127 ();
 sg13g2_decap_8 FILLER_27_155 ();
 sg13g2_decap_8 FILLER_27_162 ();
 sg13g2_decap_4 FILLER_27_169 ();
 sg13g2_fill_1 FILLER_27_173 ();
 sg13g2_decap_4 FILLER_27_206 ();
 sg13g2_fill_1 FILLER_27_210 ();
 sg13g2_fill_1 FILLER_27_221 ();
 sg13g2_decap_8 FILLER_27_235 ();
 sg13g2_decap_8 FILLER_27_242 ();
 sg13g2_decap_8 FILLER_27_249 ();
 sg13g2_fill_2 FILLER_27_256 ();
 sg13g2_fill_2 FILLER_27_266 ();
 sg13g2_fill_1 FILLER_27_268 ();
 sg13g2_fill_2 FILLER_27_282 ();
 sg13g2_decap_8 FILLER_27_288 ();
 sg13g2_decap_8 FILLER_27_295 ();
 sg13g2_decap_8 FILLER_27_302 ();
 sg13g2_decap_4 FILLER_27_309 ();
 sg13g2_fill_1 FILLER_27_313 ();
 sg13g2_decap_8 FILLER_27_321 ();
 sg13g2_decap_4 FILLER_27_328 ();
 sg13g2_fill_2 FILLER_27_332 ();
 sg13g2_fill_2 FILLER_27_342 ();
 sg13g2_fill_1 FILLER_27_360 ();
 sg13g2_decap_8 FILLER_27_370 ();
 sg13g2_decap_4 FILLER_27_377 ();
 sg13g2_fill_1 FILLER_27_381 ();
 sg13g2_decap_8 FILLER_27_388 ();
 sg13g2_decap_4 FILLER_27_395 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_11 ();
 sg13g2_decap_4 FILLER_28_18 ();
 sg13g2_fill_2 FILLER_28_30 ();
 sg13g2_fill_1 FILLER_28_76 ();
 sg13g2_fill_2 FILLER_28_92 ();
 sg13g2_fill_1 FILLER_28_94 ();
 sg13g2_decap_8 FILLER_28_110 ();
 sg13g2_fill_2 FILLER_28_117 ();
 sg13g2_fill_1 FILLER_28_119 ();
 sg13g2_fill_2 FILLER_28_127 ();
 sg13g2_fill_1 FILLER_28_129 ();
 sg13g2_fill_2 FILLER_28_133 ();
 sg13g2_decap_4 FILLER_28_140 ();
 sg13g2_fill_2 FILLER_28_144 ();
 sg13g2_fill_1 FILLER_28_177 ();
 sg13g2_decap_4 FILLER_28_187 ();
 sg13g2_decap_4 FILLER_28_196 ();
 sg13g2_fill_1 FILLER_28_200 ();
 sg13g2_fill_1 FILLER_28_206 ();
 sg13g2_decap_8 FILLER_28_211 ();
 sg13g2_fill_1 FILLER_28_218 ();
 sg13g2_fill_2 FILLER_28_230 ();
 sg13g2_fill_1 FILLER_28_236 ();
 sg13g2_decap_8 FILLER_28_246 ();
 sg13g2_decap_4 FILLER_28_253 ();
 sg13g2_fill_2 FILLER_28_267 ();
 sg13g2_fill_1 FILLER_28_269 ();
 sg13g2_decap_4 FILLER_28_288 ();
 sg13g2_fill_2 FILLER_28_292 ();
 sg13g2_decap_8 FILLER_28_332 ();
 sg13g2_decap_4 FILLER_28_339 ();
 sg13g2_fill_2 FILLER_28_343 ();
 sg13g2_fill_1 FILLER_28_352 ();
 sg13g2_fill_1 FILLER_28_403 ();
 sg13g2_decap_8 FILLER_28_413 ();
 sg13g2_decap_8 FILLER_28_420 ();
 sg13g2_fill_2 FILLER_28_427 ();
 sg13g2_fill_1 FILLER_28_429 ();
 sg13g2_fill_1 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_27 ();
 sg13g2_fill_1 FILLER_29_45 ();
 sg13g2_fill_2 FILLER_29_80 ();
 sg13g2_fill_1 FILLER_29_82 ();
 sg13g2_decap_4 FILLER_29_92 ();
 sg13g2_decap_8 FILLER_29_101 ();
 sg13g2_fill_2 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_fill_1 FILLER_29_126 ();
 sg13g2_fill_1 FILLER_29_139 ();
 sg13g2_decap_8 FILLER_29_148 ();
 sg13g2_decap_4 FILLER_29_155 ();
 sg13g2_decap_8 FILLER_29_163 ();
 sg13g2_fill_2 FILLER_29_170 ();
 sg13g2_fill_1 FILLER_29_172 ();
 sg13g2_fill_2 FILLER_29_187 ();
 sg13g2_fill_1 FILLER_29_198 ();
 sg13g2_fill_1 FILLER_29_211 ();
 sg13g2_fill_1 FILLER_29_216 ();
 sg13g2_fill_2 FILLER_29_222 ();
 sg13g2_decap_8 FILLER_29_250 ();
 sg13g2_decap_8 FILLER_29_257 ();
 sg13g2_fill_2 FILLER_29_264 ();
 sg13g2_fill_1 FILLER_29_266 ();
 sg13g2_decap_8 FILLER_29_277 ();
 sg13g2_decap_8 FILLER_29_284 ();
 sg13g2_decap_8 FILLER_29_291 ();
 sg13g2_fill_1 FILLER_29_298 ();
 sg13g2_decap_8 FILLER_29_303 ();
 sg13g2_decap_8 FILLER_29_310 ();
 sg13g2_decap_8 FILLER_29_317 ();
 sg13g2_fill_2 FILLER_29_324 ();
 sg13g2_fill_1 FILLER_29_326 ();
 sg13g2_fill_1 FILLER_29_336 ();
 sg13g2_fill_1 FILLER_29_348 ();
 sg13g2_fill_1 FILLER_29_352 ();
 sg13g2_decap_4 FILLER_29_373 ();
 sg13g2_decap_8 FILLER_29_381 ();
 sg13g2_decap_4 FILLER_29_388 ();
 sg13g2_decap_8 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_29_415 ();
 sg13g2_decap_8 FILLER_29_422 ();
 sg13g2_fill_1 FILLER_29_429 ();
 sg13g2_fill_2 FILLER_30_30 ();
 sg13g2_fill_2 FILLER_30_41 ();
 sg13g2_fill_1 FILLER_30_54 ();
 sg13g2_fill_2 FILLER_30_69 ();
 sg13g2_fill_1 FILLER_30_71 ();
 sg13g2_fill_2 FILLER_30_79 ();
 sg13g2_fill_1 FILLER_30_81 ();
 sg13g2_decap_4 FILLER_30_87 ();
 sg13g2_fill_2 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_123 ();
 sg13g2_decap_4 FILLER_30_130 ();
 sg13g2_fill_2 FILLER_30_134 ();
 sg13g2_decap_8 FILLER_30_141 ();
 sg13g2_decap_4 FILLER_30_148 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_4 FILLER_30_173 ();
 sg13g2_fill_2 FILLER_30_177 ();
 sg13g2_fill_1 FILLER_30_188 ();
 sg13g2_fill_1 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_237 ();
 sg13g2_fill_2 FILLER_30_257 ();
 sg13g2_decap_8 FILLER_30_289 ();
 sg13g2_fill_1 FILLER_30_296 ();
 sg13g2_decap_8 FILLER_30_301 ();
 sg13g2_decap_4 FILLER_30_308 ();
 sg13g2_decap_8 FILLER_30_329 ();
 sg13g2_decap_8 FILLER_30_336 ();
 sg13g2_fill_2 FILLER_30_383 ();
 sg13g2_fill_2 FILLER_30_389 ();
 sg13g2_fill_2 FILLER_30_396 ();
 sg13g2_fill_1 FILLER_30_398 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_11 ();
 sg13g2_decap_4 FILLER_31_18 ();
 sg13g2_fill_2 FILLER_31_22 ();
 sg13g2_decap_4 FILLER_31_37 ();
 sg13g2_fill_1 FILLER_31_41 ();
 sg13g2_fill_1 FILLER_31_66 ();
 sg13g2_decap_8 FILLER_31_72 ();
 sg13g2_decap_8 FILLER_31_79 ();
 sg13g2_decap_8 FILLER_31_86 ();
 sg13g2_decap_4 FILLER_31_93 ();
 sg13g2_fill_2 FILLER_31_97 ();
 sg13g2_decap_8 FILLER_31_108 ();
 sg13g2_decap_8 FILLER_31_115 ();
 sg13g2_decap_4 FILLER_31_122 ();
 sg13g2_fill_2 FILLER_31_126 ();
 sg13g2_fill_1 FILLER_31_141 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_decap_4 FILLER_31_182 ();
 sg13g2_decap_4 FILLER_31_197 ();
 sg13g2_decap_8 FILLER_31_206 ();
 sg13g2_decap_8 FILLER_31_213 ();
 sg13g2_decap_4 FILLER_31_220 ();
 sg13g2_fill_1 FILLER_31_224 ();
 sg13g2_decap_8 FILLER_31_239 ();
 sg13g2_decap_8 FILLER_31_246 ();
 sg13g2_fill_1 FILLER_31_253 ();
 sg13g2_decap_8 FILLER_31_271 ();
 sg13g2_decap_8 FILLER_31_278 ();
 sg13g2_fill_2 FILLER_31_285 ();
 sg13g2_fill_1 FILLER_31_287 ();
 sg13g2_decap_4 FILLER_31_318 ();
 sg13g2_decap_4 FILLER_31_327 ();
 sg13g2_fill_1 FILLER_31_331 ();
 sg13g2_fill_1 FILLER_31_336 ();
 sg13g2_decap_4 FILLER_31_344 ();
 sg13g2_fill_2 FILLER_31_348 ();
 sg13g2_fill_2 FILLER_31_361 ();
 sg13g2_fill_1 FILLER_31_363 ();
 sg13g2_fill_2 FILLER_31_370 ();
 sg13g2_decap_8 FILLER_31_378 ();
 sg13g2_fill_1 FILLER_31_385 ();
 sg13g2_decap_4 FILLER_31_403 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_31_413 ();
 sg13g2_decap_8 FILLER_31_420 ();
 sg13g2_fill_2 FILLER_31_427 ();
 sg13g2_fill_1 FILLER_31_429 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_fill_2 FILLER_32_21 ();
 sg13g2_fill_2 FILLER_32_34 ();
 sg13g2_decap_8 FILLER_32_69 ();
 sg13g2_decap_8 FILLER_32_76 ();
 sg13g2_decap_8 FILLER_32_83 ();
 sg13g2_decap_4 FILLER_32_90 ();
 sg13g2_fill_1 FILLER_32_94 ();
 sg13g2_decap_4 FILLER_32_130 ();
 sg13g2_fill_1 FILLER_32_134 ();
 sg13g2_decap_4 FILLER_32_145 ();
 sg13g2_fill_1 FILLER_32_149 ();
 sg13g2_decap_4 FILLER_32_154 ();
 sg13g2_fill_2 FILLER_32_195 ();
 sg13g2_decap_4 FILLER_32_203 ();
 sg13g2_fill_2 FILLER_32_207 ();
 sg13g2_fill_1 FILLER_32_213 ();
 sg13g2_fill_2 FILLER_32_219 ();
 sg13g2_fill_1 FILLER_32_226 ();
 sg13g2_fill_2 FILLER_32_237 ();
 sg13g2_fill_1 FILLER_32_251 ();
 sg13g2_fill_1 FILLER_32_265 ();
 sg13g2_fill_1 FILLER_32_270 ();
 sg13g2_decap_8 FILLER_32_275 ();
 sg13g2_fill_2 FILLER_32_282 ();
 sg13g2_fill_2 FILLER_32_314 ();
 sg13g2_fill_2 FILLER_32_336 ();
 sg13g2_fill_1 FILLER_32_338 ();
 sg13g2_fill_1 FILLER_32_348 ();
 sg13g2_decap_4 FILLER_32_376 ();
 sg13g2_fill_1 FILLER_32_380 ();
 sg13g2_decap_8 FILLER_32_401 ();
 sg13g2_fill_2 FILLER_32_408 ();
 sg13g2_fill_1 FILLER_32_410 ();
 sg13g2_decap_4 FILLER_32_415 ();
 sg13g2_fill_1 FILLER_32_419 ();
 sg13g2_decap_4 FILLER_32_425 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_fill_1 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_27 ();
 sg13g2_fill_1 FILLER_33_34 ();
 sg13g2_fill_1 FILLER_33_40 ();
 sg13g2_fill_1 FILLER_33_50 ();
 sg13g2_decap_4 FILLER_33_69 ();
 sg13g2_fill_1 FILLER_33_73 ();
 sg13g2_decap_8 FILLER_33_78 ();
 sg13g2_decap_4 FILLER_33_85 ();
 sg13g2_decap_8 FILLER_33_93 ();
 sg13g2_decap_8 FILLER_33_100 ();
 sg13g2_decap_4 FILLER_33_107 ();
 sg13g2_decap_8 FILLER_33_115 ();
 sg13g2_decap_8 FILLER_33_122 ();
 sg13g2_decap_4 FILLER_33_143 ();
 sg13g2_fill_2 FILLER_33_147 ();
 sg13g2_fill_1 FILLER_33_154 ();
 sg13g2_fill_2 FILLER_33_167 ();
 sg13g2_decap_4 FILLER_33_194 ();
 sg13g2_fill_2 FILLER_33_198 ();
 sg13g2_decap_4 FILLER_33_205 ();
 sg13g2_fill_1 FILLER_33_209 ();
 sg13g2_decap_8 FILLER_33_216 ();
 sg13g2_decap_8 FILLER_33_223 ();
 sg13g2_fill_1 FILLER_33_240 ();
 sg13g2_decap_8 FILLER_33_245 ();
 sg13g2_fill_2 FILLER_33_252 ();
 sg13g2_decap_8 FILLER_33_285 ();
 sg13g2_fill_1 FILLER_33_292 ();
 sg13g2_decap_8 FILLER_33_297 ();
 sg13g2_fill_2 FILLER_33_304 ();
 sg13g2_fill_1 FILLER_33_306 ();
 sg13g2_fill_1 FILLER_33_318 ();
 sg13g2_fill_1 FILLER_33_323 ();
 sg13g2_decap_4 FILLER_33_344 ();
 sg13g2_decap_4 FILLER_33_358 ();
 sg13g2_decap_8 FILLER_33_367 ();
 sg13g2_decap_4 FILLER_33_374 ();
 sg13g2_fill_2 FILLER_33_378 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_9 ();
 sg13g2_fill_1 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_18 ();
 sg13g2_fill_2 FILLER_34_25 ();
 sg13g2_decap_8 FILLER_34_61 ();
 sg13g2_fill_1 FILLER_34_68 ();
 sg13g2_fill_2 FILLER_34_79 ();
 sg13g2_fill_1 FILLER_34_81 ();
 sg13g2_fill_2 FILLER_34_108 ();
 sg13g2_decap_8 FILLER_34_146 ();
 sg13g2_decap_4 FILLER_34_161 ();
 sg13g2_fill_1 FILLER_34_165 ();
 sg13g2_decap_4 FILLER_34_175 ();
 sg13g2_fill_1 FILLER_34_179 ();
 sg13g2_fill_1 FILLER_34_196 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_8 FILLER_34_222 ();
 sg13g2_fill_1 FILLER_34_229 ();
 sg13g2_decap_4 FILLER_34_235 ();
 sg13g2_fill_1 FILLER_34_247 ();
 sg13g2_fill_1 FILLER_34_266 ();
 sg13g2_decap_8 FILLER_34_285 ();
 sg13g2_decap_8 FILLER_34_292 ();
 sg13g2_decap_8 FILLER_34_299 ();
 sg13g2_fill_1 FILLER_34_306 ();
 sg13g2_fill_1 FILLER_34_311 ();
 sg13g2_decap_4 FILLER_34_317 ();
 sg13g2_decap_8 FILLER_34_333 ();
 sg13g2_fill_2 FILLER_34_340 ();
 sg13g2_decap_8 FILLER_34_346 ();
 sg13g2_decap_4 FILLER_34_353 ();
 sg13g2_fill_1 FILLER_34_369 ();
 sg13g2_decap_4 FILLER_34_375 ();
 sg13g2_fill_2 FILLER_34_379 ();
 sg13g2_fill_1 FILLER_34_385 ();
 sg13g2_decap_8 FILLER_34_390 ();
 sg13g2_fill_2 FILLER_34_397 ();
 sg13g2_fill_1 FILLER_34_429 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_39 ();
 sg13g2_decap_4 FILLER_35_46 ();
 sg13g2_fill_2 FILLER_35_50 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_fill_2 FILLER_35_63 ();
 sg13g2_fill_1 FILLER_35_65 ();
 sg13g2_decap_8 FILLER_35_110 ();
 sg13g2_decap_4 FILLER_35_121 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_fill_1 FILLER_35_170 ();
 sg13g2_fill_2 FILLER_35_177 ();
 sg13g2_fill_1 FILLER_35_179 ();
 sg13g2_decap_4 FILLER_35_184 ();
 sg13g2_fill_1 FILLER_35_192 ();
 sg13g2_decap_8 FILLER_35_224 ();
 sg13g2_decap_8 FILLER_35_231 ();
 sg13g2_decap_8 FILLER_35_238 ();
 sg13g2_decap_4 FILLER_35_254 ();
 sg13g2_fill_1 FILLER_35_258 ();
 sg13g2_fill_2 FILLER_35_263 ();
 sg13g2_fill_1 FILLER_35_265 ();
 sg13g2_fill_1 FILLER_35_292 ();
 sg13g2_fill_1 FILLER_35_319 ();
 sg13g2_fill_1 FILLER_35_346 ();
 sg13g2_fill_2 FILLER_35_373 ();
 sg13g2_decap_4 FILLER_35_405 ();
 sg13g2_fill_1 FILLER_35_409 ();
 sg13g2_fill_2 FILLER_35_414 ();
 sg13g2_fill_1 FILLER_35_416 ();
 sg13g2_decap_8 FILLER_35_422 ();
 sg13g2_fill_1 FILLER_35_429 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_71 ();
 sg13g2_decap_8 FILLER_36_78 ();
 sg13g2_decap_8 FILLER_36_94 ();
 sg13g2_fill_2 FILLER_36_127 ();
 sg13g2_decap_4 FILLER_36_133 ();
 sg13g2_fill_2 FILLER_36_137 ();
 sg13g2_fill_1 FILLER_36_144 ();
 sg13g2_fill_1 FILLER_36_148 ();
 sg13g2_fill_2 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_160 ();
 sg13g2_decap_4 FILLER_36_167 ();
 sg13g2_fill_2 FILLER_36_179 ();
 sg13g2_fill_1 FILLER_36_181 ();
 sg13g2_fill_2 FILLER_36_186 ();
 sg13g2_fill_1 FILLER_36_188 ();
 sg13g2_decap_8 FILLER_36_219 ();
 sg13g2_decap_8 FILLER_36_226 ();
 sg13g2_decap_4 FILLER_36_233 ();
 sg13g2_fill_1 FILLER_36_237 ();
 sg13g2_decap_8 FILLER_36_269 ();
 sg13g2_decap_8 FILLER_36_276 ();
 sg13g2_fill_1 FILLER_36_283 ();
 sg13g2_decap_8 FILLER_36_288 ();
 sg13g2_decap_4 FILLER_36_295 ();
 sg13g2_fill_2 FILLER_36_299 ();
 sg13g2_fill_2 FILLER_36_305 ();
 sg13g2_fill_1 FILLER_36_307 ();
 sg13g2_fill_1 FILLER_36_311 ();
 sg13g2_fill_1 FILLER_36_315 ();
 sg13g2_decap_8 FILLER_36_321 ();
 sg13g2_fill_2 FILLER_36_332 ();
 sg13g2_fill_2 FILLER_36_339 ();
 sg13g2_fill_1 FILLER_36_341 ();
 sg13g2_decap_4 FILLER_36_350 ();
 sg13g2_decap_4 FILLER_36_358 ();
 sg13g2_fill_1 FILLER_36_362 ();
 sg13g2_decap_8 FILLER_36_368 ();
 sg13g2_decap_4 FILLER_36_375 ();
 sg13g2_fill_2 FILLER_36_389 ();
 sg13g2_fill_1 FILLER_36_391 ();
 sg13g2_fill_2 FILLER_36_402 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_fill_2 FILLER_37_91 ();
 sg13g2_fill_1 FILLER_37_93 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_fill_1 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_110 ();
 sg13g2_fill_1 FILLER_37_117 ();
 sg13g2_fill_2 FILLER_37_181 ();
 sg13g2_decap_4 FILLER_37_209 ();
 sg13g2_decap_4 FILLER_37_218 ();
 sg13g2_fill_2 FILLER_37_229 ();
 sg13g2_fill_1 FILLER_37_231 ();
 sg13g2_fill_2 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_decap_8 FILLER_37_406 ();
 sg13g2_decap_8 FILLER_37_413 ();
 sg13g2_decap_8 FILLER_37_420 ();
 sg13g2_fill_2 FILLER_37_427 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_fill_1 FILLER_38_141 ();
 sg13g2_fill_1 FILLER_38_146 ();
 sg13g2_fill_1 FILLER_38_151 ();
 sg13g2_fill_1 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_201 ();
 sg13g2_decap_4 FILLER_38_216 ();
 sg13g2_fill_2 FILLER_38_224 ();
 sg13g2_fill_1 FILLER_38_234 ();
 sg13g2_fill_1 FILLER_38_239 ();
 sg13g2_fill_1 FILLER_38_244 ();
 sg13g2_fill_2 FILLER_38_264 ();
 sg13g2_decap_4 FILLER_38_270 ();
 sg13g2_fill_1 FILLER_38_274 ();
 sg13g2_decap_8 FILLER_38_279 ();
 sg13g2_decap_8 FILLER_38_286 ();
 sg13g2_decap_8 FILLER_38_297 ();
 sg13g2_decap_8 FILLER_38_304 ();
 sg13g2_decap_8 FILLER_38_311 ();
 sg13g2_decap_8 FILLER_38_322 ();
 sg13g2_decap_8 FILLER_38_329 ();
 sg13g2_decap_4 FILLER_38_336 ();
 sg13g2_fill_1 FILLER_38_340 ();
 sg13g2_fill_2 FILLER_38_349 ();
 sg13g2_decap_4 FILLER_38_355 ();
 sg13g2_fill_2 FILLER_38_371 ();
 sg13g2_fill_2 FILLER_38_388 ();
 sg13g2_fill_1 FILLER_38_390 ();
 sg13g2_fill_2 FILLER_38_395 ();
 sg13g2_decap_8 FILLER_38_402 ();
 sg13g2_fill_2 FILLER_38_409 ();
 sg13g2_decap_8 FILLER_38_415 ();
 sg13g2_decap_8 FILLER_38_422 ();
 sg13g2_fill_1 FILLER_38_429 ();
endmodule
