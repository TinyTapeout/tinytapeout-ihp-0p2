module tt_um_phansel_laplace_lut (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire clknet_0_clk;
 wire net221;
 wire \chars_remaining[0] ;
 wire \chars_remaining[1] ;
 wire \chars_remaining[2] ;
 wire \chars_remaining[3] ;
 wire \chars_remaining[4] ;
 wire \chars_remaining[5] ;
 wire \chars_remaining[6] ;
 wire \chars_remaining[7] ;
 wire \chars_remaining[8] ;
 wire \chars_remaining[9] ;
 wire clk_buffered;
 wire \clk_picker.clk_slow ;
 wire \clk_picker.counter[0] ;
 wire \clk_picker.counter[10] ;
 wire \clk_picker.counter[11] ;
 wire \clk_picker.counter[12] ;
 wire \clk_picker.counter[13] ;
 wire \clk_picker.counter[14] ;
 wire \clk_picker.counter[15] ;
 wire \clk_picker.counter[16] ;
 wire \clk_picker.counter[17] ;
 wire \clk_picker.counter[18] ;
 wire \clk_picker.counter[19] ;
 wire \clk_picker.counter[1] ;
 wire \clk_picker.counter[20] ;
 wire \clk_picker.counter[21] ;
 wire \clk_picker.counter[22] ;
 wire \clk_picker.counter[23] ;
 wire \clk_picker.counter[24] ;
 wire \clk_picker.counter[25] ;
 wire \clk_picker.counter[2] ;
 wire \clk_picker.counter[3] ;
 wire \clk_picker.counter[4] ;
 wire \clk_picker.counter[5] ;
 wire \clk_picker.counter[6] ;
 wire \clk_picker.counter[7] ;
 wire \clk_picker.counter[8] ;
 wire \clk_picker.counter[9] ;
 wire \line_mapper_1.pointer_addr[0] ;
 wire \line_mapper_1.pointer_addr[10] ;
 wire \line_mapper_1.pointer_addr[11] ;
 wire \line_mapper_1.pointer_addr[12] ;
 wire \line_mapper_1.pointer_addr[13] ;
 wire \line_mapper_1.pointer_addr[14] ;
 wire \line_mapper_1.pointer_addr[15] ;
 wire \line_mapper_1.pointer_addr[1] ;
 wire \line_mapper_1.pointer_addr[2] ;
 wire \line_mapper_1.pointer_addr[3] ;
 wire \line_mapper_1.pointer_addr[4] ;
 wire \line_mapper_1.pointer_addr[5] ;
 wire \line_mapper_1.pointer_addr[6] ;
 wire \line_mapper_1.pointer_addr[7] ;
 wire \line_mapper_1.pointer_addr[8] ;
 wire \line_mapper_1.pointer_addr[9] ;
 wire \mem_addr[0] ;
 wire \mem_addr[1] ;
 wire \mem_addr[2] ;
 wire \mem_addr[3] ;
 wire \mem_addr[4] ;
 wire \mem_addr[5] ;
 wire \mem_addr[6] ;
 wire \mem_addr[7] ;
 wire \mem_addr[8] ;
 wire \memory_1.mem_addr[9] ;
 wire \transformer_1.started ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_level_0_1_10_clk;
 wire clknet_level_1_1_11_clk;
 wire clknet_level_2_1_12_clk;
 wire clknet_level_0_1_23_clk;
 wire clknet_level_1_1_24_clk;
 wire clknet_level_2_1_25_clk;
 wire clknet_level_0_1_36_clk;
 wire clknet_level_1_1_37_clk;
 wire clknet_level_2_1_38_clk;
 wire clknet_level_0_1_49_clk;
 wire clknet_level_1_1_410_clk;
 wire clknet_level_2_1_411_clk;
 wire clknet_0_clk_buffered;
 wire clknet_3_0__leaf_clk_buffered;
 wire clknet_3_1__leaf_clk_buffered;
 wire clknet_3_2__leaf_clk_buffered;
 wire clknet_3_3__leaf_clk_buffered;
 wire clknet_3_4__leaf_clk_buffered;
 wire clknet_3_5__leaf_clk_buffered;
 wire clknet_3_6__leaf_clk_buffered;
 wire clknet_3_7__leaf_clk_buffered;

 sg13g2_buf_8 _3120_ (.A(\mem_addr[2] ),
    .X(_0725_));
 sg13g2_inv_2 _3121_ (.Y(_0736_),
    .A(_0725_));
 sg13g2_buf_8 _3122_ (.A(_0736_),
    .X(_0746_));
 sg13g2_buf_8 _3123_ (.A(net190),
    .X(_0757_));
 sg13g2_buf_8 _3124_ (.A(\mem_addr[1] ),
    .X(_0768_));
 sg13g2_inv_4 _3125_ (.A(_0768_),
    .Y(_0779_));
 sg13g2_buf_1 _3126_ (.A(_0779_),
    .X(_0790_));
 sg13g2_nand2_1 _3127_ (.Y(_0801_),
    .A(net158),
    .B(net189));
 sg13g2_buf_4 _3128_ (.X(_0812_),
    .A(\mem_addr[3] ));
 sg13g2_inv_2 _3129_ (.Y(_0823_),
    .A(_0812_));
 sg13g2_buf_8 _3130_ (.A(_0823_),
    .X(_0834_));
 sg13g2_buf_8 _3131_ (.A(net188),
    .X(_0845_));
 sg13g2_buf_8 _3132_ (.A(net157),
    .X(_0856_));
 sg13g2_buf_8 _3133_ (.A(_0725_),
    .X(_0867_));
 sg13g2_buf_16 _3134_ (.X(_0878_),
    .A(\mem_addr[0] ));
 sg13g2_buf_8 _3135_ (.A(_0878_),
    .X(_0889_));
 sg13g2_nand2_1 _3136_ (.Y(_0900_),
    .A(net208),
    .B(net207));
 sg13g2_buf_1 _3137_ (.A(_0900_),
    .X(_0910_));
 sg13g2_nand3_1 _3138_ (.B(net111),
    .C(net156),
    .A(_0801_),
    .Y(_0921_));
 sg13g2_buf_4 _3139_ (.X(_0932_),
    .A(_0037_));
 sg13g2_buf_2 _3140_ (.A(_0932_),
    .X(_0943_));
 sg13g2_nor2_1 _3141_ (.A(_0768_),
    .B(_0878_),
    .Y(_0954_));
 sg13g2_buf_2 _3142_ (.A(_0954_),
    .X(_0965_));
 sg13g2_buf_1 _3143_ (.A(_0965_),
    .X(_0976_));
 sg13g2_nor2_2 _3144_ (.A(net206),
    .B(_0976_),
    .Y(_0987_));
 sg13g2_buf_8 _3145_ (.A(_0812_),
    .X(_0998_));
 sg13g2_buf_8 _3146_ (.A(net205),
    .X(_1009_));
 sg13g2_buf_8 _3147_ (.A(net187),
    .X(_1020_));
 sg13g2_nand2_1 _3148_ (.Y(_1031_),
    .A(_0987_),
    .B(net154));
 sg13g2_buf_2 _3149_ (.A(\mem_addr[4] ),
    .X(_1042_));
 sg13g2_buf_8 _3150_ (.A(\mem_addr[5] ),
    .X(_1053_));
 sg13g2_inv_1 _3151_ (.Y(_1064_),
    .A(net210));
 sg13g2_nor2_1 _3152_ (.A(_1042_),
    .B(_1064_),
    .Y(_1074_));
 sg13g2_buf_2 _3153_ (.A(_1074_),
    .X(_1085_));
 sg13g2_inv_2 _3154_ (.Y(_1096_),
    .A(_1085_));
 sg13g2_buf_2 _3155_ (.A(_1096_),
    .X(_1107_));
 sg13g2_a21oi_1 _3156_ (.A1(_0921_),
    .A2(_1031_),
    .Y(_1118_),
    .B1(net64));
 sg13g2_inv_4 _3157_ (.A(_0878_),
    .Y(_1129_));
 sg13g2_nand2_1 _3158_ (.Y(_1140_),
    .A(net190),
    .B(_1129_));
 sg13g2_buf_4 _3159_ (.X(_1151_),
    .A(_1140_));
 sg13g2_buf_2 _3160_ (.A(_0032_),
    .X(_1162_));
 sg13g2_nand2_1 _3161_ (.Y(_1173_),
    .A(net208),
    .B(_1162_));
 sg13g2_buf_4 _3162_ (.X(_1184_),
    .A(_1173_));
 sg13g2_nand2_1 _3163_ (.Y(_1195_),
    .A(_1151_),
    .B(_1184_));
 sg13g2_buf_8 _3164_ (.A(_0768_),
    .X(_1205_));
 sg13g2_nor2_2 _3165_ (.A(net208),
    .B(net204),
    .Y(_1216_));
 sg13g2_nor2_2 _3166_ (.A(net205),
    .B(_1216_),
    .Y(_1227_));
 sg13g2_nand2_2 _3167_ (.Y(_1238_),
    .A(_1195_),
    .B(_1227_));
 sg13g2_buf_8 _3168_ (.A(net204),
    .X(_1249_));
 sg13g2_buf_8 _3169_ (.A(net207),
    .X(_1260_));
 sg13g2_a21oi_2 _3170_ (.B1(net206),
    .Y(_1271_),
    .A2(net185),
    .A1(net186));
 sg13g2_buf_1 _3171_ (.A(net205),
    .X(_1282_));
 sg13g2_nand2_2 _3172_ (.Y(_1293_),
    .A(_1271_),
    .B(_1282_));
 sg13g2_nand2_1 _3173_ (.Y(_1304_),
    .A(_1238_),
    .B(_1293_));
 sg13g2_nand2_1 _3174_ (.Y(_1315_),
    .A(_1042_),
    .B(net210));
 sg13g2_buf_2 _3175_ (.A(_1315_),
    .X(_1326_));
 sg13g2_inv_1 _3176_ (.Y(_1336_),
    .A(_1326_));
 sg13g2_buf_1 _3177_ (.A(_1336_),
    .X(_1347_));
 sg13g2_nand2_1 _3178_ (.Y(_1358_),
    .A(_1304_),
    .B(net110));
 sg13g2_buf_2 _3179_ (.A(\mem_addr[6] ),
    .X(_1369_));
 sg13g2_buf_2 _3180_ (.A(net209),
    .X(_1380_));
 sg13g2_nand2_1 _3181_ (.Y(_1391_),
    .A(_1358_),
    .B(net203));
 sg13g2_nor2_1 _3182_ (.A(_1118_),
    .B(_1391_),
    .Y(_1402_));
 sg13g2_xnor2_1 _3183_ (.Y(_1413_),
    .A(net204),
    .B(_0878_));
 sg13g2_buf_8 _3184_ (.A(net208),
    .X(_1424_));
 sg13g2_buf_8 _3185_ (.A(_1424_),
    .X(_1435_));
 sg13g2_nand2_1 _3186_ (.Y(_1446_),
    .A(_1413_),
    .B(net153));
 sg13g2_inv_1 _3187_ (.Y(_1457_),
    .A(_1162_));
 sg13g2_nor2_1 _3188_ (.A(net208),
    .B(_1457_),
    .Y(_1467_));
 sg13g2_buf_2 _3189_ (.A(_1467_),
    .X(_1478_));
 sg13g2_nor2_1 _3190_ (.A(net157),
    .B(_1478_),
    .Y(_1489_));
 sg13g2_nand2_1 _3191_ (.Y(_1500_),
    .A(_1446_),
    .B(_1489_));
 sg13g2_buf_8 _3192_ (.A(net188),
    .X(_1511_));
 sg13g2_buf_1 _3193_ (.A(net152),
    .X(_1522_));
 sg13g2_inv_2 _3194_ (.Y(_1533_),
    .A(_1042_));
 sg13g2_buf_8 _3195_ (.A(_1533_),
    .X(_1544_));
 sg13g2_buf_1 _3196_ (.A(net182),
    .X(_1555_));
 sg13g2_a21oi_1 _3197_ (.A1(_0987_),
    .A2(net109),
    .Y(_1566_),
    .B1(net151));
 sg13g2_nand2_1 _3198_ (.Y(_1577_),
    .A(_1500_),
    .B(_1566_));
 sg13g2_buf_8 _3199_ (.A(_1129_),
    .X(_1588_));
 sg13g2_nor2_1 _3200_ (.A(_0725_),
    .B(_0779_),
    .Y(_1599_));
 sg13g2_buf_2 _3201_ (.A(_1599_),
    .X(_1609_));
 sg13g2_nor2_1 _3202_ (.A(net181),
    .B(_1609_),
    .Y(_1620_));
 sg13g2_buf_1 _3203_ (.A(net151),
    .X(_1631_));
 sg13g2_nand2_1 _3204_ (.Y(_1642_),
    .A(_0812_),
    .B(_0725_));
 sg13g2_buf_4 _3205_ (.X(_1653_),
    .A(_1642_));
 sg13g2_nand3_1 _3206_ (.B(net108),
    .C(_1653_),
    .A(_1620_),
    .Y(_1664_));
 sg13g2_nand2_1 _3207_ (.Y(_1675_),
    .A(_1577_),
    .B(_1664_));
 sg13g2_buf_1 _3208_ (.A(_1064_),
    .X(_1685_));
 sg13g2_buf_2 _3209_ (.A(net180),
    .X(_1696_));
 sg13g2_buf_1 _3210_ (.A(net150),
    .X(_1707_));
 sg13g2_nand2_1 _3211_ (.Y(_1718_),
    .A(_1675_),
    .B(net107));
 sg13g2_nand2_1 _3212_ (.Y(_1729_),
    .A(_1402_),
    .B(_1718_));
 sg13g2_buf_2 _3213_ (.A(_1042_),
    .X(_1740_));
 sg13g2_buf_1 _3214_ (.A(net202),
    .X(_1751_));
 sg13g2_nand2_1 _3215_ (.Y(_1762_),
    .A(_0768_),
    .B(_0878_));
 sg13g2_buf_8 _3216_ (.A(_1762_),
    .X(_1773_));
 sg13g2_nand2_1 _3217_ (.Y(_1784_),
    .A(net178),
    .B(net190));
 sg13g2_buf_4 _3218_ (.X(_1795_),
    .A(_1784_));
 sg13g2_nor2_2 _3219_ (.A(net188),
    .B(_1795_),
    .Y(_1805_));
 sg13g2_nor2_1 _3220_ (.A(net179),
    .B(_1805_),
    .Y(_1816_));
 sg13g2_nand2_1 _3221_ (.Y(_1827_),
    .A(net188),
    .B(net204));
 sg13g2_buf_8 _3222_ (.A(_1827_),
    .X(_1838_));
 sg13g2_inv_4 _3223_ (.A(_0932_),
    .Y(_1848_));
 sg13g2_nand2_2 _3224_ (.Y(_1859_),
    .A(net201),
    .B(net185));
 sg13g2_nor2_2 _3225_ (.A(net106),
    .B(_1859_),
    .Y(_1869_));
 sg13g2_inv_2 _3226_ (.Y(_1880_),
    .A(_1869_));
 sg13g2_nand2_1 _3227_ (.Y(_1890_),
    .A(_1816_),
    .B(_1880_));
 sg13g2_nand2_1 _3228_ (.Y(_1901_),
    .A(_0725_),
    .B(net204));
 sg13g2_buf_2 _3229_ (.A(_1901_),
    .X(_1911_));
 sg13g2_nand2_2 _3230_ (.Y(_1921_),
    .A(_1911_),
    .B(_0834_));
 sg13g2_nor2_2 _3231_ (.A(net185),
    .B(_1921_),
    .Y(_1930_));
 sg13g2_nand2_1 _3232_ (.Y(_1938_),
    .A(_1216_),
    .B(_0834_));
 sg13g2_buf_2 _3233_ (.A(_1938_),
    .X(_1948_));
 sg13g2_nand2_1 _3234_ (.Y(_1958_),
    .A(_1948_),
    .B(net202));
 sg13g2_nor2_2 _3235_ (.A(_1930_),
    .B(_1958_),
    .Y(_1968_));
 sg13g2_inv_1 _3236_ (.Y(_1976_),
    .A(_1968_));
 sg13g2_nand2_1 _3237_ (.Y(_1987_),
    .A(net205),
    .B(_1042_));
 sg13g2_buf_4 _3238_ (.X(_1998_),
    .A(_1987_));
 sg13g2_nand3_1 _3239_ (.B(net186),
    .C(net207),
    .A(net183),
    .Y(_2009_));
 sg13g2_buf_4 _3240_ (.X(_2020_),
    .A(_2009_));
 sg13g2_nand2_2 _3241_ (.Y(_2031_),
    .A(_1795_),
    .B(_2020_));
 sg13g2_nor2_1 _3242_ (.A(net209),
    .B(net180),
    .Y(_2042_));
 sg13g2_buf_1 _3243_ (.A(_2042_),
    .X(_2053_));
 sg13g2_o21ai_1 _3244_ (.B1(net105),
    .Y(_2064_),
    .A1(_1998_),
    .A2(_2031_));
 sg13g2_a21oi_1 _3245_ (.A1(_1890_),
    .A2(_1976_),
    .Y(_2075_),
    .B1(_2064_));
 sg13g2_nand2_2 _3246_ (.Y(_2086_),
    .A(_1413_),
    .B(net158));
 sg13g2_nand2_2 _3247_ (.Y(_2097_),
    .A(net178),
    .B(net183));
 sg13g2_nand3_1 _3248_ (.B(net152),
    .C(_2097_),
    .A(_2086_),
    .Y(_2108_));
 sg13g2_buf_2 _3249_ (.A(_2108_),
    .X(_2119_));
 sg13g2_nor2_1 _3250_ (.A(net210),
    .B(net209),
    .Y(_2130_));
 sg13g2_buf_2 _3251_ (.A(_2130_),
    .X(_2141_));
 sg13g2_nand2_1 _3252_ (.Y(_2151_),
    .A(_2119_),
    .B(_2141_));
 sg13g2_buf_1 _3253_ (.A(net202),
    .X(_2162_));
 sg13g2_buf_1 _3254_ (.A(net177),
    .X(_2173_));
 sg13g2_nand2_1 _3255_ (.Y(_2183_),
    .A(_0812_),
    .B(_0878_));
 sg13g2_buf_1 _3256_ (.A(_2183_),
    .X(_2193_));
 sg13g2_nor2_2 _3257_ (.A(net153),
    .B(net176),
    .Y(_2203_));
 sg13g2_nand2_1 _3258_ (.Y(_2212_),
    .A(_1216_),
    .B(net205));
 sg13g2_buf_4 _3259_ (.X(_2221_),
    .A(_2212_));
 sg13g2_inv_1 _3260_ (.Y(_2230_),
    .A(_2221_));
 sg13g2_nor2_2 _3261_ (.A(_2203_),
    .B(_2230_),
    .Y(_2239_));
 sg13g2_nand2_1 _3262_ (.Y(_2248_),
    .A(_0779_),
    .B(_0812_));
 sg13g2_buf_1 _3263_ (.A(_2248_),
    .X(_2257_));
 sg13g2_xnor2_1 _3264_ (.Y(_2266_),
    .A(net183),
    .B(net207));
 sg13g2_buf_4 _3265_ (.X(_2273_),
    .A(_2266_));
 sg13g2_nor2_2 _3266_ (.A(net148),
    .B(_2273_),
    .Y(_2279_));
 sg13g2_nor2_1 _3267_ (.A(net177),
    .B(_2279_),
    .Y(_2289_));
 sg13g2_a21oi_1 _3268_ (.A1(net149),
    .A2(_2239_),
    .Y(_2299_),
    .B1(_2289_));
 sg13g2_nor2_1 _3269_ (.A(_2151_),
    .B(_2299_),
    .Y(_2308_));
 sg13g2_nor2_1 _3270_ (.A(_2075_),
    .B(_2308_),
    .Y(_2317_));
 sg13g2_nand2_1 _3271_ (.Y(_2325_),
    .A(_1729_),
    .B(_2317_));
 sg13g2_buf_1 _3272_ (.A(\mem_addr[7] ),
    .X(_2332_));
 sg13g2_inv_1 _3273_ (.Y(_2341_),
    .A(_2332_));
 sg13g2_buf_2 _3274_ (.A(_2341_),
    .X(_2351_));
 sg13g2_buf_2 _3275_ (.A(net175),
    .X(_2360_));
 sg13g2_nand2_1 _3276_ (.Y(_2369_),
    .A(_2325_),
    .B(net147));
 sg13g2_nor2_1 _3277_ (.A(net209),
    .B(_2341_),
    .Y(_2372_));
 sg13g2_buf_2 _3278_ (.A(_2372_),
    .X(_2373_));
 sg13g2_inv_1 _3279_ (.Y(_2374_),
    .A(_2373_));
 sg13g2_buf_1 _3280_ (.A(_2374_),
    .X(_2375_));
 sg13g2_buf_2 _3281_ (.A(_0036_),
    .X(_2376_));
 sg13g2_nand2_1 _3282_ (.Y(_2377_),
    .A(net205),
    .B(_2376_));
 sg13g2_inv_1 _3283_ (.Y(_2378_),
    .A(_2377_));
 sg13g2_nand2_2 _3284_ (.Y(_2379_),
    .A(net178),
    .B(net201));
 sg13g2_nor3_1 _3285_ (.A(_2378_),
    .B(net64),
    .C(_2379_),
    .Y(_2380_));
 sg13g2_nor2_1 _3286_ (.A(_1053_),
    .B(net182),
    .Y(_2381_));
 sg13g2_buf_1 _3287_ (.A(_2381_),
    .X(_2382_));
 sg13g2_inv_2 _3288_ (.Y(_2383_),
    .A(net104));
 sg13g2_buf_2 _3289_ (.A(net62),
    .X(_2384_));
 sg13g2_nand2_1 _3290_ (.Y(_2385_),
    .A(_0812_),
    .B(net204));
 sg13g2_buf_2 _3291_ (.A(_2385_),
    .X(_2386_));
 sg13g2_inv_2 _3292_ (.Y(_2387_),
    .A(net146));
 sg13g2_nor2_1 _3293_ (.A(net103),
    .B(_2203_),
    .Y(_2388_));
 sg13g2_nor2_1 _3294_ (.A(net31),
    .B(_2388_),
    .Y(_2389_));
 sg13g2_buf_1 _3295_ (.A(_1326_),
    .X(_2390_));
 sg13g2_nor2_1 _3296_ (.A(_0889_),
    .B(net190),
    .Y(_2391_));
 sg13g2_buf_4 _3297_ (.X(_2392_),
    .A(_2391_));
 sg13g2_nor2_1 _3298_ (.A(net146),
    .B(_2392_),
    .Y(_2393_));
 sg13g2_nor2_2 _3299_ (.A(_2203_),
    .B(_2393_),
    .Y(_2394_));
 sg13g2_nor2_1 _3300_ (.A(net145),
    .B(_2394_),
    .Y(_2395_));
 sg13g2_nor4_1 _3301_ (.A(net63),
    .B(_2380_),
    .C(_2389_),
    .D(_2395_),
    .Y(_2396_));
 sg13g2_inv_1 _3302_ (.Y(_2397_),
    .A(_0038_));
 sg13g2_nor2_1 _3303_ (.A(net208),
    .B(_2397_),
    .Y(_2398_));
 sg13g2_inv_2 _3304_ (.Y(_2399_),
    .A(_2398_));
 sg13g2_nand2_1 _3305_ (.Y(_2400_),
    .A(_2097_),
    .B(net144));
 sg13g2_buf_8 _3306_ (.A(net184),
    .X(_2401_));
 sg13g2_buf_1 _3307_ (.A(net143),
    .X(_2402_));
 sg13g2_nand2_1 _3308_ (.Y(_2403_),
    .A(_2400_),
    .B(net102));
 sg13g2_nor2_1 _3309_ (.A(_1042_),
    .B(net210),
    .Y(_2404_));
 sg13g2_buf_2 _3310_ (.A(_2404_),
    .X(_2405_));
 sg13g2_inv_1 _3311_ (.Y(_2406_),
    .A(_2405_));
 sg13g2_buf_1 _3312_ (.A(_2406_),
    .X(_2407_));
 sg13g2_buf_2 _3313_ (.A(net101),
    .X(_2408_));
 sg13g2_a21o_1 _3314_ (.A2(_1238_),
    .A1(_2403_),
    .B1(net61),
    .X(_2409_));
 sg13g2_nor2_1 _3315_ (.A(_0725_),
    .B(_0878_),
    .Y(_2410_));
 sg13g2_buf_2 _3316_ (.A(_2410_),
    .X(_2411_));
 sg13g2_nand2_1 _3317_ (.Y(_2412_),
    .A(_2411_),
    .B(net189));
 sg13g2_buf_1 _3318_ (.A(_2412_),
    .X(_2413_));
 sg13g2_nand2_1 _3319_ (.Y(_2414_),
    .A(net100),
    .B(_2020_));
 sg13g2_buf_1 _3320_ (.A(_0856_),
    .X(_2415_));
 sg13g2_buf_2 _3321_ (.A(net60),
    .X(_2416_));
 sg13g2_buf_1 _3322_ (.A(net202),
    .X(_2417_));
 sg13g2_buf_1 _3323_ (.A(_2417_),
    .X(_2418_));
 sg13g2_buf_1 _3324_ (.A(net142),
    .X(_2419_));
 sg13g2_nand3_1 _3325_ (.B(net30),
    .C(_2419_),
    .A(_2414_),
    .Y(_2420_));
 sg13g2_nand3_1 _3326_ (.B(_2409_),
    .C(_2420_),
    .A(_2396_),
    .Y(_2421_));
 sg13g2_nand2_1 _3327_ (.Y(_2422_),
    .A(_2369_),
    .B(_2421_));
 sg13g2_buf_4 _3328_ (.X(_2423_),
    .A(\mem_addr[8] ));
 sg13g2_buf_1 _3329_ (.A(_2423_),
    .X(_2424_));
 sg13g2_nand2_1 _3330_ (.Y(_2425_),
    .A(_2422_),
    .B(net200));
 sg13g2_buf_1 _3331_ (.A(net181),
    .X(_2426_));
 sg13g2_nand4_1 _3332_ (.B(_1911_),
    .C(net152),
    .A(_0801_),
    .Y(_2427_),
    .D(net141));
 sg13g2_buf_1 _3333_ (.A(_2427_),
    .X(_2428_));
 sg13g2_nor2_2 _3334_ (.A(_2386_),
    .B(_1859_),
    .Y(_2429_));
 sg13g2_inv_2 _3335_ (.Y(_2430_),
    .A(_2429_));
 sg13g2_a21oi_1 _3336_ (.A1(_2428_),
    .A2(_2430_),
    .Y(_2431_),
    .B1(net101));
 sg13g2_nand2_1 _3337_ (.Y(_2432_),
    .A(net190),
    .B(_1205_));
 sg13g2_buf_2 _3338_ (.A(_2432_),
    .X(_2433_));
 sg13g2_nand2_1 _3339_ (.Y(_2434_),
    .A(net189),
    .B(net183));
 sg13g2_buf_1 _3340_ (.A(_2434_),
    .X(_2435_));
 sg13g2_nand2_2 _3341_ (.Y(_2436_),
    .A(_2433_),
    .B(net98));
 sg13g2_buf_2 _3342_ (.A(net184),
    .X(_2437_));
 sg13g2_nand3_1 _3343_ (.B(net140),
    .C(net141),
    .A(_2436_),
    .Y(_2438_));
 sg13g2_nor2_1 _3344_ (.A(_0867_),
    .B(net181),
    .Y(_2439_));
 sg13g2_buf_4 _3345_ (.X(_2440_),
    .A(_2439_));
 sg13g2_nor2_2 _3346_ (.A(_0812_),
    .B(_1205_),
    .Y(_2441_));
 sg13g2_buf_2 _3347_ (.A(_2441_),
    .X(_2442_));
 sg13g2_nand2_1 _3348_ (.Y(_2443_),
    .A(_2440_),
    .B(_2442_));
 sg13g2_buf_2 _3349_ (.A(_2443_),
    .X(_2444_));
 sg13g2_buf_1 _3350_ (.A(_1326_),
    .X(_2445_));
 sg13g2_a21oi_1 _3351_ (.A1(_2438_),
    .A2(_2444_),
    .Y(_2446_),
    .B1(net138));
 sg13g2_nor2_1 _3352_ (.A(_2431_),
    .B(_2446_),
    .Y(_2447_));
 sg13g2_nand2_1 _3353_ (.Y(_2448_),
    .A(net183),
    .B(_0038_));
 sg13g2_buf_1 _3354_ (.A(_2448_),
    .X(_2449_));
 sg13g2_nor2_2 _3355_ (.A(_1009_),
    .B(net97),
    .Y(_2450_));
 sg13g2_nand2_1 _3356_ (.Y(_2451_),
    .A(net188),
    .B(net207));
 sg13g2_buf_1 _3357_ (.A(_2451_),
    .X(_2452_));
 sg13g2_nor2_2 _3358_ (.A(_2433_),
    .B(net96),
    .Y(_2453_));
 sg13g2_nor2_1 _3359_ (.A(_2450_),
    .B(_2453_),
    .Y(_2454_));
 sg13g2_inv_1 _3360_ (.Y(_2455_),
    .A(_2393_));
 sg13g2_a21oi_1 _3361_ (.A1(_2454_),
    .A2(_2455_),
    .Y(_2456_),
    .B1(net64));
 sg13g2_inv_2 _3362_ (.Y(_2457_),
    .A(_0965_));
 sg13g2_buf_1 _3363_ (.A(_2457_),
    .X(_2458_));
 sg13g2_nand3_1 _3364_ (.B(_2458_),
    .C(net104),
    .A(_1805_),
    .Y(_2459_));
 sg13g2_inv_2 _3365_ (.Y(_2460_),
    .A(_1369_));
 sg13g2_nand2_2 _3366_ (.Y(_2461_),
    .A(net104),
    .B(_0845_));
 sg13g2_nor2_2 _3367_ (.A(net100),
    .B(_2461_),
    .Y(_2462_));
 sg13g2_nor2_1 _3368_ (.A(_2460_),
    .B(_2462_),
    .Y(_2463_));
 sg13g2_nand2_1 _3369_ (.Y(_2464_),
    .A(_2459_),
    .B(_2463_));
 sg13g2_nor2_1 _3370_ (.A(_2456_),
    .B(_2464_),
    .Y(_2465_));
 sg13g2_nand2_1 _3371_ (.Y(_2466_),
    .A(_2447_),
    .B(_2465_));
 sg13g2_nor2_2 _3372_ (.A(net152),
    .B(net156),
    .Y(_2467_));
 sg13g2_xnor2_1 _3373_ (.Y(_2468_),
    .A(net208),
    .B(net186));
 sg13g2_buf_2 _3374_ (.A(_2468_),
    .X(_2469_));
 sg13g2_nor2_2 _3375_ (.A(_2452_),
    .B(_2469_),
    .Y(_2470_));
 sg13g2_nor2_1 _3376_ (.A(_2467_),
    .B(_2470_),
    .Y(_2471_));
 sg13g2_nor2_1 _3377_ (.A(net62),
    .B(_2471_),
    .Y(_2472_));
 sg13g2_nand2_1 _3378_ (.Y(_2473_),
    .A(net190),
    .B(net207));
 sg13g2_nand2_1 _3379_ (.Y(_2474_),
    .A(_2473_),
    .B(net188));
 sg13g2_buf_1 _3380_ (.A(_2474_),
    .X(_2475_));
 sg13g2_nand2_1 _3381_ (.Y(_2476_),
    .A(_1129_),
    .B(_0725_));
 sg13g2_buf_2 _3382_ (.A(_2476_),
    .X(_2477_));
 sg13g2_nand2_2 _3383_ (.Y(_2478_),
    .A(net137),
    .B(net187));
 sg13g2_nand3_1 _3384_ (.B(_2478_),
    .C(_1085_),
    .A(net59),
    .Y(_2479_));
 sg13g2_buf_2 _3385_ (.A(_2460_),
    .X(_2480_));
 sg13g2_nor2_1 _3386_ (.A(_1042_),
    .B(_2376_),
    .Y(_2481_));
 sg13g2_buf_2 _3387_ (.A(_2481_),
    .X(_2482_));
 sg13g2_nand3_1 _3388_ (.B(net150),
    .C(_2482_),
    .A(_0987_),
    .Y(_2483_));
 sg13g2_nand3_1 _3389_ (.B(net173),
    .C(_2483_),
    .A(_2479_),
    .Y(_2484_));
 sg13g2_nor2_1 _3390_ (.A(_2472_),
    .B(_2484_),
    .Y(_2485_));
 sg13g2_nand2_1 _3391_ (.Y(_2486_),
    .A(_0965_),
    .B(net183));
 sg13g2_buf_8 _3392_ (.A(_2486_),
    .X(_2487_));
 sg13g2_inv_1 _3393_ (.Y(_2488_),
    .A(_1478_));
 sg13g2_nand2_1 _3394_ (.Y(_2489_),
    .A(net94),
    .B(_2488_));
 sg13g2_buf_8 _3395_ (.A(net157),
    .X(_2490_));
 sg13g2_buf_8 _3396_ (.A(net93),
    .X(_2491_));
 sg13g2_nand2_1 _3397_ (.Y(_2492_),
    .A(_2489_),
    .B(net58));
 sg13g2_nor2_1 _3398_ (.A(net204),
    .B(_0736_),
    .Y(_2493_));
 sg13g2_buf_2 _3399_ (.A(_2493_),
    .X(_2494_));
 sg13g2_buf_1 _3400_ (.A(net187),
    .X(_2495_));
 sg13g2_nand2_2 _3401_ (.Y(_2496_),
    .A(_2494_),
    .B(net136));
 sg13g2_a21o_1 _3402_ (.A2(_2496_),
    .A1(_2492_),
    .B1(net138),
    .X(_2497_));
 sg13g2_nand2_1 _3403_ (.Y(_2498_),
    .A(_2485_),
    .B(_2497_));
 sg13g2_nand2_1 _3404_ (.Y(_2499_),
    .A(_2466_),
    .B(_2498_));
 sg13g2_nand2_1 _3405_ (.Y(_2500_),
    .A(_2499_),
    .B(net147));
 sg13g2_a21oi_2 _3406_ (.B1(net190),
    .Y(_2501_),
    .A2(net185),
    .A1(net186));
 sg13g2_nand2_1 _3407_ (.Y(_2502_),
    .A(_2501_),
    .B(_2457_));
 sg13g2_buf_1 _3408_ (.A(_2502_),
    .X(_2503_));
 sg13g2_nand2_1 _3409_ (.Y(_2504_),
    .A(net57),
    .B(net100));
 sg13g2_buf_1 _3410_ (.A(net154),
    .X(_2505_));
 sg13g2_buf_1 _3411_ (.A(net92),
    .X(_2506_));
 sg13g2_nand2_1 _3412_ (.Y(_2507_),
    .A(_2504_),
    .B(net56));
 sg13g2_buf_1 _3413_ (.A(net182),
    .X(_2508_));
 sg13g2_buf_1 _3414_ (.A(net135),
    .X(_2509_));
 sg13g2_buf_1 _3415_ (.A(net91),
    .X(_2510_));
 sg13g2_inv_1 _3416_ (.Y(_2511_),
    .A(_1838_));
 sg13g2_buf_1 _3417_ (.A(_2511_),
    .X(_2512_));
 sg13g2_buf_2 _3418_ (.A(_2473_),
    .X(_2513_));
 sg13g2_nand2_1 _3419_ (.Y(_2514_),
    .A(net29),
    .B(net90));
 sg13g2_nand3_1 _3420_ (.B(net55),
    .C(_2514_),
    .A(_2507_),
    .Y(_2515_));
 sg13g2_buf_1 _3421_ (.A(net210),
    .X(_2516_));
 sg13g2_buf_1 _3422_ (.A(_2516_),
    .X(_2517_));
 sg13g2_buf_1 _3423_ (.A(net135),
    .X(_2518_));
 sg13g2_nor2_2 _3424_ (.A(net187),
    .B(_1911_),
    .Y(_2519_));
 sg13g2_inv_2 _3425_ (.Y(_2520_),
    .A(_1031_));
 sg13g2_nor3_1 _3426_ (.A(net89),
    .B(_2519_),
    .C(_2520_),
    .Y(_2521_));
 sg13g2_nor2_1 _3427_ (.A(net172),
    .B(_2521_),
    .Y(_2522_));
 sg13g2_nand2_1 _3428_ (.Y(_2523_),
    .A(_2515_),
    .B(_2522_));
 sg13g2_nand2_2 _3429_ (.Y(_2524_),
    .A(_0779_),
    .B(_0878_));
 sg13g2_nand2_2 _3430_ (.Y(_2525_),
    .A(_2524_),
    .B(net201));
 sg13g2_nand2_2 _3431_ (.Y(_2526_),
    .A(_2411_),
    .B(net205));
 sg13g2_nand2_1 _3432_ (.Y(_2527_),
    .A(_1347_),
    .B(_2386_));
 sg13g2_a21oi_1 _3433_ (.A1(_2525_),
    .A2(_2526_),
    .Y(_2528_),
    .B1(_2527_));
 sg13g2_a21oi_2 _3434_ (.B1(net181),
    .Y(_2529_),
    .A2(net153),
    .A1(net206));
 sg13g2_nand2_2 _3435_ (.Y(_2530_),
    .A(_2529_),
    .B(_2512_));
 sg13g2_nand3_1 _3436_ (.B(net208),
    .C(net186),
    .A(_0812_),
    .Y(_2531_));
 sg13g2_buf_2 _3437_ (.A(_2531_),
    .X(_2532_));
 sg13g2_buf_1 _3438_ (.A(_1096_),
    .X(_2533_));
 sg13g2_a21oi_1 _3439_ (.A1(_2530_),
    .A2(_2532_),
    .Y(_2534_),
    .B1(net54));
 sg13g2_nor3_1 _3440_ (.A(_2375_),
    .B(_2528_),
    .C(_2534_),
    .Y(_2535_));
 sg13g2_inv_1 _3441_ (.Y(_2536_),
    .A(_1958_));
 sg13g2_nor2_2 _3442_ (.A(net157),
    .B(_2379_),
    .Y(_2537_));
 sg13g2_nand2_1 _3443_ (.Y(_2538_),
    .A(_2537_),
    .B(net95));
 sg13g2_nor2_1 _3444_ (.A(net202),
    .B(_2429_),
    .Y(_2539_));
 sg13g2_nor2_1 _3445_ (.A(net96),
    .B(_1609_),
    .Y(_2540_));
 sg13g2_inv_1 _3446_ (.Y(_2541_),
    .A(_2540_));
 sg13g2_nand2_1 _3447_ (.Y(_2542_),
    .A(_2539_),
    .B(_2541_));
 sg13g2_buf_2 _3448_ (.A(net210),
    .X(_2543_));
 sg13g2_buf_1 _3449_ (.A(_2543_),
    .X(_2544_));
 sg13g2_nand2_1 _3450_ (.Y(_2545_),
    .A(_2542_),
    .B(net171));
 sg13g2_a21oi_1 _3451_ (.A1(_2536_),
    .A2(_2538_),
    .Y(_2546_),
    .B1(_2545_));
 sg13g2_nand2_1 _3452_ (.Y(_2547_),
    .A(_2221_),
    .B(net176));
 sg13g2_inv_1 _3453_ (.Y(_2548_),
    .A(_2547_));
 sg13g2_a21oi_1 _3454_ (.A1(net183),
    .A2(net186),
    .Y(_2549_),
    .B1(net205));
 sg13g2_buf_4 _3455_ (.X(_2550_),
    .A(_2549_));
 sg13g2_nand2_1 _3456_ (.Y(_2551_),
    .A(_2550_),
    .B(net100));
 sg13g2_buf_2 _3457_ (.A(_2405_),
    .X(_2552_));
 sg13g2_nand3_1 _3458_ (.B(_2551_),
    .C(net134),
    .A(_2548_),
    .Y(_2553_));
 sg13g2_buf_1 _3459_ (.A(net178),
    .X(_2554_));
 sg13g2_a21oi_1 _3460_ (.A1(net133),
    .A2(net98),
    .Y(_2555_),
    .B1(_2461_));
 sg13g2_inv_1 _3461_ (.Y(_2556_),
    .A(_2555_));
 sg13g2_buf_2 _3462_ (.A(_2332_),
    .X(_2557_));
 sg13g2_nand2_1 _3463_ (.Y(_2558_),
    .A(net209),
    .B(net197));
 sg13g2_inv_2 _3464_ (.Y(_2559_),
    .A(_2558_));
 sg13g2_nand3_1 _3465_ (.B(_2556_),
    .C(_2559_),
    .A(_2553_),
    .Y(_2560_));
 sg13g2_nor2_1 _3466_ (.A(_2546_),
    .B(_2560_),
    .Y(_2561_));
 sg13g2_a21oi_1 _3467_ (.A1(_2523_),
    .A2(_2535_),
    .Y(_2562_),
    .B1(_2561_));
 sg13g2_nand2_1 _3468_ (.Y(_2563_),
    .A(_2500_),
    .B(_2562_));
 sg13g2_inv_2 _3469_ (.Y(_2564_),
    .A(_2423_));
 sg13g2_buf_1 _3470_ (.A(_2564_),
    .X(_2565_));
 sg13g2_buf_2 _3471_ (.A(net170),
    .X(_2566_));
 sg13g2_nand2_1 _3472_ (.Y(_2567_),
    .A(_2563_),
    .B(net132));
 sg13g2_buf_2 _3473_ (.A(_1085_),
    .X(_2568_));
 sg13g2_buf_2 _3474_ (.A(net88),
    .X(_2569_));
 sg13g2_nor2_1 _3475_ (.A(net188),
    .B(_2440_),
    .Y(_2570_));
 sg13g2_buf_2 _3476_ (.A(_2570_),
    .X(_2571_));
 sg13g2_inv_1 _3477_ (.Y(_2572_),
    .A(_2571_));
 sg13g2_nor2_2 _3478_ (.A(_0965_),
    .B(_2097_),
    .Y(_2573_));
 sg13g2_nor2_1 _3479_ (.A(_2572_),
    .B(_2573_),
    .Y(_2574_));
 sg13g2_inv_1 _3480_ (.Y(_2575_),
    .A(net97));
 sg13g2_nor2_1 _3481_ (.A(_0867_),
    .B(_0965_),
    .Y(_2576_));
 sg13g2_buf_2 _3482_ (.A(_2576_),
    .X(_2577_));
 sg13g2_o21ai_1 _3483_ (.B1(net60),
    .Y(_2578_),
    .A1(_2575_),
    .A2(_2577_));
 sg13g2_buf_2 _3484_ (.A(_2578_),
    .X(_2579_));
 sg13g2_nand2b_1 _3485_ (.Y(_2580_),
    .B(_2579_),
    .A_N(_2574_));
 sg13g2_nand2_1 _3486_ (.Y(_2581_),
    .A(net90),
    .B(net137));
 sg13g2_buf_2 _3487_ (.A(_2581_),
    .X(_2582_));
 sg13g2_buf_1 _3488_ (.A(_0801_),
    .X(_2583_));
 sg13g2_nor2_1 _3489_ (.A(_0790_),
    .B(_0900_),
    .Y(_2584_));
 sg13g2_nor2_2 _3490_ (.A(_2490_),
    .B(_2584_),
    .Y(_2585_));
 sg13g2_a22oi_1 _3491_ (.Y(_2586_),
    .B1(net52),
    .B2(_2585_),
    .A2(net139),
    .A1(_2582_));
 sg13g2_nor2_1 _3492_ (.A(net145),
    .B(_2586_),
    .Y(_2587_));
 sg13g2_a21oi_1 _3493_ (.A1(net53),
    .A2(_2580_),
    .Y(_2588_),
    .B1(_2587_));
 sg13g2_buf_2 _3494_ (.A(net111),
    .X(_2589_));
 sg13g2_nand2_2 _3495_ (.Y(_2590_),
    .A(_2273_),
    .B(net51));
 sg13g2_nand2_1 _3496_ (.Y(_2591_),
    .A(net103),
    .B(_2411_));
 sg13g2_nand2_1 _3497_ (.Y(_2592_),
    .A(_2590_),
    .B(_2591_));
 sg13g2_buf_1 _3498_ (.A(net104),
    .X(_2593_));
 sg13g2_nand2_1 _3499_ (.Y(_2594_),
    .A(_2592_),
    .B(net50));
 sg13g2_buf_2 _3500_ (.A(net203),
    .X(_2595_));
 sg13g2_buf_1 _3501_ (.A(net169),
    .X(_2596_));
 sg13g2_nand2_2 _3502_ (.Y(_2597_),
    .A(net197),
    .B(_2423_));
 sg13g2_inv_2 _3503_ (.Y(_2598_),
    .A(_2597_));
 sg13g2_nand3_1 _3504_ (.B(net131),
    .C(_2598_),
    .A(_2594_),
    .Y(_2599_));
 sg13g2_buf_2 _3505_ (.A(net198),
    .X(_2600_));
 sg13g2_buf_1 _3506_ (.A(net168),
    .X(_2601_));
 sg13g2_nor2_1 _3507_ (.A(net143),
    .B(net98),
    .Y(_2602_));
 sg13g2_buf_1 _3508_ (.A(_1911_),
    .X(_2603_));
 sg13g2_nand2_1 _3509_ (.Y(_2604_),
    .A(_1489_),
    .B(net87));
 sg13g2_nand2_2 _3510_ (.Y(_2605_),
    .A(_2411_),
    .B(net93));
 sg13g2_nand3_1 _3511_ (.B(_2508_),
    .C(_2605_),
    .A(_2604_),
    .Y(_2606_));
 sg13g2_nor3_1 _3512_ (.A(net130),
    .B(_2602_),
    .C(_2606_),
    .Y(_2607_));
 sg13g2_nor2_1 _3513_ (.A(_2599_),
    .B(_2607_),
    .Y(_2608_));
 sg13g2_buf_2 _3514_ (.A(\memory_1.mem_addr[9] ),
    .X(_2609_));
 sg13g2_buf_1 _3515_ (.A(_2609_),
    .X(_2610_));
 sg13g2_a21oi_1 _3516_ (.A1(_2588_),
    .A2(_2608_),
    .Y(_2611_),
    .B1(net196));
 sg13g2_nand3_1 _3517_ (.B(_2567_),
    .C(_2611_),
    .A(_2425_),
    .Y(_2612_));
 sg13g2_a21oi_1 _3518_ (.A1(net155),
    .A2(net153),
    .Y(_2613_),
    .B1(_1609_));
 sg13g2_nand2_1 _3519_ (.Y(_2614_),
    .A(_2613_),
    .B(_2571_));
 sg13g2_buf_2 _3520_ (.A(net104),
    .X(_2615_));
 sg13g2_nor2_2 _3521_ (.A(_1009_),
    .B(_2469_),
    .Y(_2616_));
 sg13g2_inv_1 _3522_ (.Y(_2617_),
    .A(_2616_));
 sg13g2_nand3_1 _3523_ (.B(net49),
    .C(_2617_),
    .A(_2614_),
    .Y(_2618_));
 sg13g2_buf_2 _3524_ (.A(net203),
    .X(_2619_));
 sg13g2_nand2_1 _3525_ (.Y(_2620_),
    .A(_2618_),
    .B(net167));
 sg13g2_nand2_1 _3526_ (.Y(_2621_),
    .A(_2577_),
    .B(net178));
 sg13g2_buf_2 _3527_ (.A(_2621_),
    .X(_2622_));
 sg13g2_nand2_1 _3528_ (.Y(_2623_),
    .A(net137),
    .B(net188));
 sg13g2_inv_1 _3529_ (.Y(_2624_),
    .A(_2623_));
 sg13g2_nand2_2 _3530_ (.Y(_2625_),
    .A(_2622_),
    .B(_2624_));
 sg13g2_buf_1 _3531_ (.A(_2405_),
    .X(_2626_));
 sg13g2_nand2_1 _3532_ (.Y(_2627_),
    .A(_1653_),
    .B(net176));
 sg13g2_buf_1 _3533_ (.A(_2627_),
    .X(_2628_));
 sg13g2_inv_1 _3534_ (.Y(_2629_),
    .A(net86));
 sg13g2_nand3_1 _3535_ (.B(net129),
    .C(_2629_),
    .A(_2625_),
    .Y(_2630_));
 sg13g2_nor2b_1 _3536_ (.A(_2620_),
    .B_N(_2630_),
    .Y(_2631_));
 sg13g2_nor2_1 _3537_ (.A(_0932_),
    .B(net207),
    .Y(_2632_));
 sg13g2_buf_4 _3538_ (.X(_2633_),
    .A(_2632_));
 sg13g2_inv_2 _3539_ (.Y(_2634_),
    .A(_2633_));
 sg13g2_nor2_2 _3540_ (.A(net148),
    .B(_2634_),
    .Y(_2635_));
 sg13g2_nor2_1 _3541_ (.A(_0932_),
    .B(net181),
    .Y(_2636_));
 sg13g2_nand2_2 _3542_ (.Y(_2637_),
    .A(_2636_),
    .B(_2441_));
 sg13g2_inv_1 _3543_ (.Y(_2638_),
    .A(_2637_));
 sg13g2_nor2_1 _3544_ (.A(_2635_),
    .B(_2638_),
    .Y(_2639_));
 sg13g2_inv_1 _3545_ (.Y(_2640_),
    .A(_2639_));
 sg13g2_nand2_2 _3546_ (.Y(_2641_),
    .A(net184),
    .B(_1053_));
 sg13g2_nand2_2 _3547_ (.Y(_2642_),
    .A(_2637_),
    .B(net202));
 sg13g2_nand2_1 _3548_ (.Y(_2643_),
    .A(_2642_),
    .B(net199));
 sg13g2_o21ai_1 _3549_ (.B1(_2643_),
    .Y(_2644_),
    .A1(_2641_),
    .A2(_2613_));
 sg13g2_o21ai_1 _3550_ (.B1(_2644_),
    .Y(_2645_),
    .A1(_2419_),
    .A2(_2640_));
 sg13g2_buf_1 _3551_ (.A(net197),
    .X(_2646_));
 sg13g2_a21oi_1 _3552_ (.A1(_2631_),
    .A2(_2645_),
    .Y(_2647_),
    .B1(net166));
 sg13g2_nor2_1 _3553_ (.A(_0998_),
    .B(_2411_),
    .Y(_2648_));
 sg13g2_buf_1 _3554_ (.A(_2648_),
    .X(_2649_));
 sg13g2_nand2_1 _3555_ (.Y(_2650_),
    .A(net85),
    .B(_2634_));
 sg13g2_nand2_1 _3556_ (.Y(_2651_),
    .A(net86),
    .B(_2433_));
 sg13g2_nand3_1 _3557_ (.B(_2651_),
    .C(net199),
    .A(_2650_),
    .Y(_2652_));
 sg13g2_buf_1 _3558_ (.A(net179),
    .X(_2653_));
 sg13g2_buf_1 _3559_ (.A(net128),
    .X(_2654_));
 sg13g2_nand2_1 _3560_ (.Y(_2655_),
    .A(_2652_),
    .B(_2654_));
 sg13g2_nand2_1 _3561_ (.Y(_2656_),
    .A(_2622_),
    .B(net143));
 sg13g2_inv_1 _3562_ (.Y(_2657_),
    .A(_2656_));
 sg13g2_nor3_1 _3563_ (.A(net168),
    .B(_2392_),
    .C(_2657_),
    .Y(_2658_));
 sg13g2_nand2_2 _3564_ (.Y(_2659_),
    .A(net155),
    .B(net201));
 sg13g2_inv_1 _3565_ (.Y(_2660_),
    .A(net96));
 sg13g2_nor2_1 _3566_ (.A(_1751_),
    .B(_2660_),
    .Y(_2661_));
 sg13g2_o21ai_1 _3567_ (.B1(_2661_),
    .Y(_2662_),
    .A1(_2641_),
    .A2(_2659_));
 sg13g2_o21ai_1 _3568_ (.B1(_2662_),
    .Y(_2663_),
    .A1(_2655_),
    .A2(_2658_));
 sg13g2_buf_1 _3569_ (.A(net173),
    .X(_2664_));
 sg13g2_buf_2 _3570_ (.A(net127),
    .X(_2665_));
 sg13g2_nand2_1 _3571_ (.Y(_2666_),
    .A(_2663_),
    .B(net83));
 sg13g2_nand2_1 _3572_ (.Y(_2667_),
    .A(_2647_),
    .B(_2666_));
 sg13g2_nand2_1 _3573_ (.Y(_2668_),
    .A(_1129_),
    .B(net204));
 sg13g2_buf_8 _3574_ (.A(_2668_),
    .X(_2669_));
 sg13g2_nand2_1 _3575_ (.Y(_2670_),
    .A(net126),
    .B(_0746_));
 sg13g2_buf_2 _3576_ (.A(_2670_),
    .X(_2671_));
 sg13g2_nand3_1 _3577_ (.B(net183),
    .C(_1249_),
    .A(_1588_),
    .Y(_2672_));
 sg13g2_buf_1 _3578_ (.A(_2672_),
    .X(_2673_));
 sg13g2_nand2_1 _3579_ (.Y(_2674_),
    .A(_2671_),
    .B(net82));
 sg13g2_nand2_1 _3580_ (.Y(_2675_),
    .A(net181),
    .B(_0038_));
 sg13g2_nand2_1 _3581_ (.Y(_2676_),
    .A(_0932_),
    .B(net185));
 sg13g2_nand2_2 _3582_ (.Y(_2677_),
    .A(_2675_),
    .B(_2676_));
 sg13g2_nor2_2 _3583_ (.A(net111),
    .B(_2677_),
    .Y(_2678_));
 sg13g2_nor2_1 _3584_ (.A(net99),
    .B(_2678_),
    .Y(_2679_));
 sg13g2_buf_1 _3585_ (.A(net109),
    .X(_2680_));
 sg13g2_nand2_1 _3586_ (.Y(_2681_),
    .A(net48),
    .B(net206));
 sg13g2_buf_1 _3587_ (.A(_2524_),
    .X(_2682_));
 sg13g2_nand2_1 _3588_ (.Y(_2683_),
    .A(net125),
    .B(net126));
 sg13g2_buf_1 _3589_ (.A(_2683_),
    .X(_2684_));
 sg13g2_nand2b_1 _3590_ (.Y(_2685_),
    .B(net47),
    .A_N(_2681_));
 sg13g2_nor2_2 _3591_ (.A(_2376_),
    .B(net182),
    .Y(_2686_));
 sg13g2_inv_1 _3592_ (.Y(_2687_),
    .A(_2686_));
 sg13g2_buf_2 _3593_ (.A(net180),
    .X(_2688_));
 sg13g2_buf_2 _3594_ (.A(net124),
    .X(_2689_));
 sg13g2_nand2_1 _3595_ (.Y(_2690_),
    .A(_2332_),
    .B(_0033_));
 sg13g2_inv_1 _3596_ (.Y(_2691_),
    .A(_2690_));
 sg13g2_nand3_1 _3597_ (.B(net81),
    .C(_2691_),
    .A(_2687_),
    .Y(_2692_));
 sg13g2_a221oi_1 _3598_ (.B2(_2685_),
    .C1(_2692_),
    .B1(_2679_),
    .A1(net99),
    .Y(_2693_),
    .A2(_2674_));
 sg13g2_nor2_1 _3599_ (.A(net170),
    .B(_2693_),
    .Y(_2694_));
 sg13g2_inv_1 _3600_ (.Y(_2695_),
    .A(_2609_));
 sg13g2_buf_1 _3601_ (.A(net195),
    .X(_2696_));
 sg13g2_a21oi_1 _3602_ (.A1(_2667_),
    .A2(_2694_),
    .Y(_2697_),
    .B1(net165));
 sg13g2_buf_1 _3603_ (.A(net173),
    .X(_2698_));
 sg13g2_buf_1 _3604_ (.A(net123),
    .X(_2699_));
 sg13g2_a21oi_1 _3605_ (.A1(_1238_),
    .A2(_2221_),
    .Y(_2700_),
    .B1(net145));
 sg13g2_inv_2 _3606_ (.Y(_2701_),
    .A(_2482_));
 sg13g2_nor2_1 _3607_ (.A(net87),
    .B(_2701_),
    .Y(_2702_));
 sg13g2_inv_1 _3608_ (.Y(_2703_),
    .A(_2702_));
 sg13g2_buf_1 _3609_ (.A(_1413_),
    .X(_2704_));
 sg13g2_nand2_1 _3610_ (.Y(_2705_),
    .A(net122),
    .B(net86));
 sg13g2_nand3_1 _3611_ (.B(net106),
    .C(net129),
    .A(_2705_),
    .Y(_2706_));
 sg13g2_o21ai_1 _3612_ (.B1(_2706_),
    .Y(_2707_),
    .A1(net81),
    .A2(_2703_));
 sg13g2_nor3_1 _3613_ (.A(net80),
    .B(_2700_),
    .C(_2707_),
    .Y(_2708_));
 sg13g2_nand2_2 _3614_ (.Y(_2709_),
    .A(_2440_),
    .B(net189));
 sg13g2_nand2_2 _3615_ (.Y(_2710_),
    .A(_2709_),
    .B(_2672_));
 sg13g2_buf_1 _3616_ (.A(net154),
    .X(_2711_));
 sg13g2_nand2_2 _3617_ (.Y(_2712_),
    .A(_2710_),
    .B(net79));
 sg13g2_nor2_1 _3618_ (.A(net187),
    .B(_0910_),
    .Y(_2713_));
 sg13g2_nor2_1 _3619_ (.A(_1740_),
    .B(_2713_),
    .Y(_2714_));
 sg13g2_buf_2 _3620_ (.A(_2714_),
    .X(_2715_));
 sg13g2_buf_1 _3621_ (.A(net124),
    .X(_2716_));
 sg13g2_a21oi_1 _3622_ (.A1(_2712_),
    .A2(_2715_),
    .Y(_2717_),
    .B1(net78));
 sg13g2_nand3_1 _3623_ (.B(net93),
    .C(_2426_),
    .A(_2469_),
    .Y(_2718_));
 sg13g2_buf_2 _3624_ (.A(_2718_),
    .X(_2719_));
 sg13g2_nand3_1 _3625_ (.B(net84),
    .C(_2705_),
    .A(_2719_),
    .Y(_2720_));
 sg13g2_nand2_1 _3626_ (.Y(_2721_),
    .A(_2717_),
    .B(_2720_));
 sg13g2_nand2_1 _3627_ (.Y(_2722_),
    .A(_2489_),
    .B(net102));
 sg13g2_nor2_2 _3628_ (.A(net106),
    .B(_2634_),
    .Y(_2723_));
 sg13g2_nor2_1 _3629_ (.A(net128),
    .B(_2723_),
    .Y(_2724_));
 sg13g2_nand2_1 _3630_ (.Y(_2725_),
    .A(_2722_),
    .B(_2724_));
 sg13g2_nor2_1 _3631_ (.A(net155),
    .B(_2379_),
    .Y(_2726_));
 sg13g2_nand2_2 _3632_ (.Y(_2727_),
    .A(_2726_),
    .B(net60));
 sg13g2_buf_1 _3633_ (.A(net136),
    .X(_2728_));
 sg13g2_buf_1 _3634_ (.A(net151),
    .X(_2729_));
 sg13g2_a21oi_1 _3635_ (.A1(_2494_),
    .A2(net77),
    .Y(_2730_),
    .B1(net76));
 sg13g2_nand2_1 _3636_ (.Y(_2731_),
    .A(_2727_),
    .B(_2730_));
 sg13g2_buf_2 _3637_ (.A(net150),
    .X(_2732_));
 sg13g2_buf_2 _3638_ (.A(net75),
    .X(_2733_));
 sg13g2_nand3_1 _3639_ (.B(_2731_),
    .C(net46),
    .A(_2725_),
    .Y(_2734_));
 sg13g2_nand3_1 _3640_ (.B(_2734_),
    .C(net80),
    .A(_2721_),
    .Y(_2735_));
 sg13g2_buf_1 _3641_ (.A(net197),
    .X(_2736_));
 sg13g2_nand3b_1 _3642_ (.B(_2735_),
    .C(net164),
    .Y(_2737_),
    .A_N(_2708_));
 sg13g2_buf_1 _3643_ (.A(_2564_),
    .X(_2738_));
 sg13g2_inv_2 _3644_ (.Y(_2739_),
    .A(_2526_));
 sg13g2_nor2_2 _3645_ (.A(net76),
    .B(_2739_),
    .Y(_2740_));
 sg13g2_a21oi_1 _3646_ (.A1(_2740_),
    .A2(_1238_),
    .Y(_2741_),
    .B1(net78));
 sg13g2_nand2_1 _3647_ (.Y(_2742_),
    .A(_2221_),
    .B(net135));
 sg13g2_inv_1 _3648_ (.Y(_2743_),
    .A(_2742_));
 sg13g2_nor2_1 _3649_ (.A(_0998_),
    .B(_2494_),
    .Y(_2744_));
 sg13g2_buf_2 _3650_ (.A(_2744_),
    .X(_2745_));
 sg13g2_nand2_1 _3651_ (.Y(_2746_),
    .A(_2745_),
    .B(net122));
 sg13g2_inv_1 _3652_ (.Y(_2747_),
    .A(_2203_));
 sg13g2_nand3_1 _3653_ (.B(_2746_),
    .C(_2747_),
    .A(_2743_),
    .Y(_2748_));
 sg13g2_buf_1 _3654_ (.A(net169),
    .X(_2749_));
 sg13g2_a21oi_1 _3655_ (.A1(_2741_),
    .A2(_2748_),
    .Y(_2750_),
    .B1(net121));
 sg13g2_inv_2 _3656_ (.Y(_2751_),
    .A(_2193_));
 sg13g2_nand2_1 _3657_ (.Y(_2752_),
    .A(_2583_),
    .B(_2751_));
 sg13g2_buf_2 _3658_ (.A(_2729_),
    .X(_2753_));
 sg13g2_nand2_1 _3659_ (.Y(_2754_),
    .A(_2752_),
    .B(net45));
 sg13g2_nand2_1 _3660_ (.Y(_2755_),
    .A(_2502_),
    .B(_2671_));
 sg13g2_nor2_1 _3661_ (.A(net79),
    .B(_2755_),
    .Y(_2756_));
 sg13g2_inv_1 _3662_ (.Y(_2757_),
    .A(_1805_));
 sg13g2_inv_1 _3663_ (.Y(_2758_),
    .A(net87));
 sg13g2_nor2_1 _3664_ (.A(net91),
    .B(_2758_),
    .Y(_2759_));
 sg13g2_buf_1 _3665_ (.A(net198),
    .X(_2760_));
 sg13g2_a21oi_1 _3666_ (.A1(_2757_),
    .A2(_2759_),
    .Y(_2761_),
    .B1(net162));
 sg13g2_o21ai_1 _3667_ (.B1(_2761_),
    .Y(_2762_),
    .A1(_2754_),
    .A2(_2756_));
 sg13g2_nand2_1 _3668_ (.Y(_2763_),
    .A(_2750_),
    .B(_2762_));
 sg13g2_a21oi_1 _3669_ (.A1(_2571_),
    .A2(net47),
    .Y(_2764_),
    .B1(net149));
 sg13g2_nand2_1 _3670_ (.Y(_2765_),
    .A(net94),
    .B(net144));
 sg13g2_nand2_1 _3671_ (.Y(_2766_),
    .A(_2765_),
    .B(_2491_));
 sg13g2_nand2_1 _3672_ (.Y(_2767_),
    .A(_2764_),
    .B(_2766_));
 sg13g2_nand2_1 _3673_ (.Y(_2768_),
    .A(_1609_),
    .B(net51));
 sg13g2_buf_1 _3674_ (.A(net174),
    .X(_2769_));
 sg13g2_a21oi_1 _3675_ (.A1(_2768_),
    .A2(net120),
    .Y(_2770_),
    .B1(net78));
 sg13g2_nand2_1 _3676_ (.Y(_2771_),
    .A(_2767_),
    .B(_2770_));
 sg13g2_nand2_1 _3677_ (.Y(_2772_),
    .A(_2629_),
    .B(net146));
 sg13g2_nand2_1 _3678_ (.Y(_2773_),
    .A(_2772_),
    .B(net97));
 sg13g2_buf_1 _3679_ (.A(net62),
    .X(_2774_));
 sg13g2_nor2_1 _3680_ (.A(net79),
    .B(_2636_),
    .Y(_2775_));
 sg13g2_nor3_1 _3681_ (.A(net139),
    .B(net28),
    .C(_2775_),
    .Y(_2776_));
 sg13g2_a21oi_1 _3682_ (.A1(_2773_),
    .A2(_2776_),
    .Y(_2777_),
    .B1(net127));
 sg13g2_buf_8 _3683_ (.A(_2469_),
    .X(_2778_));
 sg13g2_nand2_2 _3684_ (.Y(_2779_),
    .A(net44),
    .B(net154));
 sg13g2_inv_1 _3685_ (.Y(_2780_),
    .A(_2779_));
 sg13g2_a21oi_1 _3686_ (.A1(_2020_),
    .A2(net144),
    .Y(_2781_),
    .B1(net154));
 sg13g2_buf_1 _3687_ (.A(net134),
    .X(_2782_));
 sg13g2_o21ai_1 _3688_ (.B1(_2782_),
    .Y(_2783_),
    .A1(_2780_),
    .A2(_2781_));
 sg13g2_nand3_1 _3689_ (.B(_2777_),
    .C(_2783_),
    .A(_2771_),
    .Y(_2784_));
 sg13g2_buf_1 _3690_ (.A(net147),
    .X(_2785_));
 sg13g2_nand3_1 _3691_ (.B(_2784_),
    .C(net73),
    .A(_2763_),
    .Y(_2786_));
 sg13g2_nand3_1 _3692_ (.B(net163),
    .C(_2786_),
    .A(_2737_),
    .Y(_2787_));
 sg13g2_nand2_1 _3693_ (.Y(_2788_),
    .A(_2697_),
    .B(_2787_));
 sg13g2_nand2_1 _3694_ (.Y(_0021_),
    .A(_2612_),
    .B(_2788_));
 sg13g2_nand2_2 _3695_ (.Y(_2789_),
    .A(_2529_),
    .B(net139));
 sg13g2_inv_1 _3696_ (.Y(_2790_),
    .A(_2789_));
 sg13g2_nor2_1 _3697_ (.A(_2518_),
    .B(_2790_),
    .Y(_2791_));
 sg13g2_nand2_1 _3698_ (.Y(_2792_),
    .A(_1609_),
    .B(net181));
 sg13g2_buf_2 _3699_ (.A(_2792_),
    .X(_2793_));
 sg13g2_nand2_1 _3700_ (.Y(_2794_),
    .A(_2494_),
    .B(_0889_));
 sg13g2_buf_8 _3701_ (.A(_2794_),
    .X(_2795_));
 sg13g2_nand2_2 _3702_ (.Y(_2796_),
    .A(_2793_),
    .B(net43));
 sg13g2_nand2_2 _3703_ (.Y(_2797_),
    .A(_2796_),
    .B(_2437_));
 sg13g2_a21oi_1 _3704_ (.A1(_2791_),
    .A2(_2797_),
    .Y(_2798_),
    .B1(net81));
 sg13g2_nand2_1 _3705_ (.Y(_2799_),
    .A(_2524_),
    .B(net190));
 sg13g2_buf_2 _3706_ (.A(_2799_),
    .X(_2800_));
 sg13g2_inv_1 _3707_ (.Y(_2801_),
    .A(_2800_));
 sg13g2_nor2_1 _3708_ (.A(_2801_),
    .B(_2573_),
    .Y(_2802_));
 sg13g2_nand2_2 _3709_ (.Y(_2803_),
    .A(_2802_),
    .B(net60));
 sg13g2_nand2_1 _3710_ (.Y(_2804_),
    .A(_2803_),
    .B(_2764_));
 sg13g2_nand2_1 _3711_ (.Y(_2805_),
    .A(_2798_),
    .B(_2804_));
 sg13g2_nand2_1 _3712_ (.Y(_2806_),
    .A(net98),
    .B(net133));
 sg13g2_nand2_1 _3713_ (.Y(_2807_),
    .A(_2806_),
    .B(net79));
 sg13g2_buf_1 _3714_ (.A(_1249_),
    .X(_2808_));
 sg13g2_nand2_1 _3715_ (.Y(_2809_),
    .A(net156),
    .B(net119));
 sg13g2_nand2_1 _3716_ (.Y(_2810_),
    .A(net85),
    .B(_2809_));
 sg13g2_nand2_1 _3717_ (.Y(_2811_),
    .A(_2807_),
    .B(_2810_));
 sg13g2_inv_1 _3718_ (.Y(_2812_),
    .A(net85));
 sg13g2_nand2_1 _3719_ (.Y(_2813_),
    .A(_2751_),
    .B(_1609_));
 sg13g2_o21ai_1 _3720_ (.B1(_2813_),
    .Y(_2814_),
    .A1(net47),
    .A2(_2812_));
 sg13g2_a22oi_1 _3721_ (.Y(_2815_),
    .B1(net50),
    .B2(_2814_),
    .A2(net74),
    .A1(_2811_));
 sg13g2_buf_2 _3722_ (.A(_2558_),
    .X(_2816_));
 sg13g2_a21oi_1 _3723_ (.A1(_2805_),
    .A2(_2815_),
    .Y(_2817_),
    .B1(net118));
 sg13g2_nor2_1 _3724_ (.A(net198),
    .B(_2781_),
    .Y(_2818_));
 sg13g2_a21oi_2 _3725_ (.B1(net152),
    .Y(_2819_),
    .A2(_1184_),
    .A1(_1151_));
 sg13g2_nand2_1 _3726_ (.Y(_2820_),
    .A(_2819_),
    .B(net52));
 sg13g2_nand2_1 _3727_ (.Y(_2821_),
    .A(_2818_),
    .B(_2820_));
 sg13g2_a21oi_1 _3728_ (.A1(net44),
    .A2(_2660_),
    .Y(_2822_),
    .B1(net150));
 sg13g2_a22oi_1 _3729_ (.Y(_2823_),
    .B1(_2392_),
    .B2(net103),
    .A2(net143),
    .A1(_1478_));
 sg13g2_nand2_1 _3730_ (.Y(_2824_),
    .A(_2822_),
    .B(_2823_));
 sg13g2_nand2_1 _3731_ (.Y(_2825_),
    .A(_2821_),
    .B(_2824_));
 sg13g2_buf_2 _3732_ (.A(net149),
    .X(_2826_));
 sg13g2_nand2_1 _3733_ (.Y(_2827_),
    .A(_2825_),
    .B(_2826_));
 sg13g2_nand2_1 _3734_ (.Y(_2828_),
    .A(_2470_),
    .B(net198));
 sg13g2_nand2_1 _3735_ (.Y(_2829_),
    .A(_0943_),
    .B(net119));
 sg13g2_nand2_1 _3736_ (.Y(_2830_),
    .A(net125),
    .B(_2829_));
 sg13g2_a21oi_1 _3737_ (.A1(_2830_),
    .A2(net140),
    .Y(_2831_),
    .B1(net177));
 sg13g2_nand2_1 _3738_ (.Y(_2832_),
    .A(_2828_),
    .B(_2831_));
 sg13g2_nand2_1 _3739_ (.Y(_2833_),
    .A(net125),
    .B(net153));
 sg13g2_nand2_1 _3740_ (.Y(_2834_),
    .A(_2709_),
    .B(_2833_));
 sg13g2_nand2_1 _3741_ (.Y(_2835_),
    .A(_2834_),
    .B(_2491_));
 sg13g2_nor2_1 _3742_ (.A(net199),
    .B(_2835_),
    .Y(_2836_));
 sg13g2_nor2_1 _3743_ (.A(_2832_),
    .B(_2836_),
    .Y(_2837_));
 sg13g2_nor2_1 _3744_ (.A(_2374_),
    .B(_2837_),
    .Y(_2838_));
 sg13g2_nand2_1 _3745_ (.Y(_2839_),
    .A(_2827_),
    .B(_2838_));
 sg13g2_nand2_1 _3746_ (.Y(_2840_),
    .A(_2839_),
    .B(_2423_));
 sg13g2_nor2_1 _3747_ (.A(_2817_),
    .B(_2840_),
    .Y(_2841_));
 sg13g2_inv_2 _3748_ (.Y(_2842_),
    .A(_1998_));
 sg13g2_nand3_1 _3749_ (.B(net87),
    .C(_2842_),
    .A(net122),
    .Y(_2843_));
 sg13g2_buf_1 _3750_ (.A(net58),
    .X(_2844_));
 sg13g2_nand2_1 _3751_ (.Y(_2845_),
    .A(_2400_),
    .B(net27));
 sg13g2_nand2_1 _3752_ (.Y(_2846_),
    .A(_2843_),
    .B(_2845_));
 sg13g2_nor2_1 _3753_ (.A(net119),
    .B(net90),
    .Y(_2847_));
 sg13g2_buf_4 _3754_ (.X(_2848_),
    .A(_2847_));
 sg13g2_o21ai_1 _3755_ (.B1(net140),
    .Y(_2849_),
    .A1(_2575_),
    .A2(_2848_));
 sg13g2_buf_2 _3756_ (.A(_2849_),
    .X(_2850_));
 sg13g2_nor2_1 _3757_ (.A(_2769_),
    .B(_2850_),
    .Y(_2851_));
 sg13g2_o21ai_1 _3758_ (.B1(net46),
    .Y(_2852_),
    .A1(_2846_),
    .A2(_2851_));
 sg13g2_nand2_1 _3759_ (.Y(_2853_),
    .A(_1859_),
    .B(net152));
 sg13g2_inv_2 _3760_ (.Y(_2854_),
    .A(_2441_));
 sg13g2_nand3_1 _3761_ (.B(net76),
    .C(_2854_),
    .A(_2853_),
    .Y(_2855_));
 sg13g2_nand2_1 _3762_ (.Y(_2856_),
    .A(_2436_),
    .B(net140));
 sg13g2_nand2_1 _3763_ (.Y(_2857_),
    .A(_2856_),
    .B(net199));
 sg13g2_o21ai_1 _3764_ (.B1(net123),
    .Y(_2858_),
    .A1(_2855_),
    .A2(_2857_));
 sg13g2_nand3_1 _3765_ (.B(net186),
    .C(net207),
    .A(_0746_),
    .Y(_2859_));
 sg13g2_buf_2 _3766_ (.A(_2859_),
    .X(_2860_));
 sg13g2_nand2_2 _3767_ (.Y(_2861_),
    .A(_2860_),
    .B(_1020_));
 sg13g2_o21ai_1 _3768_ (.B1(_2861_),
    .Y(_2862_),
    .A1(net77),
    .A2(_2848_));
 sg13g2_a21oi_1 _3769_ (.A1(_2862_),
    .A2(net97),
    .Y(_2863_),
    .B1(net145));
 sg13g2_nor2_1 _3770_ (.A(_2858_),
    .B(_2863_),
    .Y(_2864_));
 sg13g2_nand2_1 _3771_ (.Y(_2865_),
    .A(_2852_),
    .B(_2864_));
 sg13g2_a21oi_1 _3772_ (.A1(_2634_),
    .A2(_2682_),
    .Y(_2866_),
    .B1(_1020_));
 sg13g2_nor2_1 _3773_ (.A(net62),
    .B(_2866_),
    .Y(_2867_));
 sg13g2_nand2_1 _3774_ (.Y(_2868_),
    .A(_2867_),
    .B(_2239_));
 sg13g2_nand2_1 _3775_ (.Y(_2869_),
    .A(net43),
    .B(_2800_));
 sg13g2_nand2_1 _3776_ (.Y(_2870_),
    .A(_2869_),
    .B(net51));
 sg13g2_nor2_2 _3777_ (.A(net157),
    .B(_2392_),
    .Y(_2871_));
 sg13g2_nor2_1 _3778_ (.A(_1326_),
    .B(_2871_),
    .Y(_2872_));
 sg13g2_nand2_1 _3779_ (.Y(_2873_),
    .A(_2870_),
    .B(_2872_));
 sg13g2_nand2_1 _3780_ (.Y(_2874_),
    .A(_2868_),
    .B(_2873_));
 sg13g2_a21oi_1 _3781_ (.A1(_2745_),
    .A2(_2793_),
    .Y(_2875_),
    .B1(_2467_));
 sg13g2_o21ai_1 _3782_ (.B1(net167),
    .Y(_2876_),
    .A1(net54),
    .A2(_2875_));
 sg13g2_nor2_1 _3783_ (.A(_2874_),
    .B(_2876_),
    .Y(_2877_));
 sg13g2_nand2_1 _3784_ (.Y(_2878_),
    .A(_1805_),
    .B(_2457_));
 sg13g2_buf_4 _3785_ (.X(_2879_),
    .A(_2878_));
 sg13g2_inv_4 _3786_ (.A(_2879_),
    .Y(_2880_));
 sg13g2_nor2_1 _3787_ (.A(net56),
    .B(_2504_),
    .Y(_2881_));
 sg13g2_buf_1 _3788_ (.A(_2626_),
    .X(_2882_));
 sg13g2_o21ai_1 _3789_ (.B1(net70),
    .Y(_2883_),
    .A1(_2880_),
    .A2(_2881_));
 sg13g2_nand2_1 _3790_ (.Y(_2884_),
    .A(_2877_),
    .B(_2883_));
 sg13g2_nand3_1 _3791_ (.B(_2884_),
    .C(net73),
    .A(_2865_),
    .Y(_2885_));
 sg13g2_a21oi_1 _3792_ (.A1(_2841_),
    .A2(_2885_),
    .Y(_2886_),
    .B1(net196));
 sg13g2_nor2_2 _3793_ (.A(net186),
    .B(net181),
    .Y(_2887_));
 sg13g2_nor2_1 _3794_ (.A(_2887_),
    .B(_2671_),
    .Y(_2888_));
 sg13g2_nor2_2 _3795_ (.A(net157),
    .B(_2888_),
    .Y(_2889_));
 sg13g2_nand2_1 _3796_ (.Y(_2890_),
    .A(_2889_),
    .B(_2503_));
 sg13g2_nor2_1 _3797_ (.A(net187),
    .B(_2584_),
    .Y(_2891_));
 sg13g2_buf_2 _3798_ (.A(_2891_),
    .X(_2892_));
 sg13g2_nand2_1 _3799_ (.Y(_2893_),
    .A(_2892_),
    .B(net95));
 sg13g2_nand2_1 _3800_ (.Y(_2894_),
    .A(_2890_),
    .B(_2893_));
 sg13g2_buf_1 _3801_ (.A(net110),
    .X(_2895_));
 sg13g2_nand2_1 _3802_ (.Y(_2896_),
    .A(_2894_),
    .B(net42));
 sg13g2_nand2_1 _3803_ (.Y(_2897_),
    .A(_1271_),
    .B(_2458_));
 sg13g2_a21oi_1 _3804_ (.A1(_2897_),
    .A2(net51),
    .Y(_2898_),
    .B1(_2406_));
 sg13g2_nor2_1 _3805_ (.A(net157),
    .B(_2494_),
    .Y(_2899_));
 sg13g2_buf_2 _3806_ (.A(_2899_),
    .X(_2900_));
 sg13g2_nand2_1 _3807_ (.Y(_2901_),
    .A(_2900_),
    .B(net90));
 sg13g2_nand2_1 _3808_ (.Y(_2902_),
    .A(_2898_),
    .B(_2901_));
 sg13g2_nand2_1 _3809_ (.Y(_2903_),
    .A(_2896_),
    .B(_2902_));
 sg13g2_nand2_1 _3810_ (.Y(_2904_),
    .A(_0845_),
    .B(_1740_));
 sg13g2_buf_1 _3811_ (.A(_2904_),
    .X(_2905_));
 sg13g2_nor2_2 _3812_ (.A(_2398_),
    .B(_2573_),
    .Y(_2906_));
 sg13g2_o21ai_1 _3813_ (.B1(_2842_),
    .Y(_2907_),
    .A1(_2575_),
    .A2(_2577_));
 sg13g2_o21ai_1 _3814_ (.B1(_2907_),
    .Y(_2908_),
    .A1(net41),
    .A2(_2906_));
 sg13g2_nand2_1 _3815_ (.Y(_2909_),
    .A(_2908_),
    .B(net107));
 sg13g2_nand3_1 _3816_ (.B(net82),
    .C(_0856_),
    .A(_2671_),
    .Y(_2910_));
 sg13g2_nand2_1 _3817_ (.Y(_2911_),
    .A(_2897_),
    .B(net143));
 sg13g2_nand3_1 _3818_ (.B(_2911_),
    .C(_2568_),
    .A(_2910_),
    .Y(_2912_));
 sg13g2_nand2_1 _3819_ (.Y(_2913_),
    .A(_2909_),
    .B(_2912_));
 sg13g2_nor2_1 _3820_ (.A(_2903_),
    .B(_2913_),
    .Y(_2914_));
 sg13g2_nor2_1 _3821_ (.A(net63),
    .B(_2914_),
    .Y(_2915_));
 sg13g2_nor2_1 _3822_ (.A(net146),
    .B(_2273_),
    .Y(_2916_));
 sg13g2_nor2_1 _3823_ (.A(net174),
    .B(_2916_),
    .Y(_2917_));
 sg13g2_nand2_1 _3824_ (.Y(_2918_),
    .A(_2803_),
    .B(_2917_));
 sg13g2_a21oi_2 _3825_ (.B1(net151),
    .Y(_2919_),
    .A2(net154),
    .A1(_2726_));
 sg13g2_nand2_2 _3826_ (.Y(_2920_),
    .A(_2273_),
    .B(net139));
 sg13g2_nand2_1 _3827_ (.Y(_2921_),
    .A(_2919_),
    .B(_2920_));
 sg13g2_nand3_1 _3828_ (.B(_2921_),
    .C(net168),
    .A(_2918_),
    .Y(_2922_));
 sg13g2_nand2_1 _3829_ (.Y(_2923_),
    .A(_2854_),
    .B(net135));
 sg13g2_nor2_1 _3830_ (.A(_2923_),
    .B(_2869_),
    .Y(_2924_));
 sg13g2_a22oi_1 _3831_ (.Y(_2925_),
    .B1(net49),
    .B2(_2756_),
    .A2(_2924_),
    .A1(net107));
 sg13g2_nand2_1 _3832_ (.Y(_2926_),
    .A(_2922_),
    .B(_2925_));
 sg13g2_nand2_1 _3833_ (.Y(_2927_),
    .A(_2926_),
    .B(_2559_));
 sg13g2_nand2_1 _3834_ (.Y(_2928_),
    .A(_2927_),
    .B(net170));
 sg13g2_nor2_1 _3835_ (.A(_2915_),
    .B(_2928_),
    .Y(_2929_));
 sg13g2_o21ai_1 _3836_ (.B1(_2524_),
    .Y(_2930_),
    .A1(net201),
    .A2(net158));
 sg13g2_nor2_2 _3837_ (.A(_2490_),
    .B(_2930_),
    .Y(_2931_));
 sg13g2_nand2_1 _3838_ (.Y(_2932_),
    .A(_2931_),
    .B(net126));
 sg13g2_nand2_1 _3839_ (.Y(_2933_),
    .A(_2649_),
    .B(net87));
 sg13g2_a21oi_1 _3840_ (.A1(_2932_),
    .A2(_2933_),
    .Y(_2934_),
    .B1(net145));
 sg13g2_buf_2 _3841_ (.A(_1085_),
    .X(_2935_));
 sg13g2_nor2_1 _3842_ (.A(net203),
    .B(net69),
    .Y(_2936_));
 sg13g2_nand2_1 _3843_ (.Y(_2937_),
    .A(net43),
    .B(net144));
 sg13g2_nand2_1 _3844_ (.Y(_2938_),
    .A(_2937_),
    .B(net79));
 sg13g2_nand3_1 _3845_ (.B(_2428_),
    .C(net173),
    .A(_2938_),
    .Y(_2939_));
 sg13g2_nand2b_1 _3846_ (.Y(_2940_),
    .B(_2939_),
    .A_N(_2936_));
 sg13g2_nor2b_1 _3847_ (.A(_2934_),
    .B_N(_2940_),
    .Y(_2941_));
 sg13g2_nand2_1 _3848_ (.Y(_2942_),
    .A(net57),
    .B(_2800_));
 sg13g2_nand2_1 _3849_ (.Y(_2943_),
    .A(_2942_),
    .B(net30));
 sg13g2_nand2_1 _3850_ (.Y(_2944_),
    .A(_2919_),
    .B(_2943_));
 sg13g2_nor2_1 _3851_ (.A(net174),
    .B(_2638_),
    .Y(_2945_));
 sg13g2_nand2_1 _3852_ (.Y(_2946_),
    .A(net126),
    .B(net201));
 sg13g2_buf_2 _3853_ (.A(_2946_),
    .X(_2947_));
 sg13g2_nor2_1 _3854_ (.A(net58),
    .B(_2947_),
    .Y(_2948_));
 sg13g2_inv_1 _3855_ (.Y(_2949_),
    .A(_2948_));
 sg13g2_a21oi_1 _3856_ (.A1(_2945_),
    .A2(_2949_),
    .Y(_2950_),
    .B1(_2517_));
 sg13g2_nand2_1 _3857_ (.Y(_2951_),
    .A(_2944_),
    .B(_2950_));
 sg13g2_a21oi_1 _3858_ (.A1(_2941_),
    .A2(_2951_),
    .Y(_2952_),
    .B1(net164));
 sg13g2_nand2_1 _3859_ (.Y(_2953_),
    .A(net71),
    .B(net94));
 sg13g2_nor2_1 _3860_ (.A(net30),
    .B(_2953_),
    .Y(_2954_));
 sg13g2_a21oi_1 _3861_ (.A1(_2503_),
    .A2(_2433_),
    .Y(_2955_),
    .B1(_2506_));
 sg13g2_o21ai_1 _3862_ (.B1(net53),
    .Y(_2956_),
    .A1(_2954_),
    .A2(_2955_));
 sg13g2_buf_1 _3863_ (.A(net167),
    .X(_2957_));
 sg13g2_nor2_2 _3864_ (.A(net184),
    .B(_1795_),
    .Y(_2958_));
 sg13g2_nand2_2 _3865_ (.Y(_2959_),
    .A(_2958_),
    .B(net95));
 sg13g2_nor2_2 _3866_ (.A(net185),
    .B(_1653_),
    .Y(_2960_));
 sg13g2_nor2_1 _3867_ (.A(net103),
    .B(_2960_),
    .Y(_2961_));
 sg13g2_a21o_1 _3868_ (.A2(_2961_),
    .A1(_2959_),
    .B1(_2390_),
    .X(_2962_));
 sg13g2_buf_1 _3869_ (.A(net101),
    .X(_2963_));
 sg13g2_nand2_1 _3870_ (.Y(_2964_),
    .A(_1911_),
    .B(net187));
 sg13g2_inv_1 _3871_ (.Y(_2965_),
    .A(_2964_));
 sg13g2_nor2_1 _3872_ (.A(net40),
    .B(_2965_),
    .Y(_2966_));
 sg13g2_nand2_2 _3873_ (.Y(_2967_),
    .A(_2273_),
    .B(net189));
 sg13g2_buf_2 _3874_ (.A(net49),
    .X(_2968_));
 sg13g2_nor2_2 _3875_ (.A(_1838_),
    .B(_2392_),
    .Y(_2969_));
 sg13g2_inv_2 _3876_ (.Y(_2970_),
    .A(_2969_));
 sg13g2_nand2_1 _3877_ (.Y(_2971_),
    .A(_2970_),
    .B(net148));
 sg13g2_a22oi_1 _3878_ (.Y(_2972_),
    .B1(net26),
    .B2(_2971_),
    .A2(_2967_),
    .A1(_2966_));
 sg13g2_nand4_1 _3879_ (.B(net117),
    .C(_2962_),
    .A(_2956_),
    .Y(_2973_),
    .D(_2972_));
 sg13g2_nand2_1 _3880_ (.Y(_2974_),
    .A(_2952_),
    .B(_2973_));
 sg13g2_nand2_1 _3881_ (.Y(_2975_),
    .A(_2929_),
    .B(_2974_));
 sg13g2_nand2_1 _3882_ (.Y(_2976_),
    .A(_2886_),
    .B(_2975_));
 sg13g2_a21oi_2 _3883_ (.B1(_2450_),
    .Y(_2977_),
    .A2(net95),
    .A1(_2958_));
 sg13g2_nand2_1 _3884_ (.Y(_2978_),
    .A(_2020_),
    .B(net144));
 sg13g2_nand2_1 _3885_ (.Y(_2979_),
    .A(_2978_),
    .B(net102));
 sg13g2_nand3_1 _3886_ (.B(net84),
    .C(_2979_),
    .A(_2977_),
    .Y(_2980_));
 sg13g2_nor2_1 _3887_ (.A(net176),
    .B(net44),
    .Y(_2981_));
 sg13g2_inv_1 _3888_ (.Y(_2982_),
    .A(_2981_));
 sg13g2_nor2_1 _3889_ (.A(net179),
    .B(_2519_),
    .Y(_2983_));
 sg13g2_a21oi_1 _3890_ (.A1(_2982_),
    .A2(_2983_),
    .Y(_2984_),
    .B1(net162));
 sg13g2_nand2_1 _3891_ (.Y(_2985_),
    .A(_2980_),
    .B(_2984_));
 sg13g2_a21oi_2 _3892_ (.B1(net154),
    .Y(_2986_),
    .A2(net201),
    .A1(net155));
 sg13g2_nor2_1 _3893_ (.A(_2533_),
    .B(_2986_),
    .Y(_2987_));
 sg13g2_nand2_1 _3894_ (.Y(_2988_),
    .A(net94),
    .B(net90));
 sg13g2_nand2_1 _3895_ (.Y(_2989_),
    .A(_2988_),
    .B(net56));
 sg13g2_buf_1 _3896_ (.A(net110),
    .X(_2990_));
 sg13g2_buf_1 _3897_ (.A(net39),
    .X(_2991_));
 sg13g2_nor2_2 _3898_ (.A(net187),
    .B(_2887_),
    .Y(_2992_));
 sg13g2_nand2_1 _3899_ (.Y(_2993_),
    .A(_2992_),
    .B(net158));
 sg13g2_nand2_1 _3900_ (.Y(_2994_),
    .A(_2993_),
    .B(_2455_));
 sg13g2_a22oi_1 _3901_ (.Y(_2995_),
    .B1(net25),
    .B2(_2994_),
    .A2(_2989_),
    .A1(_2987_));
 sg13g2_a21oi_1 _3902_ (.A1(_2985_),
    .A2(_2995_),
    .Y(_2996_),
    .B1(net63));
 sg13g2_buf_8 _3903_ (.A(_1151_),
    .X(_2997_));
 sg13g2_nor2_2 _3904_ (.A(net106),
    .B(net38),
    .Y(_2998_));
 sg13g2_nor2_1 _3905_ (.A(_2998_),
    .B(_2723_),
    .Y(_2999_));
 sg13g2_nand2_1 _3906_ (.Y(_3000_),
    .A(_2999_),
    .B(_2221_));
 sg13g2_nand2_1 _3907_ (.Y(_3001_),
    .A(_2579_),
    .B(_2979_));
 sg13g2_a22oi_1 _3908_ (.Y(_3002_),
    .B1(net53),
    .B2(_3001_),
    .A2(_3000_),
    .A1(net50));
 sg13g2_nand2_2 _3909_ (.Y(_3003_),
    .A(_1609_),
    .B(net136));
 sg13g2_nand2_1 _3910_ (.Y(_3004_),
    .A(_2530_),
    .B(_3003_));
 sg13g2_nand2_2 _3911_ (.Y(_3005_),
    .A(_1948_),
    .B(net96));
 sg13g2_nor2_1 _3912_ (.A(net40),
    .B(_3005_),
    .Y(_3006_));
 sg13g2_nand2_1 _3913_ (.Y(_3007_),
    .A(_2622_),
    .B(net137));
 sg13g2_nand2_2 _3914_ (.Y(_3008_),
    .A(_3007_),
    .B(net92));
 sg13g2_a22oi_1 _3915_ (.Y(_3009_),
    .B1(_3006_),
    .B2(_3008_),
    .A2(_3004_),
    .A1(net42));
 sg13g2_a21oi_1 _3916_ (.A1(_3002_),
    .A2(_3009_),
    .Y(_3010_),
    .B1(net118));
 sg13g2_nor3_1 _3917_ (.A(net200),
    .B(_2996_),
    .C(_3010_),
    .Y(_3011_));
 sg13g2_nand2_1 _3918_ (.Y(_3012_),
    .A(_2582_),
    .B(_2442_));
 sg13g2_nor2_2 _3919_ (.A(net157),
    .B(_2633_),
    .Y(_3013_));
 sg13g2_nand2_2 _3920_ (.Y(_3014_),
    .A(_2397_),
    .B(_1260_));
 sg13g2_nand2_1 _3921_ (.Y(_3015_),
    .A(_3013_),
    .B(_3014_));
 sg13g2_a21oi_1 _3922_ (.A1(_3012_),
    .A2(_3015_),
    .Y(_3016_),
    .B1(_2408_));
 sg13g2_nand3_1 _3923_ (.B(net100),
    .C(net60),
    .A(net82),
    .Y(_3017_));
 sg13g2_nor2_2 _3924_ (.A(net111),
    .B(_1620_),
    .Y(_3018_));
 sg13g2_inv_1 _3925_ (.Y(_3019_),
    .A(_3018_));
 sg13g2_and3_1 _3926_ (.X(_3020_),
    .A(_3017_),
    .B(net50),
    .C(_3019_));
 sg13g2_nor3_1 _3927_ (.A(net121),
    .B(_3016_),
    .C(_3020_),
    .Y(_3021_));
 sg13g2_buf_1 _3928_ (.A(_1631_),
    .X(_3022_));
 sg13g2_buf_1 _3929_ (.A(net37),
    .X(_3023_));
 sg13g2_nand2_1 _3930_ (.Y(_3024_),
    .A(_2796_),
    .B(_1522_));
 sg13g2_buf_2 _3931_ (.A(_3024_),
    .X(_3025_));
 sg13g2_nand2_1 _3932_ (.Y(_3026_),
    .A(_2751_),
    .B(net98));
 sg13g2_nand2_1 _3933_ (.Y(_3027_),
    .A(_3025_),
    .B(_3026_));
 sg13g2_nor2_1 _3934_ (.A(net184),
    .B(_2379_),
    .Y(_3028_));
 sg13g2_nor2_2 _3935_ (.A(net148),
    .B(_1151_),
    .Y(_3029_));
 sg13g2_nor2_2 _3936_ (.A(net202),
    .B(_3029_),
    .Y(_3030_));
 sg13g2_nand2b_1 _3937_ (.Y(_3031_),
    .B(_3030_),
    .A_N(_2635_));
 sg13g2_nor2_1 _3938_ (.A(_3028_),
    .B(_3031_),
    .Y(_3032_));
 sg13g2_nor2_1 _3939_ (.A(_2689_),
    .B(_3032_),
    .Y(_3033_));
 sg13g2_o21ai_1 _3940_ (.B1(_3033_),
    .Y(_3034_),
    .A1(_3023_),
    .A2(_3027_));
 sg13g2_nand2_1 _3941_ (.Y(_3035_),
    .A(_3021_),
    .B(_3034_));
 sg13g2_inv_1 _3942_ (.Y(_3036_),
    .A(_1930_));
 sg13g2_nand3_1 _3943_ (.B(net55),
    .C(_3036_),
    .A(_2850_),
    .Y(_3037_));
 sg13g2_a21oi_1 _3944_ (.A1(_2530_),
    .A2(_2769_),
    .Y(_3038_),
    .B1(_2716_));
 sg13g2_buf_1 _3945_ (.A(_2460_),
    .X(_3039_));
 sg13g2_buf_1 _3946_ (.A(net161),
    .X(_3040_));
 sg13g2_a21oi_1 _3947_ (.A1(_3037_),
    .A2(_3038_),
    .Y(_3041_),
    .B1(_3040_));
 sg13g2_nand2_1 _3948_ (.Y(_3042_),
    .A(_2086_),
    .B(_2745_));
 sg13g2_buf_8 _3949_ (.A(_3042_),
    .X(_3043_));
 sg13g2_nand2_1 _3950_ (.Y(_3044_),
    .A(net44),
    .B(_2751_));
 sg13g2_nand2_1 _3951_ (.Y(_3045_),
    .A(_3043_),
    .B(_3044_));
 sg13g2_a21oi_2 _3952_ (.B1(_2519_),
    .Y(_3046_),
    .A2(_1478_),
    .A1(net111));
 sg13g2_nor2_1 _3953_ (.A(net152),
    .B(_2809_),
    .Y(_3047_));
 sg13g2_inv_1 _3954_ (.Y(_3048_),
    .A(_3047_));
 sg13g2_nand3_1 _3955_ (.B(_3048_),
    .C(_2496_),
    .A(_3046_),
    .Y(_3049_));
 sg13g2_a22oi_1 _3956_ (.Y(_0088_),
    .B1(net70),
    .B2(_3049_),
    .A2(net26),
    .A1(_3045_));
 sg13g2_nand2_1 _3957_ (.Y(_0089_),
    .A(_3041_),
    .B(_0088_));
 sg13g2_buf_2 _3958_ (.A(net147),
    .X(_0090_));
 sg13g2_nand3_1 _3959_ (.B(_0089_),
    .C(net68),
    .A(_3035_),
    .Y(_0091_));
 sg13g2_nand2_1 _3960_ (.Y(_0092_),
    .A(_3011_),
    .B(_0091_));
 sg13g2_nand2_2 _3961_ (.Y(_0093_),
    .A(_2965_),
    .B(net122));
 sg13g2_a21oi_1 _3962_ (.A1(_3012_),
    .A2(_0093_),
    .Y(_0094_),
    .B1(net31));
 sg13g2_nor3_1 _3963_ (.A(_1096_),
    .B(_2577_),
    .C(_2478_),
    .Y(_0095_));
 sg13g2_nand2_1 _3964_ (.Y(_0096_),
    .A(_2745_),
    .B(_2683_));
 sg13g2_nor2_1 _3965_ (.A(_2417_),
    .B(_0096_),
    .Y(_0097_));
 sg13g2_nor2_1 _3966_ (.A(_0095_),
    .B(_0097_),
    .Y(_0098_));
 sg13g2_nand2_1 _3967_ (.Y(_0099_),
    .A(_2675_),
    .B(_0910_));
 sg13g2_nand2_2 _3968_ (.Y(_0100_),
    .A(_0099_),
    .B(net136));
 sg13g2_nor2_1 _3969_ (.A(_2406_),
    .B(_0100_),
    .Y(_0101_));
 sg13g2_nor2_1 _3970_ (.A(net203),
    .B(_0101_),
    .Y(_0102_));
 sg13g2_nand2_1 _3971_ (.Y(_0103_),
    .A(_0098_),
    .B(_0102_));
 sg13g2_a21oi_1 _3972_ (.A1(_2850_),
    .A2(_3025_),
    .Y(_0104_),
    .B1(net145));
 sg13g2_nor3_1 _3973_ (.A(_0094_),
    .B(_0103_),
    .C(_0104_),
    .Y(_0105_));
 sg13g2_nor2_1 _3974_ (.A(_2646_),
    .B(_0105_),
    .Y(_0106_));
 sg13g2_nand2_1 _3975_ (.Y(_0107_),
    .A(_2673_),
    .B(_0801_));
 sg13g2_nand2_1 _3976_ (.Y(_0108_),
    .A(net43),
    .B(net86));
 sg13g2_o21ai_1 _3977_ (.B1(_0108_),
    .Y(_0109_),
    .A1(net77),
    .A2(_0107_));
 sg13g2_buf_1 _3978_ (.A(net108),
    .X(_0110_));
 sg13g2_nand2_1 _3979_ (.Y(_0111_),
    .A(_0109_),
    .B(net36));
 sg13g2_nor2_2 _3980_ (.A(_1424_),
    .B(_1773_),
    .Y(_0112_));
 sg13g2_nor3_1 _3981_ (.A(net155),
    .B(_1998_),
    .C(_0112_),
    .Y(_0113_));
 sg13g2_nor2_1 _3982_ (.A(net41),
    .B(_2897_),
    .Y(_0114_));
 sg13g2_nor3_1 _3983_ (.A(net173),
    .B(_0113_),
    .C(_0114_),
    .Y(_0115_));
 sg13g2_nand2_1 _3984_ (.Y(_0116_),
    .A(_0111_),
    .B(_0115_));
 sg13g2_nand2_1 _3985_ (.Y(_0117_),
    .A(net180),
    .B(\mem_addr[6] ));
 sg13g2_buf_2 _3986_ (.A(_0117_),
    .X(_0118_));
 sg13g2_nand2_1 _3987_ (.Y(_0119_),
    .A(_0116_),
    .B(_0118_));
 sg13g2_nand3_1 _3988_ (.B(net38),
    .C(_1653_),
    .A(net57),
    .Y(_0120_));
 sg13g2_a22oi_1 _3989_ (.Y(_0121_),
    .B1(net70),
    .B2(_3027_),
    .A2(_2593_),
    .A1(_0120_));
 sg13g2_nand2_1 _3990_ (.Y(_0122_),
    .A(_0119_),
    .B(_0121_));
 sg13g2_nand2_1 _3991_ (.Y(_0123_),
    .A(_0106_),
    .B(_0122_));
 sg13g2_nand2_1 _3992_ (.Y(_0124_),
    .A(_2793_),
    .B(net156));
 sg13g2_nand2_1 _3993_ (.Y(_0125_),
    .A(_0124_),
    .B(net56));
 sg13g2_nand2_1 _3994_ (.Y(_0126_),
    .A(_0125_),
    .B(_2854_));
 sg13g2_buf_1 _3995_ (.A(_0035_),
    .X(_0127_));
 sg13g2_inv_2 _3996_ (.Y(_0128_),
    .A(_0127_));
 sg13g2_nor3_1 _3997_ (.A(net130),
    .B(_0128_),
    .C(_2690_),
    .Y(_0129_));
 sg13g2_a21oi_1 _3998_ (.A1(_0126_),
    .A2(_0129_),
    .Y(_0130_),
    .B1(_2565_));
 sg13g2_a21oi_1 _3999_ (.A1(_0123_),
    .A2(_0130_),
    .Y(_0131_),
    .B1(net165));
 sg13g2_nand2_1 _4000_ (.Y(_0132_),
    .A(_0092_),
    .B(_0131_));
 sg13g2_nand2_1 _4001_ (.Y(_0022_),
    .A(_2976_),
    .B(_0132_));
 sg13g2_nand2_1 _4002_ (.Y(_0133_),
    .A(net71),
    .B(_2673_));
 sg13g2_nor2_2 _4003_ (.A(net111),
    .B(_0133_),
    .Y(_0134_));
 sg13g2_nand2_1 _4004_ (.Y(_0135_),
    .A(_2683_),
    .B(_2550_));
 sg13g2_nand2_1 _4005_ (.Y(_0136_),
    .A(_0135_),
    .B(_2405_));
 sg13g2_nor2_1 _4006_ (.A(_0134_),
    .B(_0136_),
    .Y(_0137_));
 sg13g2_nand2_1 _4007_ (.Y(_0138_),
    .A(_2397_),
    .B(_1588_));
 sg13g2_nand2_1 _4008_ (.Y(_0139_),
    .A(_0138_),
    .B(_1859_));
 sg13g2_nand2_1 _4009_ (.Y(_0140_),
    .A(_0139_),
    .B(net93));
 sg13g2_nand2_1 _4010_ (.Y(_0141_),
    .A(_0140_),
    .B(_1336_));
 sg13g2_inv_2 _4011_ (.Y(_0142_),
    .A(net148));
 sg13g2_nor2_2 _4012_ (.A(_0142_),
    .B(net86),
    .Y(_0143_));
 sg13g2_nor2_1 _4013_ (.A(_0757_),
    .B(_2683_),
    .Y(_0144_));
 sg13g2_nor2_2 _4014_ (.A(_0143_),
    .B(_0144_),
    .Y(_0145_));
 sg13g2_nor2_1 _4015_ (.A(_0141_),
    .B(_0145_),
    .Y(_0146_));
 sg13g2_nor2_1 _4016_ (.A(_0137_),
    .B(_0146_),
    .Y(_0147_));
 sg13g2_nor2_2 _4017_ (.A(_2495_),
    .B(_2513_),
    .Y(_0148_));
 sg13g2_nand2_2 _4018_ (.Y(_0149_),
    .A(_2469_),
    .B(_1260_));
 sg13g2_nand2_2 _4019_ (.Y(_0150_),
    .A(_0149_),
    .B(_2547_));
 sg13g2_nand2b_1 _4020_ (.Y(_0151_),
    .B(_0150_),
    .A_N(_0148_));
 sg13g2_nand2_1 _4021_ (.Y(_0152_),
    .A(_0151_),
    .B(net88));
 sg13g2_inv_1 _4022_ (.Y(_0153_),
    .A(net126));
 sg13g2_nor3_1 _4023_ (.A(net109),
    .B(_0153_),
    .C(_2848_),
    .Y(_0154_));
 sg13g2_nor2_1 _4024_ (.A(net62),
    .B(_0154_),
    .Y(_0155_));
 sg13g2_nand2_1 _4025_ (.Y(_0156_),
    .A(_3007_),
    .B(_2550_));
 sg13g2_nand2_1 _4026_ (.Y(_0157_),
    .A(_0155_),
    .B(_0156_));
 sg13g2_nand3_1 _4027_ (.B(_0152_),
    .C(_0157_),
    .A(_0147_),
    .Y(_0158_));
 sg13g2_nand2_1 _4028_ (.Y(_0159_),
    .A(_0158_),
    .B(net131));
 sg13g2_nand2_2 _4029_ (.Y(_0160_),
    .A(_2710_),
    .B(net109));
 sg13g2_buf_1 _4030_ (.A(net149),
    .X(_0161_));
 sg13g2_nand3_1 _4031_ (.B(net67),
    .C(net176),
    .A(_0160_),
    .Y(_0162_));
 sg13g2_inv_2 _4032_ (.Y(_0163_),
    .A(net105));
 sg13g2_a21oi_1 _4033_ (.A1(_0108_),
    .A2(_2715_),
    .Y(_0164_),
    .B1(net35));
 sg13g2_buf_1 _4034_ (.A(_2141_),
    .X(_0165_));
 sg13g2_nor2_1 _4035_ (.A(net182),
    .B(_3029_),
    .Y(_0166_));
 sg13g2_buf_2 _4036_ (.A(_0166_),
    .X(_0167_));
 sg13g2_a21oi_2 _4037_ (.B1(net155),
    .Y(_0168_),
    .A2(_1435_),
    .A1(net206));
 sg13g2_nand3_1 _4038_ (.B(net51),
    .C(net133),
    .A(_0168_),
    .Y(_0169_));
 sg13g2_o21ai_1 _4039_ (.B1(_0169_),
    .Y(_0170_),
    .A1(_0167_),
    .A2(_1816_));
 sg13g2_a22oi_1 _4040_ (.Y(_0171_),
    .B1(net115),
    .B2(_0170_),
    .A2(_0164_),
    .A1(_0162_));
 sg13g2_nand2_1 _4041_ (.Y(_0172_),
    .A(_0159_),
    .B(_0171_));
 sg13g2_nand2_1 _4042_ (.Y(_0173_),
    .A(_0172_),
    .B(net68));
 sg13g2_nand2_2 _4043_ (.Y(_0174_),
    .A(_2871_),
    .B(_2436_));
 sg13g2_nand2_1 _4044_ (.Y(_0175_),
    .A(_2525_),
    .B(net93));
 sg13g2_nand2_1 _4045_ (.Y(_0176_),
    .A(_0174_),
    .B(_0175_));
 sg13g2_nand2_1 _4046_ (.Y(_0177_),
    .A(_0176_),
    .B(_2509_));
 sg13g2_nand2_1 _4047_ (.Y(_0178_),
    .A(net122),
    .B(net137));
 sg13g2_nand2_1 _4048_ (.Y(_0179_),
    .A(_0178_),
    .B(_2842_));
 sg13g2_a21oi_1 _4049_ (.A1(_0177_),
    .A2(_0179_),
    .Y(_0180_),
    .B1(net81));
 sg13g2_buf_8 _4050_ (.A(_2086_),
    .X(_0181_));
 sg13g2_nand3_1 _4051_ (.B(net79),
    .C(net43),
    .A(_0181_),
    .Y(_0182_));
 sg13g2_nand3_1 _4052_ (.B(net129),
    .C(_0140_),
    .A(_0182_),
    .Y(_0183_));
 sg13g2_nand2_1 _4053_ (.Y(_0184_),
    .A(_2819_),
    .B(_1696_));
 sg13g2_nand2_1 _4054_ (.Y(_0185_),
    .A(_2273_),
    .B(_1227_));
 sg13g2_nand2_1 _4055_ (.Y(_0186_),
    .A(_0184_),
    .B(_0185_));
 sg13g2_nand2_1 _4056_ (.Y(_0187_),
    .A(_0186_),
    .B(net142));
 sg13g2_nand2_1 _4057_ (.Y(_0188_),
    .A(_0183_),
    .B(_0187_));
 sg13g2_nor2_1 _4058_ (.A(_0180_),
    .B(_0188_),
    .Y(_0189_));
 sg13g2_nor2_1 _4059_ (.A(net63),
    .B(_0189_),
    .Y(_0190_));
 sg13g2_a21oi_1 _4060_ (.A1(net43),
    .A2(net85),
    .Y(_0191_),
    .B1(net150));
 sg13g2_nand2_1 _4061_ (.Y(_0192_),
    .A(_3008_),
    .B(_0191_));
 sg13g2_nor2_1 _4062_ (.A(net198),
    .B(_3005_),
    .Y(_0193_));
 sg13g2_o21ai_1 _4063_ (.B1(_0193_),
    .Y(_0194_),
    .A1(net48),
    .A2(_2674_));
 sg13g2_nand2_1 _4064_ (.Y(_0195_),
    .A(_0192_),
    .B(_0194_));
 sg13g2_nand2_1 _4065_ (.Y(_0196_),
    .A(_0195_),
    .B(net24));
 sg13g2_nand2_1 _4066_ (.Y(_0197_),
    .A(net137),
    .B(_0790_));
 sg13g2_inv_1 _4067_ (.Y(_0198_),
    .A(_0197_));
 sg13g2_nor2_1 _4068_ (.A(_2475_),
    .B(_0198_),
    .Y(_0199_));
 sg13g2_nor3_1 _4069_ (.A(net28),
    .B(_0199_),
    .C(_2574_),
    .Y(_0200_));
 sg13g2_a21oi_1 _4070_ (.A1(_2571_),
    .A2(net82),
    .Y(_0201_),
    .B1(net150));
 sg13g2_nand2_1 _4071_ (.Y(_0202_),
    .A(_0201_),
    .B(_1968_));
 sg13g2_nand2_1 _4072_ (.Y(_0203_),
    .A(_0202_),
    .B(_2559_));
 sg13g2_nor2_1 _4073_ (.A(_0200_),
    .B(_0203_),
    .Y(_0204_));
 sg13g2_nand2_1 _4074_ (.Y(_0205_),
    .A(_0196_),
    .B(_0204_));
 sg13g2_nand2_1 _4075_ (.Y(_0206_),
    .A(_0205_),
    .B(_2423_));
 sg13g2_nor2_1 _4076_ (.A(_0190_),
    .B(_0206_),
    .Y(_0207_));
 sg13g2_nand2_1 _4077_ (.Y(_0208_),
    .A(_0173_),
    .B(_0207_));
 sg13g2_inv_1 _4078_ (.Y(_0209_),
    .A(_0143_));
 sg13g2_nand2_1 _4079_ (.Y(_0210_),
    .A(_0209_),
    .B(_1446_));
 sg13g2_nand2_1 _4080_ (.Y(_0211_),
    .A(_2967_),
    .B(net60));
 sg13g2_nand2_1 _4081_ (.Y(_0212_),
    .A(_0210_),
    .B(_0211_));
 sg13g2_nand2_1 _4082_ (.Y(_0213_),
    .A(_0212_),
    .B(net129));
 sg13g2_nor2_1 _4083_ (.A(_1511_),
    .B(_0976_),
    .Y(_0214_));
 sg13g2_nand2_1 _4084_ (.Y(_0215_),
    .A(_0149_),
    .B(_0214_));
 sg13g2_nand2_1 _4085_ (.Y(_0216_),
    .A(_2835_),
    .B(_0215_));
 sg13g2_nand2_1 _4086_ (.Y(_0217_),
    .A(_0216_),
    .B(net49));
 sg13g2_nand2_1 _4087_ (.Y(_0218_),
    .A(_0213_),
    .B(_0217_));
 sg13g2_nand2_2 _4088_ (.Y(_0219_),
    .A(_2812_),
    .B(net106));
 sg13g2_buf_1 _4089_ (.A(net177),
    .X(_0220_));
 sg13g2_a21oi_2 _4090_ (.B1(net114),
    .Y(_0221_),
    .A2(net156),
    .A1(_0219_));
 sg13g2_nand2_1 _4091_ (.Y(_0222_),
    .A(net34),
    .B(net87));
 sg13g2_nand2_1 _4092_ (.Y(_0223_),
    .A(_0222_),
    .B(_2402_));
 sg13g2_nor2_1 _4093_ (.A(net60),
    .B(net44),
    .Y(_0224_));
 sg13g2_nor2_1 _4094_ (.A(_1544_),
    .B(_2511_),
    .Y(_0225_));
 sg13g2_inv_1 _4095_ (.Y(_0226_),
    .A(_2467_));
 sg13g2_nand2_1 _4096_ (.Y(_0227_),
    .A(_0225_),
    .B(_0226_));
 sg13g2_o21ai_1 _4097_ (.B1(net171),
    .Y(_0228_),
    .A1(_0224_),
    .A2(_0227_));
 sg13g2_a21oi_1 _4098_ (.A1(_0221_),
    .A2(_0223_),
    .Y(_0229_),
    .B1(_0228_));
 sg13g2_nor2_1 _4099_ (.A(_0218_),
    .B(_0229_),
    .Y(_0230_));
 sg13g2_nor2_1 _4100_ (.A(net63),
    .B(_0230_),
    .Y(_0231_));
 sg13g2_nor2_1 _4101_ (.A(_2407_),
    .B(_2678_),
    .Y(_0232_));
 sg13g2_nand2_1 _4102_ (.Y(_0233_),
    .A(_2624_),
    .B(_2709_));
 sg13g2_buf_2 _4103_ (.A(_0233_),
    .X(_0234_));
 sg13g2_a21oi_1 _4104_ (.A1(_2752_),
    .A2(_2605_),
    .Y(_0235_),
    .B1(_1326_));
 sg13g2_a21oi_1 _4105_ (.A1(_0232_),
    .A2(_0234_),
    .Y(_0236_),
    .B1(_0235_));
 sg13g2_nand2_1 _4106_ (.Y(_0237_),
    .A(_2428_),
    .B(_2430_));
 sg13g2_nand2_1 _4107_ (.Y(_0238_),
    .A(_0237_),
    .B(net49));
 sg13g2_nand3_1 _4108_ (.B(_2495_),
    .C(net141),
    .A(_2778_),
    .Y(_0239_));
 sg13g2_nand2_1 _4109_ (.Y(_0240_),
    .A(net43),
    .B(net85));
 sg13g2_nand2_1 _4110_ (.Y(_0241_),
    .A(_0239_),
    .B(_0240_));
 sg13g2_nand2_1 _4111_ (.Y(_0242_),
    .A(_0241_),
    .B(net88));
 sg13g2_nand3_1 _4112_ (.B(_0238_),
    .C(_0242_),
    .A(_0236_),
    .Y(_0243_));
 sg13g2_nand2_1 _4113_ (.Y(_0244_),
    .A(_0243_),
    .B(_2559_));
 sg13g2_nand2_1 _4114_ (.Y(_0245_),
    .A(_0244_),
    .B(net170));
 sg13g2_nor2_1 _4115_ (.A(_0231_),
    .B(_0245_),
    .Y(_0246_));
 sg13g2_a21oi_1 _4116_ (.A1(_0099_),
    .A2(net143),
    .Y(_0247_),
    .B1(net135));
 sg13g2_nand2_1 _4117_ (.Y(_0248_),
    .A(_0247_),
    .B(_2910_));
 sg13g2_a21oi_1 _4118_ (.A1(_2529_),
    .A2(_0142_),
    .Y(_0249_),
    .B1(_2162_));
 sg13g2_nand2_2 _4119_ (.Y(_0250_),
    .A(_2582_),
    .B(_1227_));
 sg13g2_nand2_1 _4120_ (.Y(_0251_),
    .A(_0249_),
    .B(_0250_));
 sg13g2_nand3_1 _4121_ (.B(_0251_),
    .C(net168),
    .A(_0248_),
    .Y(_0252_));
 sg13g2_nand2_1 _4122_ (.Y(_0253_),
    .A(_2965_),
    .B(_0197_));
 sg13g2_nand3_1 _4123_ (.B(_0149_),
    .C(net104),
    .A(_0253_),
    .Y(_0254_));
 sg13g2_and2_1 _4124_ (.A(_0254_),
    .B(_2483_),
    .X(_0255_));
 sg13g2_nand2_1 _4125_ (.Y(_0256_),
    .A(_0252_),
    .B(_0255_));
 sg13g2_nand2_1 _4126_ (.Y(_0257_),
    .A(_0256_),
    .B(net80));
 sg13g2_inv_1 _4127_ (.Y(_0258_),
    .A(_2031_));
 sg13g2_a21oi_1 _4128_ (.A1(_0258_),
    .A2(net48),
    .Y(_0259_),
    .B1(net114));
 sg13g2_nand2_2 _4129_ (.Y(_0260_),
    .A(_2526_),
    .B(net146));
 sg13g2_nor2_1 _4130_ (.A(net75),
    .B(_0260_),
    .Y(_0261_));
 sg13g2_o21ai_1 _4131_ (.B1(_0261_),
    .Y(_0262_),
    .A1(_1968_),
    .A2(_0259_));
 sg13g2_o21ai_1 _4132_ (.B1(_2688_),
    .Y(_0263_),
    .A1(_2905_),
    .A2(net34));
 sg13g2_nor2_1 _4133_ (.A(net141),
    .B(_2494_),
    .Y(_0264_));
 sg13g2_o21ai_1 _4134_ (.B1(net135),
    .Y(_0265_),
    .A1(net29),
    .A2(_0264_));
 sg13g2_nor2_2 _4135_ (.A(_2964_),
    .B(net122),
    .Y(_0266_));
 sg13g2_nand2_1 _4136_ (.Y(_0267_),
    .A(_0266_),
    .B(net177));
 sg13g2_nand2_1 _4137_ (.Y(_0268_),
    .A(_0265_),
    .B(_0267_));
 sg13g2_nor2_1 _4138_ (.A(_0263_),
    .B(_0268_),
    .Y(_0269_));
 sg13g2_nor2_1 _4139_ (.A(net123),
    .B(_0269_),
    .Y(_0270_));
 sg13g2_nand2_1 _4140_ (.Y(_0271_),
    .A(_0262_),
    .B(_0270_));
 sg13g2_nand2_1 _4141_ (.Y(_0272_),
    .A(_0257_),
    .B(_0271_));
 sg13g2_nand2_1 _4142_ (.Y(_0273_),
    .A(_0272_),
    .B(net68));
 sg13g2_nand2_1 _4143_ (.Y(_0274_),
    .A(_0246_),
    .B(_0273_));
 sg13g2_nand3_1 _4144_ (.B(_0274_),
    .C(net165),
    .A(_0208_),
    .Y(_0275_));
 sg13g2_nand2_1 _4145_ (.Y(_0276_),
    .A(_2532_),
    .B(net176));
 sg13g2_nand2_1 _4146_ (.Y(_0277_),
    .A(_0149_),
    .B(_0276_));
 sg13g2_nand2_2 _4147_ (.Y(_0278_),
    .A(_2930_),
    .B(_1511_));
 sg13g2_nand3_1 _4148_ (.B(_0278_),
    .C(_0220_),
    .A(_0277_),
    .Y(_0279_));
 sg13g2_nand2_1 _4149_ (.Y(_0280_),
    .A(_0279_),
    .B(_0177_));
 sg13g2_nand2_1 _4150_ (.Y(_0281_),
    .A(_0280_),
    .B(net46));
 sg13g2_inv_1 _4151_ (.Y(_0282_),
    .A(_0260_));
 sg13g2_nand2_1 _4152_ (.Y(_0283_),
    .A(_2660_),
    .B(net52));
 sg13g2_a21oi_1 _4153_ (.A1(_0282_),
    .A2(_0283_),
    .Y(_0284_),
    .B1(net138));
 sg13g2_nand2_1 _4154_ (.Y(_0285_),
    .A(_2900_),
    .B(_2997_));
 sg13g2_a21oi_1 _4155_ (.A1(_2617_),
    .A2(_0285_),
    .Y(_0286_),
    .B1(_2533_));
 sg13g2_nor3_1 _4156_ (.A(net127),
    .B(_0284_),
    .C(_0286_),
    .Y(_0287_));
 sg13g2_a21oi_1 _4157_ (.A1(_0281_),
    .A2(_0287_),
    .Y(_0288_),
    .B1(net166));
 sg13g2_nand2_2 _4158_ (.Y(_0289_),
    .A(_0900_),
    .B(_1911_));
 sg13g2_o21ai_1 _4159_ (.B1(_2506_),
    .Y(_0290_),
    .A1(_1478_),
    .A2(_0289_));
 sg13g2_nand2_1 _4160_ (.Y(_0291_),
    .A(_2119_),
    .B(_0290_));
 sg13g2_nand2_1 _4161_ (.Y(_0292_),
    .A(_2890_),
    .B(_3012_));
 sg13g2_a22oi_1 _4162_ (.Y(_0293_),
    .B1(net26),
    .B2(_0292_),
    .A2(_2882_),
    .A1(_0291_));
 sg13g2_buf_1 _4163_ (.A(net64),
    .X(_0294_));
 sg13g2_a21oi_1 _4164_ (.A1(_2119_),
    .A2(_2572_),
    .Y(_0295_),
    .B1(net23));
 sg13g2_nand2_1 _4165_ (.Y(_0296_),
    .A(_2830_),
    .B(_2589_));
 sg13g2_nand2_1 _4166_ (.Y(_0297_),
    .A(_0174_),
    .B(_0296_));
 sg13g2_a21oi_1 _4167_ (.A1(_0297_),
    .A2(_2895_),
    .Y(_0298_),
    .B1(_2595_));
 sg13g2_nor2b_1 _4168_ (.A(_0295_),
    .B_N(_0298_),
    .Y(_0299_));
 sg13g2_nand2_1 _4169_ (.Y(_0300_),
    .A(_0293_),
    .B(_0299_));
 sg13g2_nand2_1 _4170_ (.Y(_0301_),
    .A(_0288_),
    .B(_0300_));
 sg13g2_a21oi_2 _4171_ (.B1(net149),
    .Y(_0302_),
    .A2(_2633_),
    .A1(net103));
 sg13g2_nand2_2 _4172_ (.Y(_0303_),
    .A(_2691_),
    .B(_0034_));
 sg13g2_a221oi_1 _4173_ (.B2(_0302_),
    .C1(_0303_),
    .B1(_0169_),
    .A1(_0167_),
    .Y(_0304_),
    .A2(_1880_));
 sg13g2_nor2_1 _4174_ (.A(net170),
    .B(_0304_),
    .Y(_0305_));
 sg13g2_a21oi_1 _4175_ (.A1(_0301_),
    .A2(_0305_),
    .Y(_0306_),
    .B1(net165));
 sg13g2_a21oi_1 _4176_ (.A1(_2803_),
    .A2(_0285_),
    .Y(_0307_),
    .B1(net23));
 sg13g2_a21oi_1 _4177_ (.A1(_2746_),
    .A2(_2747_),
    .Y(_0308_),
    .B1(net28));
 sg13g2_inv_1 _4178_ (.Y(_0309_),
    .A(_2960_));
 sg13g2_nand3b_1 _4179_ (.B(net134),
    .C(_0309_),
    .Y(_0310_),
    .A_N(_2470_));
 sg13g2_nand2_1 _4180_ (.Y(_0311_),
    .A(_2440_),
    .B(net177));
 sg13g2_o21ai_1 _4181_ (.B1(_0311_),
    .Y(_0312_),
    .A1(_1998_),
    .A2(net47));
 sg13g2_nand2_1 _4182_ (.Y(_0313_),
    .A(_0312_),
    .B(net171));
 sg13g2_nand3b_1 _4183_ (.B(_0310_),
    .C(_0313_),
    .Y(_0314_),
    .A_N(_0308_));
 sg13g2_nor2_1 _4184_ (.A(_0307_),
    .B(_0314_),
    .Y(_0315_));
 sg13g2_nor2_1 _4185_ (.A(net118),
    .B(_0315_),
    .Y(_0316_));
 sg13g2_nor2_1 _4186_ (.A(net200),
    .B(_0316_),
    .Y(_0317_));
 sg13g2_nand2_1 _4187_ (.Y(_0318_),
    .A(_2086_),
    .B(net140));
 sg13g2_nand2_1 _4188_ (.Y(_0319_),
    .A(_2704_),
    .B(_2550_));
 sg13g2_nand2_1 _4189_ (.Y(_0320_),
    .A(_0318_),
    .B(_0319_));
 sg13g2_nor2_2 _4190_ (.A(net29),
    .B(_2713_),
    .Y(_0321_));
 sg13g2_o21ai_1 _4191_ (.B1(_0321_),
    .Y(_0322_),
    .A1(_2494_),
    .A2(_0143_));
 sg13g2_a22oi_1 _4192_ (.Y(_0323_),
    .B1(net25),
    .B2(_0322_),
    .A2(net53),
    .A1(_0320_));
 sg13g2_a21oi_2 _4193_ (.B1(_2589_),
    .Y(_0324_),
    .A2(net94),
    .A1(_2622_));
 sg13g2_o21ai_1 _4194_ (.B1(_2968_),
    .Y(_0325_),
    .A1(_2955_),
    .A2(_0324_));
 sg13g2_buf_1 _4195_ (.A(_2711_),
    .X(_0326_));
 sg13g2_nor2_1 _4196_ (.A(net33),
    .B(_2525_),
    .Y(_0327_));
 sg13g2_o21ai_1 _4197_ (.B1(net70),
    .Y(_0328_),
    .A1(_0327_),
    .A2(_2948_));
 sg13g2_nand3_1 _4198_ (.B(_0325_),
    .C(_0328_),
    .A(_0323_),
    .Y(_0329_));
 sg13g2_nand2_1 _4199_ (.Y(_0330_),
    .A(_0329_),
    .B(_2373_));
 sg13g2_nand3_1 _4200_ (.B(_2895_),
    .C(_0174_),
    .A(_2870_),
    .Y(_0331_));
 sg13g2_nand2_2 _4201_ (.Y(_0332_),
    .A(net87),
    .B(net141));
 sg13g2_nand2_1 _4202_ (.Y(_0333_),
    .A(_2892_),
    .B(_0332_));
 sg13g2_buf_2 _4203_ (.A(net69),
    .X(_0334_));
 sg13g2_nand3_1 _4204_ (.B(_0333_),
    .C(net32),
    .A(_0150_),
    .Y(_0335_));
 sg13g2_a21oi_1 _4205_ (.A1(_0331_),
    .A2(_0335_),
    .Y(_0336_),
    .B1(_2596_));
 sg13g2_inv_1 _4206_ (.Y(_0337_),
    .A(_2141_));
 sg13g2_buf_1 _4207_ (.A(_0337_),
    .X(_0338_));
 sg13g2_nand2_1 _4208_ (.Y(_0339_),
    .A(_2671_),
    .B(_2947_));
 sg13g2_nor2_1 _4209_ (.A(net48),
    .B(_0339_),
    .Y(_0340_));
 sg13g2_nand2_1 _4210_ (.Y(_0341_),
    .A(_0234_),
    .B(net114));
 sg13g2_nor2_1 _4211_ (.A(_0340_),
    .B(_0341_),
    .Y(_0342_));
 sg13g2_nor2_1 _4212_ (.A(net66),
    .B(_0342_),
    .Y(_0343_));
 sg13g2_nand2_1 _4213_ (.Y(_0344_),
    .A(_2436_),
    .B(net141));
 sg13g2_nand2_1 _4214_ (.Y(_0345_),
    .A(_3018_),
    .B(_0344_));
 sg13g2_nor2_2 _4215_ (.A(_1216_),
    .B(net59),
    .Y(_0346_));
 sg13g2_nand2_1 _4216_ (.Y(_0347_),
    .A(_0346_),
    .B(_2947_));
 sg13g2_nand3_1 _4217_ (.B(_0347_),
    .C(_3023_),
    .A(_0345_),
    .Y(_0348_));
 sg13g2_a21oi_1 _4218_ (.A1(_0343_),
    .A2(_0348_),
    .Y(_0349_),
    .B1(net166));
 sg13g2_nand2_2 _4219_ (.Y(_0350_),
    .A(_2800_),
    .B(_2525_));
 sg13g2_nand2_1 _4220_ (.Y(_0351_),
    .A(_0350_),
    .B(net27));
 sg13g2_nor2_1 _4221_ (.A(_1751_),
    .B(_2751_),
    .Y(_0352_));
 sg13g2_nand2_1 _4222_ (.Y(_0353_),
    .A(_0351_),
    .B(_0352_));
 sg13g2_nand2_1 _4223_ (.Y(_0354_),
    .A(_2616_),
    .B(net95));
 sg13g2_nand2_1 _4224_ (.Y(_0355_),
    .A(_0354_),
    .B(_0167_));
 sg13g2_nand3_1 _4225_ (.B(_0355_),
    .C(net130),
    .A(_0353_),
    .Y(_0356_));
 sg13g2_nor2_1 _4226_ (.A(net101),
    .B(_0266_),
    .Y(_0357_));
 sg13g2_a21oi_1 _4227_ (.A1(_2969_),
    .A2(net104),
    .Y(_0358_),
    .B1(net173));
 sg13g2_nand2_1 _4228_ (.Y(_0359_),
    .A(_1795_),
    .B(_1184_));
 sg13g2_nor2_2 _4229_ (.A(_2543_),
    .B(_1998_),
    .Y(_0360_));
 sg13g2_nand2_1 _4230_ (.Y(_0361_),
    .A(_0359_),
    .B(_0360_));
 sg13g2_nand2_1 _4231_ (.Y(_0362_),
    .A(_0358_),
    .B(_0361_));
 sg13g2_a21oi_1 _4232_ (.A1(_0160_),
    .A2(_0357_),
    .Y(_0363_),
    .B1(_0362_));
 sg13g2_nand2_1 _4233_ (.Y(_0364_),
    .A(_0356_),
    .B(_0363_));
 sg13g2_nand3b_1 _4234_ (.B(_0349_),
    .C(_0364_),
    .Y(_0365_),
    .A_N(_0336_));
 sg13g2_nand3_1 _4235_ (.B(_0330_),
    .C(_0365_),
    .A(_0317_),
    .Y(_0366_));
 sg13g2_nand2_1 _4236_ (.Y(_0367_),
    .A(_0306_),
    .B(_0366_));
 sg13g2_nand2_1 _4237_ (.Y(_0023_),
    .A(_0275_),
    .B(_0367_));
 sg13g2_nor2_1 _4238_ (.A(net128),
    .B(_2602_),
    .Y(_0368_));
 sg13g2_a21oi_1 _4239_ (.A1(_0150_),
    .A2(_0368_),
    .Y(_0369_),
    .B1(net162));
 sg13g2_nand2_2 _4240_ (.Y(_0370_),
    .A(_2086_),
    .B(net97));
 sg13g2_nand2_1 _4241_ (.Y(_0371_),
    .A(_0370_),
    .B(net27));
 sg13g2_inv_1 _4242_ (.Y(_0372_),
    .A(_2813_));
 sg13g2_nor2_1 _4243_ (.A(net37),
    .B(_0372_),
    .Y(_0373_));
 sg13g2_nand2_1 _4244_ (.Y(_0374_),
    .A(_0371_),
    .B(_0373_));
 sg13g2_nand2_1 _4245_ (.Y(_0375_),
    .A(_0369_),
    .B(_0374_));
 sg13g2_nand2_1 _4246_ (.Y(_0376_),
    .A(net126),
    .B(net153));
 sg13g2_nand2_1 _4247_ (.Y(_0377_),
    .A(_0376_),
    .B(_2488_));
 sg13g2_nand2_1 _4248_ (.Y(_0378_),
    .A(_0377_),
    .B(net27));
 sg13g2_nand3_1 _4249_ (.B(_2614_),
    .C(net45),
    .A(_0378_),
    .Y(_0379_));
 sg13g2_nand3_1 _4250_ (.B(net198),
    .C(_2020_),
    .A(_0276_),
    .Y(_0380_));
 sg13g2_nand2_1 _4251_ (.Y(_0381_),
    .A(_0380_),
    .B(_2643_));
 sg13g2_nand2_1 _4252_ (.Y(_0382_),
    .A(_0379_),
    .B(_0381_));
 sg13g2_a21oi_1 _4253_ (.A1(_0375_),
    .A2(_0382_),
    .Y(_0383_),
    .B1(_2816_));
 sg13g2_nor2_1 _4254_ (.A(_1326_),
    .B(_0260_),
    .Y(_0384_));
 sg13g2_nand2_1 _4255_ (.Y(_0385_),
    .A(_0160_),
    .B(_0384_));
 sg13g2_nand2_1 _4256_ (.Y(_0386_),
    .A(_0385_),
    .B(_2373_));
 sg13g2_nand2_2 _4257_ (.Y(_0387_),
    .A(_2582_),
    .B(net29));
 sg13g2_nand2_1 _4258_ (.Y(_0388_),
    .A(_2582_),
    .B(_0214_));
 sg13g2_nand3_1 _4259_ (.B(_0388_),
    .C(_2935_),
    .A(_0387_),
    .Y(_0389_));
 sg13g2_nor2b_1 _4260_ (.A(_0386_),
    .B_N(_0389_),
    .Y(_0390_));
 sg13g2_a21oi_1 _4261_ (.A1(_0214_),
    .A2(_1859_),
    .Y(_0391_),
    .B1(net174));
 sg13g2_nand2_1 _4262_ (.Y(_0392_),
    .A(_3043_),
    .B(_0391_));
 sg13g2_nand2_1 _4263_ (.Y(_0393_),
    .A(net144),
    .B(_2477_));
 sg13g2_nand2_1 _4264_ (.Y(_0394_),
    .A(_0393_),
    .B(_2745_));
 sg13g2_nor2_1 _4265_ (.A(_1555_),
    .B(_2387_),
    .Y(_0395_));
 sg13g2_nand2_1 _4266_ (.Y(_0396_),
    .A(_0394_),
    .B(_0395_));
 sg13g2_nand2_1 _4267_ (.Y(_0397_),
    .A(_0392_),
    .B(_0396_));
 sg13g2_nand2_1 _4268_ (.Y(_0398_),
    .A(_0397_),
    .B(net46));
 sg13g2_nand2_1 _4269_ (.Y(_0399_),
    .A(_0390_),
    .B(_0398_));
 sg13g2_nand2_1 _4270_ (.Y(_0400_),
    .A(_0399_),
    .B(_2423_));
 sg13g2_nor2_1 _4271_ (.A(_0383_),
    .B(_0400_),
    .Y(_0401_));
 sg13g2_nand2_1 _4272_ (.Y(_0402_),
    .A(_2833_),
    .B(_2399_));
 sg13g2_nand2_1 _4273_ (.Y(_0403_),
    .A(_0402_),
    .B(net27));
 sg13g2_inv_1 _4274_ (.Y(_0404_),
    .A(_2525_));
 sg13g2_nand2_2 _4275_ (.Y(_0405_),
    .A(_0404_),
    .B(net79));
 sg13g2_a21oi_1 _4276_ (.A1(_0403_),
    .A2(_0405_),
    .Y(_0406_),
    .B1(net23));
 sg13g2_a21oi_1 _4277_ (.A1(_3043_),
    .A2(_0277_),
    .Y(_0407_),
    .B1(net145));
 sg13g2_nor2_1 _4278_ (.A(_0406_),
    .B(_0407_),
    .Y(_0408_));
 sg13g2_nand2_1 _4279_ (.Y(_0409_),
    .A(_2889_),
    .B(_2097_));
 sg13g2_nand2_1 _4280_ (.Y(_0410_),
    .A(_0409_),
    .B(_2977_));
 sg13g2_nand2_1 _4281_ (.Y(_0411_),
    .A(_0410_),
    .B(_2882_));
 sg13g2_nand3_1 _4282_ (.B(_2416_),
    .C(_2413_),
    .A(net57),
    .Y(_0412_));
 sg13g2_nand2_1 _4283_ (.Y(_0413_),
    .A(_0412_),
    .B(_0100_));
 sg13g2_nand2_1 _4284_ (.Y(_0414_),
    .A(_0413_),
    .B(_2968_));
 sg13g2_nand3_1 _4285_ (.B(_0411_),
    .C(_0414_),
    .A(_0408_),
    .Y(_0415_));
 sg13g2_nor2_1 _4286_ (.A(_2646_),
    .B(_2665_),
    .Y(_0416_));
 sg13g2_nand2_1 _4287_ (.Y(_0417_),
    .A(_0415_),
    .B(_0416_));
 sg13g2_inv_1 _4288_ (.Y(_0418_),
    .A(_2900_));
 sg13g2_nand3_1 _4289_ (.B(net37),
    .C(_0418_),
    .A(net34),
    .Y(_0419_));
 sg13g2_nand2_1 _4290_ (.Y(_0420_),
    .A(_2988_),
    .B(_2842_));
 sg13g2_nor2_1 _4291_ (.A(net184),
    .B(_1544_),
    .Y(_0421_));
 sg13g2_buf_2 _4292_ (.A(_0421_),
    .X(_0422_));
 sg13g2_nand2_1 _4293_ (.Y(_0423_),
    .A(_0178_),
    .B(_0422_));
 sg13g2_nand3_1 _4294_ (.B(_0420_),
    .C(_0423_),
    .A(_0419_),
    .Y(_0424_));
 sg13g2_nand2_1 _4295_ (.Y(_0425_),
    .A(_0424_),
    .B(_0165_));
 sg13g2_a21oi_1 _4296_ (.A1(_1609_),
    .A2(net141),
    .Y(_0426_),
    .B1(_2575_));
 sg13g2_nor2_1 _4297_ (.A(net33),
    .B(_0426_),
    .Y(_0427_));
 sg13g2_nand2_1 _4298_ (.Y(_0428_),
    .A(net103),
    .B(_1162_));
 sg13g2_nand2_1 _4299_ (.Y(_0429_),
    .A(_2730_),
    .B(_0428_));
 sg13g2_nand2_1 _4300_ (.Y(_0430_),
    .A(_2871_),
    .B(_2860_));
 sg13g2_a21oi_1 _4301_ (.A1(_2724_),
    .A2(_0430_),
    .Y(_0431_),
    .B1(net35));
 sg13g2_o21ai_1 _4302_ (.B1(_0431_),
    .Y(_0432_),
    .A1(_0427_),
    .A2(_0429_));
 sg13g2_nand2_1 _4303_ (.Y(_0433_),
    .A(_0425_),
    .B(_0432_));
 sg13g2_nand2_1 _4304_ (.Y(_0434_),
    .A(_0433_),
    .B(_2785_));
 sg13g2_nand3_1 _4305_ (.B(_0417_),
    .C(_0434_),
    .A(_0401_),
    .Y(_0435_));
 sg13g2_nand2_1 _4306_ (.Y(_0436_),
    .A(_0370_),
    .B(_2842_));
 sg13g2_a21oi_1 _4307_ (.A1(_2983_),
    .A2(_3003_),
    .Y(_0437_),
    .B1(net35));
 sg13g2_nor2_2 _4308_ (.A(_0932_),
    .B(net178),
    .Y(_0438_));
 sg13g2_inv_1 _4309_ (.Y(_0439_),
    .A(_0438_));
 sg13g2_nand3_1 _4310_ (.B(net114),
    .C(_0439_),
    .A(_2986_),
    .Y(_0440_));
 sg13g2_nand3_1 _4311_ (.B(_0437_),
    .C(_0440_),
    .A(_0436_),
    .Y(_0441_));
 sg13g2_nand2_1 _4312_ (.Y(_0442_),
    .A(_0441_),
    .B(net175));
 sg13g2_nand3_1 _4313_ (.B(net111),
    .C(net158),
    .A(_2669_),
    .Y(_0443_));
 sg13g2_nand2_1 _4314_ (.Y(_0444_),
    .A(_0443_),
    .B(_2430_));
 sg13g2_a21oi_1 _4315_ (.A1(_0444_),
    .A2(net134),
    .Y(_0445_),
    .B1(_2480_));
 sg13g2_nand3_1 _4316_ (.B(net77),
    .C(net97),
    .A(_2622_),
    .Y(_0446_));
 sg13g2_nand2_1 _4317_ (.Y(_0447_),
    .A(_0446_),
    .B(_2867_));
 sg13g2_nand2_1 _4318_ (.Y(_0448_),
    .A(_0445_),
    .B(_0447_));
 sg13g2_nor2b_1 _4319_ (.A(_0107_),
    .B_N(_2992_),
    .Y(_0449_));
 sg13g2_nor2_1 _4320_ (.A(net114),
    .B(_0449_),
    .Y(_0450_));
 sg13g2_nand2_1 _4321_ (.Y(_0451_),
    .A(_2942_),
    .B(net56));
 sg13g2_nor2_1 _4322_ (.A(_2641_),
    .B(net90),
    .Y(_0452_));
 sg13g2_nor2_2 _4323_ (.A(net182),
    .B(_2453_),
    .Y(_0453_));
 sg13g2_nor2_1 _4324_ (.A(net150),
    .B(_0453_),
    .Y(_0454_));
 sg13g2_nor2_1 _4325_ (.A(_0452_),
    .B(_0454_),
    .Y(_0455_));
 sg13g2_a21oi_1 _4326_ (.A1(_0450_),
    .A2(_0451_),
    .Y(_0456_),
    .B1(_0455_));
 sg13g2_nor2_1 _4327_ (.A(_0448_),
    .B(_0456_),
    .Y(_0457_));
 sg13g2_nor2_1 _4328_ (.A(_0442_),
    .B(_0457_),
    .Y(_0458_));
 sg13g2_nand3_1 _4329_ (.B(net72),
    .C(_0405_),
    .A(_2119_),
    .Y(_0459_));
 sg13g2_nor2_1 _4330_ (.A(net149),
    .B(_2537_),
    .Y(_0460_));
 sg13g2_nand2_1 _4331_ (.Y(_0461_),
    .A(_0460_),
    .B(_2920_));
 sg13g2_nand2_1 _4332_ (.Y(_0462_),
    .A(_0459_),
    .B(_0461_));
 sg13g2_nand2_1 _4333_ (.Y(_0463_),
    .A(_0462_),
    .B(net115));
 sg13g2_nand2_1 _4334_ (.Y(_0464_),
    .A(_0458_),
    .B(_0463_));
 sg13g2_nand2_1 _4335_ (.Y(_0465_),
    .A(_3043_),
    .B(_2879_));
 sg13g2_a21oi_1 _4336_ (.A1(_1948_),
    .A2(_2532_),
    .Y(_0466_),
    .B1(_0294_));
 sg13g2_a21oi_1 _4337_ (.A1(_0465_),
    .A2(_2991_),
    .Y(_0467_),
    .B1(_0466_));
 sg13g2_nand2_1 _4338_ (.Y(_0468_),
    .A(_0987_),
    .B(net111));
 sg13g2_a21o_1 _4339_ (.A2(_0468_),
    .A1(_0215_),
    .B1(_2408_),
    .X(_0469_));
 sg13g2_nand3_1 _4340_ (.B(net136),
    .C(net178),
    .A(_0168_),
    .Y(_0470_));
 sg13g2_nand2_1 _4341_ (.Y(_0471_),
    .A(_2778_),
    .B(net109));
 sg13g2_nand2_1 _4342_ (.Y(_0472_),
    .A(_0470_),
    .B(_0471_));
 sg13g2_nand2_1 _4343_ (.Y(_0473_),
    .A(_0472_),
    .B(net26));
 sg13g2_nand3_1 _4344_ (.B(_0469_),
    .C(_0473_),
    .A(_0467_),
    .Y(_0474_));
 sg13g2_nand2_1 _4345_ (.Y(_0475_),
    .A(_0474_),
    .B(_2373_));
 sg13g2_nor2_1 _4346_ (.A(_1151_),
    .B(_2854_),
    .Y(_0476_));
 sg13g2_buf_2 _4347_ (.A(_0476_),
    .X(_0477_));
 sg13g2_nand2_2 _4348_ (.Y(_0478_),
    .A(_0477_),
    .B(net182));
 sg13g2_o21ai_1 _4349_ (.B1(_0478_),
    .Y(_0479_),
    .A1(_1998_),
    .A2(_2634_));
 sg13g2_nor2_1 _4350_ (.A(_2450_),
    .B(_2916_),
    .Y(_0480_));
 sg13g2_nor2_1 _4351_ (.A(net120),
    .B(_0480_),
    .Y(_0481_));
 sg13g2_nand2_1 _4352_ (.Y(_0482_),
    .A(net210),
    .B(net209));
 sg13g2_buf_2 _4353_ (.A(_0482_),
    .X(_0483_));
 sg13g2_nor2_1 _4354_ (.A(net175),
    .B(net160),
    .Y(_0484_));
 sg13g2_o21ai_1 _4355_ (.B1(_0484_),
    .Y(_0485_),
    .A1(_0479_),
    .A2(_0481_));
 sg13g2_nand2_1 _4356_ (.Y(_0486_),
    .A(_0485_),
    .B(_2564_));
 sg13g2_nand2_2 _4357_ (.Y(_0487_),
    .A(net34),
    .B(_2900_));
 sg13g2_nand2_1 _4358_ (.Y(_0488_),
    .A(_0487_),
    .B(_2715_));
 sg13g2_a21oi_1 _4359_ (.A1(_0185_),
    .A2(net120),
    .Y(_0489_),
    .B1(net162));
 sg13g2_a22oi_1 _4360_ (.Y(_0490_),
    .B1(_0488_),
    .B2(_0489_),
    .A2(_2790_),
    .A1(net25));
 sg13g2_nor2_1 _4361_ (.A(net118),
    .B(_0490_),
    .Y(_0491_));
 sg13g2_nor2_1 _4362_ (.A(_0486_),
    .B(_0491_),
    .Y(_0492_));
 sg13g2_nand3_1 _4363_ (.B(_0475_),
    .C(_0492_),
    .A(_0464_),
    .Y(_0493_));
 sg13g2_nand3_1 _4364_ (.B(_0493_),
    .C(net165),
    .A(_0435_),
    .Y(_0494_));
 sg13g2_nand2_1 _4365_ (.Y(_0495_),
    .A(net100),
    .B(_1184_));
 sg13g2_nand2_1 _4366_ (.Y(_0496_),
    .A(_0495_),
    .B(net60));
 sg13g2_a21oi_1 _4367_ (.A1(_2289_),
    .A2(_0496_),
    .Y(_0497_),
    .B1(net75));
 sg13g2_nand2_1 _4368_ (.Y(_0498_),
    .A(_2538_),
    .B(_2993_));
 sg13g2_nand2_1 _4369_ (.Y(_0499_),
    .A(_0498_),
    .B(_0220_));
 sg13g2_nand2_1 _4370_ (.Y(_0500_),
    .A(_0497_),
    .B(_0499_));
 sg13g2_nor2_1 _4371_ (.A(_2577_),
    .B(_2623_),
    .Y(_0501_));
 sg13g2_nor2_1 _4372_ (.A(_0266_),
    .B(_0501_),
    .Y(_0502_));
 sg13g2_nor2_1 _4373_ (.A(net28),
    .B(_0502_),
    .Y(_0503_));
 sg13g2_nand2_1 _4374_ (.Y(_0504_),
    .A(_2801_),
    .B(net143));
 sg13g2_a21oi_1 _4375_ (.A1(_2959_),
    .A2(_0504_),
    .Y(_0505_),
    .B1(net101));
 sg13g2_nor2_1 _4376_ (.A(_0503_),
    .B(_0505_),
    .Y(_0506_));
 sg13g2_nand2_1 _4377_ (.Y(_0507_),
    .A(_0500_),
    .B(_0506_));
 sg13g2_nand2_1 _4378_ (.Y(_0508_),
    .A(_0507_),
    .B(net80));
 sg13g2_nor2_1 _4379_ (.A(net142),
    .B(_2960_),
    .Y(_0509_));
 sg13g2_nor2_1 _4380_ (.A(net47),
    .B(_2812_),
    .Y(_0510_));
 sg13g2_inv_1 _4381_ (.Y(_0511_),
    .A(net160));
 sg13g2_o21ai_1 _4382_ (.B1(net113),
    .Y(_0512_),
    .A1(net37),
    .A2(_0510_));
 sg13g2_a21oi_1 _4383_ (.A1(_2977_),
    .A2(_0509_),
    .Y(_0513_),
    .B1(_0512_));
 sg13g2_nand2_2 _4384_ (.Y(_0514_),
    .A(_2414_),
    .B(net136));
 sg13g2_nand2_1 _4385_ (.Y(_0515_),
    .A(_0514_),
    .B(net128));
 sg13g2_inv_2 _4386_ (.Y(_0516_),
    .A(_2119_));
 sg13g2_nor2_1 _4387_ (.A(_0515_),
    .B(_0516_),
    .Y(_0517_));
 sg13g2_nand2_1 _4388_ (.Y(_0518_),
    .A(_0282_),
    .B(net108));
 sg13g2_nor2_1 _4389_ (.A(net77),
    .B(_0258_),
    .Y(_0519_));
 sg13g2_inv_1 _4390_ (.Y(_0520_),
    .A(_0118_));
 sg13g2_buf_2 _4391_ (.A(_0520_),
    .X(_0521_));
 sg13g2_o21ai_1 _4392_ (.B1(net22),
    .Y(_0522_),
    .A1(_0518_),
    .A2(_0519_));
 sg13g2_nor2_1 _4393_ (.A(_0517_),
    .B(_0522_),
    .Y(_0523_));
 sg13g2_nor2_1 _4394_ (.A(_0513_),
    .B(_0523_),
    .Y(_0524_));
 sg13g2_nand2_1 _4395_ (.Y(_0525_),
    .A(_0508_),
    .B(_0524_));
 sg13g2_nand2_1 _4396_ (.Y(_0526_),
    .A(_0525_),
    .B(net68));
 sg13g2_nor2_2 _4397_ (.A(net184),
    .B(net158),
    .Y(_0527_));
 sg13g2_inv_1 _4398_ (.Y(_0528_),
    .A(_0527_));
 sg13g2_a21oi_1 _4399_ (.A1(_2478_),
    .A2(_0528_),
    .Y(_0529_),
    .B1(net64));
 sg13g2_buf_2 _4400_ (.A(_2376_),
    .X(_0530_));
 sg13g2_nor2_1 _4401_ (.A(net194),
    .B(_1326_),
    .Y(_0531_));
 sg13g2_buf_1 _4402_ (.A(_0531_),
    .X(_0532_));
 sg13g2_inv_1 _4403_ (.Y(_0533_),
    .A(net65));
 sg13g2_nor2_1 _4404_ (.A(_0533_),
    .B(_2755_),
    .Y(_0534_));
 sg13g2_nor3_1 _4405_ (.A(net167),
    .B(_0529_),
    .C(_0534_),
    .Y(_0535_));
 sg13g2_inv_1 _4406_ (.Y(_0536_),
    .A(_2585_));
 sg13g2_a21oi_1 _4407_ (.A1(_0536_),
    .A2(_2715_),
    .Y(_0537_),
    .B1(net162));
 sg13g2_nor2_1 _4408_ (.A(net89),
    .B(_2547_),
    .Y(_0538_));
 sg13g2_nand2_1 _4409_ (.Y(_0539_),
    .A(_0169_),
    .B(_0538_));
 sg13g2_nand2_1 _4410_ (.Y(_0540_),
    .A(_0537_),
    .B(_0539_));
 sg13g2_a21oi_1 _4411_ (.A1(_0535_),
    .A2(_0540_),
    .Y(_0541_),
    .B1(net147));
 sg13g2_nand2_1 _4412_ (.Y(_0542_),
    .A(_0402_),
    .B(net77));
 sg13g2_nand2_1 _4413_ (.Y(_0543_),
    .A(_0542_),
    .B(net36));
 sg13g2_a21oi_1 _4414_ (.A1(net34),
    .A2(net57),
    .Y(_0544_),
    .B1(net33));
 sg13g2_a21oi_1 _4415_ (.A1(_2999_),
    .A2(_0167_),
    .Y(_0545_),
    .B1(net162));
 sg13g2_o21ai_1 _4416_ (.B1(_0545_),
    .Y(_0546_),
    .A1(_0543_),
    .A2(_0544_));
 sg13g2_nand2_1 _4417_ (.Y(_0547_),
    .A(net153),
    .B(_2376_));
 sg13g2_inv_1 _4418_ (.Y(_0548_),
    .A(_0547_));
 sg13g2_o21ai_1 _4419_ (.B1(net110),
    .Y(_0549_),
    .A1(_0548_),
    .A2(_2801_));
 sg13g2_nand2_1 _4420_ (.Y(_0550_),
    .A(_0549_),
    .B(net169));
 sg13g2_a21oi_1 _4421_ (.A1(_0514_),
    .A2(_2789_),
    .Y(_0551_),
    .B1(net23));
 sg13g2_nor2_1 _4422_ (.A(_0550_),
    .B(_0551_),
    .Y(_0552_));
 sg13g2_nand2_1 _4423_ (.Y(_0553_),
    .A(_0546_),
    .B(_0552_));
 sg13g2_a21oi_1 _4424_ (.A1(_0541_),
    .A2(_0553_),
    .Y(_0554_),
    .B1(net200));
 sg13g2_nand2_1 _4425_ (.Y(_0555_),
    .A(_0526_),
    .B(_0554_));
 sg13g2_nand2_1 _4426_ (.Y(_0556_),
    .A(_0376_),
    .B(net144));
 sg13g2_nand3_1 _4427_ (.B(net92),
    .C(net150),
    .A(_0556_),
    .Y(_0557_));
 sg13g2_nand2_1 _4428_ (.Y(_0558_),
    .A(net59),
    .B(net106));
 sg13g2_a21oi_1 _4429_ (.A1(net52),
    .A2(net156),
    .Y(_0559_),
    .B1(_2641_));
 sg13g2_nor2_1 _4430_ (.A(_0558_),
    .B(_0559_),
    .Y(_0560_));
 sg13g2_nand2_1 _4431_ (.Y(_0561_),
    .A(_0557_),
    .B(_0560_));
 sg13g2_nand2_1 _4432_ (.Y(_0562_),
    .A(_0561_),
    .B(net36));
 sg13g2_nand2_2 _4433_ (.Y(_0563_),
    .A(_1795_),
    .B(net97));
 sg13g2_nand2_1 _4434_ (.Y(_0564_),
    .A(_0563_),
    .B(net136));
 sg13g2_nand2_1 _4435_ (.Y(_0565_),
    .A(net95),
    .B(net158));
 sg13g2_nand2_1 _4436_ (.Y(_0566_),
    .A(_0565_),
    .B(net58));
 sg13g2_nand2_1 _4437_ (.Y(_0567_),
    .A(_0564_),
    .B(_0566_));
 sg13g2_inv_1 _4438_ (.Y(_0568_),
    .A(_1948_));
 sg13g2_nor3_1 _4439_ (.A(_0568_),
    .B(net62),
    .C(_2678_),
    .Y(_0569_));
 sg13g2_a21oi_1 _4440_ (.A1(_0567_),
    .A2(net39),
    .Y(_0570_),
    .B1(_0569_));
 sg13g2_nand2_1 _4441_ (.Y(_0571_),
    .A(_0562_),
    .B(_0570_));
 sg13g2_nand2_1 _4442_ (.Y(_0572_),
    .A(_0571_),
    .B(net80));
 sg13g2_nand2_1 _4443_ (.Y(_0573_),
    .A(_2502_),
    .B(_2433_));
 sg13g2_nand2_1 _4444_ (.Y(_0574_),
    .A(_0573_),
    .B(_2842_));
 sg13g2_o21ai_1 _4445_ (.B1(net89),
    .Y(_0575_),
    .A1(_0112_),
    .A2(_1869_));
 sg13g2_nor2_1 _4446_ (.A(net137),
    .B(net41),
    .Y(_0576_));
 sg13g2_inv_1 _4447_ (.Y(_0577_),
    .A(_0576_));
 sg13g2_nand3_1 _4448_ (.B(_0575_),
    .C(_0577_),
    .A(_0574_),
    .Y(_0578_));
 sg13g2_nand2_1 _4449_ (.Y(_0579_),
    .A(_2435_),
    .B(net152));
 sg13g2_nor2_1 _4450_ (.A(_0112_),
    .B(_0579_),
    .Y(_0580_));
 sg13g2_nand2_1 _4451_ (.Y(_0581_),
    .A(_0395_),
    .B(_0226_));
 sg13g2_o21ai_1 _4452_ (.B1(net22),
    .Y(_0582_),
    .A1(_0580_),
    .A2(_0581_));
 sg13g2_nor2_1 _4453_ (.A(_2162_),
    .B(_0527_),
    .Y(_0583_));
 sg13g2_nand2_1 _4454_ (.Y(_0584_),
    .A(_2911_),
    .B(_0583_));
 sg13g2_nor2b_1 _4455_ (.A(_0582_),
    .B_N(_0584_),
    .Y(_0585_));
 sg13g2_a21oi_1 _4456_ (.A1(_0578_),
    .A2(net113),
    .Y(_0586_),
    .B1(_0585_));
 sg13g2_nand2_1 _4457_ (.Y(_0587_),
    .A(_0572_),
    .B(_0586_));
 sg13g2_nand2_1 _4458_ (.Y(_0588_),
    .A(_0587_),
    .B(net68));
 sg13g2_nand3_1 _4459_ (.B(net52),
    .C(_0422_),
    .A(net82),
    .Y(_0589_));
 sg13g2_o21ai_1 _4460_ (.B1(_0589_),
    .Y(_0590_),
    .A1(net99),
    .A2(_2977_));
 sg13g2_inv_1 _4461_ (.Y(_0591_),
    .A(_0303_));
 sg13g2_a21oi_1 _4462_ (.A1(_0590_),
    .A2(_0591_),
    .Y(_0592_),
    .B1(net163));
 sg13g2_nand2_1 _4463_ (.Y(_0593_),
    .A(_0588_),
    .B(_0592_));
 sg13g2_nand3_1 _4464_ (.B(_0593_),
    .C(net196),
    .A(_0555_),
    .Y(_0594_));
 sg13g2_nand2_1 _4465_ (.Y(_0024_),
    .A(_0494_),
    .B(_0594_));
 sg13g2_a21oi_1 _4466_ (.A1(_1773_),
    .A2(_0757_),
    .Y(_0595_),
    .B1(_1282_));
 sg13g2_inv_1 _4467_ (.Y(_0596_),
    .A(_0289_));
 sg13g2_nand2_2 _4468_ (.Y(_0597_),
    .A(_0595_),
    .B(_0596_));
 sg13g2_nor2_2 _4469_ (.A(_1653_),
    .B(net178),
    .Y(_0598_));
 sg13g2_inv_1 _4470_ (.Y(_0599_),
    .A(_0598_));
 sg13g2_nor2_2 _4471_ (.A(_2460_),
    .B(_2406_),
    .Y(_0600_));
 sg13g2_nand3_1 _4472_ (.B(_0599_),
    .C(_0600_),
    .A(_0597_),
    .Y(_0601_));
 sg13g2_inv_1 _4473_ (.Y(_0602_),
    .A(_2376_));
 sg13g2_nand2_1 _4474_ (.Y(_0603_),
    .A(_2848_),
    .B(net193));
 sg13g2_nor2_2 _4475_ (.A(net151),
    .B(_0118_),
    .Y(_0604_));
 sg13g2_a21oi_1 _4476_ (.A1(_0603_),
    .A2(_0604_),
    .Y(_0605_),
    .B1(_2423_));
 sg13g2_nand2_1 _4477_ (.Y(_0606_),
    .A(_0601_),
    .B(_0605_));
 sg13g2_nor2_2 _4478_ (.A(net206),
    .B(net125),
    .Y(_0607_));
 sg13g2_nand2_1 _4479_ (.Y(_0608_),
    .A(_0607_),
    .B(net193));
 sg13g2_nand2_2 _4480_ (.Y(_0609_),
    .A(_2633_),
    .B(net119));
 sg13g2_nor2_1 _4481_ (.A(net194),
    .B(_0609_),
    .Y(_0610_));
 sg13g2_nor2_1 _4482_ (.A(net108),
    .B(_0610_),
    .Y(_0611_));
 sg13g2_a21oi_1 _4483_ (.A1(net37),
    .A2(_0608_),
    .Y(_0612_),
    .B1(_0611_));
 sg13g2_nor2_1 _4484_ (.A(net66),
    .B(_0612_),
    .Y(_0613_));
 sg13g2_nor2_1 _4485_ (.A(_0606_),
    .B(_0613_),
    .Y(_0614_));
 sg13g2_nor2_1 _4486_ (.A(net138),
    .B(_2640_),
    .Y(_0615_));
 sg13g2_nand2_2 _4487_ (.Y(_0616_),
    .A(_2887_),
    .B(net201));
 sg13g2_nand2_2 _4488_ (.Y(_0617_),
    .A(_0616_),
    .B(net136));
 sg13g2_nand2_2 _4489_ (.Y(_0618_),
    .A(_2659_),
    .B(net51));
 sg13g2_a21oi_1 _4490_ (.A1(_0617_),
    .A2(_0618_),
    .Y(_0619_),
    .B1(net54));
 sg13g2_o21ai_1 _4491_ (.B1(net116),
    .Y(_0620_),
    .A1(_0615_),
    .A2(_0619_));
 sg13g2_nor2_1 _4492_ (.A(net184),
    .B(_0112_),
    .Y(_0621_));
 sg13g2_inv_2 _4493_ (.Y(_0622_),
    .A(_0621_));
 sg13g2_nand3_1 _4494_ (.B(net45),
    .C(_0143_),
    .A(_0622_),
    .Y(_0623_));
 sg13g2_nand2_1 _4495_ (.Y(_0624_),
    .A(_2953_),
    .B(_2686_));
 sg13g2_nand3_1 _4496_ (.B(net113),
    .C(_0624_),
    .A(_0623_),
    .Y(_0625_));
 sg13g2_nand3_1 _4497_ (.B(_0620_),
    .C(_0625_),
    .A(_0614_),
    .Y(_0626_));
 sg13g2_nand2_2 _4498_ (.Y(_0627_),
    .A(_1795_),
    .B(net93));
 sg13g2_nor2_2 _4499_ (.A(_1271_),
    .B(_0627_),
    .Y(_0628_));
 sg13g2_nand2_2 _4500_ (.Y(_0629_),
    .A(net139),
    .B(_2633_));
 sg13g2_a21oi_1 _4501_ (.A1(net108),
    .A2(_0128_),
    .Y(_0630_),
    .B1(net124));
 sg13g2_nand2_1 _4502_ (.Y(_0631_),
    .A(_2848_),
    .B(net194));
 sg13g2_a22oi_1 _4503_ (.Y(_0632_),
    .B1(_0630_),
    .B2(_0631_),
    .A2(_0629_),
    .A1(net134));
 sg13g2_o21ai_1 _4504_ (.B1(_0632_),
    .Y(_0633_),
    .A1(net31),
    .A2(_0628_));
 sg13g2_nand2_1 _4505_ (.Y(_0634_),
    .A(_0633_),
    .B(net121));
 sg13g2_a22oi_1 _4506_ (.Y(_0635_),
    .B1(_2701_),
    .B2(_0608_),
    .A2(net89),
    .A1(_0149_));
 sg13g2_nor2_1 _4507_ (.A(net35),
    .B(_0635_),
    .Y(_0636_));
 sg13g2_nand2_1 _4508_ (.Y(_0637_),
    .A(_2710_),
    .B(net194));
 sg13g2_a21oi_1 _4509_ (.A1(net76),
    .A2(_0128_),
    .Y(_0638_),
    .B1(_0337_));
 sg13g2_a21oi_1 _4510_ (.A1(_0637_),
    .A2(_0638_),
    .Y(_0639_),
    .B1(_2564_));
 sg13g2_nor2b_1 _4511_ (.A(_0636_),
    .B_N(_0639_),
    .Y(_0640_));
 sg13g2_nand2_1 _4512_ (.Y(_0641_),
    .A(_0634_),
    .B(_0640_));
 sg13g2_nand2_1 _4513_ (.Y(_0642_),
    .A(_0626_),
    .B(_0641_));
 sg13g2_nand2_1 _4514_ (.Y(_0643_),
    .A(_0642_),
    .B(net68));
 sg13g2_nor3_2 _4515_ (.A(net177),
    .B(_0142_),
    .C(_3013_),
    .Y(_0644_));
 sg13g2_a21o_1 _4516_ (.A2(_0618_),
    .A1(_0644_),
    .B1(net160),
    .X(_0645_));
 sg13g2_nor2_1 _4517_ (.A(net206),
    .B(net126),
    .Y(_0646_));
 sg13g2_o21ai_1 _4518_ (.B1(_0646_),
    .Y(_0647_),
    .A1(_0422_),
    .A2(_2482_));
 sg13g2_nand2_2 _4519_ (.Y(_0648_),
    .A(_0609_),
    .B(net93));
 sg13g2_nand2_1 _4520_ (.Y(_0649_),
    .A(_0617_),
    .B(_0648_));
 sg13g2_nand2_1 _4521_ (.Y(_0650_),
    .A(net180),
    .B(_0128_));
 sg13g2_buf_2 _4522_ (.A(_0650_),
    .X(_0651_));
 sg13g2_a21oi_1 _4523_ (.A1(net101),
    .A2(_0651_),
    .Y(_0652_),
    .B1(net169));
 sg13g2_a22oi_1 _4524_ (.Y(_0653_),
    .B1(_0649_),
    .B2(_0652_),
    .A2(net105),
    .A1(_0647_));
 sg13g2_nand2_1 _4525_ (.Y(_0654_),
    .A(_0603_),
    .B(net91));
 sg13g2_inv_1 _4526_ (.Y(_0655_),
    .A(_2998_));
 sg13g2_nand2_1 _4527_ (.Y(_0656_),
    .A(_0655_),
    .B(net149));
 sg13g2_nand2_1 _4528_ (.Y(_0657_),
    .A(_0654_),
    .B(_0656_));
 sg13g2_nand2_1 _4529_ (.Y(_0658_),
    .A(_0657_),
    .B(net22));
 sg13g2_nand3_1 _4530_ (.B(_0653_),
    .C(_0658_),
    .A(_0645_),
    .Y(_0659_));
 sg13g2_nand2_1 _4531_ (.Y(_0660_),
    .A(_0659_),
    .B(_2565_));
 sg13g2_nand2_1 _4532_ (.Y(_0661_),
    .A(_0339_),
    .B(net128));
 sg13g2_nand2_1 _4533_ (.Y(_0662_),
    .A(net174),
    .B(net194));
 sg13g2_nand2_1 _4534_ (.Y(_0663_),
    .A(_0661_),
    .B(_0662_));
 sg13g2_nand2_1 _4535_ (.Y(_0664_),
    .A(net71),
    .B(_2377_));
 sg13g2_o21ai_1 _4536_ (.B1(net161),
    .Y(_0665_),
    .A1(net64),
    .A2(_0664_));
 sg13g2_nor2_1 _4537_ (.A(_0663_),
    .B(_0665_),
    .Y(_0666_));
 sg13g2_nand2_1 _4538_ (.Y(_0667_),
    .A(_2862_),
    .B(net74));
 sg13g2_a21oi_1 _4539_ (.A1(_0666_),
    .A2(_0667_),
    .Y(_0668_),
    .B1(_2564_));
 sg13g2_nand2_2 _4540_ (.Y(_0669_),
    .A(_0609_),
    .B(_2401_));
 sg13g2_o21ai_1 _4541_ (.B1(_0669_),
    .Y(_0670_),
    .A1(_0438_),
    .A2(_0618_));
 sg13g2_nand2_1 _4542_ (.Y(_0671_),
    .A(_0670_),
    .B(net32));
 sg13g2_nor3_1 _4543_ (.A(net101),
    .B(_2378_),
    .C(_0607_),
    .Y(_0672_));
 sg13g2_nand2_2 _4544_ (.Y(_0673_),
    .A(_0629_),
    .B(net179));
 sg13g2_nor2_1 _4545_ (.A(net171),
    .B(_0673_),
    .Y(_0674_));
 sg13g2_nor2_1 _4546_ (.A(_0672_),
    .B(_0674_),
    .Y(_0675_));
 sg13g2_a21oi_1 _4547_ (.A1(_0608_),
    .A2(net42),
    .Y(_0676_),
    .B1(net127));
 sg13g2_nand3_1 _4548_ (.B(_0675_),
    .C(_0676_),
    .A(_0671_),
    .Y(_0677_));
 sg13g2_nand2_1 _4549_ (.Y(_0678_),
    .A(_0668_),
    .B(_0677_));
 sg13g2_nand3_1 _4550_ (.B(_0678_),
    .C(net164),
    .A(_0660_),
    .Y(_0679_));
 sg13g2_a21oi_1 _4551_ (.A1(_0643_),
    .A2(_0679_),
    .Y(_0680_),
    .B1(net196));
 sg13g2_nor2_1 _4552_ (.A(net133),
    .B(_0547_),
    .Y(_0681_));
 sg13g2_nand2_1 _4553_ (.Y(_0682_),
    .A(_0565_),
    .B(_2097_));
 sg13g2_nand2_1 _4554_ (.Y(_0683_),
    .A(_0682_),
    .B(_2844_));
 sg13g2_a22oi_1 _4555_ (.Y(_0684_),
    .B1(_0644_),
    .B2(_0683_),
    .A2(_0681_),
    .A1(net84));
 sg13g2_nand2_1 _4556_ (.Y(_0685_),
    .A(_0597_),
    .B(_3022_));
 sg13g2_nand2_1 _4557_ (.Y(_0686_),
    .A(_2768_),
    .B(net114));
 sg13g2_a21oi_1 _4558_ (.A1(_0685_),
    .A2(_0686_),
    .Y(_0687_),
    .B1(net160));
 sg13g2_a21oi_1 _4559_ (.A1(_0684_),
    .A2(net22),
    .Y(_0688_),
    .B1(_0687_));
 sg13g2_nor2_1 _4560_ (.A(net64),
    .B(_2723_),
    .Y(_0689_));
 sg13g2_nand3_1 _4561_ (.B(_2444_),
    .C(_2405_),
    .A(_2591_),
    .Y(_0690_));
 sg13g2_nor2b_1 _4562_ (.A(_0689_),
    .B_N(_0690_),
    .Y(_0691_));
 sg13g2_o21ai_1 _4563_ (.B1(_2861_),
    .Y(_0692_),
    .A1(net92),
    .A2(_0607_));
 sg13g2_nand2_1 _4564_ (.Y(_0693_),
    .A(_0692_),
    .B(net39));
 sg13g2_o21ai_1 _4565_ (.B1(net49),
    .Y(_0694_),
    .A1(net194),
    .A2(_0350_));
 sg13g2_nand3_1 _4566_ (.B(_0693_),
    .C(_0694_),
    .A(_0691_),
    .Y(_0695_));
 sg13g2_nand2_1 _4567_ (.Y(_0696_),
    .A(_0695_),
    .B(net116));
 sg13g2_nand2_1 _4568_ (.Y(_0697_),
    .A(_0688_),
    .B(_0696_));
 sg13g2_nand2_1 _4569_ (.Y(_0698_),
    .A(_0697_),
    .B(net68));
 sg13g2_nor2_1 _4570_ (.A(net61),
    .B(_2892_),
    .Y(_0699_));
 sg13g2_nand2_1 _4571_ (.Y(_0700_),
    .A(net100),
    .B(net193));
 sg13g2_nand3_1 _4572_ (.B(net55),
    .C(_2532_),
    .A(_2444_),
    .Y(_0701_));
 sg13g2_a221oi_1 _4573_ (.B2(_0701_),
    .C1(net118),
    .B1(_0454_),
    .A1(_0699_),
    .Y(_0702_),
    .A2(_0700_));
 sg13g2_nand2_1 _4574_ (.Y(_0703_),
    .A(_2273_),
    .B(net119));
 sg13g2_nand2_1 _4575_ (.Y(_0704_),
    .A(_0703_),
    .B(net92));
 sg13g2_a21oi_1 _4576_ (.A1(_0704_),
    .A2(_0618_),
    .Y(_0705_),
    .B1(net54));
 sg13g2_nand2_1 _4577_ (.Y(_0706_),
    .A(_0599_),
    .B(net128));
 sg13g2_nor3_1 _4578_ (.A(net107),
    .B(_0477_),
    .C(_0706_),
    .Y(_0707_));
 sg13g2_nor2_1 _4579_ (.A(net62),
    .B(_2638_),
    .Y(_0708_));
 sg13g2_nor2_1 _4580_ (.A(_0530_),
    .B(_0607_),
    .Y(_0709_));
 sg13g2_o21ai_1 _4581_ (.B1(net134),
    .Y(_0710_),
    .A1(_2892_),
    .A2(_0709_));
 sg13g2_nand2b_1 _4582_ (.Y(_0711_),
    .B(_0710_),
    .A_N(_0708_));
 sg13g2_nor3_1 _4583_ (.A(_0705_),
    .B(_0707_),
    .C(_0711_),
    .Y(_0712_));
 sg13g2_nor2_1 _4584_ (.A(net63),
    .B(_0712_),
    .Y(_0713_));
 sg13g2_nor2_1 _4585_ (.A(_0702_),
    .B(_0713_),
    .Y(_0714_));
 sg13g2_nand2_1 _4586_ (.Y(_0715_),
    .A(_0698_),
    .B(_0714_));
 sg13g2_nor2_2 _4587_ (.A(net179),
    .B(_2998_),
    .Y(_0716_));
 sg13g2_a22oi_1 _4588_ (.Y(_0717_),
    .B1(_0716_),
    .B2(_0514_),
    .A2(_2637_),
    .A1(net42));
 sg13g2_nand3b_1 _4589_ (.B(_0717_),
    .C(net80),
    .Y(_0718_),
    .A_N(_0674_));
 sg13g2_nand2_1 _4590_ (.Y(_0719_),
    .A(_0692_),
    .B(net24));
 sg13g2_nor2_1 _4591_ (.A(net146),
    .B(_1151_),
    .Y(_0720_));
 sg13g2_nor2_2 _4592_ (.A(net151),
    .B(_0720_),
    .Y(_0721_));
 sg13g2_nand2_1 _4593_ (.Y(_0722_),
    .A(_2719_),
    .B(_0721_));
 sg13g2_nand3_1 _4594_ (.B(_0722_),
    .C(net22),
    .A(_0719_),
    .Y(_0723_));
 sg13g2_nand2_1 _4595_ (.Y(_0724_),
    .A(_0664_),
    .B(net32));
 sg13g2_o21ai_1 _4596_ (.B1(_0724_),
    .Y(_0726_),
    .A1(_2793_),
    .A2(_0533_));
 sg13g2_nor2_1 _4597_ (.A(net197),
    .B(_2564_),
    .Y(_0727_));
 sg13g2_buf_2 _4598_ (.A(_0727_),
    .X(_0728_));
 sg13g2_inv_1 _4599_ (.Y(_0729_),
    .A(net112));
 sg13g2_a21oi_1 _4600_ (.A1(_0726_),
    .A2(net131),
    .Y(_0730_),
    .B1(_0729_));
 sg13g2_nand3_1 _4601_ (.B(_0723_),
    .C(_0730_),
    .A(_0718_),
    .Y(_0731_));
 sg13g2_nand2_1 _4602_ (.Y(_0732_),
    .A(net115),
    .B(_0127_));
 sg13g2_o21ai_1 _4603_ (.B1(_2598_),
    .Y(_0733_),
    .A1(_0732_),
    .A2(_0631_));
 sg13g2_nand3_1 _4604_ (.B(net196),
    .C(_0733_),
    .A(_0731_),
    .Y(_0734_));
 sg13g2_a21oi_1 _4605_ (.A1(_0715_),
    .A2(net132),
    .Y(_0735_),
    .B1(_0734_));
 sg13g2_nor2_1 _4606_ (.A(_0680_),
    .B(_0735_),
    .Y(_0025_));
 sg13g2_nor2_1 _4607_ (.A(_1631_),
    .B(_0580_),
    .Y(_0737_));
 sg13g2_o21ai_1 _4608_ (.B1(_0737_),
    .Y(_0738_),
    .A1(_2392_),
    .A2(_2656_));
 sg13g2_nor3_1 _4609_ (.A(net179),
    .B(net103),
    .C(_3013_),
    .Y(_0739_));
 sg13g2_a21oi_1 _4610_ (.A1(_0739_),
    .A2(_3046_),
    .Y(_0740_),
    .B1(net173));
 sg13g2_nand2_1 _4611_ (.Y(_0741_),
    .A(_0738_),
    .B(_0740_));
 sg13g2_nand2_1 _4612_ (.Y(_0742_),
    .A(_0596_),
    .B(net144));
 sg13g2_nand2_1 _4613_ (.Y(_0743_),
    .A(_0742_),
    .B(_2401_));
 sg13g2_inv_1 _4614_ (.Y(_0744_),
    .A(_0477_));
 sg13g2_nand2_1 _4615_ (.Y(_0745_),
    .A(_0743_),
    .B(_0744_));
 sg13g2_nand3_1 _4616_ (.B(net142),
    .C(net161),
    .A(_0745_),
    .Y(_0747_));
 sg13g2_nor2_2 _4617_ (.A(net174),
    .B(net209),
    .Y(_0748_));
 sg13g2_nand3_1 _4618_ (.B(_2719_),
    .C(_0748_),
    .A(_2712_),
    .Y(_0749_));
 sg13g2_nand3_1 _4619_ (.B(_0747_),
    .C(_0749_),
    .A(_0741_),
    .Y(_0750_));
 sg13g2_nand2_1 _4620_ (.Y(_0751_),
    .A(_0750_),
    .B(net46));
 sg13g2_a21oi_1 _4621_ (.A1(_2489_),
    .A2(_2402_),
    .Y(_0752_),
    .B1(net142));
 sg13g2_nand2_1 _4622_ (.Y(_0753_),
    .A(_2616_),
    .B(_2682_));
 sg13g2_o21ai_1 _4623_ (.B1(net113),
    .Y(_0754_),
    .A1(net89),
    .A2(net29));
 sg13g2_a21oi_1 _4624_ (.A1(_0752_),
    .A2(_0753_),
    .Y(_0755_),
    .B1(_0754_));
 sg13g2_nand2_1 _4625_ (.Y(_0756_),
    .A(_0468_),
    .B(_0669_));
 sg13g2_nor2_1 _4626_ (.A(_1107_),
    .B(_2678_),
    .Y(_0758_));
 sg13g2_a22oi_1 _4627_ (.Y(_0759_),
    .B1(_0758_),
    .B2(_3025_),
    .A2(net110),
    .A1(_0756_));
 sg13g2_nor2_1 _4628_ (.A(net167),
    .B(_0759_),
    .Y(_0760_));
 sg13g2_nor3_1 _4629_ (.A(_2557_),
    .B(_0755_),
    .C(_0760_),
    .Y(_0761_));
 sg13g2_nand2_1 _4630_ (.Y(_0762_),
    .A(_0751_),
    .B(_0761_));
 sg13g2_a21oi_1 _4631_ (.A1(_0096_),
    .A2(_2526_),
    .Y(_0763_),
    .B1(net31));
 sg13g2_nor2_1 _4632_ (.A(_2844_),
    .B(_2031_),
    .Y(_0764_));
 sg13g2_nor3_1 _4633_ (.A(net40),
    .B(_2616_),
    .C(_0764_),
    .Y(_0765_));
 sg13g2_nor3_1 _4634_ (.A(_2816_),
    .B(_0763_),
    .C(_0765_),
    .Y(_0766_));
 sg13g2_nand3_1 _4635_ (.B(net55),
    .C(_2901_),
    .A(_0683_),
    .Y(_0767_));
 sg13g2_a21oi_1 _4636_ (.A1(_2728_),
    .A2(_0943_),
    .Y(_0769_),
    .B1(_2729_));
 sg13g2_a21oi_1 _4637_ (.A1(_0627_),
    .A2(_0769_),
    .Y(_0770_),
    .B1(net81));
 sg13g2_nand2_1 _4638_ (.Y(_0771_),
    .A(_0767_),
    .B(_0770_));
 sg13g2_nand3_1 _4639_ (.B(net72),
    .C(_2853_),
    .A(_0125_),
    .Y(_0772_));
 sg13g2_a21oi_1 _4640_ (.A1(_0669_),
    .A2(_0583_),
    .Y(_0773_),
    .B1(_2733_));
 sg13g2_nand2_1 _4641_ (.Y(_0774_),
    .A(_0772_),
    .B(_0773_));
 sg13g2_o21ai_1 _4642_ (.B1(_2779_),
    .Y(_0775_),
    .A1(net33),
    .A2(_2888_));
 sg13g2_o21ai_1 _4643_ (.B1(_2373_),
    .Y(_0776_),
    .A1(net172),
    .A2(_2855_));
 sg13g2_a21oi_1 _4644_ (.A1(net26),
    .A2(_0775_),
    .Y(_0777_),
    .B1(_0776_));
 sg13g2_a22oi_1 _4645_ (.Y(_0778_),
    .B1(_0774_),
    .B2(_0777_),
    .A2(_0771_),
    .A1(_0766_));
 sg13g2_nand2_1 _4646_ (.Y(_0780_),
    .A(_0762_),
    .B(_0778_));
 sg13g2_nand2_1 _4647_ (.Y(_0781_),
    .A(_0780_),
    .B(net132));
 sg13g2_nand3_1 _4648_ (.B(_2433_),
    .C(_1522_),
    .A(net95),
    .Y(_0782_));
 sg13g2_a21oi_1 _4649_ (.A1(_0644_),
    .A2(_0782_),
    .Y(_0783_),
    .B1(_0118_));
 sg13g2_inv_1 _4650_ (.Y(_0784_),
    .A(net59));
 sg13g2_nand2_1 _4651_ (.Y(_0785_),
    .A(_0784_),
    .B(net94));
 sg13g2_nand3_1 _4652_ (.B(net120),
    .C(_0785_),
    .A(_0487_),
    .Y(_0786_));
 sg13g2_nor4_1 _4653_ (.A(net36),
    .B(_0337_),
    .C(_2453_),
    .D(_2520_),
    .Y(_0787_));
 sg13g2_a21oi_1 _4654_ (.A1(_0783_),
    .A2(_0786_),
    .Y(_0788_),
    .B1(_0787_));
 sg13g2_nand3_1 _4655_ (.B(_0514_),
    .C(net110),
    .A(_3017_),
    .Y(_0789_));
 sg13g2_inv_1 _4656_ (.Y(_0791_),
    .A(_1653_));
 sg13g2_o21ai_1 _4657_ (.B1(net69),
    .Y(_0792_),
    .A1(_0791_),
    .A2(_2806_));
 sg13g2_nand2_1 _4658_ (.Y(_0793_),
    .A(_0789_),
    .B(_0792_));
 sg13g2_nand2_1 _4659_ (.Y(_0794_),
    .A(_0793_),
    .B(net121));
 sg13g2_nand2_1 _4660_ (.Y(_0795_),
    .A(_1948_),
    .B(net182));
 sg13g2_nor2_1 _4661_ (.A(_0795_),
    .B(_2916_),
    .Y(_0796_));
 sg13g2_inv_1 _4662_ (.Y(_0797_),
    .A(_2532_));
 sg13g2_nor3_1 _4663_ (.A(net75),
    .B(_0797_),
    .C(_0673_),
    .Y(_0798_));
 sg13g2_o21ai_1 _4664_ (.B1(net116),
    .Y(_0799_),
    .A1(_0796_),
    .A2(_0798_));
 sg13g2_nand3_1 _4665_ (.B(_0794_),
    .C(_0799_),
    .A(_0788_),
    .Y(_0800_));
 sg13g2_nand2_1 _4666_ (.Y(_0802_),
    .A(_0800_),
    .B(net73));
 sg13g2_nor2_1 _4667_ (.A(_2467_),
    .B(_2880_),
    .Y(_0803_));
 sg13g2_nand2_1 _4668_ (.Y(_0804_),
    .A(_0803_),
    .B(_1921_));
 sg13g2_a21oi_1 _4669_ (.A1(_0804_),
    .A2(_0129_),
    .Y(_0805_),
    .B1(net170));
 sg13g2_a21oi_1 _4670_ (.A1(_0802_),
    .A2(_0805_),
    .Y(_0806_),
    .B1(_2696_));
 sg13g2_nand2_1 _4671_ (.Y(_0807_),
    .A(_0781_),
    .B(_0806_));
 sg13g2_nand2_2 _4672_ (.Y(_0808_),
    .A(_2020_),
    .B(net109));
 sg13g2_nand2_1 _4673_ (.Y(_0809_),
    .A(_0743_),
    .B(_0808_));
 sg13g2_nand3_1 _4674_ (.B(net161),
    .C(net88),
    .A(_0809_),
    .Y(_0810_));
 sg13g2_nor2_1 _4675_ (.A(_0163_),
    .B(_0673_),
    .Y(_0811_));
 sg13g2_nand2_1 _4676_ (.Y(_0813_),
    .A(_0409_),
    .B(_0811_));
 sg13g2_nand2_1 _4677_ (.Y(_0814_),
    .A(_0810_),
    .B(_0813_));
 sg13g2_a21oi_1 _4678_ (.A1(_2945_),
    .A2(_1653_),
    .Y(_0815_),
    .B1(_0337_));
 sg13g2_nor2_1 _4679_ (.A(net151),
    .B(_0797_),
    .Y(_0816_));
 sg13g2_nand2_1 _4680_ (.Y(_0817_),
    .A(_3025_),
    .B(_0816_));
 sg13g2_nand2_1 _4681_ (.Y(_0818_),
    .A(_0815_),
    .B(_0817_));
 sg13g2_nor2b_1 _4682_ (.A(_0814_),
    .B_N(_0818_),
    .Y(_0819_));
 sg13g2_nand2b_1 _4683_ (.Y(_0820_),
    .B(_0816_),
    .A_N(_3028_));
 sg13g2_nand2_1 _4684_ (.Y(_0821_),
    .A(_2606_),
    .B(_0820_));
 sg13g2_nand2_1 _4685_ (.Y(_0822_),
    .A(_0821_),
    .B(_1707_));
 sg13g2_nor2_1 _4686_ (.A(_1096_),
    .B(_0598_),
    .Y(_0824_));
 sg13g2_nand2_2 _4687_ (.Y(_0825_),
    .A(_1795_),
    .B(net154));
 sg13g2_nand2_1 _4688_ (.Y(_0826_),
    .A(_0825_),
    .B(_2444_));
 sg13g2_a22oi_1 _4689_ (.Y(_0827_),
    .B1(net39),
    .B2(_0826_),
    .A2(_0824_),
    .A1(_0471_));
 sg13g2_nand2_1 _4690_ (.Y(_0828_),
    .A(_0822_),
    .B(_0827_));
 sg13g2_nand2_1 _4691_ (.Y(_0829_),
    .A(_0828_),
    .B(net131));
 sg13g2_nand2_1 _4692_ (.Y(_0830_),
    .A(_0819_),
    .B(_0829_));
 sg13g2_nand2_1 _4693_ (.Y(_0831_),
    .A(_0830_),
    .B(_0090_));
 sg13g2_nand2_1 _4694_ (.Y(_0832_),
    .A(_0563_),
    .B(net51));
 sg13g2_nand2_1 _4695_ (.Y(_0833_),
    .A(net103),
    .B(_2633_));
 sg13g2_and3_1 _4696_ (.X(_0835_),
    .A(_0832_),
    .B(net72),
    .C(_0833_));
 sg13g2_o21ai_1 _4697_ (.B1(_2601_),
    .Y(_0836_),
    .A1(_0346_),
    .A2(_0518_));
 sg13g2_o21ai_1 _4698_ (.B1(net169),
    .Y(_0837_),
    .A1(net168),
    .A2(_0589_));
 sg13g2_nand2_2 _4699_ (.Y(_0838_),
    .A(_2967_),
    .B(net92));
 sg13g2_nand2_1 _4700_ (.Y(_0839_),
    .A(_2414_),
    .B(net27));
 sg13g2_a21oi_1 _4701_ (.A1(_0838_),
    .A2(_0839_),
    .Y(_0840_),
    .B1(net61));
 sg13g2_nor2_1 _4702_ (.A(_0837_),
    .B(_0840_),
    .Y(_0841_));
 sg13g2_o21ai_1 _4703_ (.B1(_0841_),
    .Y(_0842_),
    .A1(_0835_),
    .A2(_0836_));
 sg13g2_a21o_1 _4704_ (.A2(_0785_),
    .A1(_2656_),
    .B1(net61),
    .X(_0843_));
 sg13g2_a22oi_1 _4705_ (.Y(_0844_),
    .B1(_1848_),
    .B2(_0142_),
    .A2(_1457_),
    .A1(_2387_));
 sg13g2_nor2_1 _4706_ (.A(_2445_),
    .B(_2453_),
    .Y(_0846_));
 sg13g2_nand2_1 _4707_ (.Y(_0847_),
    .A(_2854_),
    .B(net158));
 sg13g2_nand2_1 _4708_ (.Y(_0848_),
    .A(_2392_),
    .B(net58));
 sg13g2_nand3_1 _4709_ (.B(_0848_),
    .C(net69),
    .A(_0847_),
    .Y(_0849_));
 sg13g2_nand2_1 _4710_ (.Y(_0850_),
    .A(_0849_),
    .B(_2698_));
 sg13g2_a21oi_1 _4711_ (.A1(_0844_),
    .A2(_0846_),
    .Y(_0851_),
    .B1(_0850_));
 sg13g2_nand2_1 _4712_ (.Y(_0852_),
    .A(_0742_),
    .B(_2416_));
 sg13g2_nand2_1 _4713_ (.Y(_0853_),
    .A(_0852_),
    .B(_2861_));
 sg13g2_nand2_1 _4714_ (.Y(_0854_),
    .A(_0853_),
    .B(net26));
 sg13g2_nand3_1 _4715_ (.B(_0851_),
    .C(_0854_),
    .A(_0843_),
    .Y(_0855_));
 sg13g2_nand3_1 _4716_ (.B(_0855_),
    .C(net164),
    .A(_0842_),
    .Y(_0857_));
 sg13g2_nand3_1 _4717_ (.B(_0857_),
    .C(_2738_),
    .A(_0831_),
    .Y(_0858_));
 sg13g2_inv_1 _4718_ (.Y(_0859_),
    .A(_0470_));
 sg13g2_o21ai_1 _4719_ (.B1(net99),
    .Y(_0860_),
    .A1(_0568_),
    .A2(_0859_));
 sg13g2_nand3_1 _4720_ (.B(net24),
    .C(_2920_),
    .A(_0514_),
    .Y(_0861_));
 sg13g2_a21oi_1 _4721_ (.A1(_0860_),
    .A2(_0861_),
    .Y(_0862_),
    .B1(net66));
 sg13g2_inv_1 _4722_ (.Y(_0863_),
    .A(_0716_));
 sg13g2_o21ai_1 _4723_ (.B1(net114),
    .Y(_0864_),
    .A1(_0548_),
    .A2(_2801_));
 sg13g2_o21ai_1 _4724_ (.B1(_0864_),
    .Y(_0865_),
    .A1(_2279_),
    .A2(_0863_));
 sg13g2_nor2_2 _4725_ (.A(net202),
    .B(_0482_),
    .Y(_0866_));
 sg13g2_inv_1 _4726_ (.Y(_0868_),
    .A(_0866_));
 sg13g2_nor2b_1 _4727_ (.A(_0510_),
    .B_N(_2861_),
    .Y(_0869_));
 sg13g2_o21ai_1 _4728_ (.B1(_2598_),
    .Y(_0870_),
    .A1(_0868_),
    .A2(_0869_));
 sg13g2_a21oi_1 _4729_ (.A1(_0865_),
    .A2(net22),
    .Y(_0871_),
    .B1(_0870_));
 sg13g2_nand2_1 _4730_ (.Y(_0872_),
    .A(_0259_),
    .B(_0704_));
 sg13g2_a21oi_1 _4731_ (.A1(_0487_),
    .A2(_2536_),
    .Y(_0873_),
    .B1(net35));
 sg13g2_nand2_1 _4732_ (.Y(_0874_),
    .A(_0872_),
    .B(_0873_));
 sg13g2_a21o_1 _4733_ (.A2(_2496_),
    .A1(_0832_),
    .B1(net37),
    .X(_0875_));
 sg13g2_nand2b_1 _4734_ (.Y(_0876_),
    .B(net113),
    .A_N(_0875_));
 sg13g2_nand3_1 _4735_ (.B(_0874_),
    .C(_0876_),
    .A(_0871_),
    .Y(_0877_));
 sg13g2_nor2_1 _4736_ (.A(_0862_),
    .B(_0877_),
    .Y(_0879_));
 sg13g2_nand3_1 _4737_ (.B(_0669_),
    .C(net39),
    .A(_2967_),
    .Y(_0880_));
 sg13g2_o21ai_1 _4738_ (.B1(net88),
    .Y(_0881_),
    .A1(_0438_),
    .A2(_2775_));
 sg13g2_a21oi_1 _4739_ (.A1(_0880_),
    .A2(_0881_),
    .Y(_0882_),
    .B1(net127));
 sg13g2_nand2_1 _4740_ (.Y(_0883_),
    .A(_2970_),
    .B(net149));
 sg13g2_nor2_1 _4741_ (.A(net174),
    .B(_0548_),
    .Y(_0884_));
 sg13g2_a21oi_1 _4742_ (.A1(_2622_),
    .A2(_0884_),
    .Y(_0885_),
    .B1(_0118_));
 sg13g2_o21ai_1 _4743_ (.B1(_0885_),
    .Y(_0886_),
    .A1(_0134_),
    .A2(_0883_));
 sg13g2_nand2_1 _4744_ (.Y(_0887_),
    .A(_0886_),
    .B(_0728_));
 sg13g2_nor2_1 _4745_ (.A(_0882_),
    .B(_0887_),
    .Y(_0888_));
 sg13g2_a21oi_1 _4746_ (.A1(_2978_),
    .A2(_2482_),
    .Y(_0890_),
    .B1(net107));
 sg13g2_nand2_1 _4747_ (.Y(_0891_),
    .A(_0875_),
    .B(_0890_));
 sg13g2_nand2_1 _4748_ (.Y(_0892_),
    .A(net124),
    .B(net193));
 sg13g2_a21oi_1 _4749_ (.A1(_2677_),
    .A2(net142),
    .Y(_0893_),
    .B1(_0892_));
 sg13g2_nand2_1 _4750_ (.Y(_0894_),
    .A(_0563_),
    .B(net36));
 sg13g2_a21oi_1 _4751_ (.A1(_0893_),
    .A2(_0894_),
    .Y(_0895_),
    .B1(net167));
 sg13g2_nand2_1 _4752_ (.Y(_0896_),
    .A(_0891_),
    .B(_0895_));
 sg13g2_a21oi_1 _4753_ (.A1(_0888_),
    .A2(_0896_),
    .Y(_0897_),
    .B1(_2609_));
 sg13g2_nor2b_1 _4754_ (.A(_0879_),
    .B_N(_0897_),
    .Y(_0898_));
 sg13g2_nand2_1 _4755_ (.Y(_0899_),
    .A(_0858_),
    .B(_0898_));
 sg13g2_nand2_1 _4756_ (.Y(_0026_),
    .A(_0807_),
    .B(_0899_));
 sg13g2_nand2_1 _4757_ (.Y(_0901_),
    .A(_0573_),
    .B(net58));
 sg13g2_nand2_1 _4758_ (.Y(_0902_),
    .A(_0901_),
    .B(_0470_));
 sg13g2_nand2_1 _4759_ (.Y(_0903_),
    .A(_0902_),
    .B(net42));
 sg13g2_a21oi_1 _4760_ (.A1(_3036_),
    .A2(_1948_),
    .Y(_0904_),
    .B1(net101));
 sg13g2_nor2_1 _4761_ (.A(_1685_),
    .B(_2378_),
    .Y(_0905_));
 sg13g2_nand3_1 _4762_ (.B(net135),
    .C(_0905_),
    .A(_0563_),
    .Y(_0906_));
 sg13g2_nand2_1 _4763_ (.Y(_0907_),
    .A(_2603_),
    .B(net146));
 sg13g2_nand2_1 _4764_ (.Y(_0908_),
    .A(_0907_),
    .B(net104));
 sg13g2_nand2_1 _4765_ (.Y(_0909_),
    .A(_0906_),
    .B(_0908_));
 sg13g2_nor2_1 _4766_ (.A(_0904_),
    .B(_0909_),
    .Y(_0911_));
 sg13g2_nand2_1 _4767_ (.Y(_0912_),
    .A(_0903_),
    .B(_0911_));
 sg13g2_nand2_1 _4768_ (.Y(_0913_),
    .A(_0912_),
    .B(net121));
 sg13g2_o21ai_1 _4769_ (.B1(_0564_),
    .Y(_0914_),
    .A1(net155),
    .A2(_0622_));
 sg13g2_nor2_2 _4770_ (.A(_0127_),
    .B(net180),
    .Y(_0915_));
 sg13g2_nand2_1 _4771_ (.Y(_0916_),
    .A(_0915_),
    .B(_2460_));
 sg13g2_inv_1 _4772_ (.Y(_0917_),
    .A(_0916_));
 sg13g2_nor2_1 _4773_ (.A(net140),
    .B(_2947_),
    .Y(_0918_));
 sg13g2_nor2_1 _4774_ (.A(_3047_),
    .B(_0918_),
    .Y(_0919_));
 sg13g2_a21oi_1 _4775_ (.A1(_0919_),
    .A2(net84),
    .Y(_0920_),
    .B1(_0716_));
 sg13g2_a22oi_1 _4776_ (.Y(_0922_),
    .B1(net115),
    .B2(_0920_),
    .A2(_0917_),
    .A1(_0914_));
 sg13g2_nand2_1 _4777_ (.Y(_0923_),
    .A(_0913_),
    .B(_0922_));
 sg13g2_nand2_1 _4778_ (.Y(_0924_),
    .A(_0923_),
    .B(net73));
 sg13g2_nor2_1 _4779_ (.A(net107),
    .B(_0673_),
    .Y(_0925_));
 sg13g2_inv_1 _4780_ (.Y(_0926_),
    .A(_0648_));
 sg13g2_nor2_1 _4781_ (.A(_0598_),
    .B(_0926_),
    .Y(_0927_));
 sg13g2_a22oi_1 _4782_ (.Y(_0928_),
    .B1(net50),
    .B2(_0927_),
    .A2(_0825_),
    .A1(_0925_));
 sg13g2_o21ai_1 _4783_ (.B1(net32),
    .Y(_0929_),
    .A1(net85),
    .A2(_2429_));
 sg13g2_a21oi_1 _4784_ (.A1(_0928_),
    .A2(_0929_),
    .Y(_0930_),
    .B1(net118));
 sg13g2_nand2_1 _4785_ (.Y(_0931_),
    .A(_0803_),
    .B(_0250_));
 sg13g2_nand2_1 _4786_ (.Y(_0933_),
    .A(_0931_),
    .B(net53));
 sg13g2_nor2_1 _4787_ (.A(_2537_),
    .B(_1805_),
    .Y(_0934_));
 sg13g2_nand2_1 _4788_ (.Y(_0935_),
    .A(_0934_),
    .B(_2810_));
 sg13g2_a21oi_1 _4789_ (.A1(_0935_),
    .A2(net74),
    .Y(_0936_),
    .B1(_2462_));
 sg13g2_a21oi_1 _4790_ (.A1(_0933_),
    .A2(_0936_),
    .Y(_0937_),
    .B1(net63));
 sg13g2_nor2_1 _4791_ (.A(_0930_),
    .B(_0937_),
    .Y(_0938_));
 sg13g2_nand2_1 _4792_ (.Y(_0939_),
    .A(_0924_),
    .B(_0938_));
 sg13g2_nor2_1 _4793_ (.A(net128),
    .B(_0372_),
    .Y(_0940_));
 sg13g2_o21ai_1 _4794_ (.B1(_0940_),
    .Y(_0941_),
    .A1(_0326_),
    .A2(_2031_));
 sg13g2_nand2_1 _4795_ (.Y(_0942_),
    .A(net193),
    .B(net198));
 sg13g2_o21ai_1 _4796_ (.B1(net54),
    .Y(_0944_),
    .A1(_0942_),
    .A2(_0607_));
 sg13g2_a21oi_1 _4797_ (.A1(_0351_),
    .A2(_2856_),
    .Y(_0945_),
    .B1(_2963_));
 sg13g2_a21oi_1 _4798_ (.A1(_0941_),
    .A2(_0944_),
    .Y(_0946_),
    .B1(_0945_));
 sg13g2_nor3_1 _4799_ (.A(net180),
    .B(net193),
    .C(_0128_),
    .Y(_0947_));
 sg13g2_inv_1 _4800_ (.Y(_0948_),
    .A(_0947_));
 sg13g2_nor2_1 _4801_ (.A(net203),
    .B(_0948_),
    .Y(_0949_));
 sg13g2_nand4_1 _4802_ (.B(_1948_),
    .C(_2605_),
    .A(_2430_),
    .Y(_0950_),
    .D(net120));
 sg13g2_nand2_1 _4803_ (.Y(_0951_),
    .A(_2854_),
    .B(net96));
 sg13g2_nand2_1 _4804_ (.Y(_0952_),
    .A(_0951_),
    .B(_2795_));
 sg13g2_a21oi_1 _4805_ (.A1(_0739_),
    .A2(_0952_),
    .Y(_0953_),
    .B1(net66));
 sg13g2_a22oi_1 _4806_ (.Y(_0955_),
    .B1(_0950_),
    .B2(_0953_),
    .A2(_0949_),
    .A1(_0339_));
 sg13g2_o21ai_1 _4807_ (.B1(_0955_),
    .Y(_0956_),
    .A1(net83),
    .A2(_0946_));
 sg13g2_nand2_1 _4808_ (.Y(_0957_),
    .A(_0956_),
    .B(net112));
 sg13g2_a21oi_2 _4809_ (.B1(net174),
    .Y(_0958_),
    .A2(net86),
    .A1(net44));
 sg13g2_nor2_1 _4810_ (.A(_2564_),
    .B(_0303_),
    .Y(_0959_));
 sg13g2_inv_1 _4811_ (.Y(_0960_),
    .A(_0959_));
 sg13g2_a221oi_1 _4812_ (.B2(_2959_),
    .C1(_0960_),
    .B1(_0958_),
    .A1(_2740_),
    .Y(_0961_),
    .A2(_0321_));
 sg13g2_nor2_1 _4813_ (.A(net195),
    .B(_0961_),
    .Y(_0962_));
 sg13g2_nand2_1 _4814_ (.Y(_0963_),
    .A(_0957_),
    .B(_0962_));
 sg13g2_a21oi_1 _4815_ (.A1(_0939_),
    .A2(_2566_),
    .Y(_0964_),
    .B1(_0963_));
 sg13g2_a21oi_1 _4816_ (.A1(_1968_),
    .A2(_2807_),
    .Y(_0966_),
    .B1(net81));
 sg13g2_nand2_1 _4817_ (.Y(_0967_),
    .A(_0371_),
    .B(_0460_));
 sg13g2_nand2_1 _4818_ (.Y(_0968_),
    .A(_0966_),
    .B(_0967_));
 sg13g2_nand3_1 _4819_ (.B(net94),
    .C(net27),
    .A(net71),
    .Y(_0969_));
 sg13g2_a21oi_1 _4820_ (.A1(_0969_),
    .A2(_1293_),
    .Y(_0970_),
    .B1(net40));
 sg13g2_nor2_2 _4821_ (.A(net198),
    .B(_2687_),
    .Y(_0971_));
 sg13g2_inv_1 _4822_ (.Y(_0972_),
    .A(_2947_));
 sg13g2_a21oi_1 _4823_ (.A1(_0971_),
    .A2(_0972_),
    .Y(_0973_),
    .B1(net203));
 sg13g2_nor2b_1 _4824_ (.A(_0970_),
    .B_N(_0973_),
    .Y(_0974_));
 sg13g2_nand2_1 _4825_ (.Y(_0975_),
    .A(_0968_),
    .B(_0974_));
 sg13g2_nand2_2 _4826_ (.Y(_0977_),
    .A(_0142_),
    .B(_2411_));
 sg13g2_a21oi_1 _4827_ (.A1(_0321_),
    .A2(_0977_),
    .Y(_0978_),
    .B1(net54));
 sg13g2_nand2_1 _4828_ (.Y(_0979_),
    .A(_0703_),
    .B(net65));
 sg13g2_nand2_1 _4829_ (.Y(_0980_),
    .A(_0979_),
    .B(net169));
 sg13g2_nor2_1 _4830_ (.A(_0978_),
    .B(_0980_),
    .Y(_0981_));
 sg13g2_nand2_1 _4831_ (.Y(_0982_),
    .A(_2800_),
    .B(net97));
 sg13g2_nand2_1 _4832_ (.Y(_0983_),
    .A(_0982_),
    .B(_2842_));
 sg13g2_nand2_1 _4833_ (.Y(_0984_),
    .A(_0983_),
    .B(_2703_));
 sg13g2_nand2_1 _4834_ (.Y(_0985_),
    .A(_0984_),
    .B(net46));
 sg13g2_nand2_1 _4835_ (.Y(_0986_),
    .A(_2881_),
    .B(net50));
 sg13g2_nand3_1 _4836_ (.B(_0985_),
    .C(_0986_),
    .A(_0981_),
    .Y(_0988_));
 sg13g2_nand3_1 _4837_ (.B(_0988_),
    .C(net147),
    .A(_0975_),
    .Y(_0989_));
 sg13g2_nand2_1 _4838_ (.Y(_0990_),
    .A(_1446_),
    .B(_2399_));
 sg13g2_nand2_1 _4839_ (.Y(_0991_),
    .A(_0990_),
    .B(net56));
 sg13g2_nand3_1 _4840_ (.B(net67),
    .C(_0354_),
    .A(_0991_),
    .Y(_0992_));
 sg13g2_a21oi_1 _4841_ (.A1(_0919_),
    .A2(net45),
    .Y(_0993_),
    .B1(net172));
 sg13g2_nand2_1 _4842_ (.Y(_0994_),
    .A(_0992_),
    .B(_0993_));
 sg13g2_a21oi_2 _4843_ (.B1(_2450_),
    .Y(_0995_),
    .A2(net139),
    .A1(_2440_));
 sg13g2_nand3_1 _4844_ (.B(net67),
    .C(_0995_),
    .A(_2932_),
    .Y(_0996_));
 sg13g2_a22oi_1 _4845_ (.Y(_0997_),
    .B1(net86),
    .B2(net44),
    .A2(_1478_),
    .A1(net27));
 sg13g2_a21oi_1 _4846_ (.A1(net47),
    .A2(_0527_),
    .Y(_0999_),
    .B1(_2653_));
 sg13g2_a21oi_1 _4847_ (.A1(_0997_),
    .A2(_0999_),
    .Y(_1000_),
    .B1(net78));
 sg13g2_nand2_1 _4848_ (.Y(_1001_),
    .A(_0996_),
    .B(_1000_));
 sg13g2_nand2_1 _4849_ (.Y(_1002_),
    .A(_0994_),
    .B(_1001_));
 sg13g2_nand2_1 _4850_ (.Y(_1003_),
    .A(_1002_),
    .B(_2559_));
 sg13g2_nand2_1 _4851_ (.Y(_1004_),
    .A(_2948_),
    .B(net125));
 sg13g2_nor3_1 _4852_ (.A(net36),
    .B(net168),
    .C(_2745_),
    .Y(_1005_));
 sg13g2_nand3_1 _4853_ (.B(net82),
    .C(net48),
    .A(net71),
    .Y(_1006_));
 sg13g2_nand2_1 _4854_ (.Y(_1007_),
    .A(_1006_),
    .B(_0167_));
 sg13g2_inv_1 _4855_ (.Y(_1008_),
    .A(_0795_));
 sg13g2_a21oi_1 _4856_ (.A1(_1008_),
    .A2(_2705_),
    .Y(_1010_),
    .B1(net78));
 sg13g2_a22oi_1 _4857_ (.Y(_1011_),
    .B1(_1007_),
    .B2(_1010_),
    .A2(_1005_),
    .A1(_1004_));
 sg13g2_nor2_1 _4858_ (.A(net210),
    .B(_0478_),
    .Y(_1012_));
 sg13g2_inv_2 _4859_ (.Y(_1013_),
    .A(_1012_));
 sg13g2_nand2_1 _4860_ (.Y(_1014_),
    .A(_1011_),
    .B(_1013_));
 sg13g2_nand2_1 _4861_ (.Y(_1015_),
    .A(_1014_),
    .B(_2373_));
 sg13g2_nand3_1 _4862_ (.B(_1003_),
    .C(_1015_),
    .A(_0989_),
    .Y(_1016_));
 sg13g2_nand3_1 _4863_ (.B(_2727_),
    .C(_2654_),
    .A(_2850_),
    .Y(_1017_));
 sg13g2_nand2_1 _4864_ (.Y(_1018_),
    .A(_0350_),
    .B(_0951_));
 sg13g2_nand3_1 _4865_ (.B(_2753_),
    .C(_2591_),
    .A(_1018_),
    .Y(_1019_));
 sg13g2_nand3_1 _4866_ (.B(_1019_),
    .C(_2733_),
    .A(_1017_),
    .Y(_1021_));
 sg13g2_a21oi_1 _4867_ (.A1(_0150_),
    .A2(_2727_),
    .Y(_1022_),
    .B1(_2390_));
 sg13g2_nand2_1 _4868_ (.Y(_1023_),
    .A(_0240_),
    .B(_2935_));
 sg13g2_o21ai_1 _4869_ (.B1(_2698_),
    .Y(_1024_),
    .A1(_1023_),
    .A2(_2657_));
 sg13g2_nor2_1 _4870_ (.A(_1022_),
    .B(_1024_),
    .Y(_1025_));
 sg13g2_nand2_1 _4871_ (.Y(_1026_),
    .A(_1021_),
    .B(_1025_));
 sg13g2_nand2_1 _4872_ (.Y(_1027_),
    .A(_0438_),
    .B(_0602_));
 sg13g2_nand3_1 _4873_ (.B(net65),
    .C(net98),
    .A(_2793_),
    .Y(_1028_));
 sg13g2_o21ai_1 _4874_ (.B1(_1028_),
    .Y(_1029_),
    .A1(net28),
    .A2(_1027_));
 sg13g2_nand2_1 _4875_ (.Y(_1030_),
    .A(_1013_),
    .B(net169));
 sg13g2_nor2_1 _4876_ (.A(_1029_),
    .B(_1030_),
    .Y(_1032_));
 sg13g2_nand2_1 _4877_ (.Y(_1033_),
    .A(_2592_),
    .B(net53));
 sg13g2_a21oi_1 _4878_ (.A1(_1032_),
    .A2(_1033_),
    .Y(_1034_),
    .B1(_2597_));
 sg13g2_a21oi_1 _4879_ (.A1(_1026_),
    .A2(_1034_),
    .Y(_1035_),
    .B1(_2609_));
 sg13g2_nor2_1 _4880_ (.A(net122),
    .B(net59),
    .Y(_1036_));
 sg13g2_nor3_1 _4881_ (.A(net91),
    .B(_2279_),
    .C(_1036_),
    .Y(_1037_));
 sg13g2_nand2_1 _4882_ (.Y(_1038_),
    .A(_2571_),
    .B(net44));
 sg13g2_nand2_1 _4883_ (.Y(_1039_),
    .A(_1038_),
    .B(net108));
 sg13g2_a21oi_1 _4884_ (.A1(_0350_),
    .A2(_0951_),
    .Y(_1040_),
    .B1(_1039_));
 sg13g2_nor3_1 _4885_ (.A(_2760_),
    .B(_1037_),
    .C(_1040_),
    .Y(_1041_));
 sg13g2_a21oi_1 _4886_ (.A1(_2797_),
    .A2(_0135_),
    .Y(_1043_),
    .B1(_2445_));
 sg13g2_nand2_1 _4887_ (.Y(_1044_),
    .A(net71),
    .B(_1184_));
 sg13g2_nor2_2 _4888_ (.A(net180),
    .B(_2701_),
    .Y(_1045_));
 sg13g2_a21oi_1 _4889_ (.A1(_1044_),
    .A2(_1045_),
    .Y(_1046_),
    .B1(_3039_));
 sg13g2_nand2b_1 _4890_ (.Y(_1047_),
    .B(_1046_),
    .A_N(_1043_));
 sg13g2_nor2_1 _4891_ (.A(_1041_),
    .B(_1047_),
    .Y(_1048_));
 sg13g2_nor2_1 _4892_ (.A(_0729_),
    .B(_1048_),
    .Y(_1049_));
 sg13g2_nor2_1 _4893_ (.A(net140),
    .B(net95),
    .Y(_1050_));
 sg13g2_nor2_1 _4894_ (.A(_0264_),
    .B(_1050_),
    .Y(_1051_));
 sg13g2_a21oi_1 _4895_ (.A1(_1051_),
    .A2(_0110_),
    .Y(_1052_),
    .B1(net169));
 sg13g2_nand3_1 _4896_ (.B(net133),
    .C(_0422_),
    .A(_2577_),
    .Y(_1054_));
 sg13g2_a21oi_1 _4897_ (.A1(_1052_),
    .A2(_1054_),
    .Y(_1055_),
    .B1(_2141_));
 sg13g2_nand3_1 _4898_ (.B(net109),
    .C(_2554_),
    .A(_2487_),
    .Y(_1056_));
 sg13g2_nor2_1 _4899_ (.A(_2513_),
    .B(net148),
    .Y(_1057_));
 sg13g2_nor2_1 _4900_ (.A(net179),
    .B(_1057_),
    .Y(_1058_));
 sg13g2_a21oi_1 _4901_ (.A1(_1056_),
    .A2(_1058_),
    .Y(_1059_),
    .B1(net172));
 sg13g2_nand3_1 _4902_ (.B(net67),
    .C(_0418_),
    .A(_2579_),
    .Y(_1060_));
 sg13g2_a22oi_1 _4903_ (.Y(_1061_),
    .B1(_1059_),
    .B2(_1060_),
    .A2(_0324_),
    .A1(net25));
 sg13g2_nand2b_1 _4904_ (.Y(_1062_),
    .B(_1061_),
    .A_N(_1055_));
 sg13g2_nand2_1 _4905_ (.Y(_1063_),
    .A(_1049_),
    .B(_1062_));
 sg13g2_nand2_1 _4906_ (.Y(_1065_),
    .A(_1035_),
    .B(_1063_));
 sg13g2_a21oi_1 _4907_ (.A1(_1016_),
    .A2(net132),
    .Y(_1066_),
    .B1(_1065_));
 sg13g2_nor2_1 _4908_ (.A(_0964_),
    .B(_1066_),
    .Y(_0027_));
 sg13g2_nand3_1 _4909_ (.B(_2727_),
    .C(net84),
    .A(_0838_),
    .Y(_1067_));
 sg13g2_a21oi_1 _4910_ (.A1(_2743_),
    .A2(_0808_),
    .Y(_1068_),
    .B1(net162));
 sg13g2_nand2_1 _4911_ (.Y(_1069_),
    .A(_1067_),
    .B(_1068_));
 sg13g2_o21ai_1 _4912_ (.B1(net25),
    .Y(_1070_),
    .A1(_2723_),
    .A2(_0145_));
 sg13g2_nor2_1 _4913_ (.A(_1685_),
    .B(_0795_),
    .Y(_1071_));
 sg13g2_nand2b_1 _4914_ (.Y(_1072_),
    .B(_1071_),
    .A_N(_2772_));
 sg13g2_nand4_1 _4915_ (.B(_1070_),
    .C(net80),
    .A(_1069_),
    .Y(_1073_),
    .D(_1072_));
 sg13g2_a21oi_1 _4916_ (.A1(_0234_),
    .A2(_0977_),
    .Y(_1075_),
    .B1(net23));
 sg13g2_nand3_1 _4917_ (.B(net38),
    .C(net65),
    .A(net57),
    .Y(_1076_));
 sg13g2_nor2_1 _4918_ (.A(_0651_),
    .B(_1027_),
    .Y(_1077_));
 sg13g2_nor2_1 _4919_ (.A(_2480_),
    .B(_1077_),
    .Y(_1078_));
 sg13g2_nand3b_1 _4920_ (.B(_1076_),
    .C(_1078_),
    .Y(_1079_),
    .A_N(_1075_));
 sg13g2_a21oi_1 _4921_ (.A1(_1073_),
    .A2(_1079_),
    .Y(_1080_),
    .B1(_2597_));
 sg13g2_nand2_1 _4922_ (.Y(_1081_),
    .A(_2477_),
    .B(net133));
 sg13g2_a22oi_1 _4923_ (.Y(_1082_),
    .B1(_2552_),
    .B2(_2892_),
    .A2(_1081_),
    .A1(_1045_));
 sg13g2_inv_1 _4924_ (.Y(_1083_),
    .A(_2642_));
 sg13g2_nand3_1 _4925_ (.B(_2779_),
    .C(net199),
    .A(_1083_),
    .Y(_1084_));
 sg13g2_a21oi_1 _4926_ (.A1(_1082_),
    .A2(_1084_),
    .Y(_1086_),
    .B1(net123));
 sg13g2_a221oi_1 _4927_ (.B2(_0627_),
    .C1(_0338_),
    .B1(_3030_),
    .A1(_2789_),
    .Y(_1087_),
    .A2(net120));
 sg13g2_nand2_1 _4928_ (.Y(_1088_),
    .A(_0438_),
    .B(_2482_));
 sg13g2_inv_1 _4929_ (.Y(_1089_),
    .A(_1088_));
 sg13g2_a21oi_1 _4930_ (.A1(net77),
    .A2(_2800_),
    .Y(_1090_),
    .B1(_1958_));
 sg13g2_o21ai_1 _4931_ (.B1(_0521_),
    .Y(_1091_),
    .A1(_1089_),
    .A2(_1090_));
 sg13g2_nand2_1 _4932_ (.Y(_1092_),
    .A(_1091_),
    .B(net112));
 sg13g2_nor3_1 _4933_ (.A(_1086_),
    .B(_1087_),
    .C(_1092_),
    .Y(_1093_));
 sg13g2_o21ai_1 _4934_ (.B1(_0394_),
    .Y(_1094_),
    .A1(_2680_),
    .A2(_2848_));
 sg13g2_a22oi_1 _4935_ (.Y(_1095_),
    .B1(_2568_),
    .B2(_1094_),
    .A2(_0360_),
    .A1(_0565_));
 sg13g2_nand2_1 _4936_ (.Y(_1097_),
    .A(_0428_),
    .B(_2496_));
 sg13g2_o21ai_1 _4937_ (.B1(net42),
    .Y(_1098_),
    .A1(_0477_),
    .A2(_1097_));
 sg13g2_nand2_1 _4938_ (.Y(_1099_),
    .A(_1095_),
    .B(_1098_));
 sg13g2_nand2_1 _4939_ (.Y(_1100_),
    .A(_1099_),
    .B(_2699_));
 sg13g2_nand2_1 _4940_ (.Y(_1101_),
    .A(_1093_),
    .B(_1100_));
 sg13g2_nand2_1 _4941_ (.Y(_1102_),
    .A(_1101_),
    .B(net195));
 sg13g2_nor2_1 _4942_ (.A(_1080_),
    .B(_1102_),
    .Y(_1103_));
 sg13g2_nor2_2 _4943_ (.A(net179),
    .B(_0477_),
    .Y(_1104_));
 sg13g2_nor2_1 _4944_ (.A(_2577_),
    .B(_2478_),
    .Y(_1105_));
 sg13g2_nor2_1 _4945_ (.A(_2642_),
    .B(_1105_),
    .Y(_1106_));
 sg13g2_nor2_1 _4946_ (.A(_1104_),
    .B(_1106_),
    .Y(_1108_));
 sg13g2_nand2_1 _4947_ (.Y(_1109_),
    .A(net94),
    .B(net133));
 sg13g2_a21o_1 _4948_ (.A2(_2482_),
    .A1(_1109_),
    .B1(_0576_),
    .X(_1110_));
 sg13g2_a22oi_1 _4949_ (.Y(_1111_),
    .B1(_2053_),
    .B2(_1110_),
    .A2(_2141_),
    .A1(_1108_));
 sg13g2_nor3_1 _4950_ (.A(_2518_),
    .B(_2512_),
    .C(_0148_),
    .Y(_1112_));
 sg13g2_nand2_1 _4951_ (.Y(_1113_),
    .A(_1112_),
    .B(_1004_));
 sg13g2_nand2_1 _4952_ (.Y(_1114_),
    .A(_2992_),
    .B(net82));
 sg13g2_nand3_1 _4953_ (.B(_1114_),
    .C(_2753_),
    .A(_1038_),
    .Y(_1115_));
 sg13g2_nand3_1 _4954_ (.B(_1115_),
    .C(_0511_),
    .A(_1113_),
    .Y(_1116_));
 sg13g2_a22oi_1 _4955_ (.Y(_1117_),
    .B1(_0321_),
    .B2(_0769_),
    .A2(_2964_),
    .A1(_2715_));
 sg13g2_nand2_1 _4956_ (.Y(_1119_),
    .A(_1117_),
    .B(_0521_));
 sg13g2_nand3_1 _4957_ (.B(_1116_),
    .C(_1119_),
    .A(_1111_),
    .Y(_1120_));
 sg13g2_nand2_1 _4958_ (.Y(_1121_),
    .A(_1120_),
    .B(_2736_));
 sg13g2_a21oi_1 _4959_ (.A1(_0743_),
    .A2(_3043_),
    .Y(_1122_),
    .B1(net61));
 sg13g2_nor2_1 _4960_ (.A(net28),
    .B(_0226_),
    .Y(_1123_));
 sg13g2_inv_1 _4961_ (.Y(_1124_),
    .A(_2462_));
 sg13g2_nand2_1 _4962_ (.Y(_1125_),
    .A(_1124_),
    .B(net173));
 sg13g2_a21oi_1 _4963_ (.A1(_1293_),
    .A2(_2681_),
    .Y(_1126_),
    .B1(net138));
 sg13g2_nor3_1 _4964_ (.A(_1123_),
    .B(_1125_),
    .C(_1126_),
    .Y(_1127_));
 sg13g2_nor3_1 _4965_ (.A(net56),
    .B(_2411_),
    .C(_0289_),
    .Y(_1128_));
 sg13g2_o21ai_1 _4966_ (.B1(net53),
    .Y(_1130_),
    .A1(_2520_),
    .A2(_1128_));
 sg13g2_nand3b_1 _4967_ (.B(_1127_),
    .C(_1130_),
    .Y(_1131_),
    .A_N(_1122_));
 sg13g2_nand2_1 _4968_ (.Y(_1132_),
    .A(_2901_),
    .B(_2444_));
 sg13g2_a22oi_1 _4969_ (.Y(_1133_),
    .B1(net50),
    .B2(_1132_),
    .A2(_0532_),
    .A1(_0264_));
 sg13g2_o21ai_1 _4970_ (.B1(net32),
    .Y(_1134_),
    .A1(_2470_),
    .A2(_2880_));
 sg13g2_a21oi_2 _4971_ (.B1(_2460_),
    .Y(_1135_),
    .A2(net124),
    .A1(_1089_));
 sg13g2_nand3_1 _4972_ (.B(_1134_),
    .C(_1135_),
    .A(_1133_),
    .Y(_1136_));
 sg13g2_nand3_1 _4973_ (.B(_2785_),
    .C(_1136_),
    .A(_1131_),
    .Y(_1137_));
 sg13g2_nand3_1 _4974_ (.B(_1137_),
    .C(_2738_),
    .A(_1121_),
    .Y(_1138_));
 sg13g2_nand2_1 _4975_ (.Y(_1139_),
    .A(_1103_),
    .B(_1138_));
 sg13g2_a21oi_1 _4976_ (.A1(net52),
    .A2(net185),
    .Y(_1141_),
    .B1(net108));
 sg13g2_nand3_1 _4977_ (.B(_2856_),
    .C(net176),
    .A(_1141_),
    .Y(_1142_));
 sg13g2_nand3_1 _4978_ (.B(net89),
    .C(_0848_),
    .A(_2239_),
    .Y(_1143_));
 sg13g2_nand3_1 _4979_ (.B(_1143_),
    .C(_2760_),
    .A(_1142_),
    .Y(_1144_));
 sg13g2_nor2_1 _4980_ (.A(_1555_),
    .B(_1869_),
    .Y(_1145_));
 sg13g2_o21ai_1 _4981_ (.B1(_1145_),
    .Y(_1146_),
    .A1(_0198_),
    .A2(_2572_));
 sg13g2_a21oi_1 _4982_ (.A1(_0443_),
    .A2(net89),
    .Y(_1147_),
    .B1(_2544_));
 sg13g2_nand2_1 _4983_ (.Y(_1148_),
    .A(_1146_),
    .B(_1147_));
 sg13g2_a21oi_1 _4984_ (.A1(_1144_),
    .A2(_1148_),
    .Y(_1149_),
    .B1(_3040_));
 sg13g2_nor3_1 _4985_ (.A(net66),
    .B(net41),
    .C(_2947_),
    .Y(_1150_));
 sg13g2_a21oi_1 _4986_ (.A1(_2843_),
    .A2(_0478_),
    .Y(_1152_),
    .B1(net66));
 sg13g2_a21oi_1 _4987_ (.A1(_0333_),
    .A2(_0309_),
    .Y(_1153_),
    .B1(_0916_));
 sg13g2_nor4_1 _4988_ (.A(net197),
    .B(_1150_),
    .C(_1152_),
    .D(_1153_),
    .Y(_1154_));
 sg13g2_nand2b_1 _4989_ (.Y(_1155_),
    .B(_1154_),
    .A_N(_1149_));
 sg13g2_nand2_1 _4990_ (.Y(_1156_),
    .A(_0556_),
    .B(net30));
 sg13g2_nand3_1 _4991_ (.B(_0161_),
    .C(_2221_),
    .A(_1156_),
    .Y(_1157_));
 sg13g2_inv_1 _4992_ (.Y(_1158_),
    .A(net156));
 sg13g2_nor2_1 _4993_ (.A(net106),
    .B(_1158_),
    .Y(_1159_));
 sg13g2_inv_1 _4994_ (.Y(_1160_),
    .A(_1159_));
 sg13g2_a21oi_1 _4995_ (.A1(_1160_),
    .A2(net45),
    .Y(_1161_),
    .B1(net160));
 sg13g2_a21oi_1 _4996_ (.A1(_1157_),
    .A2(_1161_),
    .Y(_1163_),
    .B1(net175));
 sg13g2_nand2_1 _4997_ (.Y(_1164_),
    .A(net34),
    .B(net57));
 sg13g2_nand2_1 _4998_ (.Y(_1165_),
    .A(_1164_),
    .B(net102));
 sg13g2_nand2_1 _4999_ (.Y(_1166_),
    .A(_1165_),
    .B(_1880_));
 sg13g2_inv_2 _5000_ (.Y(_1167_),
    .A(_0651_));
 sg13g2_nand3_1 _5001_ (.B(_2749_),
    .C(_1167_),
    .A(_1166_),
    .Y(_1168_));
 sg13g2_inv_1 _5002_ (.Y(_1169_),
    .A(_0175_));
 sg13g2_o21ai_1 _5003_ (.B1(net172),
    .Y(_1170_),
    .A1(_0266_),
    .A2(_1169_));
 sg13g2_nand2_1 _5004_ (.Y(_1171_),
    .A(_0099_),
    .B(net58));
 sg13g2_nand3_1 _5005_ (.B(_0825_),
    .C(_2716_),
    .A(_1171_),
    .Y(_1172_));
 sg13g2_nand3_1 _5006_ (.B(_0748_),
    .C(_1172_),
    .A(_1170_),
    .Y(_1174_));
 sg13g2_nand3_1 _5007_ (.B(_1168_),
    .C(_1174_),
    .A(_1163_),
    .Y(_1175_));
 sg13g2_nand2_1 _5008_ (.Y(_1176_),
    .A(_1155_),
    .B(_1175_));
 sg13g2_nand2_1 _5009_ (.Y(_1177_),
    .A(_1176_),
    .B(net132));
 sg13g2_inv_1 _5010_ (.Y(_1178_),
    .A(_2678_));
 sg13g2_a221oi_1 _5011_ (.B2(_2740_),
    .C1(_0303_),
    .B1(_0901_),
    .A1(_1178_),
    .Y(_1179_),
    .A2(_1104_));
 sg13g2_nor2_1 _5012_ (.A(net163),
    .B(_1179_),
    .Y(_1180_));
 sg13g2_a21oi_1 _5013_ (.A1(_0495_),
    .A2(_0326_),
    .Y(_1181_),
    .B1(_2642_));
 sg13g2_nand2_1 _5014_ (.Y(_1182_),
    .A(_0368_),
    .B(_2747_));
 sg13g2_nand3b_1 _5015_ (.B(net130),
    .C(_1182_),
    .Y(_1183_),
    .A_N(_1181_));
 sg13g2_nand3_1 _5016_ (.B(_2782_),
    .C(_2651_),
    .A(_2625_),
    .Y(_1185_));
 sg13g2_nand3_1 _5017_ (.B(net117),
    .C(_1185_),
    .A(_1183_),
    .Y(_1186_));
 sg13g2_nor3_1 _5018_ (.A(net171),
    .B(net41),
    .C(net52),
    .Y(_1187_));
 sg13g2_nor3_1 _5019_ (.A(net75),
    .B(_0128_),
    .C(_0808_),
    .Y(_1188_));
 sg13g2_a21oi_1 _5020_ (.A1(_0100_),
    .A2(net96),
    .Y(_1189_),
    .B1(net40));
 sg13g2_nor3_1 _5021_ (.A(_1187_),
    .B(_1188_),
    .C(_1189_),
    .Y(_1190_));
 sg13g2_a21oi_1 _5022_ (.A1(_1190_),
    .A2(net80),
    .Y(_1191_),
    .B1(net166));
 sg13g2_nand2_1 _5023_ (.Y(_1192_),
    .A(_1186_),
    .B(_1191_));
 sg13g2_a21oi_1 _5024_ (.A1(_1180_),
    .A2(_1192_),
    .Y(_1193_),
    .B1(net165));
 sg13g2_nand2_1 _5025_ (.Y(_1194_),
    .A(_1177_),
    .B(_1193_));
 sg13g2_nand2_1 _5026_ (.Y(_0028_),
    .A(_1139_),
    .B(_1194_));
 sg13g2_nand3_1 _5027_ (.B(net93),
    .C(_1848_),
    .A(_1413_),
    .Y(_1196_));
 sg13g2_buf_2 _5028_ (.A(_1196_),
    .X(_1197_));
 sg13g2_nand2_1 _5029_ (.Y(_1198_),
    .A(_1197_),
    .B(_0388_));
 sg13g2_a21oi_1 _5030_ (.A1(_1198_),
    .A2(net32),
    .Y(_1199_),
    .B1(_1125_));
 sg13g2_nand2_1 _5031_ (.Y(_1200_),
    .A(_0345_),
    .B(_2789_));
 sg13g2_nand2_1 _5032_ (.Y(_1201_),
    .A(_1200_),
    .B(net74));
 sg13g2_a21oi_1 _5033_ (.A1(_1199_),
    .A2(_1201_),
    .Y(_1202_),
    .B1(net147));
 sg13g2_o21ai_1 _5034_ (.B1(net55),
    .Y(_1203_),
    .A1(net33),
    .A2(_1164_));
 sg13g2_nand2_1 _5035_ (.Y(_1204_),
    .A(_2671_),
    .B(_1184_));
 sg13g2_nand2_1 _5036_ (.Y(_1206_),
    .A(_0558_),
    .B(_1204_));
 sg13g2_a21oi_1 _5037_ (.A1(_1206_),
    .A2(_2740_),
    .Y(_1207_),
    .B1(net78));
 sg13g2_nand2_1 _5038_ (.Y(_1208_),
    .A(_1203_),
    .B(_1207_));
 sg13g2_nor3_1 _5039_ (.A(net51),
    .B(_2575_),
    .C(_2848_),
    .Y(_1209_));
 sg13g2_nor3_1 _5040_ (.A(_2550_),
    .B(_0651_),
    .C(_1209_),
    .Y(_1210_));
 sg13g2_nor2_1 _5041_ (.A(net116),
    .B(_1210_),
    .Y(_1211_));
 sg13g2_nand2_1 _5042_ (.Y(_1212_),
    .A(_1208_),
    .B(_1211_));
 sg13g2_a21oi_1 _5043_ (.A1(_1202_),
    .A2(_1212_),
    .Y(_1213_),
    .B1(net195));
 sg13g2_nand2_1 _5044_ (.Y(_1214_),
    .A(_2900_),
    .B(_2704_));
 sg13g2_nand2_1 _5045_ (.Y(_1215_),
    .A(_0597_),
    .B(_1214_));
 sg13g2_nor2_1 _5046_ (.A(_2751_),
    .B(_1096_),
    .Y(_1217_));
 sg13g2_nand2_1 _5047_ (.Y(_1218_),
    .A(_2779_),
    .B(_1217_));
 sg13g2_nor2_1 _5048_ (.A(_2866_),
    .B(_1218_),
    .Y(_1219_));
 sg13g2_a21oi_1 _5049_ (.A1(_1215_),
    .A2(net39),
    .Y(_1220_),
    .B1(_1219_));
 sg13g2_nand2_1 _5050_ (.Y(_1221_),
    .A(_2529_),
    .B(_0142_));
 sg13g2_a21oi_1 _5051_ (.A1(_1145_),
    .A2(_1221_),
    .Y(_1222_),
    .B1(net199));
 sg13g2_nand2_1 _5052_ (.Y(_1223_),
    .A(_2428_),
    .B(_2509_));
 sg13g2_nand2_1 _5053_ (.Y(_1224_),
    .A(_1222_),
    .B(_1223_));
 sg13g2_nand2_1 _5054_ (.Y(_1225_),
    .A(_1220_),
    .B(_1224_));
 sg13g2_nand2_1 _5055_ (.Y(_1226_),
    .A(_1225_),
    .B(net121));
 sg13g2_nand2_1 _5056_ (.Y(_1228_),
    .A(_0564_),
    .B(_1083_));
 sg13g2_nor2_1 _5057_ (.A(_0337_),
    .B(_1008_),
    .Y(_1229_));
 sg13g2_o21ai_1 _5058_ (.B1(_2394_),
    .Y(_1230_),
    .A1(net47),
    .A2(net59));
 sg13g2_a22oi_1 _5059_ (.Y(_1231_),
    .B1(_0917_),
    .B2(_1230_),
    .A2(_1229_),
    .A1(_1228_));
 sg13g2_nand2_1 _5060_ (.Y(_1232_),
    .A(_1226_),
    .B(_1231_));
 sg13g2_nand2_1 _5061_ (.Y(_1233_),
    .A(_1232_),
    .B(net73));
 sg13g2_a21oi_1 _5062_ (.A1(_1213_),
    .A2(_1233_),
    .Y(_1234_),
    .B1(net200));
 sg13g2_a21oi_1 _5063_ (.A1(_2879_),
    .A2(_0387_),
    .Y(_1235_),
    .B1(net23));
 sg13g2_nand2_1 _5064_ (.Y(_1236_),
    .A(_2802_),
    .B(net65));
 sg13g2_nand2_1 _5065_ (.Y(_1237_),
    .A(_1135_),
    .B(_1236_));
 sg13g2_a21oi_1 _5066_ (.A1(_0345_),
    .A2(_0655_),
    .Y(_1239_),
    .B1(net31));
 sg13g2_nor3_1 _5067_ (.A(_1235_),
    .B(_1237_),
    .C(_1239_),
    .Y(_1240_));
 sg13g2_nor2_1 _5068_ (.A(net166),
    .B(_1240_),
    .Y(_1241_));
 sg13g2_nand2_1 _5069_ (.Y(_1242_),
    .A(_2428_),
    .B(_0309_));
 sg13g2_nand2_1 _5070_ (.Y(_1243_),
    .A(_3025_),
    .B(_0226_));
 sg13g2_a22oi_1 _5071_ (.Y(_1244_),
    .B1(net53),
    .B2(_1243_),
    .A2(net25),
    .A1(_1242_));
 sg13g2_nor2_1 _5072_ (.A(net177),
    .B(_1105_),
    .Y(_1245_));
 sg13g2_a21oi_1 _5073_ (.A1(_1245_),
    .A2(_0160_),
    .Y(_1246_),
    .B1(net199));
 sg13g2_nand2_1 _5074_ (.Y(_1247_),
    .A(_2919_),
    .B(_0744_));
 sg13g2_nand2_1 _5075_ (.Y(_1248_),
    .A(_1246_),
    .B(_1247_));
 sg13g2_nand3_1 _5076_ (.B(_1248_),
    .C(net83),
    .A(_1244_),
    .Y(_1250_));
 sg13g2_nand2_1 _5077_ (.Y(_1251_),
    .A(_1241_),
    .B(_1250_));
 sg13g2_a21oi_1 _5078_ (.A1(_2712_),
    .A2(_2637_),
    .Y(_1252_),
    .B1(_0651_));
 sg13g2_inv_1 _5079_ (.Y(_1253_),
    .A(_2659_));
 sg13g2_nor2_1 _5080_ (.A(net145),
    .B(_2920_),
    .Y(_1254_));
 sg13g2_a21oi_1 _5081_ (.A1(_1253_),
    .A2(_1045_),
    .Y(_1255_),
    .B1(_1254_));
 sg13g2_nand3b_1 _5082_ (.B(net83),
    .C(_1255_),
    .Y(_1256_),
    .A_N(_1252_));
 sg13g2_a21oi_1 _5083_ (.A1(_2879_),
    .A2(_0387_),
    .Y(_1257_),
    .B1(net31));
 sg13g2_nor2_1 _5084_ (.A(net91),
    .B(_2635_),
    .Y(_1258_));
 sg13g2_a21oi_1 _5085_ (.A1(_1258_),
    .A2(_1238_),
    .Y(_1259_),
    .B1(net78));
 sg13g2_nand2_1 _5086_ (.Y(_1261_),
    .A(_2625_),
    .B(_2539_));
 sg13g2_nand2_1 _5087_ (.Y(_1262_),
    .A(_1259_),
    .B(_1261_));
 sg13g2_nand2_1 _5088_ (.Y(_1263_),
    .A(_0093_),
    .B(_2637_));
 sg13g2_a21oi_1 _5089_ (.A1(_1263_),
    .A2(net74),
    .Y(_1264_),
    .B1(net127));
 sg13g2_nand3b_1 _5090_ (.B(_1262_),
    .C(_1264_),
    .Y(_1265_),
    .A_N(_1257_));
 sg13g2_nand3_1 _5091_ (.B(_1265_),
    .C(net164),
    .A(_1256_),
    .Y(_1266_));
 sg13g2_nand3_1 _5092_ (.B(_1266_),
    .C(_2696_),
    .A(_1251_),
    .Y(_1267_));
 sg13g2_nand2_1 _5093_ (.Y(_1268_),
    .A(_1234_),
    .B(_1267_));
 sg13g2_nand2_1 _5094_ (.Y(_1269_),
    .A(net38),
    .B(_2808_));
 sg13g2_o21ai_1 _5095_ (.B1(_2719_),
    .Y(_1270_),
    .A1(_2680_),
    .A2(_1269_));
 sg13g2_nand2_1 _5096_ (.Y(_1272_),
    .A(_1270_),
    .B(net32));
 sg13g2_nand2_1 _5097_ (.Y(_1273_),
    .A(_2796_),
    .B(_0532_));
 sg13g2_nand2_1 _5098_ (.Y(_1274_),
    .A(_1272_),
    .B(_1273_));
 sg13g2_nand2_1 _5099_ (.Y(_1275_),
    .A(_1274_),
    .B(_2699_));
 sg13g2_nand2_1 _5100_ (.Y(_1276_),
    .A(_0995_),
    .B(_2539_));
 sg13g2_nand2_1 _5101_ (.Y(_1277_),
    .A(net29),
    .B(net38));
 sg13g2_nand2_1 _5102_ (.Y(_1278_),
    .A(_0721_),
    .B(_1277_));
 sg13g2_nand3_1 _5103_ (.B(_1278_),
    .C(_0520_),
    .A(_1276_),
    .Y(_1279_));
 sg13g2_nand2_1 _5104_ (.Y(_1280_),
    .A(_1279_),
    .B(net175));
 sg13g2_o21ai_1 _5105_ (.B1(net110),
    .Y(_1281_),
    .A1(_1159_),
    .A2(_2981_));
 sg13g2_inv_1 _5106_ (.Y(_1283_),
    .A(_1045_));
 sg13g2_nor2_1 _5107_ (.A(_2947_),
    .B(_1283_),
    .Y(_1284_));
 sg13g2_nand2_1 _5108_ (.Y(_1285_),
    .A(_1284_),
    .B(net125));
 sg13g2_a21oi_1 _5109_ (.A1(_1281_),
    .A2(_1285_),
    .Y(_1286_),
    .B1(_2664_));
 sg13g2_nor2_1 _5110_ (.A(_1280_),
    .B(_1286_),
    .Y(_1287_));
 sg13g2_nand2_1 _5111_ (.Y(_1288_),
    .A(_2802_),
    .B(net102));
 sg13g2_nand3_1 _5112_ (.B(_2826_),
    .C(_3025_),
    .A(_1288_),
    .Y(_1289_));
 sg13g2_o21ai_1 _5113_ (.B1(_2983_),
    .Y(_1290_),
    .A1(net33),
    .A2(net34));
 sg13g2_nand3_1 _5114_ (.B(_1290_),
    .C(_0165_),
    .A(_1289_),
    .Y(_1291_));
 sg13g2_nand3_1 _5115_ (.B(_1287_),
    .C(_1291_),
    .A(_1275_),
    .Y(_1292_));
 sg13g2_and3_1 _5116_ (.X(_1294_),
    .A(net38),
    .B(_2686_),
    .C(_3014_));
 sg13g2_a21oi_1 _5117_ (.A1(_1206_),
    .A2(_2221_),
    .Y(_1295_),
    .B1(net67));
 sg13g2_nor2_1 _5118_ (.A(_0034_),
    .B(net161),
    .Y(_1296_));
 sg13g2_o21ai_1 _5119_ (.B1(_1296_),
    .Y(_1297_),
    .A1(_1294_),
    .A2(_1295_));
 sg13g2_nor2_1 _5120_ (.A(net76),
    .B(_0926_),
    .Y(_1298_));
 sg13g2_nand2_1 _5121_ (.Y(_1299_),
    .A(_1298_),
    .B(_0150_));
 sg13g2_o21ai_1 _5122_ (.B1(_1299_),
    .Y(_1300_),
    .A1(net67),
    .A2(_2530_));
 sg13g2_nand2_1 _5123_ (.Y(_1301_),
    .A(_1300_),
    .B(net105));
 sg13g2_a22oi_1 _5124_ (.Y(_1302_),
    .B1(_3030_),
    .B2(_0995_),
    .A2(_0609_),
    .A1(_0721_));
 sg13g2_a21oi_1 _5125_ (.A1(_1302_),
    .A2(_2141_),
    .Y(_1303_),
    .B1(net175));
 sg13g2_nand3_1 _5126_ (.B(_1301_),
    .C(_1303_),
    .A(_1297_),
    .Y(_1305_));
 sg13g2_nand2_1 _5127_ (.Y(_1306_),
    .A(_1292_),
    .B(_1305_));
 sg13g2_nand2_1 _5128_ (.Y(_1307_),
    .A(_1306_),
    .B(net165));
 sg13g2_inv_1 _5129_ (.Y(_1308_),
    .A(_2450_));
 sg13g2_nand3_1 _5130_ (.B(_1308_),
    .C(_0453_),
    .A(_1288_),
    .Y(_1309_));
 sg13g2_a21oi_1 _5131_ (.A1(_1197_),
    .A2(_2743_),
    .Y(_1310_),
    .B1(net81));
 sg13g2_nand2_1 _5132_ (.Y(_1311_),
    .A(_1309_),
    .B(_1310_));
 sg13g2_inv_1 _5133_ (.Y(_1312_),
    .A(_0199_));
 sg13g2_nand3b_1 _5134_ (.B(net74),
    .C(_1312_),
    .Y(_1313_),
    .A_N(_1209_));
 sg13g2_nand3_1 _5135_ (.B(net117),
    .C(_1313_),
    .A(_1311_),
    .Y(_1314_));
 sg13g2_nor3_1 _5136_ (.A(net107),
    .B(_0128_),
    .C(_2590_),
    .Y(_1316_));
 sg13g2_o21ai_1 _5137_ (.B1(net161),
    .Y(_1317_),
    .A1(net38),
    .A2(_2461_));
 sg13g2_nand2_1 _5138_ (.Y(_1318_),
    .A(_2582_),
    .B(net143));
 sg13g2_a21oi_1 _5139_ (.A1(_0096_),
    .A2(_1318_),
    .Y(_1319_),
    .B1(net40));
 sg13g2_nor3_1 _5140_ (.A(_1316_),
    .B(_1317_),
    .C(_1319_),
    .Y(_1320_));
 sg13g2_nor2_1 _5141_ (.A(net166),
    .B(_1320_),
    .Y(_1321_));
 sg13g2_nand2_1 _5142_ (.Y(_1322_),
    .A(_1314_),
    .B(_1321_));
 sg13g2_nor2_1 _5143_ (.A(_2739_),
    .B(_0656_),
    .Y(_1323_));
 sg13g2_a21oi_1 _5144_ (.A1(_0124_),
    .A2(net193),
    .Y(_1324_),
    .B1(net99));
 sg13g2_nor3_1 _5145_ (.A(_0303_),
    .B(_1323_),
    .C(_1324_),
    .Y(_1325_));
 sg13g2_nor2_1 _5146_ (.A(net195),
    .B(_1325_),
    .Y(_1327_));
 sg13g2_a21oi_1 _5147_ (.A1(_1322_),
    .A2(_1327_),
    .Y(_1328_),
    .B1(net132));
 sg13g2_nand2_1 _5148_ (.Y(_1329_),
    .A(_1307_),
    .B(_1328_));
 sg13g2_nand2_1 _5149_ (.Y(_0029_),
    .A(_1268_),
    .B(_1329_));
 sg13g2_nor2_1 _5150_ (.A(_2508_),
    .B(_2960_),
    .Y(_1330_));
 sg13g2_a21oi_1 _5151_ (.A1(_2492_),
    .A2(_1330_),
    .Y(_1331_),
    .B1(net124));
 sg13g2_nand2_1 _5152_ (.Y(_1332_),
    .A(_2471_),
    .B(net91));
 sg13g2_nand2_1 _5153_ (.Y(_1333_),
    .A(_1331_),
    .B(_1332_));
 sg13g2_nand3_1 _5154_ (.B(net127),
    .C(_1333_),
    .A(_1248_),
    .Y(_1334_));
 sg13g2_o21ai_1 _5155_ (.B1(net50),
    .Y(_1335_),
    .A1(_1930_),
    .A2(_0145_));
 sg13g2_nand2_1 _5156_ (.Y(_1337_),
    .A(_0825_),
    .B(_1085_));
 sg13g2_nor2_1 _5157_ (.A(net79),
    .B(_1044_),
    .Y(_1338_));
 sg13g2_nor2_1 _5158_ (.A(_1337_),
    .B(_1338_),
    .Y(_1339_));
 sg13g2_nand3_1 _5159_ (.B(net43),
    .C(_0531_),
    .A(net34),
    .Y(_1340_));
 sg13g2_nor2b_1 _5160_ (.A(_1339_),
    .B_N(_1340_),
    .Y(_1341_));
 sg13g2_nand3_1 _5161_ (.B(_1341_),
    .C(_1135_),
    .A(_1335_),
    .Y(_1342_));
 sg13g2_nand2_1 _5162_ (.Y(_1343_),
    .A(_1334_),
    .B(_1342_));
 sg13g2_nand2_1 _5163_ (.Y(_1344_),
    .A(_1343_),
    .B(_2360_));
 sg13g2_nor2_1 _5164_ (.A(net140),
    .B(_1162_),
    .Y(_1345_));
 sg13g2_nor3_1 _5165_ (.A(net76),
    .B(_0483_),
    .C(_1345_),
    .Y(_1346_));
 sg13g2_a21o_1 _5166_ (.A2(_1346_),
    .A1(_2394_),
    .B1(_2351_),
    .X(_1348_));
 sg13g2_o21ai_1 _5167_ (.B1(_0250_),
    .Y(_1349_),
    .A1(net48),
    .A2(_0332_));
 sg13g2_and2_1 _5168_ (.A(_1349_),
    .B(_0604_),
    .X(_1350_));
 sg13g2_nand2_1 _5169_ (.Y(_1351_),
    .A(_2897_),
    .B(net48));
 sg13g2_nand2_1 _5170_ (.Y(_1352_),
    .A(_1489_),
    .B(net137));
 sg13g2_nand3_1 _5171_ (.B(_0600_),
    .C(_1352_),
    .A(_1351_),
    .Y(_1353_));
 sg13g2_inv_1 _5172_ (.Y(_1354_),
    .A(_3005_));
 sg13g2_nand2_1 _5173_ (.Y(_1355_),
    .A(_1354_),
    .B(_3044_));
 sg13g2_nand2_1 _5174_ (.Y(_1356_),
    .A(_1355_),
    .B(_0866_));
 sg13g2_nand2_1 _5175_ (.Y(_1357_),
    .A(_1353_),
    .B(_1356_));
 sg13g2_nor3_1 _5176_ (.A(_1348_),
    .B(_1350_),
    .C(_1357_),
    .Y(_1359_));
 sg13g2_nand2_1 _5177_ (.Y(_1360_),
    .A(_0234_),
    .B(_0167_));
 sg13g2_nand2_1 _5178_ (.Y(_1361_),
    .A(_1008_),
    .B(_1293_));
 sg13g2_nand3_1 _5179_ (.B(_1361_),
    .C(net171),
    .A(_1360_),
    .Y(_1362_));
 sg13g2_nand2_1 _5180_ (.Y(_1363_),
    .A(_1318_),
    .B(_0468_));
 sg13g2_a21oi_1 _5181_ (.A1(_1363_),
    .A2(net49),
    .Y(_1364_),
    .B1(_1012_));
 sg13g2_nand2_1 _5182_ (.Y(_1365_),
    .A(_1362_),
    .B(_1364_));
 sg13g2_nand2_1 _5183_ (.Y(_1366_),
    .A(_1365_),
    .B(net116));
 sg13g2_a21oi_1 _5184_ (.A1(_1359_),
    .A2(_1366_),
    .Y(_1367_),
    .B1(_2424_));
 sg13g2_nand2_1 _5185_ (.Y(_1368_),
    .A(_1344_),
    .B(_1367_));
 sg13g2_inv_1 _5186_ (.Y(_1370_),
    .A(_2519_));
 sg13g2_nand3_1 _5187_ (.B(_1370_),
    .C(_0184_),
    .A(_0380_),
    .Y(_1371_));
 sg13g2_nor2_1 _5188_ (.A(_1369_),
    .B(net76),
    .Y(_1372_));
 sg13g2_nor2_1 _5189_ (.A(net75),
    .B(_3005_),
    .Y(_1373_));
 sg13g2_nand2_1 _5190_ (.Y(_1374_),
    .A(net96),
    .B(_1696_));
 sg13g2_o21ai_1 _5191_ (.B1(_0748_),
    .Y(_1375_),
    .A1(_1374_),
    .A2(_2739_));
 sg13g2_a21oi_1 _5192_ (.A1(_2879_),
    .A2(_1373_),
    .Y(_1376_),
    .B1(_1375_));
 sg13g2_a21oi_1 _5193_ (.A1(_1371_),
    .A2(_1372_),
    .Y(_1377_),
    .B1(_1376_));
 sg13g2_o21ai_1 _5194_ (.B1(net69),
    .Y(_1378_),
    .A1(_2739_),
    .A2(_3005_));
 sg13g2_nand3_1 _5195_ (.B(_1013_),
    .C(_1340_),
    .A(_1378_),
    .Y(_1379_));
 sg13g2_nand2_1 _5196_ (.Y(_1381_),
    .A(_1379_),
    .B(net121));
 sg13g2_a21oi_1 _5197_ (.A1(_1377_),
    .A2(_1381_),
    .Y(_1382_),
    .B1(_2597_));
 sg13g2_a21oi_1 _5198_ (.A1(_2871_),
    .A2(_2583_),
    .Y(_1383_),
    .B1(net108));
 sg13g2_nand2_1 _5199_ (.Y(_1384_),
    .A(_1383_),
    .B(_2959_));
 sg13g2_nand2_1 _5200_ (.Y(_1385_),
    .A(_3046_),
    .B(_0352_));
 sg13g2_nand3_1 _5201_ (.B(_2600_),
    .C(_1385_),
    .A(_1384_),
    .Y(_1386_));
 sg13g2_nor2_1 _5202_ (.A(net135),
    .B(_0784_),
    .Y(_1387_));
 sg13g2_nand2_1 _5203_ (.Y(_1388_),
    .A(_1387_),
    .B(_1318_));
 sg13g2_nand2_1 _5204_ (.Y(_1389_),
    .A(_0234_),
    .B(_1058_));
 sg13g2_nand3_1 _5205_ (.B(_1389_),
    .C(net75),
    .A(_1388_),
    .Y(_1390_));
 sg13g2_nand3_1 _5206_ (.B(_2664_),
    .C(_1390_),
    .A(_1386_),
    .Y(_1392_));
 sg13g2_nand2_1 _5207_ (.Y(_1393_),
    .A(_1354_),
    .B(net128));
 sg13g2_a21oi_1 _5208_ (.A1(_0514_),
    .A2(_2661_),
    .Y(_1394_),
    .B1(net199));
 sg13g2_o21ai_1 _5209_ (.B1(_1394_),
    .Y(_1395_),
    .A1(_0324_),
    .A2(_1393_));
 sg13g2_nand2_1 _5210_ (.Y(_1396_),
    .A(net52),
    .B(_2437_));
 sg13g2_nand2_1 _5211_ (.Y(_1397_),
    .A(_0332_),
    .B(_1336_));
 sg13g2_a21oi_1 _5212_ (.A1(_0808_),
    .A2(_1396_),
    .Y(_1398_),
    .B1(_1397_));
 sg13g2_nor3_1 _5213_ (.A(net161),
    .B(_1284_),
    .C(_1398_),
    .Y(_1399_));
 sg13g2_nand2_1 _5214_ (.Y(_1400_),
    .A(_1395_),
    .B(_1399_));
 sg13g2_nand2_1 _5215_ (.Y(_1401_),
    .A(_1392_),
    .B(_1400_));
 sg13g2_nor2_1 _5216_ (.A(_0729_),
    .B(_1401_),
    .Y(_1403_));
 sg13g2_nor2_1 _5217_ (.A(_1382_),
    .B(_1403_),
    .Y(_1404_));
 sg13g2_nand2_1 _5218_ (.Y(_1405_),
    .A(_1368_),
    .B(_1404_));
 sg13g2_nand2_1 _5219_ (.Y(_1406_),
    .A(_1405_),
    .B(net165));
 sg13g2_nand2_1 _5220_ (.Y(_1407_),
    .A(_2684_),
    .B(_2649_));
 sg13g2_a21oi_1 _5221_ (.A1(_3019_),
    .A2(_1407_),
    .Y(_1408_),
    .B1(net61));
 sg13g2_o21ai_1 _5222_ (.B1(net88),
    .Y(_1409_),
    .A1(_0276_),
    .A2(_0918_));
 sg13g2_nand2_1 _5223_ (.Y(_1410_),
    .A(_1409_),
    .B(_1124_));
 sg13g2_o21ai_1 _5224_ (.B1(_2373_),
    .Y(_1411_),
    .A1(_1408_),
    .A2(_1410_));
 sg13g2_nand2_1 _5225_ (.Y(_1412_),
    .A(_1411_),
    .B(net170));
 sg13g2_nor2b_1 _5226_ (.A(_0449_),
    .B_N(_0833_),
    .Y(_1414_));
 sg13g2_nand2_1 _5227_ (.Y(_1415_),
    .A(_0791_),
    .B(net133));
 sg13g2_nor2_1 _5228_ (.A(net138),
    .B(_2440_),
    .Y(_1416_));
 sg13g2_nand2_1 _5229_ (.Y(_1417_),
    .A(_1880_),
    .B(net148));
 sg13g2_a22oi_1 _5230_ (.Y(_1418_),
    .B1(_1167_),
    .B2(_1417_),
    .A2(_1416_),
    .A1(_1415_));
 sg13g2_o21ai_1 _5231_ (.B1(_1418_),
    .Y(_1419_),
    .A1(net23),
    .A2(_1414_));
 sg13g2_nand2_1 _5232_ (.Y(_1420_),
    .A(_1419_),
    .B(_2559_));
 sg13g2_nor2b_1 _5233_ (.A(_1412_),
    .B_N(_1420_),
    .Y(_1421_));
 sg13g2_nand3b_1 _5234_ (.B(_2747_),
    .C(_3003_),
    .Y(_1422_),
    .A_N(_0501_));
 sg13g2_a21oi_1 _5235_ (.A1(_1422_),
    .A2(_0915_),
    .Y(_1423_),
    .B1(_2749_));
 sg13g2_nor2b_1 _5236_ (.A(_2819_),
    .B_N(_3003_),
    .Y(_1425_));
 sg13g2_nand3_1 _5237_ (.B(_0161_),
    .C(_2727_),
    .A(_1425_),
    .Y(_1426_));
 sg13g2_a21oi_1 _5238_ (.A1(_2605_),
    .A2(net45),
    .Y(_1427_),
    .B1(net162));
 sg13g2_nand2_1 _5239_ (.Y(_1428_),
    .A(_1426_),
    .B(_1427_));
 sg13g2_nand4_1 _5240_ (.B(net67),
    .C(net176),
    .A(_0597_),
    .Y(_1429_),
    .D(net113));
 sg13g2_nand2_1 _5241_ (.Y(_1430_),
    .A(_1429_),
    .B(_2351_));
 sg13g2_a21oi_1 _5242_ (.A1(_1423_),
    .A2(_1428_),
    .Y(_1431_),
    .B1(_1430_));
 sg13g2_nand2_1 _5243_ (.Y(_1432_),
    .A(_0393_),
    .B(_2900_));
 sg13g2_a22oi_1 _5244_ (.Y(_1433_),
    .B1(_1145_),
    .B2(_1432_),
    .A2(net45),
    .A1(_3036_));
 sg13g2_nand2_1 _5245_ (.Y(_1434_),
    .A(_2571_),
    .B(_2603_));
 sg13g2_nand3_1 _5246_ (.B(_2993_),
    .C(_0334_),
    .A(_1434_),
    .Y(_1436_));
 sg13g2_o21ai_1 _5247_ (.B1(_1436_),
    .Y(_1437_),
    .A1(_2601_),
    .A2(_1433_));
 sg13g2_nand2_1 _5248_ (.Y(_1438_),
    .A(_1437_),
    .B(net117));
 sg13g2_nand2_1 _5249_ (.Y(_1439_),
    .A(_1431_),
    .B(_1438_));
 sg13g2_nand2_1 _5250_ (.Y(_1440_),
    .A(_1421_),
    .B(_1439_));
 sg13g2_o21ai_1 _5251_ (.B1(_2579_),
    .Y(_1441_),
    .A1(net30),
    .A2(_0426_));
 sg13g2_nand2_1 _5252_ (.Y(_1442_),
    .A(_1441_),
    .B(net70));
 sg13g2_nand2_1 _5253_ (.Y(_1443_),
    .A(_1312_),
    .B(_2743_));
 sg13g2_nand2_1 _5254_ (.Y(_1444_),
    .A(net38),
    .B(net126));
 sg13g2_nor2_1 _5255_ (.A(net91),
    .B(_0527_),
    .Y(_1445_));
 sg13g2_o21ai_1 _5256_ (.B1(_1445_),
    .Y(_1447_),
    .A1(net139),
    .A2(_1444_));
 sg13g2_nand3_1 _5257_ (.B(net130),
    .C(_1447_),
    .A(_1443_),
    .Y(_1448_));
 sg13g2_nand3_1 _5258_ (.B(_1448_),
    .C(_2596_),
    .A(_1442_),
    .Y(_1449_));
 sg13g2_o21ai_1 _5259_ (.B1(net70),
    .Y(_1450_),
    .A1(_2889_),
    .A2(_0516_));
 sg13g2_a21oi_1 _5260_ (.A1(net156),
    .A2(_2800_),
    .Y(_1451_),
    .B1(_0948_));
 sg13g2_nor2_1 _5261_ (.A(_1451_),
    .B(_1317_),
    .Y(_1452_));
 sg13g2_nand2_1 _5262_ (.Y(_1453_),
    .A(_1450_),
    .B(_1452_));
 sg13g2_nand3_1 _5263_ (.B(_1453_),
    .C(net73),
    .A(_1449_),
    .Y(_1454_));
 sg13g2_a221oi_1 _5264_ (.B2(_2685_),
    .C1(_2692_),
    .B1(_0302_),
    .A1(net99),
    .Y(_1455_),
    .A2(_0616_));
 sg13g2_nor2_1 _5265_ (.A(net163),
    .B(_1455_),
    .Y(_1456_));
 sg13g2_nand2_1 _5266_ (.Y(_1458_),
    .A(_1454_),
    .B(_1456_));
 sg13g2_nand3_1 _5267_ (.B(_1458_),
    .C(net196),
    .A(_1440_),
    .Y(_1459_));
 sg13g2_nand2_1 _5268_ (.Y(_0017_),
    .A(_1406_),
    .B(_1459_));
 sg13g2_nand3_1 _5269_ (.B(_2415_),
    .C(_2405_),
    .A(_2765_),
    .Y(_1460_));
 sg13g2_nand3_1 _5270_ (.B(net100),
    .C(_2382_),
    .A(_0648_),
    .Y(_1461_));
 sg13g2_nand2_1 _5271_ (.Y(_1462_),
    .A(_1460_),
    .B(_1461_));
 sg13g2_inv_1 _5272_ (.Y(_1463_),
    .A(_2765_));
 sg13g2_nand2_1 _5273_ (.Y(_1464_),
    .A(_1463_),
    .B(_2505_));
 sg13g2_nand2_1 _5274_ (.Y(_1465_),
    .A(_1464_),
    .B(_1071_));
 sg13g2_nor2b_1 _5275_ (.A(_1462_),
    .B_N(_1465_),
    .Y(_1466_));
 sg13g2_nand2b_1 _5276_ (.Y(_1468_),
    .B(_2911_),
    .A_N(_0346_));
 sg13g2_nand2_1 _5277_ (.Y(_1469_),
    .A(_1468_),
    .B(net42));
 sg13g2_nand2_1 _5278_ (.Y(_1470_),
    .A(_1466_),
    .B(_1469_));
 sg13g2_nand2_1 _5279_ (.Y(_1471_),
    .A(_1470_),
    .B(net131));
 sg13g2_nand2_1 _5280_ (.Y(_1472_),
    .A(_0808_),
    .B(_2629_));
 sg13g2_nand3_1 _5281_ (.B(net72),
    .C(net148),
    .A(_1197_),
    .Y(_1473_));
 sg13g2_a22oi_1 _5282_ (.Y(_1474_),
    .B1(_1229_),
    .B2(_1473_),
    .A2(_1472_),
    .A1(_0917_));
 sg13g2_nand2_1 _5283_ (.Y(_1475_),
    .A(_1471_),
    .B(_1474_));
 sg13g2_nand2_1 _5284_ (.Y(_1476_),
    .A(_1475_),
    .B(net68));
 sg13g2_a21oi_1 _5285_ (.A1(_0439_),
    .A2(net106),
    .Y(_1477_),
    .B1(net54));
 sg13g2_a21oi_1 _5286_ (.A1(_2879_),
    .A2(_0995_),
    .Y(_1479_),
    .B1(net138));
 sg13g2_nand2_1 _5287_ (.Y(_1480_),
    .A(_3018_),
    .B(_2793_));
 sg13g2_a21oi_1 _5288_ (.A1(_1480_),
    .A2(_1880_),
    .Y(_1481_),
    .B1(_0651_));
 sg13g2_nor3_1 _5289_ (.A(_1477_),
    .B(_1479_),
    .C(_1481_),
    .Y(_1482_));
 sg13g2_nor2_1 _5290_ (.A(net118),
    .B(_1482_),
    .Y(_1483_));
 sg13g2_nand2_1 _5291_ (.Y(_1484_),
    .A(_1480_),
    .B(_1277_));
 sg13g2_a21oi_1 _5292_ (.A1(_1484_),
    .A2(net32),
    .Y(_1485_),
    .B1(_2462_));
 sg13g2_nand2_1 _5293_ (.Y(_1486_),
    .A(_0990_),
    .B(net30));
 sg13g2_nand2_1 _5294_ (.Y(_1487_),
    .A(_1486_),
    .B(_2807_));
 sg13g2_nand2_1 _5295_ (.Y(_1488_),
    .A(_1487_),
    .B(net70));
 sg13g2_a21oi_1 _5296_ (.A1(_1485_),
    .A2(_1488_),
    .Y(_1490_),
    .B1(net63));
 sg13g2_nor2_1 _5297_ (.A(_1483_),
    .B(_1490_),
    .Y(_1491_));
 sg13g2_nand2_1 _5298_ (.Y(_1492_),
    .A(_1476_),
    .B(_1491_));
 sg13g2_nand2_1 _5299_ (.Y(_1493_),
    .A(_1492_),
    .B(net132));
 sg13g2_o21ai_1 _5300_ (.B1(_2552_),
    .Y(_1494_),
    .A1(_2965_),
    .A2(_0621_));
 sg13g2_nand2_1 _5301_ (.Y(_1495_),
    .A(_0239_),
    .B(_0453_));
 sg13g2_nand2_1 _5302_ (.Y(_1496_),
    .A(_0940_),
    .B(_0283_));
 sg13g2_nand3_1 _5303_ (.B(_1496_),
    .C(_2517_),
    .A(_1495_),
    .Y(_1497_));
 sg13g2_o21ai_1 _5304_ (.B1(_1497_),
    .Y(_1498_),
    .A1(_1050_),
    .A2(_1494_));
 sg13g2_nand2_1 _5305_ (.Y(_1499_),
    .A(_1498_),
    .B(_2957_));
 sg13g2_nor2_1 _5306_ (.A(_3022_),
    .B(_2430_),
    .Y(_1501_));
 sg13g2_nand3_1 _5307_ (.B(net55),
    .C(net146),
    .A(_2444_),
    .Y(_1502_));
 sg13g2_nand3b_1 _5308_ (.B(_1502_),
    .C(_1054_),
    .Y(_1503_),
    .A_N(_1501_));
 sg13g2_a22oi_1 _5309_ (.Y(_1504_),
    .B1(net115),
    .B2(_1503_),
    .A2(_0949_),
    .A1(_2967_));
 sg13g2_nand2_1 _5310_ (.Y(_1505_),
    .A(_1499_),
    .B(_1504_));
 sg13g2_a21oi_1 _5311_ (.A1(_2879_),
    .A2(_2970_),
    .Y(_1506_),
    .B1(net31));
 sg13g2_nand3_1 _5312_ (.B(net200),
    .C(_2691_),
    .A(_1506_),
    .Y(_1507_));
 sg13g2_nand2_1 _5313_ (.Y(_1508_),
    .A(_1507_),
    .B(net196));
 sg13g2_a21oi_1 _5314_ (.A1(_1505_),
    .A2(net112),
    .Y(_1509_),
    .B1(_1508_));
 sg13g2_a21oi_1 _5315_ (.A1(_0542_),
    .A2(_2590_),
    .Y(_1510_),
    .B1(net61));
 sg13g2_nor2_1 _5316_ (.A(_2173_),
    .B(_2550_),
    .Y(_1512_));
 sg13g2_a21oi_1 _5317_ (.A1(_0405_),
    .A2(_1512_),
    .Y(_1513_),
    .B1(_1707_));
 sg13g2_nor2_1 _5318_ (.A(net92),
    .B(_0139_),
    .Y(_1514_));
 sg13g2_nor2_1 _5319_ (.A(net89),
    .B(_1514_),
    .Y(_1515_));
 sg13g2_nand2_1 _5320_ (.Y(_1516_),
    .A(_1515_),
    .B(_0277_));
 sg13g2_nand2_1 _5321_ (.Y(_1517_),
    .A(_1513_),
    .B(_1516_));
 sg13g2_a21oi_1 _5322_ (.A1(_0971_),
    .A2(_0404_),
    .Y(_1518_),
    .B1(net167));
 sg13g2_nand3b_1 _5323_ (.B(_1517_),
    .C(_1518_),
    .Y(_1519_),
    .A_N(_1510_));
 sg13g2_nor3_1 _5324_ (.A(net96),
    .B(_2774_),
    .C(_2436_),
    .Y(_1520_));
 sg13g2_nand2_1 _5325_ (.Y(_1521_),
    .A(_0610_),
    .B(_2405_));
 sg13g2_nand3_1 _5326_ (.B(net65),
    .C(net98),
    .A(net122),
    .Y(_1523_));
 sg13g2_nand2_1 _5327_ (.Y(_1524_),
    .A(_1521_),
    .B(_1523_));
 sg13g2_nor2_1 _5328_ (.A(net189),
    .B(_2440_),
    .Y(_1525_));
 sg13g2_a21o_1 _5329_ (.A2(_0360_),
    .A1(_1525_),
    .B1(net161),
    .X(_1526_));
 sg13g2_nor3_1 _5330_ (.A(_1520_),
    .B(_1524_),
    .C(_1526_),
    .Y(_1527_));
 sg13g2_nand2b_1 _5331_ (.Y(_1528_),
    .B(_3025_),
    .A_N(_1057_));
 sg13g2_nand2_1 _5332_ (.Y(_1529_),
    .A(_1528_),
    .B(_2569_));
 sg13g2_nand2_1 _5333_ (.Y(_1530_),
    .A(_1527_),
    .B(_1529_));
 sg13g2_a21oi_1 _5334_ (.A1(_1519_),
    .A2(_1530_),
    .Y(_1531_),
    .B1(_2736_));
 sg13g2_nand3_1 _5335_ (.B(net82),
    .C(net109),
    .A(_0197_),
    .Y(_1532_));
 sg13g2_a21oi_1 _5336_ (.A1(_1532_),
    .A2(_0239_),
    .Y(_1534_),
    .B1(_0868_));
 sg13g2_nor3_1 _5337_ (.A(net209),
    .B(_0651_),
    .C(_2986_),
    .Y(_1535_));
 sg13g2_nand2_1 _5338_ (.Y(_1536_),
    .A(_0439_),
    .B(net71));
 sg13g2_nor2_1 _5339_ (.A(_1998_),
    .B(_0482_),
    .Y(_1537_));
 sg13g2_nand2_1 _5340_ (.Y(_1538_),
    .A(_1536_),
    .B(_1537_));
 sg13g2_nand2_1 _5341_ (.Y(_1539_),
    .A(_1538_),
    .B(net197));
 sg13g2_a21oi_1 _5342_ (.A1(_1535_),
    .A2(_0838_),
    .Y(_1540_),
    .B1(_1539_));
 sg13g2_nand2b_1 _5343_ (.Y(_1541_),
    .B(_1540_),
    .A_N(_1534_));
 sg13g2_nand2_1 _5344_ (.Y(_1542_),
    .A(_1536_),
    .B(_2482_));
 sg13g2_o21ai_1 _5345_ (.B1(_1542_),
    .Y(_1543_),
    .A1(net41),
    .A2(_2659_));
 sg13g2_nand2_1 _5346_ (.Y(_1545_),
    .A(_1543_),
    .B(net105));
 sg13g2_nor2b_1 _5347_ (.A(_1541_),
    .B_N(_1545_),
    .Y(_1546_));
 sg13g2_a21o_1 _5348_ (.A2(_0140_),
    .A1(_2394_),
    .B1(_2774_),
    .X(_1547_));
 sg13g2_nand2_1 _5349_ (.Y(_1548_),
    .A(_2671_),
    .B(_2449_));
 sg13g2_nand2_1 _5350_ (.Y(_1549_),
    .A(_1548_),
    .B(_2505_));
 sg13g2_nand2_1 _5351_ (.Y(_1550_),
    .A(_1549_),
    .B(_1197_));
 sg13g2_nand2_1 _5352_ (.Y(_1551_),
    .A(_1550_),
    .B(net129));
 sg13g2_o21ai_1 _5353_ (.B1(_1347_),
    .Y(_1552_),
    .A1(net29),
    .A2(_0148_));
 sg13g2_nand3_1 _5354_ (.B(_1551_),
    .C(_1552_),
    .A(_1547_),
    .Y(_1553_));
 sg13g2_nand2_1 _5355_ (.Y(_1554_),
    .A(_1553_),
    .B(net121));
 sg13g2_nand2_1 _5356_ (.Y(_1556_),
    .A(_1546_),
    .B(_1554_));
 sg13g2_nand2_1 _5357_ (.Y(_1557_),
    .A(_1556_),
    .B(net163));
 sg13g2_nor2_1 _5358_ (.A(_1531_),
    .B(_1557_),
    .Y(_1558_));
 sg13g2_nand2_1 _5359_ (.Y(_1559_),
    .A(_0197_),
    .B(net58));
 sg13g2_nand2_1 _5360_ (.Y(_1560_),
    .A(_0504_),
    .B(_1559_));
 sg13g2_nor2_1 _5361_ (.A(_1269_),
    .B(_1283_),
    .Y(_1561_));
 sg13g2_a21oi_1 _5362_ (.A1(_1560_),
    .A2(_2615_),
    .Y(_1562_),
    .B1(_1561_));
 sg13g2_inv_1 _5363_ (.Y(_1563_),
    .A(_0278_));
 sg13g2_nor2_1 _5364_ (.A(net91),
    .B(_1563_),
    .Y(_1564_));
 sg13g2_a21oi_1 _5365_ (.A1(_2613_),
    .A2(net77),
    .Y(_1565_),
    .B1(net124));
 sg13g2_nand2_1 _5366_ (.Y(_1567_),
    .A(_1564_),
    .B(_1565_));
 sg13g2_nand2_1 _5367_ (.Y(_1568_),
    .A(_1562_),
    .B(_1567_));
 sg13g2_nand2_1 _5368_ (.Y(_1569_),
    .A(_1568_),
    .B(net131));
 sg13g2_inv_1 _5369_ (.Y(_1570_),
    .A(_2931_));
 sg13g2_nand2_1 _5370_ (.Y(_1571_),
    .A(_2937_),
    .B(_2415_));
 sg13g2_nand2_1 _5371_ (.Y(_1572_),
    .A(_1570_),
    .B(_1571_));
 sg13g2_nand2_1 _5372_ (.Y(_1573_),
    .A(_1572_),
    .B(net88));
 sg13g2_a21oi_1 _5373_ (.A1(_2628_),
    .A2(_3014_),
    .Y(_1574_),
    .B1(_0477_));
 sg13g2_nand2b_1 _5374_ (.Y(_1575_),
    .B(net39),
    .A_N(_1574_));
 sg13g2_nand2_1 _5375_ (.Y(_1576_),
    .A(_1573_),
    .B(_1575_));
 sg13g2_nand2_1 _5376_ (.Y(_1578_),
    .A(_1576_),
    .B(net116));
 sg13g2_nor4_1 _5377_ (.A(_2418_),
    .B(_0118_),
    .C(_0142_),
    .D(_3013_),
    .Y(_1579_));
 sg13g2_inv_1 _5378_ (.Y(_1580_),
    .A(_0628_));
 sg13g2_nand2_1 _5379_ (.Y(_1581_),
    .A(_0247_),
    .B(_2444_));
 sg13g2_nand2_1 _5380_ (.Y(_1582_),
    .A(net85),
    .B(net125));
 sg13g2_a21oi_1 _5381_ (.A1(_3030_),
    .A2(_1582_),
    .Y(_1583_),
    .B1(_0338_));
 sg13g2_a22oi_1 _5382_ (.Y(_1584_),
    .B1(_1581_),
    .B2(_1583_),
    .A2(_1580_),
    .A1(_1579_));
 sg13g2_nand3_1 _5383_ (.B(_1578_),
    .C(_1584_),
    .A(_1569_),
    .Y(_1585_));
 sg13g2_nand2_1 _5384_ (.Y(_1586_),
    .A(_1585_),
    .B(net112));
 sg13g2_nand2_1 _5385_ (.Y(_1587_),
    .A(_0225_),
    .B(_2853_));
 sg13g2_inv_1 _5386_ (.Y(_1589_),
    .A(_1587_));
 sg13g2_a21oi_1 _5387_ (.A1(_1589_),
    .A2(_2982_),
    .Y(_1590_),
    .B1(_2732_));
 sg13g2_nand2_1 _5388_ (.Y(_1591_),
    .A(_1532_),
    .B(_0977_));
 sg13g2_nand2_1 _5389_ (.Y(_1592_),
    .A(_1591_),
    .B(_0110_));
 sg13g2_nand2_1 _5390_ (.Y(_1593_),
    .A(_1590_),
    .B(_1592_));
 sg13g2_nor2_1 _5391_ (.A(net171),
    .B(_3028_),
    .Y(_1594_));
 sg13g2_nor2_1 _5392_ (.A(_2958_),
    .B(_2742_),
    .Y(_1595_));
 sg13g2_a22oi_1 _5393_ (.Y(_1596_),
    .B1(_1594_),
    .B2(_1595_),
    .A2(_2388_),
    .A1(_0708_));
 sg13g2_nand2_1 _5394_ (.Y(_1597_),
    .A(_1593_),
    .B(_1596_));
 sg13g2_nand2_1 _5395_ (.Y(_1598_),
    .A(_1597_),
    .B(_2665_));
 sg13g2_nand2_1 _5396_ (.Y(_1600_),
    .A(_0921_),
    .B(_2221_));
 sg13g2_nand2_1 _5397_ (.Y(_1601_),
    .A(_1600_),
    .B(net69));
 sg13g2_nand2_1 _5398_ (.Y(_1602_),
    .A(_1601_),
    .B(_1078_));
 sg13g2_a21oi_1 _5399_ (.A1(_0370_),
    .A2(net65),
    .Y(_1603_),
    .B1(_1602_));
 sg13g2_nor2_1 _5400_ (.A(_2597_),
    .B(_1603_),
    .Y(_1604_));
 sg13g2_a21oi_1 _5401_ (.A1(_1598_),
    .A2(_1604_),
    .Y(_1605_),
    .B1(_2609_));
 sg13g2_nand2_1 _5402_ (.Y(_1606_),
    .A(_1586_),
    .B(_1605_));
 sg13g2_nor2_1 _5403_ (.A(_1558_),
    .B(_1606_),
    .Y(_1607_));
 sg13g2_a21oi_1 _5404_ (.A1(_1493_),
    .A2(_1509_),
    .Y(_0018_),
    .B1(_1607_));
 sg13g2_nand3_1 _5405_ (.B(net120),
    .C(_0618_),
    .A(_0934_),
    .Y(_1608_));
 sg13g2_nand2_1 _5406_ (.Y(_1610_),
    .A(_2453_),
    .B(net45));
 sg13g2_nand3_1 _5407_ (.B(net130),
    .C(_1610_),
    .A(_1608_),
    .Y(_1611_));
 sg13g2_o21ai_1 _5408_ (.B1(net46),
    .Y(_1612_),
    .A1(_0127_),
    .A2(_0603_));
 sg13g2_nand2_1 _5409_ (.Y(_1613_),
    .A(_1611_),
    .B(_1612_));
 sg13g2_nor2_1 _5410_ (.A(net48),
    .B(_0168_),
    .Y(_1614_));
 sg13g2_nand2_1 _5411_ (.Y(_1615_),
    .A(_1614_),
    .B(net67));
 sg13g2_nand3_1 _5412_ (.B(_2141_),
    .C(_0478_),
    .A(_1615_),
    .Y(_1616_));
 sg13g2_nand2_1 _5413_ (.Y(_1617_),
    .A(_2861_),
    .B(_0128_));
 sg13g2_o21ai_1 _5414_ (.B1(net105),
    .Y(_1618_),
    .A1(_0219_),
    .A2(_1617_));
 sg13g2_nand3_1 _5415_ (.B(_1618_),
    .C(_2360_),
    .A(_1616_),
    .Y(_1619_));
 sg13g2_a21oi_1 _5416_ (.A1(_1613_),
    .A2(net117),
    .Y(_1621_),
    .B1(_1619_));
 sg13g2_nand3_1 _5417_ (.B(_0673_),
    .C(net168),
    .A(_0863_),
    .Y(_1622_));
 sg13g2_a21oi_1 _5418_ (.A1(_0681_),
    .A2(_1167_),
    .Y(_1623_),
    .B1(net123));
 sg13g2_nand2_1 _5419_ (.Y(_1624_),
    .A(_1622_),
    .B(_1623_));
 sg13g2_o21ai_1 _5420_ (.B1(net105),
    .Y(_1625_),
    .A1(_2892_),
    .A2(_0134_));
 sg13g2_o21ai_1 _5421_ (.B1(_2936_),
    .Y(_1626_),
    .A1(_2701_),
    .A2(net71));
 sg13g2_nand3_1 _5422_ (.B(_1625_),
    .C(_1626_),
    .A(_1624_),
    .Y(_1627_));
 sg13g2_o21ai_1 _5423_ (.B1(net163),
    .Y(_1628_),
    .A1(net73),
    .A2(_1627_));
 sg13g2_nor2_1 _5424_ (.A(_1621_),
    .B(_1628_),
    .Y(_1629_));
 sg13g2_o21ai_1 _5425_ (.B1(_0454_),
    .Y(_1630_),
    .A1(net72),
    .A2(_0681_));
 sg13g2_a21oi_1 _5426_ (.A1(_1563_),
    .A2(net74),
    .Y(_1632_),
    .B1(net127));
 sg13g2_a221oi_1 _5427_ (.B2(_2635_),
    .C1(net167),
    .B1(net74),
    .A1(_2998_),
    .Y(_1633_),
    .A2(net55));
 sg13g2_a21oi_1 _5428_ (.A1(_1630_),
    .A2(_1632_),
    .Y(_1634_),
    .B1(_1633_));
 sg13g2_nand2b_1 _5429_ (.Y(_1635_),
    .B(net112),
    .A_N(_1634_));
 sg13g2_nor2_1 _5430_ (.A(_2701_),
    .B(_1204_),
    .Y(_1636_));
 sg13g2_a21oi_1 _5431_ (.A1(_2727_),
    .A2(_2757_),
    .Y(_1637_),
    .B1(net36));
 sg13g2_o21ai_1 _5432_ (.B1(net115),
    .Y(_1638_),
    .A1(_1636_),
    .A2(_1637_));
 sg13g2_nand2_1 _5433_ (.Y(_1639_),
    .A(_1638_),
    .B(_2598_));
 sg13g2_nand3_1 _5434_ (.B(_2610_),
    .C(_1639_),
    .A(_1635_),
    .Y(_1640_));
 sg13g2_nor2_1 _5435_ (.A(_1629_),
    .B(_1640_),
    .Y(_1641_));
 sg13g2_a21oi_1 _5436_ (.A1(_1006_),
    .A2(_2861_),
    .Y(_1643_),
    .B1(net55));
 sg13g2_a21oi_1 _5437_ (.A1(net24),
    .A2(_0599_),
    .Y(_1644_),
    .B1(_1643_));
 sg13g2_nor2_1 _5438_ (.A(net114),
    .B(_0219_),
    .Y(_1645_));
 sg13g2_o21ai_1 _5439_ (.B1(net171),
    .Y(_1646_),
    .A1(_2687_),
    .A2(_0616_));
 sg13g2_a21oi_1 _5440_ (.A1(_1645_),
    .A2(_0934_),
    .Y(_1647_),
    .B1(_1646_));
 sg13g2_nand2_1 _5441_ (.Y(_1648_),
    .A(_1253_),
    .B(net193));
 sg13g2_a21oi_1 _5442_ (.A1(_1648_),
    .A2(net49),
    .Y(_1649_),
    .B1(net203));
 sg13g2_o21ai_1 _5443_ (.B1(_1649_),
    .Y(_1650_),
    .A1(net40),
    .A2(_0628_));
 sg13g2_nor2_1 _5444_ (.A(_1647_),
    .B(_1650_),
    .Y(_1651_));
 sg13g2_a21oi_1 _5445_ (.A1(_1644_),
    .A2(net113),
    .Y(_1652_),
    .B1(_1651_));
 sg13g2_a21oi_1 _5446_ (.A1(_0278_),
    .A2(net24),
    .Y(_1654_),
    .B1(_0118_));
 sg13g2_nand2_1 _5447_ (.Y(_1655_),
    .A(_1580_),
    .B(_0721_));
 sg13g2_a21oi_1 _5448_ (.A1(_1654_),
    .A2(_1655_),
    .Y(_1656_),
    .B1(_0729_));
 sg13g2_a21oi_1 _5449_ (.A1(_1652_),
    .A2(_1656_),
    .Y(_1657_),
    .B1(_2609_));
 sg13g2_nand3_1 _5450_ (.B(_0706_),
    .C(net172),
    .A(_0654_),
    .Y(_1658_));
 sg13g2_a21oi_1 _5451_ (.A1(_0610_),
    .A2(_1167_),
    .Y(_1659_),
    .B1(net123));
 sg13g2_o21ai_1 _5452_ (.B1(net129),
    .Y(_1660_),
    .A1(net194),
    .A2(_0682_));
 sg13g2_nor2_1 _5453_ (.A(_0824_),
    .B(_0611_),
    .Y(_1661_));
 sg13g2_nand2_1 _5454_ (.Y(_1662_),
    .A(_1660_),
    .B(_1661_));
 sg13g2_a22oi_1 _5455_ (.Y(_1663_),
    .B1(net116),
    .B2(_1662_),
    .A2(_1659_),
    .A1(_1658_));
 sg13g2_nand2_1 _5456_ (.Y(_1665_),
    .A(_1663_),
    .B(net147));
 sg13g2_nor3_1 _5457_ (.A(net28),
    .B(_0720_),
    .C(_2723_),
    .Y(_1666_));
 sg13g2_nor2_1 _5458_ (.A(net40),
    .B(_1614_),
    .Y(_1667_));
 sg13g2_nor4_1 _5459_ (.A(net175),
    .B(_0033_),
    .C(_1666_),
    .D(_1667_),
    .Y(_1668_));
 sg13g2_a21oi_1 _5460_ (.A1(_0628_),
    .A2(net37),
    .Y(_1669_),
    .B1(net107));
 sg13g2_o21ai_1 _5461_ (.B1(_1669_),
    .Y(_1670_),
    .A1(net24),
    .A2(_0347_));
 sg13g2_a21oi_1 _5462_ (.A1(_1668_),
    .A2(_1670_),
    .Y(_1671_),
    .B1(_2423_));
 sg13g2_nand2_1 _5463_ (.Y(_1672_),
    .A(_1665_),
    .B(_1671_));
 sg13g2_nand2_1 _5464_ (.Y(_1673_),
    .A(_1657_),
    .B(_1672_));
 sg13g2_nor2_1 _5465_ (.A(net142),
    .B(_2772_),
    .Y(_1674_));
 sg13g2_a22oi_1 _5466_ (.Y(_1676_),
    .B1(_0622_),
    .B2(_1674_),
    .A2(_2686_),
    .A1(_1253_));
 sg13g2_nor2b_1 _5467_ (.A(_1676_),
    .B_N(_1296_),
    .Y(_1677_));
 sg13g2_nand2_1 _5468_ (.Y(_1678_),
    .A(_2710_),
    .B(_2686_));
 sg13g2_a21oi_1 _5469_ (.A1(_1669_),
    .A2(_1678_),
    .Y(_1679_),
    .B1(net131));
 sg13g2_nor3_1 _5470_ (.A(net72),
    .B(_3029_),
    .C(_1563_),
    .Y(_1680_));
 sg13g2_o21ai_1 _5471_ (.B1(net115),
    .Y(_1681_),
    .A1(_0663_),
    .A2(_1680_));
 sg13g2_o21ai_1 _5472_ (.B1(_1681_),
    .Y(_1682_),
    .A1(_1677_),
    .A2(_1679_));
 sg13g2_nand2_1 _5473_ (.Y(_1683_),
    .A(_1682_),
    .B(_2598_));
 sg13g2_nor2b_1 _5474_ (.A(_1673_),
    .B_N(_1683_),
    .Y(_1684_));
 sg13g2_nor2_1 _5475_ (.A(_1641_),
    .B(_1684_),
    .Y(_0019_));
 sg13g2_inv_1 _5476_ (.Y(_1686_),
    .A(_2715_));
 sg13g2_nor2_1 _5477_ (.A(_1686_),
    .B(_2880_),
    .Y(_1687_));
 sg13g2_nand3b_1 _5478_ (.B(net172),
    .C(_0662_),
    .Y(_1688_),
    .A_N(_1141_));
 sg13g2_nand3_1 _5479_ (.B(net59),
    .C(_1167_),
    .A(_2548_),
    .Y(_1689_));
 sg13g2_o21ai_1 _5480_ (.B1(_1689_),
    .Y(_1690_),
    .A1(_1687_),
    .A2(_1688_));
 sg13g2_nand2_1 _5481_ (.Y(_1691_),
    .A(_1690_),
    .B(net117));
 sg13g2_a21oi_1 _5482_ (.A1(net90),
    .A2(_2969_),
    .Y(_1692_),
    .B1(_1039_));
 sg13g2_a21oi_1 _5483_ (.A1(_0816_),
    .A2(_0744_),
    .Y(_1693_),
    .B1(net66));
 sg13g2_nor2b_1 _5484_ (.A(_1692_),
    .B_N(_1693_),
    .Y(_1694_));
 sg13g2_nor3_1 _5485_ (.A(net72),
    .B(_2550_),
    .C(_0797_),
    .Y(_1695_));
 sg13g2_nand2_1 _5486_ (.Y(_1697_),
    .A(_0744_),
    .B(_0629_));
 sg13g2_nor3_1 _5487_ (.A(_2510_),
    .B(_2520_),
    .C(_1697_),
    .Y(_1698_));
 sg13g2_nor3_1 _5488_ (.A(net35),
    .B(_1695_),
    .C(_1698_),
    .Y(_1699_));
 sg13g2_nor2_1 _5489_ (.A(_1694_),
    .B(_1699_),
    .Y(_1700_));
 sg13g2_nand3_1 _5490_ (.B(_1700_),
    .C(_0090_),
    .A(_1691_),
    .Y(_1701_));
 sg13g2_nor2b_1 _5491_ (.A(_2848_),
    .B_N(_1184_),
    .Y(_1702_));
 sg13g2_o21ai_1 _5492_ (.B1(_1542_),
    .Y(_1703_),
    .A1(net41),
    .A2(_1702_));
 sg13g2_nand2_1 _5493_ (.Y(_1704_),
    .A(_1703_),
    .B(net130));
 sg13g2_a21oi_1 _5494_ (.A1(_2273_),
    .A2(_0360_),
    .Y(_1705_),
    .B1(_1012_));
 sg13g2_nand2_1 _5495_ (.Y(_1706_),
    .A(_1704_),
    .B(_1705_));
 sg13g2_nand2_1 _5496_ (.Y(_1708_),
    .A(_1706_),
    .B(net83));
 sg13g2_nor2_1 _5497_ (.A(net72),
    .B(_1869_),
    .Y(_1709_));
 sg13g2_nor2_1 _5498_ (.A(_2510_),
    .B(_1036_),
    .Y(_1710_));
 sg13g2_a22oi_1 _5499_ (.Y(_1711_),
    .B1(_2879_),
    .B2(_1710_),
    .A2(_1709_),
    .A1(_0093_));
 sg13g2_nor3_1 _5500_ (.A(_2418_),
    .B(net189),
    .C(_3013_),
    .Y(_1712_));
 sg13g2_nor2_1 _5501_ (.A(_1501_),
    .B(_1712_),
    .Y(_1713_));
 sg13g2_nand3_1 _5502_ (.B(_2554_),
    .C(_0422_),
    .A(_0168_),
    .Y(_1714_));
 sg13g2_a21oi_1 _5503_ (.A1(_1713_),
    .A2(_1714_),
    .Y(_1715_),
    .B1(_0483_));
 sg13g2_a21oi_1 _5504_ (.A1(_1711_),
    .A2(net22),
    .Y(_1716_),
    .B1(_1715_));
 sg13g2_nand3_1 _5505_ (.B(_1716_),
    .C(net164),
    .A(_1708_),
    .Y(_1717_));
 sg13g2_nand3_1 _5506_ (.B(_1717_),
    .C(_2566_),
    .A(_1701_),
    .Y(_1719_));
 sg13g2_nor2_1 _5507_ (.A(net28),
    .B(_2793_),
    .Y(_1720_));
 sg13g2_nand2_1 _5508_ (.Y(_1721_),
    .A(_0422_),
    .B(_2808_));
 sg13g2_nand3_1 _5509_ (.B(net189),
    .C(_0530_),
    .A(net76),
    .Y(_1722_));
 sg13g2_a21oi_1 _5510_ (.A1(_1721_),
    .A2(_1722_),
    .Y(_1723_),
    .B1(_2600_));
 sg13g2_a21oi_1 _5511_ (.A1(_1160_),
    .A2(_3003_),
    .Y(_1724_),
    .B1(net138));
 sg13g2_nor4_1 _5512_ (.A(_1561_),
    .B(_1720_),
    .C(_1723_),
    .D(_1724_),
    .Y(_1725_));
 sg13g2_nand2_1 _5513_ (.Y(_1726_),
    .A(_1725_),
    .B(_2957_));
 sg13g2_inv_1 _5514_ (.Y(_1727_),
    .A(_1104_));
 sg13g2_o21ai_1 _5515_ (.B1(net54),
    .Y(_1728_),
    .A1(net98),
    .A2(_0942_));
 sg13g2_o21ai_1 _5516_ (.B1(_1728_),
    .Y(_1730_),
    .A1(_1727_),
    .A2(_2931_));
 sg13g2_o21ai_1 _5517_ (.B1(_2593_),
    .Y(_1731_),
    .A1(_0148_),
    .A2(_2574_));
 sg13g2_nor2_1 _5518_ (.A(_2494_),
    .B(_2407_),
    .Y(_1732_));
 sg13g2_a21oi_1 _5519_ (.A1(_1732_),
    .A2(net85),
    .Y(_1733_),
    .B1(_2619_));
 sg13g2_nand3_1 _5520_ (.B(_1731_),
    .C(_1733_),
    .A(_1730_),
    .Y(_1734_));
 sg13g2_nand3_1 _5521_ (.B(_0728_),
    .C(_1734_),
    .A(_1726_),
    .Y(_1735_));
 sg13g2_a21oi_1 _5522_ (.A1(_1109_),
    .A2(net65),
    .Y(_1736_),
    .B1(_1077_));
 sg13g2_o21ai_1 _5523_ (.B1(net69),
    .Y(_1737_),
    .A1(_2969_),
    .A2(_3029_));
 sg13g2_nand2_1 _5524_ (.Y(_1738_),
    .A(_1736_),
    .B(_1737_));
 sg13g2_nand2_1 _5525_ (.Y(_1739_),
    .A(_1738_),
    .B(_2559_));
 sg13g2_nand2_1 _5526_ (.Y(_1741_),
    .A(net29),
    .B(net37));
 sg13g2_o21ai_1 _5527_ (.B1(_1741_),
    .Y(_1742_),
    .A1(_2687_),
    .A2(_2906_));
 sg13g2_nor2_1 _5528_ (.A(net175),
    .B(net35),
    .Y(_1743_));
 sg13g2_nand2_1 _5529_ (.Y(_1744_),
    .A(_1742_),
    .B(_1743_));
 sg13g2_nor2_1 _5530_ (.A(_2923_),
    .B(_3029_),
    .Y(_1745_));
 sg13g2_nor3_1 _5531_ (.A(net168),
    .B(_2374_),
    .C(_1745_),
    .Y(_1746_));
 sg13g2_o21ai_1 _5532_ (.B1(_1746_),
    .Y(_1747_),
    .A1(_2642_),
    .A2(_0859_));
 sg13g2_nand3_1 _5533_ (.B(_1744_),
    .C(_1747_),
    .A(_1739_),
    .Y(_1748_));
 sg13g2_nand2_1 _5534_ (.Y(_1749_),
    .A(_1748_),
    .B(net200));
 sg13g2_nand2_1 _5535_ (.Y(_1750_),
    .A(_1735_),
    .B(_1749_));
 sg13g2_nor2_1 _5536_ (.A(_2610_),
    .B(_1750_),
    .Y(_1752_));
 sg13g2_nor2_1 _5537_ (.A(net155),
    .B(_2501_),
    .Y(_1753_));
 sg13g2_o21ai_1 _5538_ (.B1(_1054_),
    .Y(_1754_),
    .A1(_0795_),
    .A2(_0340_));
 sg13g2_a22oi_1 _5539_ (.Y(_1755_),
    .B1(net115),
    .B2(_1754_),
    .A2(_0949_),
    .A1(_1753_));
 sg13g2_nand3_1 _5540_ (.B(_1308_),
    .C(_0453_),
    .A(_2823_),
    .Y(_1756_));
 sg13g2_a21oi_1 _5541_ (.A1(_2239_),
    .A2(_2715_),
    .Y(_1757_),
    .B1(net124));
 sg13g2_nand2_1 _5542_ (.Y(_1758_),
    .A(_1756_),
    .B(_1757_));
 sg13g2_nand2_1 _5543_ (.Y(_1759_),
    .A(_1758_),
    .B(_1494_));
 sg13g2_nand2_1 _5544_ (.Y(_1760_),
    .A(_1759_),
    .B(net131));
 sg13g2_nand2_1 _5545_ (.Y(_1761_),
    .A(_1755_),
    .B(_1760_));
 sg13g2_nand2_1 _5546_ (.Y(_1763_),
    .A(_1761_),
    .B(net112));
 sg13g2_nor2b_1 _5547_ (.A(_1637_),
    .B_N(_0478_),
    .Y(_1764_));
 sg13g2_o21ai_1 _5548_ (.B1(_1764_),
    .Y(_1765_),
    .A1(net99),
    .A2(_0803_));
 sg13g2_a21oi_1 _5549_ (.A1(_1765_),
    .A2(_0959_),
    .Y(_1766_),
    .B1(net195));
 sg13g2_nand2_1 _5550_ (.Y(_1767_),
    .A(_1763_),
    .B(_1766_));
 sg13g2_a21oi_1 _5551_ (.A1(_2803_),
    .A2(_2989_),
    .Y(_1768_),
    .B1(net61));
 sg13g2_nand2_1 _5552_ (.Y(_1769_),
    .A(_0907_),
    .B(net88));
 sg13g2_nor2b_1 _5553_ (.A(_1125_),
    .B_N(_1769_),
    .Y(_1770_));
 sg13g2_nand2b_1 _5554_ (.Y(_1771_),
    .B(_1770_),
    .A_N(_1768_));
 sg13g2_nand2_1 _5555_ (.Y(_1772_),
    .A(_3019_),
    .B(_1370_));
 sg13g2_a21oi_1 _5556_ (.A1(_1772_),
    .A2(_1167_),
    .Y(_1774_),
    .B1(net116));
 sg13g2_nor2_1 _5557_ (.A(net33),
    .B(_1444_),
    .Y(_1775_));
 sg13g2_o21ai_1 _5558_ (.B1(net42),
    .Y(_1776_),
    .A1(_1775_),
    .A2(_2880_));
 sg13g2_nand4_1 _5559_ (.B(net24),
    .C(net172),
    .A(_0168_),
    .Y(_1777_),
    .D(net194));
 sg13g2_nand3_1 _5560_ (.B(_1776_),
    .C(_1777_),
    .A(_1774_),
    .Y(_1778_));
 sg13g2_a21oi_1 _5561_ (.A1(_1771_),
    .A2(_1778_),
    .Y(_1779_),
    .B1(net73));
 sg13g2_nor2_1 _5562_ (.A(net31),
    .B(_1197_),
    .Y(_1780_));
 sg13g2_o21ai_1 _5563_ (.B1(_0915_),
    .Y(_1781_),
    .A1(_2892_),
    .A2(_0209_));
 sg13g2_nand2_1 _5564_ (.Y(_1782_),
    .A(_1781_),
    .B(net123));
 sg13g2_a21oi_1 _5565_ (.A1(_0971_),
    .A2(_2413_),
    .Y(_1783_),
    .B1(_3039_));
 sg13g2_o21ai_1 _5566_ (.B1(net39),
    .Y(_1785_),
    .A1(_0527_),
    .A2(_2900_));
 sg13g2_nand2_1 _5567_ (.Y(_1786_),
    .A(_1514_),
    .B(net134));
 sg13g2_nand3_1 _5568_ (.B(_1785_),
    .C(_1786_),
    .A(_1783_),
    .Y(_1787_));
 sg13g2_o21ai_1 _5569_ (.B1(_1787_),
    .Y(_1788_),
    .A1(_1780_),
    .A2(_1782_));
 sg13g2_nor3_1 _5570_ (.A(_2678_),
    .B(net160),
    .C(_1727_),
    .Y(_1789_));
 sg13g2_nor3_1 _5571_ (.A(_2557_),
    .B(_1789_),
    .C(_1152_),
    .Y(_1790_));
 sg13g2_nand2_1 _5572_ (.Y(_1791_),
    .A(_1788_),
    .B(_1790_));
 sg13g2_nand2_1 _5573_ (.Y(_1792_),
    .A(_1791_),
    .B(net163));
 sg13g2_nor2_1 _5574_ (.A(_1779_),
    .B(_1792_),
    .Y(_1793_));
 sg13g2_nor2_1 _5575_ (.A(_1767_),
    .B(_1793_),
    .Y(_1794_));
 sg13g2_a21oi_1 _5576_ (.A1(_1719_),
    .A2(_1752_),
    .Y(_0020_),
    .B1(_1794_));
 sg13g2_buf_1 _5577_ (.A(ui_in[0]),
    .X(_1796_));
 sg13g2_buf_2 _5578_ (.A(ui_in[3]),
    .X(_1797_));
 sg13g2_buf_1 _5579_ (.A(_1797_),
    .X(_1798_));
 sg13g2_buf_1 _5580_ (.A(ui_in[2]),
    .X(_1799_));
 sg13g2_buf_1 _5581_ (.A(ui_in[1]),
    .X(_1800_));
 sg13g2_buf_1 _5582_ (.A(_1800_),
    .X(_1801_));
 sg13g2_inv_1 _5583_ (.Y(_1802_),
    .A(net216));
 sg13g2_nor2_1 _5584_ (.A(_1799_),
    .B(_1802_),
    .Y(_1803_));
 sg13g2_nor2_1 _5585_ (.A(net217),
    .B(_1803_),
    .Y(_1804_));
 sg13g2_inv_1 _5586_ (.Y(_1806_),
    .A(net218));
 sg13g2_nand2_2 _5587_ (.Y(_1807_),
    .A(_1806_),
    .B(net216));
 sg13g2_buf_1 _5588_ (.A(_1799_),
    .X(_1808_));
 sg13g2_nand2_1 _5589_ (.Y(_1809_),
    .A(_1807_),
    .B(net215));
 sg13g2_inv_1 _5590_ (.Y(_1810_),
    .A(_1797_));
 sg13g2_nand2_1 _5591_ (.Y(_1811_),
    .A(net218),
    .B(_1800_));
 sg13g2_buf_2 _5592_ (.A(_1811_),
    .X(_1812_));
 sg13g2_inv_1 _5593_ (.Y(_1813_),
    .A(_1812_));
 sg13g2_nor2_1 _5594_ (.A(net215),
    .B(_1813_),
    .Y(_1814_));
 sg13g2_nor2_1 _5595_ (.A(net214),
    .B(_1814_),
    .Y(_1815_));
 sg13g2_a22oi_1 _5596_ (.Y(_1817_),
    .B1(_1809_),
    .B2(_1815_),
    .A2(_1804_),
    .A1(net218));
 sg13g2_buf_1 _5597_ (.A(ui_in[4]),
    .X(_1818_));
 sg13g2_nor2_1 _5598_ (.A(_1818_),
    .B(net1),
    .Y(_1819_));
 sg13g2_buf_2 _5599_ (.A(_1819_),
    .X(_1820_));
 sg13g2_inv_1 _5600_ (.Y(_1821_),
    .A(_1820_));
 sg13g2_inv_1 _5601_ (.Y(_1822_),
    .A(net1));
 sg13g2_nor2_1 _5602_ (.A(_1818_),
    .B(_1822_),
    .Y(_1823_));
 sg13g2_buf_2 _5603_ (.A(_1823_),
    .X(_1824_));
 sg13g2_nor2_2 _5604_ (.A(net216),
    .B(net215),
    .Y(_1825_));
 sg13g2_nor2_2 _5605_ (.A(net214),
    .B(_1825_),
    .Y(_1826_));
 sg13g2_inv_1 _5606_ (.Y(_1828_),
    .A(_1799_));
 sg13g2_nor2_1 _5607_ (.A(net216),
    .B(_1828_),
    .Y(_1829_));
 sg13g2_nor2_2 _5608_ (.A(_1797_),
    .B(_1829_),
    .Y(_1830_));
 sg13g2_nor2_1 _5609_ (.A(_1796_),
    .B(_1799_),
    .Y(_1831_));
 sg13g2_inv_1 _5610_ (.Y(_1832_),
    .A(_1831_));
 sg13g2_o21ai_1 _5611_ (.B1(_1832_),
    .Y(_1833_),
    .A1(_1826_),
    .A2(_1830_));
 sg13g2_inv_1 _5612_ (.Y(_1834_),
    .A(_1818_));
 sg13g2_nor2_1 _5613_ (.A(net1),
    .B(_1834_),
    .Y(_1835_));
 sg13g2_buf_2 _5614_ (.A(_1835_),
    .X(_1836_));
 sg13g2_inv_1 _5615_ (.Y(_1837_),
    .A(_1836_));
 sg13g2_nor2_1 _5616_ (.A(_1831_),
    .B(_1803_),
    .Y(_1839_));
 sg13g2_nand2_1 _5617_ (.Y(_1840_),
    .A(net218),
    .B(net215));
 sg13g2_nand2_1 _5618_ (.Y(_1841_),
    .A(_1839_),
    .B(_1840_));
 sg13g2_nor2_1 _5619_ (.A(net217),
    .B(_1841_),
    .Y(_1842_));
 sg13g2_nor3_1 _5620_ (.A(_1826_),
    .B(net192),
    .C(_1842_),
    .Y(_1843_));
 sg13g2_a21oi_1 _5621_ (.A1(_1824_),
    .A2(_1833_),
    .Y(_1844_),
    .B1(_1843_));
 sg13g2_o21ai_1 _5622_ (.B1(_1844_),
    .Y(_0000_),
    .A1(_1817_),
    .A2(_1821_));
 sg13g2_nor2_1 _5623_ (.A(net218),
    .B(_1800_),
    .Y(_1845_));
 sg13g2_buf_2 _5624_ (.A(_1845_),
    .X(_1846_));
 sg13g2_nor2_1 _5625_ (.A(_1846_),
    .B(_1813_),
    .Y(_1847_));
 sg13g2_nand2_1 _5626_ (.Y(_1849_),
    .A(_1847_),
    .B(_1832_));
 sg13g2_buf_1 _5627_ (.A(_1828_),
    .X(_1850_));
 sg13g2_nor2_1 _5628_ (.A(_1797_),
    .B(net213),
    .Y(_1851_));
 sg13g2_a21oi_1 _5629_ (.A1(_1846_),
    .A2(net214),
    .Y(_1852_),
    .B1(_1851_));
 sg13g2_inv_1 _5630_ (.Y(_1853_),
    .A(_1852_));
 sg13g2_nand2_1 _5631_ (.Y(_1854_),
    .A(_1853_),
    .B(_1812_));
 sg13g2_o21ai_1 _5632_ (.B1(_1854_),
    .Y(_1855_),
    .A1(_1810_),
    .A2(_1849_));
 sg13g2_nand2_1 _5633_ (.Y(_1856_),
    .A(_1855_),
    .B(_1836_));
 sg13g2_nand2_1 _5634_ (.Y(_1857_),
    .A(_1839_),
    .B(_1797_));
 sg13g2_nand3_1 _5635_ (.B(_1807_),
    .C(_1824_),
    .A(_1857_),
    .Y(_1858_));
 sg13g2_inv_1 _5636_ (.Y(_1860_),
    .A(_1847_));
 sg13g2_nand2_1 _5637_ (.Y(_1861_),
    .A(_1860_),
    .B(net213));
 sg13g2_inv_1 _5638_ (.Y(_1862_),
    .A(_1846_));
 sg13g2_nand2_1 _5639_ (.Y(_1863_),
    .A(_1862_),
    .B(net215));
 sg13g2_a21oi_1 _5640_ (.A1(_1862_),
    .A2(net215),
    .Y(_1864_),
    .B1(net217));
 sg13g2_a21oi_1 _5641_ (.A1(_1861_),
    .A2(_1863_),
    .Y(_1865_),
    .B1(_1864_));
 sg13g2_nand2_1 _5642_ (.Y(_1866_),
    .A(_1865_),
    .B(_1820_));
 sg13g2_nand3_1 _5643_ (.B(_1858_),
    .C(_1866_),
    .A(_1856_),
    .Y(_0007_));
 sg13g2_buf_1 _5644_ (.A(net217),
    .X(_1867_));
 sg13g2_nor2_1 _5645_ (.A(_1850_),
    .B(_1860_),
    .Y(_1868_));
 sg13g2_nor2_1 _5646_ (.A(_1798_),
    .B(_1868_),
    .Y(_1870_));
 sg13g2_nand2_1 _5647_ (.Y(_1871_),
    .A(_1807_),
    .B(_1850_));
 sg13g2_nand2_1 _5648_ (.Y(_1872_),
    .A(_1798_),
    .B(net218));
 sg13g2_inv_1 _5649_ (.Y(_1873_),
    .A(_1872_));
 sg13g2_a221oi_1 _5650_ (.B2(_1871_),
    .C1(_1873_),
    .B1(_1870_),
    .A1(_1867_),
    .Y(_1874_),
    .A2(_1825_));
 sg13g2_nor2_1 _5651_ (.A(net216),
    .B(_1806_),
    .Y(_1875_));
 sg13g2_nor2_1 _5652_ (.A(net213),
    .B(_1875_),
    .Y(_1876_));
 sg13g2_nor2_1 _5653_ (.A(_1808_),
    .B(_1807_),
    .Y(_1877_));
 sg13g2_inv_1 _5654_ (.Y(_1878_),
    .A(_1877_));
 sg13g2_nand2_1 _5655_ (.Y(_1879_),
    .A(_1878_),
    .B(net212));
 sg13g2_nor2_1 _5656_ (.A(net215),
    .B(_1806_),
    .Y(_1881_));
 sg13g2_inv_1 _5657_ (.Y(_1882_),
    .A(_1830_));
 sg13g2_o21ai_1 _5658_ (.B1(_1824_),
    .Y(_1883_),
    .A1(_1881_),
    .A2(_1882_));
 sg13g2_o21ai_1 _5659_ (.B1(_1883_),
    .Y(_1884_),
    .A1(_1821_),
    .A2(_1853_));
 sg13g2_a22oi_1 _5660_ (.Y(_1885_),
    .B1(_1879_),
    .B2(_1884_),
    .A2(_1876_),
    .A1(_1820_));
 sg13g2_o21ai_1 _5661_ (.B1(_1885_),
    .Y(_0008_),
    .A1(net192),
    .A2(_1874_));
 sg13g2_nor2_1 _5662_ (.A(net213),
    .B(_1813_),
    .Y(_1886_));
 sg13g2_a21oi_1 _5663_ (.A1(_1860_),
    .A2(net213),
    .Y(_1887_),
    .B1(_1886_));
 sg13g2_inv_1 _5664_ (.Y(_1888_),
    .A(_1814_));
 sg13g2_nand2_1 _5665_ (.Y(_1889_),
    .A(net216),
    .B(net215));
 sg13g2_nand3_1 _5666_ (.B(_1889_),
    .C(_1824_),
    .A(_1888_),
    .Y(_1891_));
 sg13g2_o21ai_1 _5667_ (.B1(_1891_),
    .Y(_1892_),
    .A1(net192),
    .A2(_1887_));
 sg13g2_nand2_1 _5668_ (.Y(_1893_),
    .A(_1892_),
    .B(net214));
 sg13g2_nor2_2 _5669_ (.A(net214),
    .B(_1846_),
    .Y(_1894_));
 sg13g2_inv_1 _5670_ (.Y(_1895_),
    .A(_1824_));
 sg13g2_a21oi_1 _5671_ (.A1(_1895_),
    .A2(net192),
    .Y(_1896_),
    .B1(_1888_));
 sg13g2_nor2b_1 _5672_ (.A(_1881_),
    .B_N(_1889_),
    .Y(_1897_));
 sg13g2_inv_1 _5673_ (.Y(_1898_),
    .A(_1886_));
 sg13g2_a22oi_1 _5674_ (.Y(_1899_),
    .B1(_1804_),
    .B2(_1898_),
    .A2(net212),
    .A1(_1897_));
 sg13g2_a22oi_1 _5675_ (.Y(_1900_),
    .B1(_1820_),
    .B2(_1899_),
    .A2(_1896_),
    .A1(_1894_));
 sg13g2_nand2_1 _5676_ (.Y(_0009_),
    .A(_1893_),
    .B(_1900_));
 sg13g2_nor2_1 _5677_ (.A(net213),
    .B(_1812_),
    .Y(_1902_));
 sg13g2_inv_1 _5678_ (.Y(_1903_),
    .A(_1902_));
 sg13g2_a22oi_1 _5679_ (.Y(_1904_),
    .B1(_1830_),
    .B2(_1878_),
    .A2(net212),
    .A1(_1903_));
 sg13g2_nor2_1 _5680_ (.A(_1875_),
    .B(_1882_),
    .Y(_1905_));
 sg13g2_nand2_1 _5681_ (.Y(_1906_),
    .A(_1894_),
    .B(_1812_));
 sg13g2_nand2_1 _5682_ (.Y(_1907_),
    .A(_1797_),
    .B(_1799_));
 sg13g2_nand2_1 _5683_ (.Y(_1908_),
    .A(_1824_),
    .B(_1907_));
 sg13g2_inv_1 _5684_ (.Y(_1909_),
    .A(_1908_));
 sg13g2_nand2_1 _5685_ (.Y(_1910_),
    .A(_1906_),
    .B(_1909_));
 sg13g2_nor2_1 _5686_ (.A(_1905_),
    .B(_1910_),
    .Y(_1912_));
 sg13g2_nand3b_1 _5687_ (.B(net214),
    .C(net218),
    .Y(_1913_),
    .A_N(_1825_));
 sg13g2_a21oi_1 _5688_ (.A1(_1913_),
    .A2(_1906_),
    .Y(_1914_),
    .B1(_1821_));
 sg13g2_nor2_1 _5689_ (.A(_1912_),
    .B(_1914_),
    .Y(_1915_));
 sg13g2_o21ai_1 _5690_ (.B1(_1915_),
    .Y(_0010_),
    .A1(net192),
    .A2(_1904_));
 sg13g2_nand2_1 _5691_ (.Y(_1916_),
    .A(_1870_),
    .B(_1839_));
 sg13g2_nand3_1 _5692_ (.B(_1836_),
    .C(_1872_),
    .A(_1916_),
    .Y(_1917_));
 sg13g2_nor2_1 _5693_ (.A(_1821_),
    .B(_1830_),
    .Y(_1918_));
 sg13g2_nand2_1 _5694_ (.Y(_1919_),
    .A(_1826_),
    .B(_1812_));
 sg13g2_nor2_1 _5695_ (.A(_1894_),
    .B(_1908_),
    .Y(_1920_));
 sg13g2_a22oi_1 _5696_ (.Y(_1922_),
    .B1(_1849_),
    .B2(_1920_),
    .A2(_1919_),
    .A1(_1918_));
 sg13g2_nand2_1 _5697_ (.Y(_0011_),
    .A(_1917_),
    .B(_1922_));
 sg13g2_nand3_1 _5698_ (.B(_1818_),
    .C(_1906_),
    .A(_1854_),
    .Y(_1923_));
 sg13g2_nor2_1 _5699_ (.A(_1801_),
    .B(_1810_),
    .Y(_1924_));
 sg13g2_nand3b_1 _5700_ (.B(_1834_),
    .C(_1889_),
    .Y(_1925_),
    .A_N(_1924_));
 sg13g2_nand3_1 _5701_ (.B(_1822_),
    .C(_1925_),
    .A(_1923_),
    .Y(_1926_));
 sg13g2_o21ai_1 _5702_ (.B1(_1920_),
    .Y(_1927_),
    .A1(_1876_),
    .A2(_1852_));
 sg13g2_nand2_1 _5703_ (.Y(_0012_),
    .A(_1926_),
    .B(_1927_));
 sg13g2_nor3_1 _5704_ (.A(net212),
    .B(_1846_),
    .C(_1902_),
    .Y(_1928_));
 sg13g2_o21ai_1 _5705_ (.B1(_1836_),
    .Y(_1929_),
    .A1(_1902_),
    .A2(_1814_));
 sg13g2_a21oi_1 _5706_ (.A1(_1846_),
    .A2(net212),
    .Y(_1931_),
    .B1(_1895_));
 sg13g2_a22oi_1 _5707_ (.Y(_1932_),
    .B1(_1863_),
    .B2(_1931_),
    .A2(_1820_),
    .A1(_1826_));
 sg13g2_o21ai_1 _5708_ (.B1(_1932_),
    .Y(_0013_),
    .A1(_1928_),
    .A2(_1929_));
 sg13g2_inv_1 _5709_ (.Y(_1933_),
    .A(_1815_));
 sg13g2_nand3_1 _5710_ (.B(net214),
    .C(net213),
    .A(_1846_),
    .Y(_1934_));
 sg13g2_nand3_1 _5711_ (.B(_1836_),
    .C(_1934_),
    .A(_1933_),
    .Y(_1935_));
 sg13g2_o21ai_1 _5712_ (.B1(_1935_),
    .Y(_0014_),
    .A1(_1864_),
    .A2(_1908_));
 sg13g2_o21ai_1 _5713_ (.B1(_1908_),
    .Y(_0015_),
    .A1(_1837_),
    .A2(_1933_));
 sg13g2_nor2_1 _5714_ (.A(net217),
    .B(_1902_),
    .Y(_1936_));
 sg13g2_inv_1 _5715_ (.Y(_1937_),
    .A(_1857_));
 sg13g2_a22oi_1 _5716_ (.Y(_1939_),
    .B1(_1898_),
    .B2(_1937_),
    .A2(_1878_),
    .A1(_1936_));
 sg13g2_nor2_1 _5717_ (.A(net218),
    .B(net213),
    .Y(_1940_));
 sg13g2_o21ai_1 _5718_ (.B1(_1909_),
    .Y(_1941_),
    .A1(_1940_),
    .A2(_1924_));
 sg13g2_xor2_1 _5719_ (.B(_1801_),
    .A(net217),
    .X(_1942_));
 sg13g2_nand3_1 _5720_ (.B(_1942_),
    .C(_1822_),
    .A(_1863_),
    .Y(_1943_));
 sg13g2_nand3_1 _5721_ (.B(_1943_),
    .C(_1837_),
    .A(_1941_),
    .Y(_1944_));
 sg13g2_o21ai_1 _5722_ (.B1(_1944_),
    .Y(_0001_),
    .A1(net192),
    .A2(_1939_));
 sg13g2_inv_1 _5723_ (.Y(_1945_),
    .A(_1803_));
 sg13g2_nand2_1 _5724_ (.Y(_1946_),
    .A(_1945_),
    .B(_1796_));
 sg13g2_a21oi_1 _5725_ (.A1(_1946_),
    .A2(_1830_),
    .Y(_1947_),
    .B1(_1873_));
 sg13g2_a21oi_1 _5726_ (.A1(_1809_),
    .A2(_1945_),
    .Y(_1949_),
    .B1(_1867_));
 sg13g2_a21oi_1 _5727_ (.A1(_1894_),
    .A2(_1889_),
    .Y(_1950_),
    .B1(net192));
 sg13g2_o21ai_1 _5728_ (.B1(_1950_),
    .Y(_1951_),
    .A1(net212),
    .A2(_1868_));
 sg13g2_o21ai_1 _5729_ (.B1(_1951_),
    .Y(_1952_),
    .A1(_1910_),
    .A2(_1949_));
 sg13g2_a21oi_1 _5730_ (.A1(_1820_),
    .A2(_1947_),
    .Y(_0002_),
    .B1(_1952_));
 sg13g2_nor2_1 _5731_ (.A(net217),
    .B(_1840_),
    .Y(_1953_));
 sg13g2_nor2_1 _5732_ (.A(_1857_),
    .B(_1868_),
    .Y(_1954_));
 sg13g2_o21ai_1 _5733_ (.B1(_1836_),
    .Y(_1955_),
    .A1(_1953_),
    .A2(_1954_));
 sg13g2_nor2_1 _5734_ (.A(_1853_),
    .B(_1937_),
    .Y(_1956_));
 sg13g2_o21ai_1 _5735_ (.B1(_1820_),
    .Y(_1957_),
    .A1(_1940_),
    .A2(_1956_));
 sg13g2_o21ai_1 _5736_ (.B1(_1920_),
    .Y(_1959_),
    .A1(_1813_),
    .A2(_1882_));
 sg13g2_nand3_1 _5737_ (.B(_1957_),
    .C(_1959_),
    .A(_1955_),
    .Y(_0003_));
 sg13g2_nand2b_1 _5738_ (.Y(_1960_),
    .B(_1870_),
    .A_N(_1825_));
 sg13g2_nand3_1 _5739_ (.B(_1834_),
    .C(_1857_),
    .A(_1960_),
    .Y(_1961_));
 sg13g2_a21oi_1 _5740_ (.A1(_1841_),
    .A2(net217),
    .Y(_1962_),
    .B1(_1851_));
 sg13g2_a21oi_1 _5741_ (.A1(_1962_),
    .A2(_1818_),
    .Y(_1963_),
    .B1(net1));
 sg13g2_nand2_1 _5742_ (.Y(_1964_),
    .A(_1961_),
    .B(_1963_));
 sg13g2_nand2_1 _5743_ (.Y(_1965_),
    .A(_1853_),
    .B(_1809_));
 sg13g2_o21ai_1 _5744_ (.B1(net212),
    .Y(_1966_),
    .A1(_1808_),
    .A2(_1812_));
 sg13g2_nand3_1 _5745_ (.B(_1824_),
    .C(_1966_),
    .A(_1965_),
    .Y(_1967_));
 sg13g2_nand2_1 _5746_ (.Y(_0004_),
    .A(_1964_),
    .B(_1967_));
 sg13g2_o21ai_1 _5747_ (.B1(net214),
    .Y(_1969_),
    .A1(net216),
    .A2(_1840_));
 sg13g2_nor2b_1 _5748_ (.A(_1894_),
    .B_N(_1969_),
    .Y(_1970_));
 sg13g2_nor2_1 _5749_ (.A(net216),
    .B(_1881_),
    .Y(_1971_));
 sg13g2_nand2_1 _5750_ (.Y(_1972_),
    .A(_1820_),
    .B(_1907_));
 sg13g2_inv_1 _5751_ (.Y(_1973_),
    .A(_1972_));
 sg13g2_a22oi_1 _5752_ (.Y(_1974_),
    .B1(_1973_),
    .B2(_1969_),
    .A2(_1971_),
    .A1(_1909_));
 sg13g2_o21ai_1 _5753_ (.B1(_1974_),
    .Y(_0005_),
    .A1(net192),
    .A2(_1970_));
 sg13g2_nand3_1 _5754_ (.B(_1846_),
    .C(net212),
    .A(_1836_),
    .Y(_1975_));
 sg13g2_o21ai_1 _5755_ (.B1(_1975_),
    .Y(_0006_),
    .A1(_1895_),
    .A2(_1965_));
 sg13g2_nand2_1 _5756_ (.Y(_1977_),
    .A(_2239_),
    .B(net120));
 sg13g2_nand2_1 _5757_ (.Y(_1978_),
    .A(_3031_),
    .B(_1977_));
 sg13g2_a21oi_1 _5758_ (.A1(_1978_),
    .A2(_0234_),
    .Y(_1979_),
    .B1(net66));
 sg13g2_nand2_1 _5759_ (.Y(_1980_),
    .A(_0359_),
    .B(_0422_));
 sg13g2_o21ai_1 _5760_ (.B1(_1980_),
    .Y(_1981_),
    .A1(net36),
    .A2(_2961_));
 sg13g2_nand2_1 _5761_ (.Y(_1982_),
    .A(_1981_),
    .B(net105));
 sg13g2_nor3_1 _5762_ (.A(_1380_),
    .B(_1107_),
    .C(_2550_),
    .Y(_1983_));
 sg13g2_nand2_1 _5763_ (.Y(_1984_),
    .A(_2890_),
    .B(_1983_));
 sg13g2_nand2_1 _5764_ (.Y(_1985_),
    .A(_0333_),
    .B(_3026_));
 sg13g2_nand2_1 _5765_ (.Y(_1986_),
    .A(_1985_),
    .B(_0600_));
 sg13g2_nand3_1 _5766_ (.B(_1984_),
    .C(_1986_),
    .A(_1982_),
    .Y(_1988_));
 sg13g2_nor2_1 _5767_ (.A(_1979_),
    .B(_1988_),
    .Y(_1989_));
 sg13g2_nand2_1 _5768_ (.Y(_1990_),
    .A(_0100_),
    .B(_0921_));
 sg13g2_nor2b_1 _5769_ (.A(_1159_),
    .B_N(_2605_),
    .Y(_1991_));
 sg13g2_nand2_1 _5770_ (.Y(_1992_),
    .A(net86),
    .B(net125));
 sg13g2_nand2_1 _5771_ (.Y(_1993_),
    .A(_1991_),
    .B(_1992_));
 sg13g2_a22oi_1 _5772_ (.Y(_1994_),
    .B1(net25),
    .B2(_1993_),
    .A2(_0334_),
    .A1(_1990_));
 sg13g2_o21ai_1 _5773_ (.B1(_0542_),
    .Y(_1995_),
    .A1(_2758_),
    .A2(net59));
 sg13g2_nand2_1 _5774_ (.Y(_1996_),
    .A(_1995_),
    .B(net26));
 sg13g2_nand2_1 _5775_ (.Y(_1997_),
    .A(_1994_),
    .B(_1996_));
 sg13g2_nand2_1 _5776_ (.Y(_1999_),
    .A(_1997_),
    .B(net117));
 sg13g2_a21oi_1 _5777_ (.A1(_1989_),
    .A2(_1999_),
    .Y(_2000_),
    .B1(_0729_));
 sg13g2_nand3b_1 _5778_ (.B(_1446_),
    .C(net90),
    .Y(_2001_),
    .A_N(_2461_));
 sg13g2_nand3_1 _5779_ (.B(_2426_),
    .C(_2615_),
    .A(_0224_),
    .Y(_2002_));
 sg13g2_nand3_1 _5780_ (.B(_2002_),
    .C(_2595_),
    .A(_2001_),
    .Y(_2003_));
 sg13g2_a22oi_1 _5781_ (.Y(_2004_),
    .B1(_2711_),
    .B2(net141),
    .A2(net119),
    .A1(_1435_));
 sg13g2_o21ai_1 _5782_ (.B1(_2004_),
    .Y(_2005_),
    .A1(net102),
    .A2(_0181_));
 sg13g2_nand2_1 _5783_ (.Y(_2006_),
    .A(_2005_),
    .B(net129));
 sg13g2_nor2b_1 _5784_ (.A(_2003_),
    .B_N(_2006_),
    .Y(_2007_));
 sg13g2_nand2b_1 _5785_ (.Y(_2008_),
    .B(_0182_),
    .A_N(_1697_));
 sg13g2_nand2_1 _5786_ (.Y(_2010_),
    .A(_1463_),
    .B(_2585_));
 sg13g2_nand2_1 _5787_ (.Y(_2011_),
    .A(_2010_),
    .B(_2910_));
 sg13g2_nor2_1 _5788_ (.A(net23),
    .B(_2011_),
    .Y(_2012_));
 sg13g2_a21oi_1 _5789_ (.A1(_2008_),
    .A2(_2991_),
    .Y(_2013_),
    .B1(_2012_));
 sg13g2_nand2_1 _5790_ (.Y(_2014_),
    .A(_2007_),
    .B(_2013_));
 sg13g2_a21oi_1 _5791_ (.A1(_2403_),
    .A2(_1160_),
    .Y(_2015_),
    .B1(_2963_));
 sg13g2_nor2_1 _5792_ (.A(net62),
    .B(_2900_),
    .Y(_2016_));
 sg13g2_a21oi_1 _5793_ (.A1(_2016_),
    .A2(_2933_),
    .Y(_2017_),
    .B1(_1380_));
 sg13g2_nor2b_1 _5794_ (.A(_2015_),
    .B_N(_2017_),
    .Y(_2018_));
 sg13g2_nand3_1 _5795_ (.B(net102),
    .C(_2997_),
    .A(net57),
    .Y(_2019_));
 sg13g2_nand2_1 _5796_ (.Y(_2021_),
    .A(_2019_),
    .B(_2514_));
 sg13g2_nand2_1 _5797_ (.Y(_2022_),
    .A(_2021_),
    .B(net25));
 sg13g2_o21ai_1 _5798_ (.B1(net102),
    .Y(_2023_),
    .A1(_1478_),
    .A2(_2501_));
 sg13g2_nand2_1 _5799_ (.Y(_2024_),
    .A(_2023_),
    .B(_2845_));
 sg13g2_nand2_1 _5800_ (.Y(_2025_),
    .A(_2024_),
    .B(_2569_));
 sg13g2_nand3_1 _5801_ (.B(_2022_),
    .C(_2025_),
    .A(_2018_),
    .Y(_2026_));
 sg13g2_nand3_1 _5802_ (.B(_2026_),
    .C(_2598_),
    .A(_2014_),
    .Y(_2027_));
 sg13g2_nand2_1 _5803_ (.Y(_2028_),
    .A(_2027_),
    .B(net195));
 sg13g2_nor2_1 _5804_ (.A(_2000_),
    .B(_2028_),
    .Y(_2029_));
 sg13g2_nand3_1 _5805_ (.B(_1197_),
    .C(net69),
    .A(_0704_),
    .Y(_2030_));
 sg13g2_nand2_1 _5806_ (.Y(_2032_),
    .A(_2030_),
    .B(_2556_));
 sg13g2_nand3_1 _5807_ (.B(_0782_),
    .C(_2526_),
    .A(_3048_),
    .Y(_2033_));
 sg13g2_nand2_1 _5808_ (.Y(_2034_),
    .A(_2033_),
    .B(net129));
 sg13g2_nand2_1 _5809_ (.Y(_2035_),
    .A(_2766_),
    .B(_1653_));
 sg13g2_nand2_1 _5810_ (.Y(_2036_),
    .A(_2035_),
    .B(_2990_));
 sg13g2_nand2_1 _5811_ (.Y(_2037_),
    .A(_2034_),
    .B(_2036_));
 sg13g2_nor2_1 _5812_ (.A(_2032_),
    .B(_2037_),
    .Y(_2038_));
 sg13g2_nor2_1 _5813_ (.A(net118),
    .B(_2038_),
    .Y(_2039_));
 sg13g2_a21oi_1 _5814_ (.A1(_2893_),
    .A2(_0100_),
    .Y(_2040_),
    .B1(_0294_));
 sg13g2_a21oi_1 _5815_ (.A1(_1425_),
    .A2(_2541_),
    .Y(_2041_),
    .B1(_2384_));
 sg13g2_nand2_1 _5816_ (.Y(_2043_),
    .A(_0234_),
    .B(_2961_));
 sg13g2_nand2_1 _5817_ (.Y(_2044_),
    .A(_2043_),
    .B(net110));
 sg13g2_nand2_1 _5818_ (.Y(_2045_),
    .A(_1114_),
    .B(_0617_));
 sg13g2_nand2_1 _5819_ (.Y(_2046_),
    .A(_2045_),
    .B(net134));
 sg13g2_nand2_1 _5820_ (.Y(_2047_),
    .A(_2044_),
    .B(_2046_));
 sg13g2_nor3_1 _5821_ (.A(_2040_),
    .B(_2041_),
    .C(_2047_),
    .Y(_2048_));
 sg13g2_nor2_1 _5822_ (.A(_2375_),
    .B(_2048_),
    .Y(_2049_));
 sg13g2_nor2_1 _5823_ (.A(_2039_),
    .B(_2049_),
    .Y(_2050_));
 sg13g2_nand3_1 _5824_ (.B(_3048_),
    .C(_2526_),
    .A(_0622_),
    .Y(_2051_));
 sg13g2_nand2_1 _5825_ (.Y(_2052_),
    .A(_2051_),
    .B(_2626_));
 sg13g2_nand2_1 _5826_ (.Y(_2054_),
    .A(_0318_),
    .B(_2617_));
 sg13g2_nand2_1 _5827_ (.Y(_2055_),
    .A(_2054_),
    .B(_2990_));
 sg13g2_nand2_1 _5828_ (.Y(_2056_),
    .A(_2052_),
    .B(_2055_));
 sg13g2_nor2_1 _5829_ (.A(net64),
    .B(_1169_),
    .Y(_2057_));
 sg13g2_nand2_1 _5830_ (.Y(_2058_),
    .A(_2057_),
    .B(_2797_));
 sg13g2_nor2_1 _5831_ (.A(_2383_),
    .B(_0346_),
    .Y(_2059_));
 sg13g2_nand2_1 _5832_ (.Y(_2060_),
    .A(_2834_),
    .B(_2728_));
 sg13g2_nand2_1 _5833_ (.Y(_2061_),
    .A(_2059_),
    .B(_2060_));
 sg13g2_nand3_1 _5834_ (.B(_2061_),
    .C(_2619_),
    .A(_2058_),
    .Y(_2062_));
 sg13g2_nor2_1 _5835_ (.A(_2056_),
    .B(_2062_),
    .Y(_2063_));
 sg13g2_nor2_1 _5836_ (.A(net166),
    .B(_2063_),
    .Y(_2065_));
 sg13g2_nand2_1 _5837_ (.Y(_2066_),
    .A(_2614_),
    .B(net84));
 sg13g2_nand2_1 _5838_ (.Y(_2067_),
    .A(_2674_),
    .B(_2992_));
 sg13g2_a21oi_1 _5839_ (.A1(_0958_),
    .A2(_2067_),
    .Y(_2068_),
    .B1(net81));
 sg13g2_o21ai_1 _5840_ (.B1(_2068_),
    .Y(_2069_),
    .A1(_2756_),
    .A2(_2066_));
 sg13g2_nand2_1 _5841_ (.Y(_2070_),
    .A(_0556_),
    .B(net92));
 sg13g2_nor2_1 _5842_ (.A(net151),
    .B(_2745_),
    .Y(_2071_));
 sg13g2_nand2_1 _5843_ (.Y(_2072_),
    .A(_2070_),
    .B(_2071_));
 sg13g2_nand2_1 _5844_ (.Y(_2073_),
    .A(_1104_),
    .B(_0833_));
 sg13g2_nand2_1 _5845_ (.Y(_2074_),
    .A(_2072_),
    .B(_2073_));
 sg13g2_nand2_1 _5846_ (.Y(_2076_),
    .A(_2074_),
    .B(net123));
 sg13g2_nand2_1 _5847_ (.Y(_2077_),
    .A(_2076_),
    .B(net35));
 sg13g2_nand2_1 _5848_ (.Y(_2078_),
    .A(_2069_),
    .B(_2077_));
 sg13g2_nand2_1 _5849_ (.Y(_2079_),
    .A(_2065_),
    .B(_2078_));
 sg13g2_nand2_1 _5850_ (.Y(_2080_),
    .A(_2050_),
    .B(_2079_));
 sg13g2_nand2_1 _5851_ (.Y(_2081_),
    .A(_2080_),
    .B(net132));
 sg13g2_a21oi_1 _5852_ (.A1(_0999_),
    .A2(_1574_),
    .Y(_2082_),
    .B1(net78));
 sg13g2_nand2_1 _5853_ (.Y(_2083_),
    .A(_1165_),
    .B(_1589_));
 sg13g2_nand2_1 _5854_ (.Y(_2084_),
    .A(_2082_),
    .B(_2083_));
 sg13g2_a21oi_1 _5855_ (.A1(_1318_),
    .A2(_1559_),
    .Y(_2085_),
    .B1(_2384_));
 sg13g2_a21oi_1 _5856_ (.A1(_2898_),
    .A2(_2010_),
    .Y(_2087_),
    .B1(_2085_));
 sg13g2_nand2_1 _5857_ (.Y(_2088_),
    .A(_2084_),
    .B(_2087_));
 sg13g2_nand2_1 _5858_ (.Y(_2089_),
    .A(_2088_),
    .B(net83));
 sg13g2_a21oi_1 _5859_ (.A1(_2394_),
    .A2(_0387_),
    .Y(_2090_),
    .B1(_0868_));
 sg13g2_nand3_1 _5860_ (.B(_2071_),
    .C(net113),
    .A(_1178_),
    .Y(_2091_));
 sg13g2_nand2_1 _5861_ (.Y(_2092_),
    .A(_2091_),
    .B(net197));
 sg13g2_nor2_1 _5862_ (.A(net41),
    .B(_1158_),
    .Y(_2093_));
 sg13g2_a22oi_1 _5863_ (.Y(_2094_),
    .B1(_0332_),
    .B2(_2093_),
    .A2(_2842_),
    .A1(_2577_));
 sg13g2_nand2_1 _5864_ (.Y(_2095_),
    .A(_0302_),
    .B(_2637_));
 sg13g2_a21oi_1 _5865_ (.A1(_2094_),
    .A2(_2095_),
    .Y(_2096_),
    .B1(_0118_));
 sg13g2_nor3_1 _5866_ (.A(_2090_),
    .B(_2092_),
    .C(_2096_),
    .Y(_2098_));
 sg13g2_a21oi_1 _5867_ (.A1(_2089_),
    .A2(_2098_),
    .Y(_2099_),
    .B1(_2424_));
 sg13g2_nor2_1 _5868_ (.A(_2257_),
    .B(_2392_),
    .Y(_2100_));
 sg13g2_nor3_1 _5869_ (.A(_2173_),
    .B(_2203_),
    .C(_2100_),
    .Y(_2101_));
 sg13g2_a21oi_1 _5870_ (.A1(_2101_),
    .A2(_2625_),
    .Y(_2102_),
    .B1(_2689_));
 sg13g2_nand3_1 _5871_ (.B(_3043_),
    .C(net84),
    .A(_2797_),
    .Y(_2103_));
 sg13g2_nand2_1 _5872_ (.Y(_2104_),
    .A(_2102_),
    .B(_2103_));
 sg13g2_nand2_1 _5873_ (.Y(_2105_),
    .A(_0223_),
    .B(_1407_));
 sg13g2_nand2_1 _5874_ (.Y(_2106_),
    .A(_2105_),
    .B(net26));
 sg13g2_nand2_1 _5875_ (.Y(_2107_),
    .A(_2019_),
    .B(_2970_));
 sg13g2_nand2_1 _5876_ (.Y(_2109_),
    .A(_2107_),
    .B(net70));
 sg13g2_nand3_1 _5877_ (.B(_2106_),
    .C(_2109_),
    .A(_2104_),
    .Y(_2110_));
 sg13g2_nand2_1 _5878_ (.Y(_2111_),
    .A(_2110_),
    .B(net83));
 sg13g2_inv_1 _5879_ (.Y(_2112_),
    .A(_0154_));
 sg13g2_nand2_1 _5880_ (.Y(_2113_),
    .A(_1204_),
    .B(net56));
 sg13g2_nand3_1 _5881_ (.B(net84),
    .C(_1991_),
    .A(_2113_),
    .Y(_2114_));
 sg13g2_nand2_1 _5882_ (.Y(_2115_),
    .A(_2114_),
    .B(net22));
 sg13g2_a21oi_1 _5883_ (.A1(_0221_),
    .A2(_2112_),
    .Y(_2116_),
    .B1(_2115_));
 sg13g2_a21oi_1 _5884_ (.A1(_0167_),
    .A2(_0387_),
    .Y(_2117_),
    .B1(net160));
 sg13g2_a21oi_1 _5885_ (.A1(net139),
    .A2(_1162_),
    .Y(_2118_),
    .B1(net142));
 sg13g2_nand3_1 _5886_ (.B(net206),
    .C(net119),
    .A(net30),
    .Y(_2120_));
 sg13g2_nand3_1 _5887_ (.B(_2118_),
    .C(_2120_),
    .A(_2548_),
    .Y(_2121_));
 sg13g2_a21oi_1 _5888_ (.A1(_2117_),
    .A2(_2121_),
    .Y(_2122_),
    .B1(net166));
 sg13g2_nor2b_1 _5889_ (.A(_2116_),
    .B_N(_2122_),
    .Y(_2123_));
 sg13g2_nand2_1 _5890_ (.Y(_2124_),
    .A(_2111_),
    .B(_2123_));
 sg13g2_nand2_1 _5891_ (.Y(_2125_),
    .A(_1056_),
    .B(_2688_));
 sg13g2_nor2_1 _5892_ (.A(_2125_),
    .B(_0324_),
    .Y(_2126_));
 sg13g2_nand3_1 _5893_ (.B(_0471_),
    .C(_2516_),
    .A(_0174_),
    .Y(_2127_));
 sg13g2_nand2_1 _5894_ (.Y(_2128_),
    .A(_2127_),
    .B(_1372_));
 sg13g2_nor2_1 _5895_ (.A(_2126_),
    .B(_2128_),
    .Y(_2129_));
 sg13g2_a22oi_1 _5896_ (.Y(_2131_),
    .B1(_2544_),
    .B2(_1097_),
    .A2(_0951_),
    .A1(_2795_));
 sg13g2_nand3_1 _5897_ (.B(_2684_),
    .C(_2732_),
    .A(_2571_),
    .Y(_2132_));
 sg13g2_inv_1 _5898_ (.Y(_2133_),
    .A(_0748_));
 sg13g2_a21oi_1 _5899_ (.A1(_2131_),
    .A2(_2132_),
    .Y(_2134_),
    .B1(_2133_));
 sg13g2_nor2_1 _5900_ (.A(_2129_),
    .B(_2134_),
    .Y(_2135_));
 sg13g2_a21oi_1 _5901_ (.A1(_0716_),
    .A2(_2651_),
    .Y(_2136_),
    .B1(net160));
 sg13g2_nand3_1 _5902_ (.B(_1171_),
    .C(_2653_),
    .A(_0285_),
    .Y(_2137_));
 sg13g2_nand2_1 _5903_ (.Y(_2138_),
    .A(_2136_),
    .B(_2137_));
 sg13g2_nand2_1 _5904_ (.Y(_2139_),
    .A(_2797_),
    .B(_3043_));
 sg13g2_nand2_1 _5905_ (.Y(_2140_),
    .A(_2139_),
    .B(_0600_));
 sg13g2_nand2_1 _5906_ (.Y(_2142_),
    .A(_2138_),
    .B(_2140_));
 sg13g2_nand3_1 _5907_ (.B(_2719_),
    .C(_0604_),
    .A(_2010_),
    .Y(_2143_));
 sg13g2_nor2b_1 _5908_ (.A(_2142_),
    .B_N(_2143_),
    .Y(_2144_));
 sg13g2_nand2_1 _5909_ (.Y(_2145_),
    .A(_2135_),
    .B(_2144_));
 sg13g2_nand2_1 _5910_ (.Y(_2146_),
    .A(_2145_),
    .B(net112));
 sg13g2_a221oi_1 _5911_ (.B2(_0958_),
    .C1(_0960_),
    .B1(_2943_),
    .A1(_0977_),
    .Y(_2147_),
    .A2(_1083_));
 sg13g2_nor2_1 _5912_ (.A(_2695_),
    .B(_2147_),
    .Y(_2148_));
 sg13g2_nand2_1 _5913_ (.Y(_2149_),
    .A(_2146_),
    .B(_2148_));
 sg13g2_a21oi_1 _5914_ (.A1(_2099_),
    .A2(_2124_),
    .Y(_2150_),
    .B1(_2149_));
 sg13g2_a21oi_1 _5915_ (.A1(_2029_),
    .A2(_2081_),
    .Y(_0016_),
    .B1(_2150_));
 sg13g2_buf_2 _5916_ (.A(\clk_picker.counter[9] ),
    .X(_2152_));
 sg13g2_nor3_1 _5917_ (.A(_2152_),
    .B(\clk_picker.counter[10] ),
    .C(\clk_picker.counter[11] ),
    .Y(_2153_));
 sg13g2_inv_1 _5918_ (.Y(_2154_),
    .A(\clk_picker.counter[7] ));
 sg13g2_inv_1 _5919_ (.Y(_2155_),
    .A(\clk_picker.counter[8] ));
 sg13g2_nand3_1 _5920_ (.B(_2154_),
    .C(_2155_),
    .A(_2153_),
    .Y(_2156_));
 sg13g2_buf_1 _5921_ (.A(\clk_picker.counter[17] ),
    .X(_2157_));
 sg13g2_nand2_1 _5922_ (.Y(_2158_),
    .A(\clk_picker.counter[12] ),
    .B(\clk_picker.counter[13] ));
 sg13g2_inv_1 _5923_ (.Y(_2159_),
    .A(_2158_));
 sg13g2_nand2_1 _5924_ (.Y(_2160_),
    .A(\clk_picker.counter[14] ),
    .B(\clk_picker.counter[15] ));
 sg13g2_inv_1 _5925_ (.Y(_2161_),
    .A(_2160_));
 sg13g2_nand4_1 _5926_ (.B(_2157_),
    .C(_2159_),
    .A(_2156_),
    .Y(_2163_),
    .D(_2161_));
 sg13g2_inv_1 _5927_ (.Y(_2164_),
    .A(\clk_picker.counter[18] ));
 sg13g2_nand2_1 _5928_ (.Y(_2165_),
    .A(\clk_picker.counter[16] ),
    .B(_2157_));
 sg13g2_nand3_1 _5929_ (.B(_2164_),
    .C(_2165_),
    .A(_2163_),
    .Y(_2166_));
 sg13g2_inv_1 _5930_ (.Y(_2167_),
    .A(\clk_picker.counter[20] ));
 sg13g2_inv_1 _5931_ (.Y(_2168_),
    .A(\clk_picker.counter[23] ));
 sg13g2_nand2_1 _5932_ (.Y(_2169_),
    .A(\clk_picker.counter[21] ),
    .B(\clk_picker.counter[22] ));
 sg13g2_nor3_1 _5933_ (.A(_2167_),
    .B(_2168_),
    .C(_2169_),
    .Y(_2170_));
 sg13g2_nand4_1 _5934_ (.B(\clk_picker.counter[19] ),
    .C(\clk_picker.counter[25] ),
    .A(_2166_),
    .Y(_2171_),
    .D(_2170_));
 sg13g2_nand2_2 _5935_ (.Y(_2172_),
    .A(\clk_picker.counter[24] ),
    .B(\clk_picker.counter[25] ));
 sg13g2_nand2_1 _5936_ (.Y(_2174_),
    .A(_2171_),
    .B(_2172_));
 sg13g2_nand2_1 _5937_ (.Y(_2175_),
    .A(_2174_),
    .B(_0030_));
 sg13g2_nand3_1 _5938_ (.B(\clk_picker.clk_slow ),
    .C(_2172_),
    .A(_2171_),
    .Y(_2176_));
 sg13g2_buf_2 _5939_ (.A(rst_n),
    .X(_2177_));
 sg13g2_inv_2 _5940_ (.Y(_2178_),
    .A(_2177_));
 sg13g2_buf_1 _5941_ (.A(_2178_),
    .X(_2179_));
 sg13g2_a21oi_1 _5942_ (.A1(_2175_),
    .A2(_2176_),
    .Y(_0040_),
    .B1(_2179_));
 sg13g2_nand3_1 _5943_ (.B(_2177_),
    .C(_2172_),
    .A(_2171_),
    .Y(_2180_));
 sg13g2_buf_2 _5944_ (.A(_2180_),
    .X(_2181_));
 sg13g2_buf_1 _5945_ (.A(_2181_),
    .X(_2182_));
 sg13g2_nor2b_1 _5946_ (.A(net21),
    .B_N(_0039_),
    .Y(_0041_));
 sg13g2_inv_1 _5947_ (.Y(_2184_),
    .A(\clk_picker.counter[10] ));
 sg13g2_inv_1 _5948_ (.Y(_2185_),
    .A(\clk_picker.counter[5] ));
 sg13g2_inv_1 _5949_ (.Y(_2186_),
    .A(\clk_picker.counter[6] ));
 sg13g2_nand2_1 _5950_ (.Y(_2187_),
    .A(\clk_picker.counter[1] ),
    .B(\clk_picker.counter[0] ));
 sg13g2_nor2b_1 _5951_ (.A(_2187_),
    .B_N(\clk_picker.counter[2] ),
    .Y(_2188_));
 sg13g2_and2_1 _5952_ (.A(_2188_),
    .B(\clk_picker.counter[3] ),
    .X(_2189_));
 sg13g2_buf_8 _5953_ (.A(_2189_),
    .X(_2190_));
 sg13g2_nand2_1 _5954_ (.Y(_2191_),
    .A(_2190_),
    .B(\clk_picker.counter[4] ));
 sg13g2_nor3_1 _5955_ (.A(_2185_),
    .B(_2186_),
    .C(_2191_),
    .Y(_2192_));
 sg13g2_nand2_1 _5956_ (.Y(_2194_),
    .A(_2192_),
    .B(\clk_picker.counter[7] ));
 sg13g2_nor2_2 _5957_ (.A(_2155_),
    .B(_2194_),
    .Y(_2195_));
 sg13g2_nand2_1 _5958_ (.Y(_2196_),
    .A(_2195_),
    .B(_2152_));
 sg13g2_xnor2_1 _5959_ (.Y(_2197_),
    .A(_2184_),
    .B(_2196_));
 sg13g2_buf_1 _5960_ (.A(_2181_),
    .X(_2198_));
 sg13g2_nor2_1 _5961_ (.A(_2197_),
    .B(net20),
    .Y(_0042_));
 sg13g2_inv_1 _5962_ (.Y(_2199_),
    .A(_2152_));
 sg13g2_nor4_1 _5963_ (.A(_2154_),
    .B(_2155_),
    .C(_2199_),
    .D(_2184_),
    .Y(_2200_));
 sg13g2_inv_1 _5964_ (.Y(_2201_),
    .A(_2200_));
 sg13g2_nor4_2 _5965_ (.A(_2185_),
    .B(_2186_),
    .C(_2201_),
    .Y(_2202_),
    .D(_2191_));
 sg13g2_xnor2_1 _5966_ (.Y(_2204_),
    .A(\clk_picker.counter[11] ),
    .B(_2202_));
 sg13g2_nor2_1 _5967_ (.A(_2204_),
    .B(net20),
    .Y(_0043_));
 sg13g2_inv_1 _5968_ (.Y(_2205_),
    .A(\clk_picker.counter[12] ));
 sg13g2_inv_2 _5969_ (.Y(_2206_),
    .A(_2194_));
 sg13g2_inv_1 _5970_ (.Y(_2207_),
    .A(\clk_picker.counter[11] ));
 sg13g2_nor4_1 _5971_ (.A(_2155_),
    .B(_2199_),
    .C(_2184_),
    .D(_2207_),
    .Y(_2208_));
 sg13g2_nand2_1 _5972_ (.Y(_2209_),
    .A(_2206_),
    .B(_2208_));
 sg13g2_xnor2_1 _5973_ (.Y(_2210_),
    .A(_2205_),
    .B(_2209_));
 sg13g2_nor2_1 _5974_ (.A(_2210_),
    .B(net20),
    .Y(_0044_));
 sg13g2_inv_1 _5975_ (.Y(_2211_),
    .A(\clk_picker.counter[13] ));
 sg13g2_nor4_1 _5976_ (.A(_2199_),
    .B(_2184_),
    .C(_2207_),
    .D(_2205_),
    .Y(_2213_));
 sg13g2_nand2_1 _5977_ (.Y(_2214_),
    .A(_2195_),
    .B(_2213_));
 sg13g2_xnor2_1 _5978_ (.Y(_2215_),
    .A(_2211_),
    .B(_2214_));
 sg13g2_nor2_1 _5979_ (.A(_2215_),
    .B(_2198_),
    .Y(_0045_));
 sg13g2_nor3_1 _5980_ (.A(_2184_),
    .B(_2207_),
    .C(_2158_),
    .Y(_2216_));
 sg13g2_inv_1 _5981_ (.Y(_2217_),
    .A(_2216_));
 sg13g2_nor2_1 _5982_ (.A(_2217_),
    .B(_2196_),
    .Y(_2218_));
 sg13g2_xnor2_1 _5983_ (.Y(_2219_),
    .A(\clk_picker.counter[14] ),
    .B(_2218_));
 sg13g2_nor2_1 _5984_ (.A(_2182_),
    .B(_2219_),
    .Y(_0046_));
 sg13g2_inv_1 _5985_ (.Y(_2220_),
    .A(\clk_picker.counter[15] ));
 sg13g2_inv_1 _5986_ (.Y(_2222_),
    .A(\clk_picker.counter[14] ));
 sg13g2_nor4_1 _5987_ (.A(_2207_),
    .B(_2205_),
    .C(_2211_),
    .D(_2222_),
    .Y(_2223_));
 sg13g2_nand2_1 _5988_ (.Y(_2224_),
    .A(_2202_),
    .B(_2223_));
 sg13g2_xnor2_1 _5989_ (.Y(_2225_),
    .A(_2220_),
    .B(_2224_));
 sg13g2_nor2_1 _5990_ (.A(_2225_),
    .B(net20),
    .Y(_0047_));
 sg13g2_nand2_1 _5991_ (.Y(_2226_),
    .A(_2159_),
    .B(_2161_));
 sg13g2_nor2_1 _5992_ (.A(_2226_),
    .B(_2209_),
    .Y(_2227_));
 sg13g2_xnor2_1 _5993_ (.Y(_2228_),
    .A(\clk_picker.counter[16] ),
    .B(_2227_));
 sg13g2_nor2_1 _5994_ (.A(_2228_),
    .B(net20),
    .Y(_0048_));
 sg13g2_inv_1 _5995_ (.Y(_2229_),
    .A(\clk_picker.counter[16] ));
 sg13g2_nor4_1 _5996_ (.A(_2211_),
    .B(_2222_),
    .C(_2220_),
    .D(_2229_),
    .Y(_2231_));
 sg13g2_nor2b_1 _5997_ (.A(_2214_),
    .B_N(_2231_),
    .Y(_2232_));
 sg13g2_xnor2_1 _5998_ (.Y(_2233_),
    .A(_2157_),
    .B(_2232_));
 sg13g2_nor2_1 _5999_ (.A(_2233_),
    .B(_2198_),
    .Y(_0049_));
 sg13g2_nor2_1 _6000_ (.A(_2165_),
    .B(_2160_),
    .Y(_2234_));
 sg13g2_nand2_1 _6001_ (.Y(_2235_),
    .A(_2218_),
    .B(_2234_));
 sg13g2_xnor2_1 _6002_ (.Y(_2236_),
    .A(_2164_),
    .B(_2235_));
 sg13g2_nor2_1 _6003_ (.A(net21),
    .B(_2236_),
    .Y(_0050_));
 sg13g2_inv_1 _6004_ (.Y(_2237_),
    .A(\clk_picker.counter[19] ));
 sg13g2_inv_1 _6005_ (.Y(_2238_),
    .A(_2157_));
 sg13g2_nor4_1 _6006_ (.A(_2220_),
    .B(_2229_),
    .C(_2238_),
    .D(_2164_),
    .Y(_2240_));
 sg13g2_nand3_1 _6007_ (.B(_2223_),
    .C(_2240_),
    .A(_2202_),
    .Y(_2241_));
 sg13g2_xnor2_1 _6008_ (.Y(_2242_),
    .A(_2237_),
    .B(_2241_));
 sg13g2_nor2_1 _6009_ (.A(_2242_),
    .B(net20),
    .Y(_0051_));
 sg13g2_inv_1 _6010_ (.Y(_2243_),
    .A(_2187_));
 sg13g2_nor2_1 _6011_ (.A(\clk_picker.counter[1] ),
    .B(\clk_picker.counter[0] ),
    .Y(_2244_));
 sg13g2_nor3_1 _6012_ (.A(_2243_),
    .B(_2244_),
    .C(net21),
    .Y(_0052_));
 sg13g2_nand2_1 _6013_ (.Y(_2245_),
    .A(\clk_picker.counter[18] ),
    .B(\clk_picker.counter[19] ));
 sg13g2_nor2_1 _6014_ (.A(_2165_),
    .B(_2245_),
    .Y(_2246_));
 sg13g2_nand2_1 _6015_ (.Y(_2247_),
    .A(_2227_),
    .B(_2246_));
 sg13g2_xnor2_1 _6016_ (.Y(_2249_),
    .A(_2167_),
    .B(_2247_));
 sg13g2_nor2_1 _6017_ (.A(net21),
    .B(_2249_),
    .Y(_0053_));
 sg13g2_inv_1 _6018_ (.Y(_2250_),
    .A(\clk_picker.counter[21] ));
 sg13g2_nor4_1 _6019_ (.A(_2238_),
    .B(_2164_),
    .C(_2237_),
    .D(_2167_),
    .Y(_2251_));
 sg13g2_nand2_1 _6020_ (.Y(_2252_),
    .A(_2232_),
    .B(_2251_));
 sg13g2_xnor2_1 _6021_ (.Y(_2253_),
    .A(_2250_),
    .B(_2252_));
 sg13g2_nor2_1 _6022_ (.A(net21),
    .B(_2253_),
    .Y(_0054_));
 sg13g2_nor2_1 _6023_ (.A(_2185_),
    .B(_2191_),
    .Y(_2254_));
 sg13g2_nor3_1 _6024_ (.A(_2167_),
    .B(_2250_),
    .C(_2245_),
    .Y(_2255_));
 sg13g2_nand4_1 _6025_ (.B(\clk_picker.counter[7] ),
    .C(\clk_picker.counter[8] ),
    .A(\clk_picker.counter[6] ),
    .Y(_2256_),
    .D(_2152_));
 sg13g2_nor2_1 _6026_ (.A(_2256_),
    .B(_2217_),
    .Y(_2258_));
 sg13g2_nand4_1 _6027_ (.B(_2255_),
    .C(_2258_),
    .A(_2254_),
    .Y(_2259_),
    .D(_2234_));
 sg13g2_xor2_1 _6028_ (.B(_2259_),
    .A(\clk_picker.counter[22] ),
    .X(_2260_));
 sg13g2_nor2_1 _6029_ (.A(_2260_),
    .B(net20),
    .Y(_0055_));
 sg13g2_nand2b_1 _6030_ (.Y(_2261_),
    .B(_2251_),
    .A_N(_2169_));
 sg13g2_nor4_1 _6031_ (.A(_2220_),
    .B(_2229_),
    .C(_2261_),
    .D(_2224_),
    .Y(_2262_));
 sg13g2_xnor2_1 _6032_ (.Y(_2263_),
    .A(\clk_picker.counter[23] ),
    .B(_2262_));
 sg13g2_nor2_1 _6033_ (.A(net21),
    .B(_2263_),
    .Y(_0056_));
 sg13g2_inv_1 _6034_ (.Y(_2264_),
    .A(\clk_picker.counter[24] ));
 sg13g2_nand3_1 _6035_ (.B(_2170_),
    .C(_2246_),
    .A(_2227_),
    .Y(_2265_));
 sg13g2_xnor2_1 _6036_ (.Y(_2267_),
    .A(_2264_),
    .B(_2265_));
 sg13g2_nor2_1 _6037_ (.A(_2182_),
    .B(_2267_),
    .Y(_0057_));
 sg13g2_nor3_1 _6038_ (.A(_2168_),
    .B(_2264_),
    .C(_2261_),
    .Y(_2268_));
 sg13g2_a21oi_1 _6039_ (.A1(_2232_),
    .A2(_2268_),
    .Y(_2269_),
    .B1(\clk_picker.counter[25] ));
 sg13g2_nor2_1 _6040_ (.A(_2269_),
    .B(net20),
    .Y(_0058_));
 sg13g2_nor2_1 _6041_ (.A(\clk_picker.counter[2] ),
    .B(_2243_),
    .Y(_2270_));
 sg13g2_nor3_1 _6042_ (.A(_2188_),
    .B(_2270_),
    .C(_2181_),
    .Y(_0059_));
 sg13g2_nor2_1 _6043_ (.A(\clk_picker.counter[3] ),
    .B(_2188_),
    .Y(_2271_));
 sg13g2_nor3_1 _6044_ (.A(_2190_),
    .B(_2271_),
    .C(_2181_),
    .Y(_0060_));
 sg13g2_xnor2_1 _6045_ (.Y(_2272_),
    .A(\clk_picker.counter[4] ),
    .B(_2190_));
 sg13g2_nor2_1 _6046_ (.A(_2272_),
    .B(net21),
    .Y(_0061_));
 sg13g2_a21oi_1 _6047_ (.A1(_2190_),
    .A2(\clk_picker.counter[4] ),
    .Y(_2274_),
    .B1(\clk_picker.counter[5] ));
 sg13g2_nor3_1 _6048_ (.A(_2254_),
    .B(_2274_),
    .C(_2181_),
    .Y(_0062_));
 sg13g2_nor2_1 _6049_ (.A(\clk_picker.counter[6] ),
    .B(_2254_),
    .Y(_2275_));
 sg13g2_nor3_1 _6050_ (.A(_2192_),
    .B(_2275_),
    .C(_2181_),
    .Y(_0063_));
 sg13g2_nor2_1 _6051_ (.A(\clk_picker.counter[7] ),
    .B(_2192_),
    .Y(_2276_));
 sg13g2_nor3_1 _6052_ (.A(_2206_),
    .B(_2276_),
    .C(_2181_),
    .Y(_0064_));
 sg13g2_nor2_1 _6053_ (.A(\clk_picker.counter[8] ),
    .B(_2206_),
    .Y(_2277_));
 sg13g2_nor3_1 _6054_ (.A(_2195_),
    .B(_2277_),
    .C(_2181_),
    .Y(_0065_));
 sg13g2_xnor2_1 _6055_ (.Y(_2278_),
    .A(_2152_),
    .B(_2195_));
 sg13g2_nor2_1 _6056_ (.A(_2278_),
    .B(net21),
    .Y(_0066_));
 sg13g2_nor2_1 _6057_ (.A(net2),
    .B(\transformer_1.started ),
    .Y(_2280_));
 sg13g2_buf_1 _6058_ (.A(_2280_),
    .X(_2281_));
 sg13g2_nor2_1 _6059_ (.A(_0031_),
    .B(net191),
    .Y(_2282_));
 sg13g2_nor3_1 _6060_ (.A(net2),
    .B(\transformer_1.started ),
    .C(\line_mapper_1.pointer_addr[10] ),
    .Y(_2283_));
 sg13g2_or2_1 _6061_ (.X(_2284_),
    .B(\chars_remaining[1] ),
    .A(\chars_remaining[2] ));
 sg13g2_nor2_1 _6062_ (.A(\chars_remaining[0] ),
    .B(_2284_),
    .Y(_2285_));
 sg13g2_inv_1 _6063_ (.Y(_2286_),
    .A(_2285_));
 sg13g2_nor4_2 _6064_ (.A(\chars_remaining[5] ),
    .B(\chars_remaining[4] ),
    .C(\chars_remaining[3] ),
    .Y(_2287_),
    .D(_2286_));
 sg13g2_nand2b_1 _6065_ (.Y(_2288_),
    .B(_2287_),
    .A_N(\chars_remaining[6] ));
 sg13g2_inv_1 _6066_ (.Y(_2290_),
    .A(\chars_remaining[8] ));
 sg13g2_nand2b_1 _6067_ (.Y(_2291_),
    .B(_2290_),
    .A_N(\chars_remaining[7] ));
 sg13g2_nor2_1 _6068_ (.A(\chars_remaining[9] ),
    .B(_2291_),
    .Y(_2292_));
 sg13g2_nor2b_1 _6069_ (.A(_2288_),
    .B_N(_2292_),
    .Y(_2293_));
 sg13g2_nor2b_1 _6070_ (.A(net191),
    .B_N(_2293_),
    .Y(_2294_));
 sg13g2_buf_1 _6071_ (.A(_2294_),
    .X(_2295_));
 sg13g2_nor4_1 _6072_ (.A(net211),
    .B(_2282_),
    .C(_2283_),
    .D(net19),
    .Y(_0067_));
 sg13g2_buf_1 _6073_ (.A(net191),
    .X(_2296_));
 sg13g2_xnor2_1 _6074_ (.Y(_2297_),
    .A(\chars_remaining[1] ),
    .B(\chars_remaining[0] ));
 sg13g2_nor2_1 _6075_ (.A(net191),
    .B(_2293_),
    .Y(_2298_));
 sg13g2_buf_2 _6076_ (.A(_2298_),
    .X(_2300_));
 sg13g2_buf_1 _6077_ (.A(_2300_),
    .X(_2301_));
 sg13g2_a22oi_1 _6078_ (.Y(_2302_),
    .B1(_2297_),
    .B2(net18),
    .A2(net159),
    .A1(\line_mapper_1.pointer_addr[11] ));
 sg13g2_nor2_1 _6079_ (.A(net211),
    .B(_2302_),
    .Y(_0068_));
 sg13g2_o21ai_1 _6080_ (.B1(\chars_remaining[2] ),
    .Y(_2303_),
    .A1(\chars_remaining[1] ),
    .A2(\chars_remaining[0] ));
 sg13g2_nand2_1 _6081_ (.Y(_2304_),
    .A(_2286_),
    .B(_2303_));
 sg13g2_a22oi_1 _6082_ (.Y(_2305_),
    .B1(_2304_),
    .B2(net18),
    .A2(net159),
    .A1(\line_mapper_1.pointer_addr[12] ));
 sg13g2_nor2_1 _6083_ (.A(net211),
    .B(_2305_),
    .Y(_0069_));
 sg13g2_nor2_1 _6084_ (.A(\chars_remaining[3] ),
    .B(_2286_),
    .Y(_2306_));
 sg13g2_nor2b_1 _6085_ (.A(_2285_),
    .B_N(\chars_remaining[3] ),
    .Y(_2307_));
 sg13g2_o21ai_1 _6086_ (.B1(_2300_),
    .Y(_2309_),
    .A1(_2306_),
    .A2(_2307_));
 sg13g2_nand2_1 _6087_ (.Y(_2310_),
    .A(net159),
    .B(\line_mapper_1.pointer_addr[13] ));
 sg13g2_a21oi_1 _6088_ (.A1(_2309_),
    .A2(_2310_),
    .Y(_0070_),
    .B1(net211));
 sg13g2_xor2_1 _6089_ (.B(_2306_),
    .A(\chars_remaining[4] ),
    .X(_2311_));
 sg13g2_a22oi_1 _6090_ (.Y(_2312_),
    .B1(_2311_),
    .B2(net18),
    .A2(net159),
    .A1(\line_mapper_1.pointer_addr[14] ));
 sg13g2_nor2_1 _6091_ (.A(net211),
    .B(_2312_),
    .Y(_0071_));
 sg13g2_nor3_1 _6092_ (.A(\chars_remaining[4] ),
    .B(\chars_remaining[3] ),
    .C(_2284_),
    .Y(_2313_));
 sg13g2_nand2_1 _6093_ (.Y(_2314_),
    .A(_2313_),
    .B(_0031_));
 sg13g2_xnor2_1 _6094_ (.Y(_2315_),
    .A(\chars_remaining[5] ),
    .B(_2314_));
 sg13g2_a22oi_1 _6095_ (.Y(_2316_),
    .B1(_2315_),
    .B2(net18),
    .A2(net159),
    .A1(\line_mapper_1.pointer_addr[15] ));
 sg13g2_nor2_1 _6096_ (.A(net211),
    .B(_2316_),
    .Y(_0072_));
 sg13g2_nor2_1 _6097_ (.A(_2178_),
    .B(net191),
    .Y(_2318_));
 sg13g2_inv_1 _6098_ (.Y(_2319_),
    .A(_2318_));
 sg13g2_xnor2_1 _6099_ (.Y(_2320_),
    .A(\chars_remaining[6] ),
    .B(_2287_));
 sg13g2_nor3_1 _6100_ (.A(_2319_),
    .B(_2293_),
    .C(_2320_),
    .Y(_0073_));
 sg13g2_or3_1 _6101_ (.A(\chars_remaining[7] ),
    .B(_2292_),
    .C(_2288_),
    .X(_2321_));
 sg13g2_buf_1 _6102_ (.A(_2321_),
    .X(_2322_));
 sg13g2_nand2_1 _6103_ (.Y(_2323_),
    .A(_2288_),
    .B(\chars_remaining[7] ));
 sg13g2_a21oi_1 _6104_ (.A1(_2322_),
    .A2(_2323_),
    .Y(_0074_),
    .B1(_2319_));
 sg13g2_o21ai_1 _6105_ (.B1(_2318_),
    .Y(_2324_),
    .A1(_2290_),
    .A2(_2322_));
 sg13g2_a21oi_1 _6106_ (.A1(_2290_),
    .A2(_2322_),
    .Y(_0075_),
    .B1(_2324_));
 sg13g2_inv_1 _6107_ (.Y(_2326_),
    .A(\chars_remaining[9] ));
 sg13g2_nor2_1 _6108_ (.A(_2291_),
    .B(_2288_),
    .Y(_2327_));
 sg13g2_nor3_1 _6109_ (.A(_2326_),
    .B(_2319_),
    .C(_2327_),
    .Y(_0076_));
 sg13g2_a22oi_1 _6110_ (.Y(_2328_),
    .B1(net185),
    .B2(net19),
    .A2(net159),
    .A1(\line_mapper_1.pointer_addr[0] ));
 sg13g2_a21oi_1 _6111_ (.A1(_2301_),
    .A2(_1162_),
    .Y(_2329_),
    .B1(_2179_));
 sg13g2_nand2_1 _6112_ (.Y(_0077_),
    .A(_2328_),
    .B(_2329_));
 sg13g2_a22oi_1 _6113_ (.Y(_2330_),
    .B1(net119),
    .B2(net19),
    .A2(_2300_),
    .A1(net47));
 sg13g2_a21oi_1 _6114_ (.A1(net159),
    .A2(\line_mapper_1.pointer_addr[1] ),
    .Y(_2331_),
    .B1(net211));
 sg13g2_nand2_1 _6115_ (.Y(_0078_),
    .A(_2330_),
    .B(_2331_));
 sg13g2_nand2_1 _6116_ (.Y(_2333_),
    .A(net19),
    .B(net153));
 sg13g2_nand2_1 _6117_ (.Y(_2334_),
    .A(net18),
    .B(_0258_));
 sg13g2_a21oi_1 _6118_ (.A1(_2296_),
    .A2(\line_mapper_1.pointer_addr[2] ),
    .Y(_2335_),
    .B1(_2178_));
 sg13g2_nand3_1 _6119_ (.B(_2334_),
    .C(_2335_),
    .A(_2333_),
    .Y(_0079_));
 sg13g2_nor2_1 _6120_ (.A(_1162_),
    .B(net87),
    .Y(_2336_));
 sg13g2_xnor2_1 _6121_ (.Y(_2337_),
    .A(net30),
    .B(_2336_));
 sg13g2_a22oi_1 _6122_ (.Y(_2338_),
    .B1(net33),
    .B2(net19),
    .A2(_2337_),
    .A1(_2300_));
 sg13g2_a21oi_1 _6123_ (.A1(_2296_),
    .A2(\line_mapper_1.pointer_addr[3] ),
    .Y(_2339_),
    .B1(_2178_));
 sg13g2_nand2_1 _6124_ (.Y(_0080_),
    .A(_2338_),
    .B(_2339_));
 sg13g2_nand2_1 _6125_ (.Y(_2340_),
    .A(net19),
    .B(net99));
 sg13g2_xnor2_1 _6126_ (.Y(_2342_),
    .A(net24),
    .B(_0598_));
 sg13g2_nand2_1 _6127_ (.Y(_2343_),
    .A(net18),
    .B(_2342_));
 sg13g2_a21oi_1 _6128_ (.A1(net191),
    .A2(\line_mapper_1.pointer_addr[4] ),
    .Y(_2344_),
    .B1(_2178_));
 sg13g2_nand3_1 _6129_ (.B(_2343_),
    .C(_2344_),
    .A(_2340_),
    .Y(_0081_));
 sg13g2_nor2_1 _6130_ (.A(_1998_),
    .B(_2020_),
    .Y(_2345_));
 sg13g2_inv_1 _6131_ (.Y(_2346_),
    .A(_2345_));
 sg13g2_nor2_1 _6132_ (.A(net75),
    .B(_2346_),
    .Y(_2347_));
 sg13g2_nand2_1 _6133_ (.Y(_2348_),
    .A(_2346_),
    .B(net46));
 sg13g2_nand3b_1 _6134_ (.B(_2300_),
    .C(_2348_),
    .Y(_2349_),
    .A_N(_2347_));
 sg13g2_nand2_1 _6135_ (.Y(_2350_),
    .A(_2295_),
    .B(net130));
 sg13g2_a21oi_1 _6136_ (.A1(net191),
    .A2(\line_mapper_1.pointer_addr[5] ),
    .Y(_2352_),
    .B1(_2178_));
 sg13g2_nand3_1 _6137_ (.B(_2350_),
    .C(_2352_),
    .A(_2349_),
    .Y(_0082_));
 sg13g2_nand2_1 _6138_ (.Y(_2353_),
    .A(_2295_),
    .B(net117));
 sg13g2_xnor2_1 _6139_ (.Y(_2354_),
    .A(net83),
    .B(_2347_));
 sg13g2_nand2_1 _6140_ (.Y(_2355_),
    .A(net18),
    .B(_2354_));
 sg13g2_a21oi_1 _6141_ (.A1(net191),
    .A2(\line_mapper_1.pointer_addr[6] ),
    .Y(_2356_),
    .B1(_2178_));
 sg13g2_nand3_1 _6142_ (.B(_2355_),
    .C(_2356_),
    .A(_2353_),
    .Y(_0083_));
 sg13g2_nand2_1 _6143_ (.Y(_2357_),
    .A(_1537_),
    .B(_2336_));
 sg13g2_xnor2_1 _6144_ (.Y(_2358_),
    .A(net164),
    .B(_2357_));
 sg13g2_a22oi_1 _6145_ (.Y(_2359_),
    .B1(net164),
    .B2(net19),
    .A2(_2358_),
    .A1(_2300_));
 sg13g2_a21oi_1 _6146_ (.A1(net159),
    .A2(\line_mapper_1.pointer_addr[7] ),
    .Y(_2361_),
    .B1(_2178_));
 sg13g2_nand2_1 _6147_ (.Y(_0084_),
    .A(_2359_),
    .B(_2361_));
 sg13g2_a22oi_1 _6148_ (.Y(_2362_),
    .B1(net200),
    .B2(net19),
    .A2(_2281_),
    .A1(\line_mapper_1.pointer_addr[8] ));
 sg13g2_nand2_1 _6149_ (.Y(_2363_),
    .A(_2347_),
    .B(_2559_));
 sg13g2_nor2_1 _6150_ (.A(net170),
    .B(_2363_),
    .Y(_2364_));
 sg13g2_nand2_1 _6151_ (.Y(_2365_),
    .A(_2363_),
    .B(net163));
 sg13g2_nand3b_1 _6152_ (.B(_2300_),
    .C(_2365_),
    .Y(_2366_),
    .A_N(_2364_));
 sg13g2_nand3_1 _6153_ (.B(_2177_),
    .C(_2366_),
    .A(_2362_),
    .Y(_0085_));
 sg13g2_a22oi_1 _6154_ (.Y(_2367_),
    .B1(net196),
    .B2(_2294_),
    .A2(_2281_),
    .A1(\line_mapper_1.pointer_addr[9] ));
 sg13g2_xnor2_1 _6155_ (.Y(_2368_),
    .A(net195),
    .B(_2364_));
 sg13g2_nand2_1 _6156_ (.Y(_2370_),
    .A(net18),
    .B(_2368_));
 sg13g2_nand3_1 _6157_ (.B(_2177_),
    .C(_2370_),
    .A(_2367_),
    .Y(_0086_));
 sg13g2_inv_1 _6158_ (.Y(_2371_),
    .A(\transformer_1.started ));
 sg13g2_a21oi_1 _6159_ (.A1(_2301_),
    .A2(_2371_),
    .Y(_0087_),
    .B1(net211));
 sg13g2_mux2_1 _6160_ (.A0(\clk_picker.clk_slow ),
    .A1(clknet_2_3__leaf_clk),
    .S(net3),
    .X(clk_buffered));
 sg13g2_buf_4 clkbuf_0_clk (.X(clknet_0_clk),
    .A(clk));
 sg13g2_tiehi _6163__221 (.L_HI(net221));
 sg13g2_buf_1 _6163_ (.A(net221),
    .X(uio_oe[0]));
 sg13g2_buf_1 _6164_ (.A(net222),
    .X(uio_oe[1]));
 sg13g2_buf_1 _6165_ (.A(net223),
    .X(uio_oe[2]));
 sg13g2_buf_1 _6166_ (.A(net224),
    .X(uio_oe[3]));
 sg13g2_buf_1 _6167_ (.A(net225),
    .X(uio_oe[4]));
 sg13g2_buf_1 _6168_ (.A(net226),
    .X(uio_oe[5]));
 sg13g2_buf_1 _6169_ (.A(net227),
    .X(uio_oe[6]));
 sg13g2_buf_1 _6170_ (.A(net228),
    .X(uio_oe[7]));
 sg13g2_buf_1 _6171_ (.A(net219),
    .X(uio_out[7]));
 sg13g2_buf_1 _6172_ (.A(net220),
    .X(uo_out[7]));
 sg13g2_dfrbp_1 \clk_picker.clk_slow$_SDFFE_PN0P_  (.CLK(clknet_level_2_1_38_clk),
    .RESET_B(net229),
    .D(_0040_),
    .Q_N(_0030_),
    .Q(\clk_picker.clk_slow ));
 sg13g2_dfrbp_1 \clk_picker.counter[0]$_SDFF_PN0_  (.CLK(clknet_level_2_1_12_clk),
    .RESET_B(net230),
    .D(_0041_),
    .Q_N(_0039_),
    .Q(\clk_picker.counter[0] ));
 sg13g2_dfrbp_1 \clk_picker.counter[10]$_SDFF_PN0_  (.CLK(clknet_level_2_1_25_clk),
    .RESET_B(net231),
    .D(_0042_),
    .Q_N(_3087_),
    .Q(\clk_picker.counter[10] ));
 sg13g2_dfrbp_1 \clk_picker.counter[11]$_SDFF_PN0_  (.CLK(clknet_level_2_1_25_clk),
    .RESET_B(net232),
    .D(_0043_),
    .Q_N(_3086_),
    .Q(\clk_picker.counter[11] ));
 sg13g2_dfrbp_1 \clk_picker.counter[12]$_SDFF_PN0_  (.CLK(clknet_level_2_1_38_clk),
    .RESET_B(net233),
    .D(_0044_),
    .Q_N(_3085_),
    .Q(\clk_picker.counter[12] ));
 sg13g2_dfrbp_1 \clk_picker.counter[13]$_SDFF_PN0_  (.CLK(clknet_level_2_1_411_clk),
    .RESET_B(net234),
    .D(_0045_),
    .Q_N(_3084_),
    .Q(\clk_picker.counter[13] ));
 sg13g2_dfrbp_1 \clk_picker.counter[14]$_SDFF_PN0_  (.CLK(clknet_level_2_1_38_clk),
    .RESET_B(net235),
    .D(_0046_),
    .Q_N(_3083_),
    .Q(\clk_picker.counter[14] ));
 sg13g2_dfrbp_1 \clk_picker.counter[15]$_SDFF_PN0_  (.CLK(clknet_level_2_1_411_clk),
    .RESET_B(net236),
    .D(_0047_),
    .Q_N(_3082_),
    .Q(\clk_picker.counter[15] ));
 sg13g2_dfrbp_1 \clk_picker.counter[16]$_SDFF_PN0_  (.CLK(clknet_level_2_1_411_clk),
    .RESET_B(net237),
    .D(_0048_),
    .Q_N(_3081_),
    .Q(\clk_picker.counter[16] ));
 sg13g2_dfrbp_1 \clk_picker.counter[17]$_SDFF_PN0_  (.CLK(clknet_level_2_1_411_clk),
    .RESET_B(net238),
    .D(_0049_),
    .Q_N(_3080_),
    .Q(\clk_picker.counter[17] ));
 sg13g2_dfrbp_1 \clk_picker.counter[18]$_SDFF_PN0_  (.CLK(clknet_level_2_1_38_clk),
    .RESET_B(net239),
    .D(_0050_),
    .Q_N(_3079_),
    .Q(\clk_picker.counter[18] ));
 sg13g2_dfrbp_1 \clk_picker.counter[19]$_SDFF_PN0_  (.CLK(clknet_level_2_1_411_clk),
    .RESET_B(net240),
    .D(_0051_),
    .Q_N(_3078_),
    .Q(\clk_picker.counter[19] ));
 sg13g2_dfrbp_1 \clk_picker.counter[1]$_SDFF_PN0_  (.CLK(clknet_level_2_1_12_clk),
    .RESET_B(net241),
    .D(_0052_),
    .Q_N(_3077_),
    .Q(\clk_picker.counter[1] ));
 sg13g2_dfrbp_1 \clk_picker.counter[20]$_SDFF_PN0_  (.CLK(clknet_level_2_1_38_clk),
    .RESET_B(net242),
    .D(_0053_),
    .Q_N(_3076_),
    .Q(\clk_picker.counter[20] ));
 sg13g2_dfrbp_1 \clk_picker.counter[21]$_SDFF_PN0_  (.CLK(clknet_level_2_1_25_clk),
    .RESET_B(net243),
    .D(_0054_),
    .Q_N(_3075_),
    .Q(\clk_picker.counter[21] ));
 sg13g2_dfrbp_1 \clk_picker.counter[22]$_SDFF_PN0_  (.CLK(clknet_level_2_1_25_clk),
    .RESET_B(net244),
    .D(_0055_),
    .Q_N(_3074_),
    .Q(\clk_picker.counter[22] ));
 sg13g2_dfrbp_1 \clk_picker.counter[23]$_SDFF_PN0_  (.CLK(clknet_level_2_1_38_clk),
    .RESET_B(net245),
    .D(_0056_),
    .Q_N(_3073_),
    .Q(\clk_picker.counter[23] ));
 sg13g2_dfrbp_1 \clk_picker.counter[24]$_SDFF_PN0_  (.CLK(clknet_level_2_1_38_clk),
    .RESET_B(net246),
    .D(_0057_),
    .Q_N(_3072_),
    .Q(\clk_picker.counter[24] ));
 sg13g2_dfrbp_1 \clk_picker.counter[25]$_SDFF_PN0_  (.CLK(clknet_level_2_1_411_clk),
    .RESET_B(net247),
    .D(_0058_),
    .Q_N(_3071_),
    .Q(\clk_picker.counter[25] ));
 sg13g2_dfrbp_1 \clk_picker.counter[2]$_SDFF_PN0_  (.CLK(clknet_level_2_1_25_clk),
    .RESET_B(net248),
    .D(_0059_),
    .Q_N(_3070_),
    .Q(\clk_picker.counter[2] ));
 sg13g2_dfrbp_1 \clk_picker.counter[3]$_SDFF_PN0_  (.CLK(clknet_level_2_1_25_clk),
    .RESET_B(net249),
    .D(_0060_),
    .Q_N(_3069_),
    .Q(\clk_picker.counter[3] ));
 sg13g2_dfrbp_1 \clk_picker.counter[4]$_SDFF_PN0_  (.CLK(clknet_level_2_1_12_clk),
    .RESET_B(net250),
    .D(_0061_),
    .Q_N(_3068_),
    .Q(\clk_picker.counter[4] ));
 sg13g2_dfrbp_1 \clk_picker.counter[5]$_SDFF_PN0_  (.CLK(clknet_level_2_1_12_clk),
    .RESET_B(net251),
    .D(_0062_),
    .Q_N(_3067_),
    .Q(\clk_picker.counter[5] ));
 sg13g2_dfrbp_1 \clk_picker.counter[6]$_SDFF_PN0_  (.CLK(clknet_level_2_1_12_clk),
    .RESET_B(net252),
    .D(_0063_),
    .Q_N(_3066_),
    .Q(\clk_picker.counter[6] ));
 sg13g2_dfrbp_1 \clk_picker.counter[7]$_SDFF_PN0_  (.CLK(clknet_level_2_1_12_clk),
    .RESET_B(net253),
    .D(_0064_),
    .Q_N(_3065_),
    .Q(\clk_picker.counter[7] ));
 sg13g2_dfrbp_1 \clk_picker.counter[8]$_SDFF_PN0_  (.CLK(clknet_level_2_1_25_clk),
    .RESET_B(net254),
    .D(_0065_),
    .Q_N(_3064_),
    .Q(\clk_picker.counter[8] ));
 sg13g2_dfrbp_1 \clk_picker.counter[9]$_SDFF_PN0_  (.CLK(clknet_level_2_1_12_clk),
    .RESET_B(net255),
    .D(_0066_),
    .Q_N(_3088_),
    .Q(\clk_picker.counter[9] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[0]$_DFF_P_  (.CLK(clknet_3_1__leaf_clk_buffered),
    .RESET_B(net256),
    .D(_0000_),
    .Q_N(_3089_),
    .Q(\line_mapper_1.pointer_addr[0] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[10]$_DFF_P_  (.CLK(clknet_3_1__leaf_clk_buffered),
    .RESET_B(net257),
    .D(_0001_),
    .Q_N(_3090_),
    .Q(\line_mapper_1.pointer_addr[10] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[11]$_DFF_P_  (.CLK(clknet_3_5__leaf_clk_buffered),
    .RESET_B(net258),
    .D(_0002_),
    .Q_N(_3091_),
    .Q(\line_mapper_1.pointer_addr[11] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[12]$_DFF_P_  (.CLK(clknet_3_0__leaf_clk_buffered),
    .RESET_B(net259),
    .D(_0003_),
    .Q_N(_3092_),
    .Q(\line_mapper_1.pointer_addr[12] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[13]$_DFF_P_  (.CLK(clknet_3_1__leaf_clk_buffered),
    .RESET_B(net260),
    .D(_0004_),
    .Q_N(_3093_),
    .Q(\line_mapper_1.pointer_addr[13] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[14]$_DFF_P_  (.CLK(clknet_3_1__leaf_clk_buffered),
    .RESET_B(net261),
    .D(_0005_),
    .Q_N(_3094_),
    .Q(\line_mapper_1.pointer_addr[14] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[15]$_DFF_P_  (.CLK(clknet_3_0__leaf_clk_buffered),
    .RESET_B(net262),
    .D(_0006_),
    .Q_N(_3095_),
    .Q(\line_mapper_1.pointer_addr[15] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[1]$_DFF_P_  (.CLK(clknet_3_4__leaf_clk_buffered),
    .RESET_B(net263),
    .D(_0007_),
    .Q_N(_3096_),
    .Q(\line_mapper_1.pointer_addr[1] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[2]$_DFF_P_  (.CLK(clknet_3_1__leaf_clk_buffered),
    .RESET_B(net264),
    .D(_0008_),
    .Q_N(_3097_),
    .Q(\line_mapper_1.pointer_addr[2] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[3]$_DFF_P_  (.CLK(clknet_3_0__leaf_clk_buffered),
    .RESET_B(net265),
    .D(_0009_),
    .Q_N(_3098_),
    .Q(\line_mapper_1.pointer_addr[3] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[4]$_DFF_P_  (.CLK(clknet_3_6__leaf_clk_buffered),
    .RESET_B(net266),
    .D(_0010_),
    .Q_N(_3099_),
    .Q(\line_mapper_1.pointer_addr[4] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[5]$_DFF_P_  (.CLK(clknet_3_4__leaf_clk_buffered),
    .RESET_B(net267),
    .D(_0011_),
    .Q_N(_3100_),
    .Q(\line_mapper_1.pointer_addr[5] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[6]$_DFF_P_  (.CLK(clknet_3_6__leaf_clk_buffered),
    .RESET_B(net268),
    .D(_0012_),
    .Q_N(_3101_),
    .Q(\line_mapper_1.pointer_addr[6] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[7]$_DFF_P_  (.CLK(clknet_3_1__leaf_clk_buffered),
    .RESET_B(net269),
    .D(_0013_),
    .Q_N(_3102_),
    .Q(\line_mapper_1.pointer_addr[7] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[8]$_DFF_P_  (.CLK(clknet_3_6__leaf_clk_buffered),
    .RESET_B(net270),
    .D(_0014_),
    .Q_N(_3103_),
    .Q(\line_mapper_1.pointer_addr[8] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[9]$_DFF_P_  (.CLK(clknet_3_4__leaf_clk_buffered),
    .RESET_B(net271),
    .D(_0015_),
    .Q_N(_3104_),
    .Q(\line_mapper_1.pointer_addr[9] ));
 sg13g2_dfrbp_1 \memory_1.dout[0]$_DFF_P_  (.CLK(clknet_3_7__leaf_clk_buffered),
    .RESET_B(net272),
    .D(_0016_),
    .Q_N(_3105_),
    .Q(net11));
 sg13g2_dfrbp_1 \memory_1.dout[10]$_DFF_P_  (.CLK(clknet_3_4__leaf_clk_buffered),
    .RESET_B(net273),
    .D(_0029_),
    .Q_N(_3106_),
    .Q(net6));
 sg13g2_dfrbp_1 \memory_1.dout[11]$_DFF_P_  (.CLK(clknet_3_5__leaf_clk_buffered),
    .RESET_B(net274),
    .D(_0017_),
    .Q_N(_3107_),
    .Q(net7));
 sg13g2_dfrbp_1 \memory_1.dout[12]$_DFF_P_  (.CLK(clknet_3_5__leaf_clk_buffered),
    .RESET_B(net275),
    .D(_0018_),
    .Q_N(_3108_),
    .Q(net8));
 sg13g2_dfrbp_1 \memory_1.dout[13]$_DFF_P_  (.CLK(clknet_3_5__leaf_clk_buffered),
    .RESET_B(net276),
    .D(_0019_),
    .Q_N(_3109_),
    .Q(net9));
 sg13g2_dfrbp_1 \memory_1.dout[14]$_DFF_P_  (.CLK(clknet_3_5__leaf_clk_buffered),
    .RESET_B(net277),
    .D(_0020_),
    .Q_N(_3110_),
    .Q(net10));
 sg13g2_dfrbp_1 \memory_1.dout[1]$_DFF_P_  (.CLK(clknet_3_4__leaf_clk_buffered),
    .RESET_B(net278),
    .D(_0021_),
    .Q_N(_3111_),
    .Q(net12));
 sg13g2_dfrbp_1 \memory_1.dout[2]$_DFF_P_  (.CLK(clknet_3_7__leaf_clk_buffered),
    .RESET_B(net279),
    .D(_0022_),
    .Q_N(_3112_),
    .Q(net13));
 sg13g2_dfrbp_1 \memory_1.dout[3]$_DFF_P_  (.CLK(clknet_3_7__leaf_clk_buffered),
    .RESET_B(net280),
    .D(_0023_),
    .Q_N(_3113_),
    .Q(net14));
 sg13g2_dfrbp_1 \memory_1.dout[4]$_DFF_P_  (.CLK(clknet_3_7__leaf_clk_buffered),
    .RESET_B(net281),
    .D(_0024_),
    .Q_N(_3114_),
    .Q(net15));
 sg13g2_dfrbp_1 \memory_1.dout[5]$_DFF_P_  (.CLK(clknet_3_7__leaf_clk_buffered),
    .RESET_B(net282),
    .D(_0025_),
    .Q_N(_3115_),
    .Q(net16));
 sg13g2_dfrbp_1 \memory_1.dout[6]$_DFF_P_  (.CLK(clknet_3_4__leaf_clk_buffered),
    .RESET_B(net283),
    .D(_0026_),
    .Q_N(_3116_),
    .Q(net17));
 sg13g2_dfrbp_1 \memory_1.dout[8]$_DFF_P_  (.CLK(clknet_3_4__leaf_clk_buffered),
    .RESET_B(net284),
    .D(_0027_),
    .Q_N(_3117_),
    .Q(net4));
 sg13g2_dfrbp_1 \memory_1.dout[9]$_DFF_P_  (.CLK(clknet_3_5__leaf_clk_buffered),
    .RESET_B(net285),
    .D(_0028_),
    .Q_N(_3063_),
    .Q(net5));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[0]$_SDFFE_PN0P_  (.CLK(clknet_3_3__leaf_clk_buffered),
    .RESET_B(net286),
    .D(_0067_),
    .Q_N(_0031_),
    .Q(\chars_remaining[0] ));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[1]$_SDFFE_PN0P_  (.CLK(clknet_3_0__leaf_clk_buffered),
    .RESET_B(net287),
    .D(_0068_),
    .Q_N(_3062_),
    .Q(\chars_remaining[1] ));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[2]$_SDFFE_PN0P_  (.CLK(clknet_3_0__leaf_clk_buffered),
    .RESET_B(net288),
    .D(_0069_),
    .Q_N(_3061_),
    .Q(\chars_remaining[2] ));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[3]$_SDFFE_PN0P_  (.CLK(clknet_3_2__leaf_clk_buffered),
    .RESET_B(net289),
    .D(_0070_),
    .Q_N(_3060_),
    .Q(\chars_remaining[3] ));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[4]$_SDFFE_PN0P_  (.CLK(clknet_3_0__leaf_clk_buffered),
    .RESET_B(net290),
    .D(_0071_),
    .Q_N(_3059_),
    .Q(\chars_remaining[4] ));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[5]$_SDFFE_PN0P_  (.CLK(clknet_3_0__leaf_clk_buffered),
    .RESET_B(net291),
    .D(_0072_),
    .Q_N(_3058_),
    .Q(\chars_remaining[5] ));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[6]$_SDFFE_PN0P_  (.CLK(clknet_3_2__leaf_clk_buffered),
    .RESET_B(net292),
    .D(_0073_),
    .Q_N(_3057_),
    .Q(\chars_remaining[6] ));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[7]$_SDFFE_PN0P_  (.CLK(clknet_3_2__leaf_clk_buffered),
    .RESET_B(net293),
    .D(_0074_),
    .Q_N(_3056_),
    .Q(\chars_remaining[7] ));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[8]$_SDFFE_PN0P_  (.CLK(clknet_3_2__leaf_clk_buffered),
    .RESET_B(net294),
    .D(_0075_),
    .Q_N(_3055_),
    .Q(\chars_remaining[8] ));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[9]$_SDFFE_PN0P_  (.CLK(clknet_3_2__leaf_clk_buffered),
    .RESET_B(net295),
    .D(_0076_),
    .Q_N(_3054_),
    .Q(\chars_remaining[9] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[0]$_SDFFE_PN1P_  (.CLK(clknet_3_3__leaf_clk_buffered),
    .RESET_B(net296),
    .D(_0077_),
    .Q_N(_0032_),
    .Q(\mem_addr[0] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[1]$_SDFFE_PN1P_  (.CLK(clknet_3_3__leaf_clk_buffered),
    .RESET_B(net297),
    .D(_0078_),
    .Q_N(_0038_),
    .Q(\mem_addr[1] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[2]$_SDFFE_PN1P_  (.CLK(clknet_3_3__leaf_clk_buffered),
    .RESET_B(net298),
    .D(_0079_),
    .Q_N(_0037_),
    .Q(\mem_addr[2] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[3]$_SDFFE_PN1P_  (.CLK(clknet_3_2__leaf_clk_buffered),
    .RESET_B(net299),
    .D(_0080_),
    .Q_N(_0036_),
    .Q(\mem_addr[3] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[4]$_SDFFE_PN1P_  (.CLK(clknet_3_7__leaf_clk_buffered),
    .RESET_B(net300),
    .D(_0081_),
    .Q_N(_0035_),
    .Q(\mem_addr[4] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[5]$_SDFFE_PN1P_  (.CLK(clknet_3_6__leaf_clk_buffered),
    .RESET_B(net301),
    .D(_0082_),
    .Q_N(_0034_),
    .Q(\mem_addr[5] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[6]$_SDFFE_PN1P_  (.CLK(clknet_3_6__leaf_clk_buffered),
    .RESET_B(net302),
    .D(_0083_),
    .Q_N(_0033_),
    .Q(\mem_addr[6] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[7]$_SDFFE_PN1P_  (.CLK(clknet_3_3__leaf_clk_buffered),
    .RESET_B(net303),
    .D(_0084_),
    .Q_N(_3053_),
    .Q(\mem_addr[7] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[8]$_SDFFE_PN1P_  (.CLK(clknet_3_3__leaf_clk_buffered),
    .RESET_B(net304),
    .D(_0085_),
    .Q_N(_3052_),
    .Q(\mem_addr[8] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[9]$_SDFFE_PN1P_  (.CLK(clknet_3_6__leaf_clk_buffered),
    .RESET_B(net305),
    .D(_0086_),
    .Q_N(_3051_),
    .Q(\memory_1.mem_addr[9] ));
 sg13g2_dfrbp_1 \transformer_1.started$_SDFFE_PN0P_  (.CLK(clknet_3_2__leaf_clk_buffered),
    .RESET_B(net306),
    .D(_0087_),
    .Q_N(_3050_),
    .Q(\transformer_1.started ));
 sg13g2_buf_1 input1 (.A(ui_in[5]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[6]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[7]),
    .X(net3));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uio_out[0]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uio_out[1]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_out[2]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[3]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[4]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[5]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[6]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[0]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[1]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[2]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[3]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[4]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[5]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[6]));
 sg13g2_buf_2 fanout18 (.A(_2301_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_2295_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_2198_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_2182_),
    .X(net21));
 sg13g2_buf_4 fanout22 (.X(net22),
    .A(_0521_));
 sg13g2_buf_2 fanout23 (.A(_0294_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_3023_),
    .X(net24));
 sg13g2_buf_4 fanout25 (.X(net25),
    .A(_2991_));
 sg13g2_buf_4 fanout26 (.X(net26),
    .A(_2968_));
 sg13g2_buf_2 fanout27 (.A(_2844_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_2774_),
    .X(net28));
 sg13g2_buf_4 fanout29 (.X(net29),
    .A(_2512_));
 sg13g2_buf_2 fanout30 (.A(_2416_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_2384_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0334_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0326_),
    .X(net33));
 sg13g2_buf_4 fanout34 (.X(net34),
    .A(_0181_));
 sg13g2_buf_2 fanout35 (.A(_0163_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0110_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_3022_),
    .X(net37));
 sg13g2_buf_4 fanout38 (.X(net38),
    .A(_2997_));
 sg13g2_buf_4 fanout39 (.X(net39),
    .A(_2990_));
 sg13g2_buf_2 fanout40 (.A(_2963_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_2905_),
    .X(net41));
 sg13g2_buf_4 fanout42 (.X(net42),
    .A(_2895_));
 sg13g2_buf_4 fanout43 (.X(net43),
    .A(_2795_));
 sg13g2_buf_4 fanout44 (.X(net44),
    .A(_2778_));
 sg13g2_buf_2 fanout45 (.A(_2753_),
    .X(net45));
 sg13g2_buf_4 fanout46 (.X(net46),
    .A(_2733_));
 sg13g2_buf_4 fanout47 (.X(net47),
    .A(_2684_));
 sg13g2_buf_2 fanout48 (.A(_2680_),
    .X(net48));
 sg13g2_buf_4 fanout49 (.X(net49),
    .A(_2615_));
 sg13g2_buf_4 fanout50 (.X(net50),
    .A(_2593_));
 sg13g2_buf_4 fanout51 (.X(net51),
    .A(_2589_));
 sg13g2_buf_2 fanout52 (.A(_2583_),
    .X(net52));
 sg13g2_buf_4 fanout53 (.X(net53),
    .A(_2569_));
 sg13g2_buf_2 fanout54 (.A(_2533_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_2510_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_2506_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_2503_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_2491_),
    .X(net58));
 sg13g2_buf_4 fanout59 (.X(net59),
    .A(_2475_));
 sg13g2_buf_4 fanout60 (.X(net60),
    .A(_2415_));
 sg13g2_buf_2 fanout61 (.A(_2408_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_2383_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_2375_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_1107_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_0532_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_0338_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_0161_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_0090_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_2935_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_2882_),
    .X(net70));
 sg13g2_buf_4 fanout71 (.X(net71),
    .A(_2860_));
 sg13g2_buf_2 fanout72 (.A(_2826_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_2785_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_2782_),
    .X(net74));
 sg13g2_buf_4 fanout75 (.X(net75),
    .A(_2732_));
 sg13g2_buf_2 fanout76 (.A(_2729_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_2728_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_2716_),
    .X(net78));
 sg13g2_buf_4 fanout79 (.X(net79),
    .A(_2711_));
 sg13g2_buf_2 fanout80 (.A(_2699_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_2689_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_2673_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_2665_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_2654_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_2649_),
    .X(net85));
 sg13g2_buf_4 fanout86 (.X(net86),
    .A(_2628_));
 sg13g2_buf_4 fanout87 (.X(net87),
    .A(_2603_));
 sg13g2_buf_2 fanout88 (.A(_2568_),
    .X(net88));
 sg13g2_buf_4 fanout89 (.X(net89),
    .A(_2518_));
 sg13g2_buf_4 fanout90 (.X(net90),
    .A(_2513_));
 sg13g2_buf_2 fanout91 (.A(_2509_),
    .X(net91));
 sg13g2_buf_4 fanout92 (.X(net92),
    .A(_2505_));
 sg13g2_buf_4 fanout93 (.X(net93),
    .A(_2490_));
 sg13g2_buf_4 fanout94 (.X(net94),
    .A(_2487_));
 sg13g2_buf_2 fanout95 (.A(_2458_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_2452_),
    .X(net96));
 sg13g2_buf_4 fanout97 (.X(net97),
    .A(_2449_));
 sg13g2_buf_4 fanout98 (.X(net98),
    .A(_2435_));
 sg13g2_buf_2 fanout99 (.A(_2419_),
    .X(net99));
 sg13g2_buf_4 fanout100 (.X(net100),
    .A(_2413_));
 sg13g2_buf_2 fanout101 (.A(_2407_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_2402_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_2387_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_2382_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_2053_),
    .X(net105));
 sg13g2_buf_4 fanout106 (.X(net106),
    .A(_1838_));
 sg13g2_buf_2 fanout107 (.A(_1707_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_1631_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_1522_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_1347_),
    .X(net110));
 sg13g2_buf_4 fanout111 (.X(net111),
    .A(_0856_));
 sg13g2_buf_2 fanout112 (.A(_0728_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_0511_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_0220_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_0165_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_3040_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_2957_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_2816_),
    .X(net118));
 sg13g2_buf_4 fanout119 (.X(net119),
    .A(_2808_));
 sg13g2_buf_2 fanout120 (.A(_2769_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_2749_),
    .X(net121));
 sg13g2_buf_4 fanout122 (.X(net122),
    .A(_2704_));
 sg13g2_buf_2 fanout123 (.A(_2698_),
    .X(net123));
 sg13g2_buf_4 fanout124 (.X(net124),
    .A(_2688_));
 sg13g2_buf_4 fanout125 (.X(net125),
    .A(_2682_));
 sg13g2_buf_4 fanout126 (.X(net126),
    .A(_2669_));
 sg13g2_buf_2 fanout127 (.A(_2664_),
    .X(net127));
 sg13g2_buf_4 fanout128 (.X(net128),
    .A(_2653_));
 sg13g2_buf_2 fanout129 (.A(_2626_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_2601_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_2596_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_2566_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_2554_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_2552_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_2508_),
    .X(net135));
 sg13g2_buf_4 fanout136 (.X(net136),
    .A(_2495_));
 sg13g2_buf_2 fanout137 (.A(_2477_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_2445_),
    .X(net138));
 sg13g2_buf_4 fanout139 (.X(net139),
    .A(_2442_));
 sg13g2_buf_2 fanout140 (.A(_2437_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_2426_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_2418_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_2401_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_2399_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_2390_),
    .X(net145));
 sg13g2_buf_4 fanout146 (.X(net146),
    .A(_2386_));
 sg13g2_buf_2 fanout147 (.A(_2360_),
    .X(net147));
 sg13g2_buf_4 fanout148 (.X(net148),
    .A(_2257_));
 sg13g2_buf_2 fanout149 (.A(_2173_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_1696_),
    .X(net150));
 sg13g2_buf_4 fanout151 (.X(net151),
    .A(_1555_));
 sg13g2_buf_2 fanout152 (.A(_1511_),
    .X(net152));
 sg13g2_buf_4 fanout153 (.X(net153),
    .A(_1435_));
 sg13g2_buf_4 fanout154 (.X(net154),
    .A(_1020_));
 sg13g2_buf_4 fanout155 (.X(net155),
    .A(_0976_));
 sg13g2_buf_2 fanout156 (.A(_0910_),
    .X(net156));
 sg13g2_buf_4 fanout157 (.X(net157),
    .A(_0845_));
 sg13g2_buf_4 fanout158 (.X(net158),
    .A(_0757_));
 sg13g2_buf_2 fanout159 (.A(_2296_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_0483_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_3039_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_2760_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_2738_),
    .X(net163));
 sg13g2_buf_4 fanout164 (.X(net164),
    .A(_2736_));
 sg13g2_buf_2 fanout165 (.A(_2696_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_2646_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_2619_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_2600_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_2595_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_2565_),
    .X(net170));
 sg13g2_buf_4 fanout171 (.X(net171),
    .A(_2544_));
 sg13g2_buf_2 fanout172 (.A(_2517_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_2480_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_2417_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_2351_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_2193_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_2162_),
    .X(net177));
 sg13g2_buf_4 fanout178 (.X(net178),
    .A(_1773_));
 sg13g2_buf_4 fanout179 (.X(net179),
    .A(_1751_));
 sg13g2_buf_2 fanout180 (.A(_1685_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_1588_),
    .X(net181));
 sg13g2_buf_4 fanout182 (.X(net182),
    .A(_1544_));
 sg13g2_buf_2 fanout183 (.A(_1424_),
    .X(net183));
 sg13g2_buf_4 fanout184 (.X(net184),
    .A(_1282_));
 sg13g2_buf_4 fanout185 (.X(net185),
    .A(_1260_));
 sg13g2_buf_2 fanout186 (.A(_1249_),
    .X(net186));
 sg13g2_buf_4 fanout187 (.X(net187),
    .A(_1009_));
 sg13g2_buf_4 fanout188 (.X(net188),
    .A(_0834_));
 sg13g2_buf_2 fanout189 (.A(_0790_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_0746_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_2281_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_1837_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_0602_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_0530_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_2695_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_2610_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_2557_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_2543_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_2516_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_2424_),
    .X(net200));
 sg13g2_buf_4 fanout201 (.X(net201),
    .A(_1848_));
 sg13g2_buf_4 fanout202 (.X(net202),
    .A(_1740_));
 sg13g2_buf_4 fanout203 (.X(net203),
    .A(_1380_));
 sg13g2_buf_2 fanout204 (.A(_1205_),
    .X(net204));
 sg13g2_buf_4 fanout205 (.X(net205),
    .A(_0998_));
 sg13g2_buf_4 fanout206 (.X(net206),
    .A(_0943_));
 sg13g2_buf_2 fanout207 (.A(_0889_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_0867_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_1369_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_1053_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_2179_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_1867_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_1850_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_1810_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_1808_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_1801_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_1798_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_1796_),
    .X(net218));
 sg13g2_tielo _6171__219 (.L_LO(net219));
 sg13g2_tielo _6172__220 (.L_LO(net220));
 sg13g2_tiehi _6164__222 (.L_HI(net222));
 sg13g2_tiehi _6165__223 (.L_HI(net223));
 sg13g2_tiehi _6166__224 (.L_HI(net224));
 sg13g2_tiehi _6167__225 (.L_HI(net225));
 sg13g2_tiehi _6168__226 (.L_HI(net226));
 sg13g2_tiehi _6169__227 (.L_HI(net227));
 sg13g2_tiehi _6170__228 (.L_HI(net228));
 sg13g2_tiehi \clk_picker.clk_slow$_SDFFE_PN0P__229  (.L_HI(net229));
 sg13g2_tiehi \clk_picker.counter[0]$_SDFF_PN0__230  (.L_HI(net230));
 sg13g2_tiehi \clk_picker.counter[10]$_SDFF_PN0__231  (.L_HI(net231));
 sg13g2_tiehi \clk_picker.counter[11]$_SDFF_PN0__232  (.L_HI(net232));
 sg13g2_tiehi \clk_picker.counter[12]$_SDFF_PN0__233  (.L_HI(net233));
 sg13g2_tiehi \clk_picker.counter[13]$_SDFF_PN0__234  (.L_HI(net234));
 sg13g2_tiehi \clk_picker.counter[14]$_SDFF_PN0__235  (.L_HI(net235));
 sg13g2_tiehi \clk_picker.counter[15]$_SDFF_PN0__236  (.L_HI(net236));
 sg13g2_tiehi \clk_picker.counter[16]$_SDFF_PN0__237  (.L_HI(net237));
 sg13g2_tiehi \clk_picker.counter[17]$_SDFF_PN0__238  (.L_HI(net238));
 sg13g2_tiehi \clk_picker.counter[18]$_SDFF_PN0__239  (.L_HI(net239));
 sg13g2_tiehi \clk_picker.counter[19]$_SDFF_PN0__240  (.L_HI(net240));
 sg13g2_tiehi \clk_picker.counter[1]$_SDFF_PN0__241  (.L_HI(net241));
 sg13g2_tiehi \clk_picker.counter[20]$_SDFF_PN0__242  (.L_HI(net242));
 sg13g2_tiehi \clk_picker.counter[21]$_SDFF_PN0__243  (.L_HI(net243));
 sg13g2_tiehi \clk_picker.counter[22]$_SDFF_PN0__244  (.L_HI(net244));
 sg13g2_tiehi \clk_picker.counter[23]$_SDFF_PN0__245  (.L_HI(net245));
 sg13g2_tiehi \clk_picker.counter[24]$_SDFF_PN0__246  (.L_HI(net246));
 sg13g2_tiehi \clk_picker.counter[25]$_SDFF_PN0__247  (.L_HI(net247));
 sg13g2_tiehi \clk_picker.counter[2]$_SDFF_PN0__248  (.L_HI(net248));
 sg13g2_tiehi \clk_picker.counter[3]$_SDFF_PN0__249  (.L_HI(net249));
 sg13g2_tiehi \clk_picker.counter[4]$_SDFF_PN0__250  (.L_HI(net250));
 sg13g2_tiehi \clk_picker.counter[5]$_SDFF_PN0__251  (.L_HI(net251));
 sg13g2_tiehi \clk_picker.counter[6]$_SDFF_PN0__252  (.L_HI(net252));
 sg13g2_tiehi \clk_picker.counter[7]$_SDFF_PN0__253  (.L_HI(net253));
 sg13g2_tiehi \clk_picker.counter[8]$_SDFF_PN0__254  (.L_HI(net254));
 sg13g2_tiehi \clk_picker.counter[9]$_SDFF_PN0__255  (.L_HI(net255));
 sg13g2_tiehi \line_mapper_1.pointer_addr[0]$_DFF_P__256  (.L_HI(net256));
 sg13g2_tiehi \line_mapper_1.pointer_addr[10]$_DFF_P__257  (.L_HI(net257));
 sg13g2_tiehi \line_mapper_1.pointer_addr[11]$_DFF_P__258  (.L_HI(net258));
 sg13g2_tiehi \line_mapper_1.pointer_addr[12]$_DFF_P__259  (.L_HI(net259));
 sg13g2_tiehi \line_mapper_1.pointer_addr[13]$_DFF_P__260  (.L_HI(net260));
 sg13g2_tiehi \line_mapper_1.pointer_addr[14]$_DFF_P__261  (.L_HI(net261));
 sg13g2_tiehi \line_mapper_1.pointer_addr[15]$_DFF_P__262  (.L_HI(net262));
 sg13g2_tiehi \line_mapper_1.pointer_addr[1]$_DFF_P__263  (.L_HI(net263));
 sg13g2_tiehi \line_mapper_1.pointer_addr[2]$_DFF_P__264  (.L_HI(net264));
 sg13g2_tiehi \line_mapper_1.pointer_addr[3]$_DFF_P__265  (.L_HI(net265));
 sg13g2_tiehi \line_mapper_1.pointer_addr[4]$_DFF_P__266  (.L_HI(net266));
 sg13g2_tiehi \line_mapper_1.pointer_addr[5]$_DFF_P__267  (.L_HI(net267));
 sg13g2_tiehi \line_mapper_1.pointer_addr[6]$_DFF_P__268  (.L_HI(net268));
 sg13g2_tiehi \line_mapper_1.pointer_addr[7]$_DFF_P__269  (.L_HI(net269));
 sg13g2_tiehi \line_mapper_1.pointer_addr[8]$_DFF_P__270  (.L_HI(net270));
 sg13g2_tiehi \line_mapper_1.pointer_addr[9]$_DFF_P__271  (.L_HI(net271));
 sg13g2_tiehi \memory_1.dout[0]$_DFF_P__272  (.L_HI(net272));
 sg13g2_tiehi \memory_1.dout[10]$_DFF_P__273  (.L_HI(net273));
 sg13g2_tiehi \memory_1.dout[11]$_DFF_P__274  (.L_HI(net274));
 sg13g2_tiehi \memory_1.dout[12]$_DFF_P__275  (.L_HI(net275));
 sg13g2_tiehi \memory_1.dout[13]$_DFF_P__276  (.L_HI(net276));
 sg13g2_tiehi \memory_1.dout[14]$_DFF_P__277  (.L_HI(net277));
 sg13g2_tiehi \memory_1.dout[1]$_DFF_P__278  (.L_HI(net278));
 sg13g2_tiehi \memory_1.dout[2]$_DFF_P__279  (.L_HI(net279));
 sg13g2_tiehi \memory_1.dout[3]$_DFF_P__280  (.L_HI(net280));
 sg13g2_tiehi \memory_1.dout[4]$_DFF_P__281  (.L_HI(net281));
 sg13g2_tiehi \memory_1.dout[5]$_DFF_P__282  (.L_HI(net282));
 sg13g2_tiehi \memory_1.dout[6]$_DFF_P__283  (.L_HI(net283));
 sg13g2_tiehi \memory_1.dout[8]$_DFF_P__284  (.L_HI(net284));
 sg13g2_tiehi \memory_1.dout[9]$_DFF_P__285  (.L_HI(net285));
 sg13g2_tiehi \transformer_1.chars_remaining[0]$_SDFFE_PN0P__286  (.L_HI(net286));
 sg13g2_tiehi \transformer_1.chars_remaining[1]$_SDFFE_PN0P__287  (.L_HI(net287));
 sg13g2_tiehi \transformer_1.chars_remaining[2]$_SDFFE_PN0P__288  (.L_HI(net288));
 sg13g2_tiehi \transformer_1.chars_remaining[3]$_SDFFE_PN0P__289  (.L_HI(net289));
 sg13g2_tiehi \transformer_1.chars_remaining[4]$_SDFFE_PN0P__290  (.L_HI(net290));
 sg13g2_tiehi \transformer_1.chars_remaining[5]$_SDFFE_PN0P__291  (.L_HI(net291));
 sg13g2_tiehi \transformer_1.chars_remaining[6]$_SDFFE_PN0P__292  (.L_HI(net292));
 sg13g2_tiehi \transformer_1.chars_remaining[7]$_SDFFE_PN0P__293  (.L_HI(net293));
 sg13g2_tiehi \transformer_1.chars_remaining[8]$_SDFFE_PN0P__294  (.L_HI(net294));
 sg13g2_tiehi \transformer_1.chars_remaining[9]$_SDFFE_PN0P__295  (.L_HI(net295));
 sg13g2_tiehi \transformer_1.mem_addr[0]$_SDFFE_PN1P__296  (.L_HI(net296));
 sg13g2_tiehi \transformer_1.mem_addr[1]$_SDFFE_PN1P__297  (.L_HI(net297));
 sg13g2_tiehi \transformer_1.mem_addr[2]$_SDFFE_PN1P__298  (.L_HI(net298));
 sg13g2_tiehi \transformer_1.mem_addr[3]$_SDFFE_PN1P__299  (.L_HI(net299));
 sg13g2_tiehi \transformer_1.mem_addr[4]$_SDFFE_PN1P__300  (.L_HI(net300));
 sg13g2_tiehi \transformer_1.mem_addr[5]$_SDFFE_PN1P__301  (.L_HI(net301));
 sg13g2_tiehi \transformer_1.mem_addr[6]$_SDFFE_PN1P__302  (.L_HI(net302));
 sg13g2_tiehi \transformer_1.mem_addr[7]$_SDFFE_PN1P__303  (.L_HI(net303));
 sg13g2_tiehi \transformer_1.mem_addr[8]$_SDFFE_PN1P__304  (.L_HI(net304));
 sg13g2_tiehi \transformer_1.mem_addr[9]$_SDFFE_PN1P__305  (.L_HI(net305));
 sg13g2_tiehi \transformer_1.started$_SDFFE_PN0P__306  (.L_HI(net306));
 sg13g2_buf_4 clkbuf_2_0__f_clk (.X(clknet_2_0__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_2_1__f_clk (.X(clknet_2_1__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_2_2__f_clk (.X(clknet_2_2__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_2_3__f_clk (.X(clknet_2_3__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_buf_8 clkbuf_level_0_1_10_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_level_0_1_10_clk));
 sg13g2_buf_8 clkbuf_level_1_1_11_clk (.A(clknet_level_0_1_10_clk),
    .X(clknet_level_1_1_11_clk));
 sg13g2_buf_8 clkbuf_level_2_1_12_clk (.A(clknet_level_1_1_11_clk),
    .X(clknet_level_2_1_12_clk));
 sg13g2_buf_8 clkbuf_level_0_1_23_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_level_0_1_23_clk));
 sg13g2_buf_8 clkbuf_level_1_1_24_clk (.A(clknet_level_0_1_23_clk),
    .X(clknet_level_1_1_24_clk));
 sg13g2_buf_8 clkbuf_level_2_1_25_clk (.A(clknet_level_1_1_24_clk),
    .X(clknet_level_2_1_25_clk));
 sg13g2_buf_8 clkbuf_level_0_1_36_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_level_0_1_36_clk));
 sg13g2_buf_8 clkbuf_level_1_1_37_clk (.A(clknet_level_0_1_36_clk),
    .X(clknet_level_1_1_37_clk));
 sg13g2_buf_8 clkbuf_level_2_1_38_clk (.A(clknet_level_1_1_37_clk),
    .X(clknet_level_2_1_38_clk));
 sg13g2_buf_8 clkbuf_level_0_1_49_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_level_0_1_49_clk));
 sg13g2_buf_8 clkbuf_level_1_1_410_clk (.A(clknet_level_0_1_49_clk),
    .X(clknet_level_1_1_410_clk));
 sg13g2_buf_8 clkbuf_level_2_1_411_clk (.A(clknet_level_1_1_410_clk),
    .X(clknet_level_2_1_411_clk));
 sg13g2_buf_4 clkload0 (.A(clknet_2_0__leaf_clk));
 sg13g2_buf_4 clkload1 (.A(clknet_2_1__leaf_clk));
 sg13g2_buf_4 clkload2 (.A(clknet_2_2__leaf_clk));
 sg13g2_buf_4 clkbuf_0_clk_buffered (.X(clknet_0_clk_buffered),
    .A(clk_buffered));
 sg13g2_buf_4 clkbuf_3_0__f_clk_buffered (.X(clknet_3_0__leaf_clk_buffered),
    .A(clknet_0_clk_buffered));
 sg13g2_buf_4 clkbuf_3_1__f_clk_buffered (.X(clknet_3_1__leaf_clk_buffered),
    .A(clknet_0_clk_buffered));
 sg13g2_buf_4 clkbuf_3_2__f_clk_buffered (.X(clknet_3_2__leaf_clk_buffered),
    .A(clknet_0_clk_buffered));
 sg13g2_buf_4 clkbuf_3_3__f_clk_buffered (.X(clknet_3_3__leaf_clk_buffered),
    .A(clknet_0_clk_buffered));
 sg13g2_buf_4 clkbuf_3_4__f_clk_buffered (.X(clknet_3_4__leaf_clk_buffered),
    .A(clknet_0_clk_buffered));
 sg13g2_buf_4 clkbuf_3_5__f_clk_buffered (.X(clknet_3_5__leaf_clk_buffered),
    .A(clknet_0_clk_buffered));
 sg13g2_buf_4 clkbuf_3_6__f_clk_buffered (.X(clknet_3_6__leaf_clk_buffered),
    .A(clknet_0_clk_buffered));
 sg13g2_buf_4 clkbuf_3_7__f_clk_buffered (.X(clknet_3_7__leaf_clk_buffered),
    .A(clknet_0_clk_buffered));
 sg13g2_inv_1 clkload3 (.A(clknet_3_1__leaf_clk_buffered));
 sg13g2_inv_1 clkload4 (.A(clknet_3_3__leaf_clk_buffered));
 sg13g2_inv_1 clkload5 (.A(clknet_3_5__leaf_clk_buffered));
 sg13g2_inv_1 clkload6 (.A(clknet_3_6__leaf_clk_buffered));
 sg13g2_inv_1 clkload7 (.A(clknet_3_7__leaf_clk_buffered));
 sg13g2_antennanp ANTENNA_1 (.A(_0003_));
 sg13g2_antennanp ANTENNA_2 (.A(_0016_));
 sg13g2_antennanp ANTENNA_3 (.A(_0018_));
 sg13g2_antennanp ANTENNA_4 (.A(_0018_));
 sg13g2_antennanp ANTENNA_5 (.A(_0021_));
 sg13g2_antennanp ANTENNA_6 (.A(_0022_));
 sg13g2_antennanp ANTENNA_7 (.A(_0023_));
 sg13g2_antennanp ANTENNA_8 (.A(_0024_));
 sg13g2_antennanp ANTENNA_9 (.A(_0025_));
 sg13g2_antennanp ANTENNA_10 (.A(_0025_));
 sg13g2_antennanp ANTENNA_11 (.A(_0026_));
 sg13g2_antennanp ANTENNA_12 (.A(_0026_));
 sg13g2_antennanp ANTENNA_13 (.A(_0027_));
 sg13g2_antennanp ANTENNA_14 (.A(_0027_));
 sg13g2_antennanp ANTENNA_15 (.A(_0028_));
 sg13g2_antennanp ANTENNA_16 (.A(_0028_));
 sg13g2_antennanp ANTENNA_17 (.A(_0038_));
 sg13g2_antennanp ANTENNA_18 (.A(_0038_));
 sg13g2_antennanp ANTENNA_19 (.A(_0038_));
 sg13g2_antennanp ANTENNA_20 (.A(_0038_));
 sg13g2_antennanp ANTENNA_21 (.A(_0038_));
 sg13g2_antennanp ANTENNA_22 (.A(_0038_));
 sg13g2_antennanp ANTENNA_23 (.A(_0038_));
 sg13g2_antennanp ANTENNA_24 (.A(_0038_));
 sg13g2_antennanp ANTENNA_25 (.A(_0038_));
 sg13g2_antennanp ANTENNA_26 (.A(_0090_));
 sg13g2_antennanp ANTENNA_27 (.A(_0090_));
 sg13g2_antennanp ANTENNA_28 (.A(_0090_));
 sg13g2_antennanp ANTENNA_29 (.A(_0100_));
 sg13g2_antennanp ANTENNA_30 (.A(_0100_));
 sg13g2_antennanp ANTENNA_31 (.A(_0100_));
 sg13g2_antennanp ANTENNA_32 (.A(_0100_));
 sg13g2_antennanp ANTENNA_33 (.A(_0100_));
 sg13g2_antennanp ANTENNA_34 (.A(_0123_));
 sg13g2_antennanp ANTENNA_35 (.A(_0123_));
 sg13g2_antennanp ANTENNA_36 (.A(_0125_));
 sg13g2_antennanp ANTENNA_37 (.A(_0125_));
 sg13g2_antennanp ANTENNA_38 (.A(_0125_));
 sg13g2_antennanp ANTENNA_39 (.A(_0150_));
 sg13g2_antennanp ANTENNA_40 (.A(_0150_));
 sg13g2_antennanp ANTENNA_41 (.A(_0150_));
 sg13g2_antennanp ANTENNA_42 (.A(_0150_));
 sg13g2_antennanp ANTENNA_43 (.A(_0150_));
 sg13g2_antennanp ANTENNA_44 (.A(_0150_));
 sg13g2_antennanp ANTENNA_45 (.A(_0150_));
 sg13g2_antennanp ANTENNA_46 (.A(_0150_));
 sg13g2_antennanp ANTENNA_47 (.A(_0150_));
 sg13g2_antennanp ANTENNA_48 (.A(_0158_));
 sg13g2_antennanp ANTENNA_49 (.A(_0160_));
 sg13g2_antennanp ANTENNA_50 (.A(_0160_));
 sg13g2_antennanp ANTENNA_51 (.A(_0160_));
 sg13g2_antennanp ANTENNA_52 (.A(_0160_));
 sg13g2_antennanp ANTENNA_53 (.A(_0165_));
 sg13g2_antennanp ANTENNA_54 (.A(_0165_));
 sg13g2_antennanp ANTENNA_55 (.A(_0165_));
 sg13g2_antennanp ANTENNA_56 (.A(_0167_));
 sg13g2_antennanp ANTENNA_57 (.A(_0167_));
 sg13g2_antennanp ANTENNA_58 (.A(_0167_));
 sg13g2_antennanp ANTENNA_59 (.A(_0167_));
 sg13g2_antennanp ANTENNA_60 (.A(_0167_));
 sg13g2_antennanp ANTENNA_61 (.A(_0167_));
 sg13g2_antennanp ANTENNA_62 (.A(_0167_));
 sg13g2_antennanp ANTENNA_63 (.A(_0167_));
 sg13g2_antennanp ANTENNA_64 (.A(_0168_));
 sg13g2_antennanp ANTENNA_65 (.A(_0168_));
 sg13g2_antennanp ANTENNA_66 (.A(_0168_));
 sg13g2_antennanp ANTENNA_67 (.A(_0168_));
 sg13g2_antennanp ANTENNA_68 (.A(_0168_));
 sg13g2_antennanp ANTENNA_69 (.A(_0168_));
 sg13g2_antennanp ANTENNA_70 (.A(_0189_));
 sg13g2_antennanp ANTENNA_71 (.A(_0230_));
 sg13g2_antennanp ANTENNA_72 (.A(_0234_));
 sg13g2_antennanp ANTENNA_73 (.A(_0234_));
 sg13g2_antennanp ANTENNA_74 (.A(_0234_));
 sg13g2_antennanp ANTENNA_75 (.A(_0234_));
 sg13g2_antennanp ANTENNA_76 (.A(_0234_));
 sg13g2_antennanp ANTENNA_77 (.A(_0234_));
 sg13g2_antennanp ANTENNA_78 (.A(_0234_));
 sg13g2_antennanp ANTENNA_79 (.A(_0234_));
 sg13g2_antennanp ANTENNA_80 (.A(_0234_));
 sg13g2_antennanp ANTENNA_81 (.A(_0234_));
 sg13g2_antennanp ANTENNA_82 (.A(_0234_));
 sg13g2_antennanp ANTENNA_83 (.A(_0234_));
 sg13g2_antennanp ANTENNA_84 (.A(_0234_));
 sg13g2_antennanp ANTENNA_85 (.A(_0234_));
 sg13g2_antennanp ANTENNA_86 (.A(_0234_));
 sg13g2_antennanp ANTENNA_87 (.A(_0250_));
 sg13g2_antennanp ANTENNA_88 (.A(_0250_));
 sg13g2_antennanp ANTENNA_89 (.A(_0250_));
 sg13g2_antennanp ANTENNA_90 (.A(_0250_));
 sg13g2_antennanp ANTENNA_91 (.A(_0250_));
 sg13g2_antennanp ANTENNA_92 (.A(_0260_));
 sg13g2_antennanp ANTENNA_93 (.A(_0260_));
 sg13g2_antennanp ANTENNA_94 (.A(_0260_));
 sg13g2_antennanp ANTENNA_95 (.A(_0260_));
 sg13g2_antennanp ANTENNA_96 (.A(_0269_));
 sg13g2_antennanp ANTENNA_97 (.A(_0301_));
 sg13g2_antennanp ANTENNA_98 (.A(_0345_));
 sg13g2_antennanp ANTENNA_99 (.A(_0345_));
 sg13g2_antennanp ANTENNA_100 (.A(_0345_));
 sg13g2_antennanp ANTENNA_101 (.A(_0345_));
 sg13g2_antennanp ANTENNA_102 (.A(_0346_));
 sg13g2_antennanp ANTENNA_103 (.A(_0346_));
 sg13g2_antennanp ANTENNA_104 (.A(_0346_));
 sg13g2_antennanp ANTENNA_105 (.A(_0346_));
 sg13g2_antennanp ANTENNA_106 (.A(_0360_));
 sg13g2_antennanp ANTENNA_107 (.A(_0360_));
 sg13g2_antennanp ANTENNA_108 (.A(_0360_));
 sg13g2_antennanp ANTENNA_109 (.A(_0360_));
 sg13g2_antennanp ANTENNA_110 (.A(_0360_));
 sg13g2_antennanp ANTENNA_111 (.A(_0387_));
 sg13g2_antennanp ANTENNA_112 (.A(_0387_));
 sg13g2_antennanp ANTENNA_113 (.A(_0387_));
 sg13g2_antennanp ANTENNA_114 (.A(_0387_));
 sg13g2_antennanp ANTENNA_115 (.A(_0387_));
 sg13g2_antennanp ANTENNA_116 (.A(_0387_));
 sg13g2_antennanp ANTENNA_117 (.A(_0435_));
 sg13g2_antennanp ANTENNA_118 (.A(_0438_));
 sg13g2_antennanp ANTENNA_119 (.A(_0438_));
 sg13g2_antennanp ANTENNA_120 (.A(_0438_));
 sg13g2_antennanp ANTENNA_121 (.A(_0438_));
 sg13g2_antennanp ANTENNA_122 (.A(_0438_));
 sg13g2_antennanp ANTENNA_123 (.A(_0438_));
 sg13g2_antennanp ANTENNA_124 (.A(_0448_));
 sg13g2_antennanp ANTENNA_125 (.A(_0474_));
 sg13g2_antennanp ANTENNA_126 (.A(_0477_));
 sg13g2_antennanp ANTENNA_127 (.A(_0477_));
 sg13g2_antennanp ANTENNA_128 (.A(_0477_));
 sg13g2_antennanp ANTENNA_129 (.A(_0477_));
 sg13g2_antennanp ANTENNA_130 (.A(_0477_));
 sg13g2_antennanp ANTENNA_131 (.A(_0477_));
 sg13g2_antennanp ANTENNA_132 (.A(_0477_));
 sg13g2_antennanp ANTENNA_133 (.A(_0490_));
 sg13g2_antennanp ANTENNA_134 (.A(_0490_));
 sg13g2_antennanp ANTENNA_135 (.A(_0507_));
 sg13g2_antennanp ANTENNA_136 (.A(_0507_));
 sg13g2_antennanp ANTENNA_137 (.A(_0511_));
 sg13g2_antennanp ANTENNA_138 (.A(_0511_));
 sg13g2_antennanp ANTENNA_139 (.A(_0521_));
 sg13g2_antennanp ANTENNA_140 (.A(_0521_));
 sg13g2_antennanp ANTENNA_141 (.A(_0521_));
 sg13g2_antennanp ANTENNA_142 (.A(_0597_));
 sg13g2_antennanp ANTENNA_143 (.A(_0597_));
 sg13g2_antennanp ANTENNA_144 (.A(_0597_));
 sg13g2_antennanp ANTENNA_145 (.A(_0597_));
 sg13g2_antennanp ANTENNA_146 (.A(_0597_));
 sg13g2_antennanp ANTENNA_147 (.A(_0598_));
 sg13g2_antennanp ANTENNA_148 (.A(_0598_));
 sg13g2_antennanp ANTENNA_149 (.A(_0598_));
 sg13g2_antennanp ANTENNA_150 (.A(_0598_));
 sg13g2_antennanp ANTENNA_151 (.A(_0598_));
 sg13g2_antennanp ANTENNA_152 (.A(_0623_));
 sg13g2_antennanp ANTENNA_153 (.A(_0780_));
 sg13g2_antennanp ANTENNA_154 (.A(_0780_));
 sg13g2_antennanp ANTENNA_155 (.A(_0800_));
 sg13g2_antennanp ANTENNA_156 (.A(_0800_));
 sg13g2_antennanp ANTENNA_157 (.A(_0824_));
 sg13g2_antennanp ANTENNA_158 (.A(_0824_));
 sg13g2_antennanp ANTENNA_159 (.A(_0824_));
 sg13g2_antennanp ANTENNA_160 (.A(_0866_));
 sg13g2_antennanp ANTENNA_161 (.A(_0866_));
 sg13g2_antennanp ANTENNA_162 (.A(_0866_));
 sg13g2_antennanp ANTENNA_163 (.A(_0878_));
 sg13g2_antennanp ANTENNA_164 (.A(_0878_));
 sg13g2_antennanp ANTENNA_165 (.A(_0878_));
 sg13g2_antennanp ANTENNA_166 (.A(_0878_));
 sg13g2_antennanp ANTENNA_167 (.A(_0878_));
 sg13g2_antennanp ANTENNA_168 (.A(_0878_));
 sg13g2_antennanp ANTENNA_169 (.A(_0878_));
 sg13g2_antennanp ANTENNA_170 (.A(_0878_));
 sg13g2_antennanp ANTENNA_171 (.A(_0878_));
 sg13g2_antennanp ANTENNA_172 (.A(_0901_));
 sg13g2_antennanp ANTENNA_173 (.A(_0901_));
 sg13g2_antennanp ANTENNA_174 (.A(_0915_));
 sg13g2_antennanp ANTENNA_175 (.A(_0915_));
 sg13g2_antennanp ANTENNA_176 (.A(_0915_));
 sg13g2_antennanp ANTENNA_177 (.A(_0990_));
 sg13g2_antennanp ANTENNA_178 (.A(_0990_));
 sg13g2_antennanp ANTENNA_179 (.A(_1002_));
 sg13g2_antennanp ANTENNA_180 (.A(_1002_));
 sg13g2_antennanp ANTENNA_181 (.A(_1071_));
 sg13g2_antennanp ANTENNA_182 (.A(_1071_));
 sg13g2_antennanp ANTENNA_183 (.A(_1071_));
 sg13g2_antennanp ANTENNA_184 (.A(_1085_));
 sg13g2_antennanp ANTENNA_185 (.A(_1085_));
 sg13g2_antennanp ANTENNA_186 (.A(_1085_));
 sg13g2_antennanp ANTENNA_187 (.A(_1085_));
 sg13g2_antennanp ANTENNA_188 (.A(_1085_));
 sg13g2_antennanp ANTENNA_189 (.A(_1151_));
 sg13g2_antennanp ANTENNA_190 (.A(_1151_));
 sg13g2_antennanp ANTENNA_191 (.A(_1151_));
 sg13g2_antennanp ANTENNA_192 (.A(_1151_));
 sg13g2_antennanp ANTENNA_193 (.A(_1151_));
 sg13g2_antennanp ANTENNA_194 (.A(_1151_));
 sg13g2_antennanp ANTENNA_195 (.A(_1151_));
 sg13g2_antennanp ANTENNA_196 (.A(_1162_));
 sg13g2_antennanp ANTENNA_197 (.A(_1162_));
 sg13g2_antennanp ANTENNA_198 (.A(_1162_));
 sg13g2_antennanp ANTENNA_199 (.A(_1162_));
 sg13g2_antennanp ANTENNA_200 (.A(_1162_));
 sg13g2_antennanp ANTENNA_201 (.A(_1162_));
 sg13g2_antennanp ANTENNA_202 (.A(_1162_));
 sg13g2_antennanp ANTENNA_203 (.A(_1162_));
 sg13g2_antennanp ANTENNA_204 (.A(_1162_));
 sg13g2_antennanp ANTENNA_205 (.A(_1162_));
 sg13g2_antennanp ANTENNA_206 (.A(_1162_));
 sg13g2_antennanp ANTENNA_207 (.A(_1199_));
 sg13g2_antennanp ANTENNA_208 (.A(_1209_));
 sg13g2_antennanp ANTENNA_209 (.A(_1209_));
 sg13g2_antennanp ANTENNA_210 (.A(_1209_));
 sg13g2_antennanp ANTENNA_211 (.A(_1225_));
 sg13g2_antennanp ANTENNA_212 (.A(_1225_));
 sg13g2_antennanp ANTENNA_213 (.A(_1292_));
 sg13g2_antennanp ANTENNA_214 (.A(_1292_));
 sg13g2_antennanp ANTENNA_215 (.A(_1319_));
 sg13g2_antennanp ANTENNA_216 (.A(_1326_));
 sg13g2_antennanp ANTENNA_217 (.A(_1326_));
 sg13g2_antennanp ANTENNA_218 (.A(_1326_));
 sg13g2_antennanp ANTENNA_219 (.A(_1326_));
 sg13g2_antennanp ANTENNA_220 (.A(_1326_));
 sg13g2_antennanp ANTENNA_221 (.A(_1326_));
 sg13g2_antennanp ANTENNA_222 (.A(_1326_));
 sg13g2_antennanp ANTENNA_223 (.A(_1326_));
 sg13g2_antennanp ANTENNA_224 (.A(_1326_));
 sg13g2_antennanp ANTENNA_225 (.A(_1326_));
 sg13g2_antennanp ANTENNA_226 (.A(_1326_));
 sg13g2_antennanp ANTENNA_227 (.A(_1326_));
 sg13g2_antennanp ANTENNA_228 (.A(_1326_));
 sg13g2_antennanp ANTENNA_229 (.A(_1326_));
 sg13g2_antennanp ANTENNA_230 (.A(_1363_));
 sg13g2_antennanp ANTENNA_231 (.A(_1411_));
 sg13g2_antennanp ANTENNA_232 (.A(_1439_));
 sg13g2_antennanp ANTENNA_233 (.A(_1470_));
 sg13g2_antennanp ANTENNA_234 (.A(_1470_));
 sg13g2_antennanp ANTENNA_235 (.A(_1519_));
 sg13g2_antennanp ANTENNA_236 (.A(_1522_));
 sg13g2_antennanp ANTENNA_237 (.A(_1522_));
 sg13g2_antennanp ANTENNA_238 (.A(_1522_));
 sg13g2_antennanp ANTENNA_239 (.A(_1531_));
 sg13g2_antennanp ANTENNA_240 (.A(_1531_));
 sg13g2_antennanp ANTENNA_241 (.A(_1532_));
 sg13g2_antennanp ANTENNA_242 (.A(_1532_));
 sg13g2_antennanp ANTENNA_243 (.A(_1532_));
 sg13g2_antennanp ANTENNA_244 (.A(_1544_));
 sg13g2_antennanp ANTENNA_245 (.A(_1544_));
 sg13g2_antennanp ANTENNA_246 (.A(_1544_));
 sg13g2_antennanp ANTENNA_247 (.A(_1553_));
 sg13g2_antennanp ANTENNA_248 (.A(_1631_));
 sg13g2_antennanp ANTENNA_249 (.A(_1631_));
 sg13g2_antennanp ANTENNA_250 (.A(_1631_));
 sg13g2_antennanp ANTENNA_251 (.A(_1685_));
 sg13g2_antennanp ANTENNA_252 (.A(_1685_));
 sg13g2_antennanp ANTENNA_253 (.A(_1685_));
 sg13g2_antennanp ANTENNA_254 (.A(_1685_));
 sg13g2_antennanp ANTENNA_255 (.A(_1696_));
 sg13g2_antennanp ANTENNA_256 (.A(_1696_));
 sg13g2_antennanp ANTENNA_257 (.A(_1696_));
 sg13g2_antennanp ANTENNA_258 (.A(_1697_));
 sg13g2_antennanp ANTENNA_259 (.A(_1697_));
 sg13g2_antennanp ANTENNA_260 (.A(_1697_));
 sg13g2_antennanp ANTENNA_261 (.A(_1707_));
 sg13g2_antennanp ANTENNA_262 (.A(_1707_));
 sg13g2_antennanp ANTENNA_263 (.A(_1707_));
 sg13g2_antennanp ANTENNA_264 (.A(_1707_));
 sg13g2_antennanp ANTENNA_265 (.A(_1707_));
 sg13g2_antennanp ANTENNA_266 (.A(_1716_));
 sg13g2_antennanp ANTENNA_267 (.A(_1716_));
 sg13g2_antennanp ANTENNA_268 (.A(_1735_));
 sg13g2_antennanp ANTENNA_269 (.A(_1735_));
 sg13g2_antennanp ANTENNA_270 (.A(_1761_));
 sg13g2_antennanp ANTENNA_271 (.A(_1761_));
 sg13g2_antennanp ANTENNA_272 (.A(_2014_));
 sg13g2_antennanp ANTENNA_273 (.A(_2014_));
 sg13g2_antennanp ANTENNA_274 (.A(_2020_));
 sg13g2_antennanp ANTENNA_275 (.A(_2020_));
 sg13g2_antennanp ANTENNA_276 (.A(_2020_));
 sg13g2_antennanp ANTENNA_277 (.A(_2020_));
 sg13g2_antennanp ANTENNA_278 (.A(_2020_));
 sg13g2_antennanp ANTENNA_279 (.A(_2020_));
 sg13g2_antennanp ANTENNA_280 (.A(_2020_));
 sg13g2_antennanp ANTENNA_281 (.A(_2037_));
 sg13g2_antennanp ANTENNA_282 (.A(_2053_));
 sg13g2_antennanp ANTENNA_283 (.A(_2053_));
 sg13g2_antennanp ANTENNA_284 (.A(_2053_));
 sg13g2_antennanp ANTENNA_285 (.A(_2097_));
 sg13g2_antennanp ANTENNA_286 (.A(_2097_));
 sg13g2_antennanp ANTENNA_287 (.A(_2097_));
 sg13g2_antennanp ANTENNA_288 (.A(_2097_));
 sg13g2_antennanp ANTENNA_289 (.A(_2097_));
 sg13g2_antennanp ANTENNA_290 (.A(_2110_));
 sg13g2_antennanp ANTENNA_291 (.A(_2112_));
 sg13g2_antennanp ANTENNA_292 (.A(_2145_));
 sg13g2_antennanp ANTENNA_293 (.A(_2171_));
 sg13g2_antennanp ANTENNA_294 (.A(_2171_));
 sg13g2_antennanp ANTENNA_295 (.A(_2171_));
 sg13g2_antennanp ANTENNA_296 (.A(_2171_));
 sg13g2_antennanp ANTENNA_297 (.A(_2171_));
 sg13g2_antennanp ANTENNA_298 (.A(_2171_));
 sg13g2_antennanp ANTENNA_299 (.A(_2171_));
 sg13g2_antennanp ANTENNA_300 (.A(_2171_));
 sg13g2_antennanp ANTENNA_301 (.A(_2171_));
 sg13g2_antennanp ANTENNA_302 (.A(_2172_));
 sg13g2_antennanp ANTENNA_303 (.A(_2172_));
 sg13g2_antennanp ANTENNA_304 (.A(_2172_));
 sg13g2_antennanp ANTENNA_305 (.A(_2172_));
 sg13g2_antennanp ANTENNA_306 (.A(_2172_));
 sg13g2_antennanp ANTENNA_307 (.A(_2172_));
 sg13g2_antennanp ANTENNA_308 (.A(_2172_));
 sg13g2_antennanp ANTENNA_309 (.A(_2172_));
 sg13g2_antennanp ANTENNA_310 (.A(_2172_));
 sg13g2_antennanp ANTENNA_311 (.A(_2257_));
 sg13g2_antennanp ANTENNA_312 (.A(_2257_));
 sg13g2_antennanp ANTENNA_313 (.A(_2408_));
 sg13g2_antennanp ANTENNA_314 (.A(_2408_));
 sg13g2_antennanp ANTENNA_315 (.A(_2408_));
 sg13g2_antennanp ANTENNA_316 (.A(_2423_));
 sg13g2_antennanp ANTENNA_317 (.A(_2423_));
 sg13g2_antennanp ANTENNA_318 (.A(_2423_));
 sg13g2_antennanp ANTENNA_319 (.A(_2423_));
 sg13g2_antennanp ANTENNA_320 (.A(_2423_));
 sg13g2_antennanp ANTENNA_321 (.A(_2423_));
 sg13g2_antennanp ANTENNA_322 (.A(_2423_));
 sg13g2_antennanp ANTENNA_323 (.A(_2423_));
 sg13g2_antennanp ANTENNA_324 (.A(_2423_));
 sg13g2_antennanp ANTENNA_325 (.A(_2429_));
 sg13g2_antennanp ANTENNA_326 (.A(_2429_));
 sg13g2_antennanp ANTENNA_327 (.A(_2429_));
 sg13g2_antennanp ANTENNA_328 (.A(_2429_));
 sg13g2_antennanp ANTENNA_329 (.A(_2429_));
 sg13g2_antennanp ANTENNA_330 (.A(_2429_));
 sg13g2_antennanp ANTENNA_331 (.A(_2429_));
 sg13g2_antennanp ANTENNA_332 (.A(_2429_));
 sg13g2_antennanp ANTENNA_333 (.A(_2430_));
 sg13g2_antennanp ANTENNA_334 (.A(_2430_));
 sg13g2_antennanp ANTENNA_335 (.A(_2430_));
 sg13g2_antennanp ANTENNA_336 (.A(_2430_));
 sg13g2_antennanp ANTENNA_337 (.A(_2430_));
 sg13g2_antennanp ANTENNA_338 (.A(_2430_));
 sg13g2_antennanp ANTENNA_339 (.A(_2444_));
 sg13g2_antennanp ANTENNA_340 (.A(_2444_));
 sg13g2_antennanp ANTENNA_341 (.A(_2444_));
 sg13g2_antennanp ANTENNA_342 (.A(_2444_));
 sg13g2_antennanp ANTENNA_343 (.A(_2444_));
 sg13g2_antennanp ANTENNA_344 (.A(_2444_));
 sg13g2_antennanp ANTENNA_345 (.A(_2444_));
 sg13g2_antennanp ANTENNA_346 (.A(_2461_));
 sg13g2_antennanp ANTENNA_347 (.A(_2461_));
 sg13g2_antennanp ANTENNA_348 (.A(_2461_));
 sg13g2_antennanp ANTENNA_349 (.A(_2461_));
 sg13g2_antennanp ANTENNA_350 (.A(_2461_));
 sg13g2_antennanp ANTENNA_351 (.A(_2467_));
 sg13g2_antennanp ANTENNA_352 (.A(_2467_));
 sg13g2_antennanp ANTENNA_353 (.A(_2467_));
 sg13g2_antennanp ANTENNA_354 (.A(_2467_));
 sg13g2_antennanp ANTENNA_355 (.A(_2467_));
 sg13g2_antennanp ANTENNA_356 (.A(_2470_));
 sg13g2_antennanp ANTENNA_357 (.A(_2470_));
 sg13g2_antennanp ANTENNA_358 (.A(_2470_));
 sg13g2_antennanp ANTENNA_359 (.A(_2470_));
 sg13g2_antennanp ANTENNA_360 (.A(_2470_));
 sg13g2_antennanp ANTENNA_361 (.A(_2478_));
 sg13g2_antennanp ANTENNA_362 (.A(_2478_));
 sg13g2_antennanp ANTENNA_363 (.A(_2478_));
 sg13g2_antennanp ANTENNA_364 (.A(_2478_));
 sg13g2_antennanp ANTENNA_365 (.A(_2478_));
 sg13g2_antennanp ANTENNA_366 (.A(_2480_));
 sg13g2_antennanp ANTENNA_367 (.A(_2480_));
 sg13g2_antennanp ANTENNA_368 (.A(_2480_));
 sg13g2_antennanp ANTENNA_369 (.A(_2480_));
 sg13g2_antennanp ANTENNA_370 (.A(_2480_));
 sg13g2_antennanp ANTENNA_371 (.A(_2482_));
 sg13g2_antennanp ANTENNA_372 (.A(_2482_));
 sg13g2_antennanp ANTENNA_373 (.A(_2482_));
 sg13g2_antennanp ANTENNA_374 (.A(_2482_));
 sg13g2_antennanp ANTENNA_375 (.A(_2482_));
 sg13g2_antennanp ANTENNA_376 (.A(_2482_));
 sg13g2_antennanp ANTENNA_377 (.A(_2482_));
 sg13g2_antennanp ANTENNA_378 (.A(_2487_));
 sg13g2_antennanp ANTENNA_379 (.A(_2487_));
 sg13g2_antennanp ANTENNA_380 (.A(_2501_));
 sg13g2_antennanp ANTENNA_381 (.A(_2501_));
 sg13g2_antennanp ANTENNA_382 (.A(_2501_));
 sg13g2_antennanp ANTENNA_383 (.A(_2501_));
 sg13g2_antennanp ANTENNA_384 (.A(_2501_));
 sg13g2_antennanp ANTENNA_385 (.A(_2501_));
 sg13g2_antennanp ANTENNA_386 (.A(_2518_));
 sg13g2_antennanp ANTENNA_387 (.A(_2518_));
 sg13g2_antennanp ANTENNA_388 (.A(_2518_));
 sg13g2_antennanp ANTENNA_389 (.A(_2518_));
 sg13g2_antennanp ANTENNA_390 (.A(_2518_));
 sg13g2_antennanp ANTENNA_391 (.A(_2518_));
 sg13g2_antennanp ANTENNA_392 (.A(_2518_));
 sg13g2_antennanp ANTENNA_393 (.A(_2518_));
 sg13g2_antennanp ANTENNA_394 (.A(_2518_));
 sg13g2_antennanp ANTENNA_395 (.A(_2520_));
 sg13g2_antennanp ANTENNA_396 (.A(_2520_));
 sg13g2_antennanp ANTENNA_397 (.A(_2520_));
 sg13g2_antennanp ANTENNA_398 (.A(_2520_));
 sg13g2_antennanp ANTENNA_399 (.A(_2520_));
 sg13g2_antennanp ANTENNA_400 (.A(_2520_));
 sg13g2_antennanp ANTENNA_401 (.A(_2530_));
 sg13g2_antennanp ANTENNA_402 (.A(_2530_));
 sg13g2_antennanp ANTENNA_403 (.A(_2530_));
 sg13g2_antennanp ANTENNA_404 (.A(_2530_));
 sg13g2_antennanp ANTENNA_405 (.A(_2530_));
 sg13g2_antennanp ANTENNA_406 (.A(_2530_));
 sg13g2_antennanp ANTENNA_407 (.A(_2532_));
 sg13g2_antennanp ANTENNA_408 (.A(_2532_));
 sg13g2_antennanp ANTENNA_409 (.A(_2532_));
 sg13g2_antennanp ANTENNA_410 (.A(_2532_));
 sg13g2_antennanp ANTENNA_411 (.A(_2532_));
 sg13g2_antennanp ANTENNA_412 (.A(_2532_));
 sg13g2_antennanp ANTENNA_413 (.A(_2532_));
 sg13g2_antennanp ANTENNA_414 (.A(_2532_));
 sg13g2_antennanp ANTENNA_415 (.A(_2532_));
 sg13g2_antennanp ANTENNA_416 (.A(_2532_));
 sg13g2_antennanp ANTENNA_417 (.A(_2537_));
 sg13g2_antennanp ANTENNA_418 (.A(_2537_));
 sg13g2_antennanp ANTENNA_419 (.A(_2537_));
 sg13g2_antennanp ANTENNA_420 (.A(_2537_));
 sg13g2_antennanp ANTENNA_421 (.A(_2552_));
 sg13g2_antennanp ANTENNA_422 (.A(_2552_));
 sg13g2_antennanp ANTENNA_423 (.A(_2552_));
 sg13g2_antennanp ANTENNA_424 (.A(_2557_));
 sg13g2_antennanp ANTENNA_425 (.A(_2557_));
 sg13g2_antennanp ANTENNA_426 (.A(_2557_));
 sg13g2_antennanp ANTENNA_427 (.A(_2573_));
 sg13g2_antennanp ANTENNA_428 (.A(_2573_));
 sg13g2_antennanp ANTENNA_429 (.A(_2573_));
 sg13g2_antennanp ANTENNA_430 (.A(_2573_));
 sg13g2_antennanp ANTENNA_431 (.A(_2574_));
 sg13g2_antennanp ANTENNA_432 (.A(_2574_));
 sg13g2_antennanp ANTENNA_433 (.A(_2574_));
 sg13g2_antennanp ANTENNA_434 (.A(_2574_));
 sg13g2_antennanp ANTENNA_435 (.A(_2577_));
 sg13g2_antennanp ANTENNA_436 (.A(_2577_));
 sg13g2_antennanp ANTENNA_437 (.A(_2577_));
 sg13g2_antennanp ANTENNA_438 (.A(_2577_));
 sg13g2_antennanp ANTENNA_439 (.A(_2577_));
 sg13g2_antennanp ANTENNA_440 (.A(_2577_));
 sg13g2_antennanp ANTENNA_441 (.A(_2577_));
 sg13g2_antennanp ANTENNA_442 (.A(_2577_));
 sg13g2_antennanp ANTENNA_443 (.A(_2585_));
 sg13g2_antennanp ANTENNA_444 (.A(_2585_));
 sg13g2_antennanp ANTENNA_445 (.A(_2585_));
 sg13g2_antennanp ANTENNA_446 (.A(_2588_));
 sg13g2_antennanp ANTENNA_447 (.A(_2595_));
 sg13g2_antennanp ANTENNA_448 (.A(_2595_));
 sg13g2_antennanp ANTENNA_449 (.A(_2595_));
 sg13g2_antennanp ANTENNA_450 (.A(_2595_));
 sg13g2_antennanp ANTENNA_451 (.A(_2595_));
 sg13g2_antennanp ANTENNA_452 (.A(_2595_));
 sg13g2_antennanp ANTENNA_453 (.A(_2596_));
 sg13g2_antennanp ANTENNA_454 (.A(_2596_));
 sg13g2_antennanp ANTENNA_455 (.A(_2596_));
 sg13g2_antennanp ANTENNA_456 (.A(_2600_));
 sg13g2_antennanp ANTENNA_457 (.A(_2600_));
 sg13g2_antennanp ANTENNA_458 (.A(_2600_));
 sg13g2_antennanp ANTENNA_459 (.A(_2601_));
 sg13g2_antennanp ANTENNA_460 (.A(_2601_));
 sg13g2_antennanp ANTENNA_461 (.A(_2601_));
 sg13g2_antennanp ANTENNA_462 (.A(_2607_));
 sg13g2_antennanp ANTENNA_463 (.A(_2607_));
 sg13g2_antennanp ANTENNA_464 (.A(_2615_));
 sg13g2_antennanp ANTENNA_465 (.A(_2615_));
 sg13g2_antennanp ANTENNA_466 (.A(_2615_));
 sg13g2_antennanp ANTENNA_467 (.A(_2615_));
 sg13g2_antennanp ANTENNA_468 (.A(_2619_));
 sg13g2_antennanp ANTENNA_469 (.A(_2619_));
 sg13g2_antennanp ANTENNA_470 (.A(_2619_));
 sg13g2_antennanp ANTENNA_471 (.A(_2619_));
 sg13g2_antennanp ANTENNA_472 (.A(_2622_));
 sg13g2_antennanp ANTENNA_473 (.A(_2622_));
 sg13g2_antennanp ANTENNA_474 (.A(_2622_));
 sg13g2_antennanp ANTENNA_475 (.A(_2622_));
 sg13g2_antennanp ANTENNA_476 (.A(_2622_));
 sg13g2_antennanp ANTENNA_477 (.A(_2622_));
 sg13g2_antennanp ANTENNA_478 (.A(_2625_));
 sg13g2_antennanp ANTENNA_479 (.A(_2625_));
 sg13g2_antennanp ANTENNA_480 (.A(_2625_));
 sg13g2_antennanp ANTENNA_481 (.A(_2625_));
 sg13g2_antennanp ANTENNA_482 (.A(_2653_));
 sg13g2_antennanp ANTENNA_483 (.A(_2653_));
 sg13g2_antennanp ANTENNA_484 (.A(_2653_));
 sg13g2_antennanp ANTENNA_485 (.A(_2659_));
 sg13g2_antennanp ANTENNA_486 (.A(_2659_));
 sg13g2_antennanp ANTENNA_487 (.A(_2659_));
 sg13g2_antennanp ANTENNA_488 (.A(_2659_));
 sg13g2_antennanp ANTENNA_489 (.A(_2659_));
 sg13g2_antennanp ANTENNA_490 (.A(_2665_));
 sg13g2_antennanp ANTENNA_491 (.A(_2665_));
 sg13g2_antennanp ANTENNA_492 (.A(_2665_));
 sg13g2_antennanp ANTENNA_493 (.A(_2665_));
 sg13g2_antennanp ANTENNA_494 (.A(_2678_));
 sg13g2_antennanp ANTENNA_495 (.A(_2678_));
 sg13g2_antennanp ANTENNA_496 (.A(_2678_));
 sg13g2_antennanp ANTENNA_497 (.A(_2678_));
 sg13g2_antennanp ANTENNA_498 (.A(_2678_));
 sg13g2_antennanp ANTENNA_499 (.A(_2678_));
 sg13g2_antennanp ANTENNA_500 (.A(_2678_));
 sg13g2_antennanp ANTENNA_501 (.A(_2681_));
 sg13g2_antennanp ANTENNA_502 (.A(_2681_));
 sg13g2_antennanp ANTENNA_503 (.A(_2719_));
 sg13g2_antennanp ANTENNA_504 (.A(_2719_));
 sg13g2_antennanp ANTENNA_505 (.A(_2719_));
 sg13g2_antennanp ANTENNA_506 (.A(_2719_));
 sg13g2_antennanp ANTENNA_507 (.A(_2719_));
 sg13g2_antennanp ANTENNA_508 (.A(_2732_));
 sg13g2_antennanp ANTENNA_509 (.A(_2732_));
 sg13g2_antennanp ANTENNA_510 (.A(_2732_));
 sg13g2_antennanp ANTENNA_511 (.A(_2732_));
 sg13g2_antennanp ANTENNA_512 (.A(_2732_));
 sg13g2_antennanp ANTENNA_513 (.A(_2733_));
 sg13g2_antennanp ANTENNA_514 (.A(_2733_));
 sg13g2_antennanp ANTENNA_515 (.A(_2733_));
 sg13g2_antennanp ANTENNA_516 (.A(_2733_));
 sg13g2_antennanp ANTENNA_517 (.A(_2739_));
 sg13g2_antennanp ANTENNA_518 (.A(_2739_));
 sg13g2_antennanp ANTENNA_519 (.A(_2739_));
 sg13g2_antennanp ANTENNA_520 (.A(_2739_));
 sg13g2_antennanp ANTENNA_521 (.A(_2745_));
 sg13g2_antennanp ANTENNA_522 (.A(_2745_));
 sg13g2_antennanp ANTENNA_523 (.A(_2745_));
 sg13g2_antennanp ANTENNA_524 (.A(_2745_));
 sg13g2_antennanp ANTENNA_525 (.A(_2745_));
 sg13g2_antennanp ANTENNA_526 (.A(_2745_));
 sg13g2_antennanp ANTENNA_527 (.A(_2745_));
 sg13g2_antennanp ANTENNA_528 (.A(_2749_));
 sg13g2_antennanp ANTENNA_529 (.A(_2749_));
 sg13g2_antennanp ANTENNA_530 (.A(_2749_));
 sg13g2_antennanp ANTENNA_531 (.A(_2749_));
 sg13g2_antennanp ANTENNA_532 (.A(_2769_));
 sg13g2_antennanp ANTENNA_533 (.A(_2769_));
 sg13g2_antennanp ANTENNA_534 (.A(_2769_));
 sg13g2_antennanp ANTENNA_535 (.A(_2769_));
 sg13g2_antennanp ANTENNA_536 (.A(_2775_));
 sg13g2_antennanp ANTENNA_537 (.A(_2775_));
 sg13g2_antennanp ANTENNA_538 (.A(_2779_));
 sg13g2_antennanp ANTENNA_539 (.A(_2779_));
 sg13g2_antennanp ANTENNA_540 (.A(_2779_));
 sg13g2_antennanp ANTENNA_541 (.A(_2779_));
 sg13g2_antennanp ANTENNA_542 (.A(_2789_));
 sg13g2_antennanp ANTENNA_543 (.A(_2789_));
 sg13g2_antennanp ANTENNA_544 (.A(_2789_));
 sg13g2_antennanp ANTENNA_545 (.A(_2789_));
 sg13g2_antennanp ANTENNA_546 (.A(_2805_));
 sg13g2_antennanp ANTENNA_547 (.A(_2805_));
 sg13g2_antennanp ANTENNA_548 (.A(_2808_));
 sg13g2_antennanp ANTENNA_549 (.A(_2808_));
 sg13g2_antennanp ANTENNA_550 (.A(_2808_));
 sg13g2_antennanp ANTENNA_551 (.A(_2808_));
 sg13g2_antennanp ANTENNA_552 (.A(_2816_));
 sg13g2_antennanp ANTENNA_553 (.A(_2816_));
 sg13g2_antennanp ANTENNA_554 (.A(_2816_));
 sg13g2_antennanp ANTENNA_555 (.A(_2816_));
 sg13g2_antennanp ANTENNA_556 (.A(_2816_));
 sg13g2_antennanp ANTENNA_557 (.A(_2816_));
 sg13g2_antennanp ANTENNA_558 (.A(_2826_));
 sg13g2_antennanp ANTENNA_559 (.A(_2826_));
 sg13g2_antennanp ANTENNA_560 (.A(_2826_));
 sg13g2_antennanp ANTENNA_561 (.A(_2826_));
 sg13g2_antennanp ANTENNA_562 (.A(_2854_));
 sg13g2_antennanp ANTENNA_563 (.A(_2854_));
 sg13g2_antennanp ANTENNA_564 (.A(_2854_));
 sg13g2_antennanp ANTENNA_565 (.A(_2854_));
 sg13g2_antennanp ANTENNA_566 (.A(_2854_));
 sg13g2_antennanp ANTENNA_567 (.A(_2854_));
 sg13g2_antennanp ANTENNA_568 (.A(_2854_));
 sg13g2_antennanp ANTENNA_569 (.A(_2854_));
 sg13g2_antennanp ANTENNA_570 (.A(_2854_));
 sg13g2_antennanp ANTENNA_571 (.A(_2854_));
 sg13g2_antennanp ANTENNA_572 (.A(_2854_));
 sg13g2_antennanp ANTENNA_573 (.A(_2854_));
 sg13g2_antennanp ANTENNA_574 (.A(_2858_));
 sg13g2_antennanp ANTENNA_575 (.A(_2858_));
 sg13g2_antennanp ANTENNA_576 (.A(_2879_));
 sg13g2_antennanp ANTENNA_577 (.A(_2879_));
 sg13g2_antennanp ANTENNA_578 (.A(_2879_));
 sg13g2_antennanp ANTENNA_579 (.A(_2879_));
 sg13g2_antennanp ANTENNA_580 (.A(_2879_));
 sg13g2_antennanp ANTENNA_581 (.A(_2879_));
 sg13g2_antennanp ANTENNA_582 (.A(_2879_));
 sg13g2_antennanp ANTENNA_583 (.A(_2879_));
 sg13g2_antennanp ANTENNA_584 (.A(_2879_));
 sg13g2_antennanp ANTENNA_585 (.A(_2879_));
 sg13g2_antennanp ANTENNA_586 (.A(_2914_));
 sg13g2_antennanp ANTENNA_587 (.A(_2931_));
 sg13g2_antennanp ANTENNA_588 (.A(_2931_));
 sg13g2_antennanp ANTENNA_589 (.A(_2931_));
 sg13g2_antennanp ANTENNA_590 (.A(_2936_));
 sg13g2_antennanp ANTENNA_591 (.A(_2936_));
 sg13g2_antennanp ANTENNA_592 (.A(_2936_));
 sg13g2_antennanp ANTENNA_593 (.A(_2957_));
 sg13g2_antennanp ANTENNA_594 (.A(_2957_));
 sg13g2_antennanp ANTENNA_595 (.A(_2957_));
 sg13g2_antennanp ANTENNA_596 (.A(_2957_));
 sg13g2_antennanp ANTENNA_597 (.A(_2967_));
 sg13g2_antennanp ANTENNA_598 (.A(_2967_));
 sg13g2_antennanp ANTENNA_599 (.A(_2967_));
 sg13g2_antennanp ANTENNA_600 (.A(_2967_));
 sg13g2_antennanp ANTENNA_601 (.A(_2967_));
 sg13g2_antennanp ANTENNA_602 (.A(_2974_));
 sg13g2_antennanp ANTENNA_603 (.A(_2977_));
 sg13g2_antennanp ANTENNA_604 (.A(_2977_));
 sg13g2_antennanp ANTENNA_605 (.A(_2977_));
 sg13g2_antennanp ANTENNA_606 (.A(_2977_));
 sg13g2_antennanp ANTENNA_607 (.A(_2977_));
 sg13g2_antennanp ANTENNA_608 (.A(_2986_));
 sg13g2_antennanp ANTENNA_609 (.A(_2986_));
 sg13g2_antennanp ANTENNA_610 (.A(_2986_));
 sg13g2_antennanp ANTENNA_611 (.A(_2986_));
 sg13g2_antennanp ANTENNA_612 (.A(_3018_));
 sg13g2_antennanp ANTENNA_613 (.A(_3018_));
 sg13g2_antennanp ANTENNA_614 (.A(_3018_));
 sg13g2_antennanp ANTENNA_615 (.A(_3018_));
 sg13g2_antennanp ANTENNA_616 (.A(_3040_));
 sg13g2_antennanp ANTENNA_617 (.A(_3040_));
 sg13g2_antennanp ANTENNA_618 (.A(_3040_));
 sg13g2_antennanp ANTENNA_619 (.A(clk));
 sg13g2_antennanp ANTENNA_620 (.A(clk));
 sg13g2_antennanp ANTENNA_621 (.A(net22));
 sg13g2_antennanp ANTENNA_622 (.A(net22));
 sg13g2_antennanp ANTENNA_623 (.A(net22));
 sg13g2_antennanp ANTENNA_624 (.A(net22));
 sg13g2_antennanp ANTENNA_625 (.A(net22));
 sg13g2_antennanp ANTENNA_626 (.A(net22));
 sg13g2_antennanp ANTENNA_627 (.A(net22));
 sg13g2_antennanp ANTENNA_628 (.A(net22));
 sg13g2_antennanp ANTENNA_629 (.A(net22));
 sg13g2_antennanp ANTENNA_630 (.A(net23));
 sg13g2_antennanp ANTENNA_631 (.A(net23));
 sg13g2_antennanp ANTENNA_632 (.A(net23));
 sg13g2_antennanp ANTENNA_633 (.A(net23));
 sg13g2_antennanp ANTENNA_634 (.A(net23));
 sg13g2_antennanp ANTENNA_635 (.A(net23));
 sg13g2_antennanp ANTENNA_636 (.A(net23));
 sg13g2_antennanp ANTENNA_637 (.A(net23));
 sg13g2_antennanp ANTENNA_638 (.A(net23));
 sg13g2_antennanp ANTENNA_639 (.A(net23));
 sg13g2_antennanp ANTENNA_640 (.A(net23));
 sg13g2_antennanp ANTENNA_641 (.A(net23));
 sg13g2_antennanp ANTENNA_642 (.A(net23));
 sg13g2_antennanp ANTENNA_643 (.A(net23));
 sg13g2_antennanp ANTENNA_644 (.A(net23));
 sg13g2_antennanp ANTENNA_645 (.A(net23));
 sg13g2_antennanp ANTENNA_646 (.A(net23));
 sg13g2_antennanp ANTENNA_647 (.A(net23));
 sg13g2_antennanp ANTENNA_648 (.A(net23));
 sg13g2_antennanp ANTENNA_649 (.A(net23));
 sg13g2_antennanp ANTENNA_650 (.A(net23));
 sg13g2_antennanp ANTENNA_651 (.A(net26));
 sg13g2_antennanp ANTENNA_652 (.A(net26));
 sg13g2_antennanp ANTENNA_653 (.A(net26));
 sg13g2_antennanp ANTENNA_654 (.A(net26));
 sg13g2_antennanp ANTENNA_655 (.A(net26));
 sg13g2_antennanp ANTENNA_656 (.A(net26));
 sg13g2_antennanp ANTENNA_657 (.A(net26));
 sg13g2_antennanp ANTENNA_658 (.A(net26));
 sg13g2_antennanp ANTENNA_659 (.A(net26));
 sg13g2_antennanp ANTENNA_660 (.A(net29));
 sg13g2_antennanp ANTENNA_661 (.A(net29));
 sg13g2_antennanp ANTENNA_662 (.A(net29));
 sg13g2_antennanp ANTENNA_663 (.A(net29));
 sg13g2_antennanp ANTENNA_664 (.A(net29));
 sg13g2_antennanp ANTENNA_665 (.A(net29));
 sg13g2_antennanp ANTENNA_666 (.A(net29));
 sg13g2_antennanp ANTENNA_667 (.A(net29));
 sg13g2_antennanp ANTENNA_668 (.A(net29));
 sg13g2_antennanp ANTENNA_669 (.A(net35));
 sg13g2_antennanp ANTENNA_670 (.A(net35));
 sg13g2_antennanp ANTENNA_671 (.A(net35));
 sg13g2_antennanp ANTENNA_672 (.A(net35));
 sg13g2_antennanp ANTENNA_673 (.A(net35));
 sg13g2_antennanp ANTENNA_674 (.A(net35));
 sg13g2_antennanp ANTENNA_675 (.A(net35));
 sg13g2_antennanp ANTENNA_676 (.A(net35));
 sg13g2_antennanp ANTENNA_677 (.A(net35));
 sg13g2_antennanp ANTENNA_678 (.A(net37));
 sg13g2_antennanp ANTENNA_679 (.A(net37));
 sg13g2_antennanp ANTENNA_680 (.A(net37));
 sg13g2_antennanp ANTENNA_681 (.A(net37));
 sg13g2_antennanp ANTENNA_682 (.A(net37));
 sg13g2_antennanp ANTENNA_683 (.A(net37));
 sg13g2_antennanp ANTENNA_684 (.A(net37));
 sg13g2_antennanp ANTENNA_685 (.A(net37));
 sg13g2_antennanp ANTENNA_686 (.A(net37));
 sg13g2_antennanp ANTENNA_687 (.A(net40));
 sg13g2_antennanp ANTENNA_688 (.A(net40));
 sg13g2_antennanp ANTENNA_689 (.A(net40));
 sg13g2_antennanp ANTENNA_690 (.A(net40));
 sg13g2_antennanp ANTENNA_691 (.A(net40));
 sg13g2_antennanp ANTENNA_692 (.A(net40));
 sg13g2_antennanp ANTENNA_693 (.A(net40));
 sg13g2_antennanp ANTENNA_694 (.A(net40));
 sg13g2_antennanp ANTENNA_695 (.A(net40));
 sg13g2_antennanp ANTENNA_696 (.A(net41));
 sg13g2_antennanp ANTENNA_697 (.A(net41));
 sg13g2_antennanp ANTENNA_698 (.A(net41));
 sg13g2_antennanp ANTENNA_699 (.A(net41));
 sg13g2_antennanp ANTENNA_700 (.A(net41));
 sg13g2_antennanp ANTENNA_701 (.A(net41));
 sg13g2_antennanp ANTENNA_702 (.A(net41));
 sg13g2_antennanp ANTENNA_703 (.A(net41));
 sg13g2_antennanp ANTENNA_704 (.A(net41));
 sg13g2_antennanp ANTENNA_705 (.A(net42));
 sg13g2_antennanp ANTENNA_706 (.A(net42));
 sg13g2_antennanp ANTENNA_707 (.A(net42));
 sg13g2_antennanp ANTENNA_708 (.A(net42));
 sg13g2_antennanp ANTENNA_709 (.A(net42));
 sg13g2_antennanp ANTENNA_710 (.A(net42));
 sg13g2_antennanp ANTENNA_711 (.A(net42));
 sg13g2_antennanp ANTENNA_712 (.A(net42));
 sg13g2_antennanp ANTENNA_713 (.A(net42));
 sg13g2_antennanp ANTENNA_714 (.A(net42));
 sg13g2_antennanp ANTENNA_715 (.A(net42));
 sg13g2_antennanp ANTENNA_716 (.A(net42));
 sg13g2_antennanp ANTENNA_717 (.A(net42));
 sg13g2_antennanp ANTENNA_718 (.A(net42));
 sg13g2_antennanp ANTENNA_719 (.A(net42));
 sg13g2_antennanp ANTENNA_720 (.A(net42));
 sg13g2_antennanp ANTENNA_721 (.A(net42));
 sg13g2_antennanp ANTENNA_722 (.A(net42));
 sg13g2_antennanp ANTENNA_723 (.A(net42));
 sg13g2_antennanp ANTENNA_724 (.A(net46));
 sg13g2_antennanp ANTENNA_725 (.A(net46));
 sg13g2_antennanp ANTENNA_726 (.A(net46));
 sg13g2_antennanp ANTENNA_727 (.A(net46));
 sg13g2_antennanp ANTENNA_728 (.A(net46));
 sg13g2_antennanp ANTENNA_729 (.A(net46));
 sg13g2_antennanp ANTENNA_730 (.A(net46));
 sg13g2_antennanp ANTENNA_731 (.A(net46));
 sg13g2_antennanp ANTENNA_732 (.A(net53));
 sg13g2_antennanp ANTENNA_733 (.A(net53));
 sg13g2_antennanp ANTENNA_734 (.A(net53));
 sg13g2_antennanp ANTENNA_735 (.A(net53));
 sg13g2_antennanp ANTENNA_736 (.A(net53));
 sg13g2_antennanp ANTENNA_737 (.A(net53));
 sg13g2_antennanp ANTENNA_738 (.A(net53));
 sg13g2_antennanp ANTENNA_739 (.A(net53));
 sg13g2_antennanp ANTENNA_740 (.A(net53));
 sg13g2_antennanp ANTENNA_741 (.A(net56));
 sg13g2_antennanp ANTENNA_742 (.A(net56));
 sg13g2_antennanp ANTENNA_743 (.A(net56));
 sg13g2_antennanp ANTENNA_744 (.A(net56));
 sg13g2_antennanp ANTENNA_745 (.A(net56));
 sg13g2_antennanp ANTENNA_746 (.A(net56));
 sg13g2_antennanp ANTENNA_747 (.A(net56));
 sg13g2_antennanp ANTENNA_748 (.A(net56));
 sg13g2_antennanp ANTENNA_749 (.A(net59));
 sg13g2_antennanp ANTENNA_750 (.A(net59));
 sg13g2_antennanp ANTENNA_751 (.A(net59));
 sg13g2_antennanp ANTENNA_752 (.A(net59));
 sg13g2_antennanp ANTENNA_753 (.A(net59));
 sg13g2_antennanp ANTENNA_754 (.A(net59));
 sg13g2_antennanp ANTENNA_755 (.A(net59));
 sg13g2_antennanp ANTENNA_756 (.A(net59));
 sg13g2_antennanp ANTENNA_757 (.A(net61));
 sg13g2_antennanp ANTENNA_758 (.A(net61));
 sg13g2_antennanp ANTENNA_759 (.A(net61));
 sg13g2_antennanp ANTENNA_760 (.A(net61));
 sg13g2_antennanp ANTENNA_761 (.A(net61));
 sg13g2_antennanp ANTENNA_762 (.A(net61));
 sg13g2_antennanp ANTENNA_763 (.A(net61));
 sg13g2_antennanp ANTENNA_764 (.A(net61));
 sg13g2_antennanp ANTENNA_765 (.A(net61));
 sg13g2_antennanp ANTENNA_766 (.A(net62));
 sg13g2_antennanp ANTENNA_767 (.A(net62));
 sg13g2_antennanp ANTENNA_768 (.A(net62));
 sg13g2_antennanp ANTENNA_769 (.A(net62));
 sg13g2_antennanp ANTENNA_770 (.A(net62));
 sg13g2_antennanp ANTENNA_771 (.A(net62));
 sg13g2_antennanp ANTENNA_772 (.A(net62));
 sg13g2_antennanp ANTENNA_773 (.A(net62));
 sg13g2_antennanp ANTENNA_774 (.A(net62));
 sg13g2_antennanp ANTENNA_775 (.A(net64));
 sg13g2_antennanp ANTENNA_776 (.A(net64));
 sg13g2_antennanp ANTENNA_777 (.A(net64));
 sg13g2_antennanp ANTENNA_778 (.A(net64));
 sg13g2_antennanp ANTENNA_779 (.A(net64));
 sg13g2_antennanp ANTENNA_780 (.A(net64));
 sg13g2_antennanp ANTENNA_781 (.A(net64));
 sg13g2_antennanp ANTENNA_782 (.A(net64));
 sg13g2_antennanp ANTENNA_783 (.A(net64));
 sg13g2_antennanp ANTENNA_784 (.A(net67));
 sg13g2_antennanp ANTENNA_785 (.A(net67));
 sg13g2_antennanp ANTENNA_786 (.A(net67));
 sg13g2_antennanp ANTENNA_787 (.A(net67));
 sg13g2_antennanp ANTENNA_788 (.A(net67));
 sg13g2_antennanp ANTENNA_789 (.A(net67));
 sg13g2_antennanp ANTENNA_790 (.A(net67));
 sg13g2_antennanp ANTENNA_791 (.A(net67));
 sg13g2_antennanp ANTENNA_792 (.A(net70));
 sg13g2_antennanp ANTENNA_793 (.A(net70));
 sg13g2_antennanp ANTENNA_794 (.A(net70));
 sg13g2_antennanp ANTENNA_795 (.A(net70));
 sg13g2_antennanp ANTENNA_796 (.A(net70));
 sg13g2_antennanp ANTENNA_797 (.A(net70));
 sg13g2_antennanp ANTENNA_798 (.A(net70));
 sg13g2_antennanp ANTENNA_799 (.A(net70));
 sg13g2_antennanp ANTENNA_800 (.A(net70));
 sg13g2_antennanp ANTENNA_801 (.A(net71));
 sg13g2_antennanp ANTENNA_802 (.A(net71));
 sg13g2_antennanp ANTENNA_803 (.A(net71));
 sg13g2_antennanp ANTENNA_804 (.A(net71));
 sg13g2_antennanp ANTENNA_805 (.A(net71));
 sg13g2_antennanp ANTENNA_806 (.A(net71));
 sg13g2_antennanp ANTENNA_807 (.A(net71));
 sg13g2_antennanp ANTENNA_808 (.A(net71));
 sg13g2_antennanp ANTENNA_809 (.A(net71));
 sg13g2_antennanp ANTENNA_810 (.A(net71));
 sg13g2_antennanp ANTENNA_811 (.A(net71));
 sg13g2_antennanp ANTENNA_812 (.A(net71));
 sg13g2_antennanp ANTENNA_813 (.A(net71));
 sg13g2_antennanp ANTENNA_814 (.A(net71));
 sg13g2_antennanp ANTENNA_815 (.A(net71));
 sg13g2_antennanp ANTENNA_816 (.A(net71));
 sg13g2_antennanp ANTENNA_817 (.A(net75));
 sg13g2_antennanp ANTENNA_818 (.A(net75));
 sg13g2_antennanp ANTENNA_819 (.A(net75));
 sg13g2_antennanp ANTENNA_820 (.A(net75));
 sg13g2_antennanp ANTENNA_821 (.A(net75));
 sg13g2_antennanp ANTENNA_822 (.A(net75));
 sg13g2_antennanp ANTENNA_823 (.A(net75));
 sg13g2_antennanp ANTENNA_824 (.A(net75));
 sg13g2_antennanp ANTENNA_825 (.A(net75));
 sg13g2_antennanp ANTENNA_826 (.A(net75));
 sg13g2_antennanp ANTENNA_827 (.A(net75));
 sg13g2_antennanp ANTENNA_828 (.A(net75));
 sg13g2_antennanp ANTENNA_829 (.A(net75));
 sg13g2_antennanp ANTENNA_830 (.A(net75));
 sg13g2_antennanp ANTENNA_831 (.A(net75));
 sg13g2_antennanp ANTENNA_832 (.A(net75));
 sg13g2_antennanp ANTENNA_833 (.A(net76));
 sg13g2_antennanp ANTENNA_834 (.A(net76));
 sg13g2_antennanp ANTENNA_835 (.A(net76));
 sg13g2_antennanp ANTENNA_836 (.A(net76));
 sg13g2_antennanp ANTENNA_837 (.A(net76));
 sg13g2_antennanp ANTENNA_838 (.A(net76));
 sg13g2_antennanp ANTENNA_839 (.A(net76));
 sg13g2_antennanp ANTENNA_840 (.A(net76));
 sg13g2_antennanp ANTENNA_841 (.A(net76));
 sg13g2_antennanp ANTENNA_842 (.A(net78));
 sg13g2_antennanp ANTENNA_843 (.A(net78));
 sg13g2_antennanp ANTENNA_844 (.A(net78));
 sg13g2_antennanp ANTENNA_845 (.A(net78));
 sg13g2_antennanp ANTENNA_846 (.A(net78));
 sg13g2_antennanp ANTENNA_847 (.A(net78));
 sg13g2_antennanp ANTENNA_848 (.A(net78));
 sg13g2_antennanp ANTENNA_849 (.A(net78));
 sg13g2_antennanp ANTENNA_850 (.A(net78));
 sg13g2_antennanp ANTENNA_851 (.A(net79));
 sg13g2_antennanp ANTENNA_852 (.A(net79));
 sg13g2_antennanp ANTENNA_853 (.A(net79));
 sg13g2_antennanp ANTENNA_854 (.A(net79));
 sg13g2_antennanp ANTENNA_855 (.A(net79));
 sg13g2_antennanp ANTENNA_856 (.A(net79));
 sg13g2_antennanp ANTENNA_857 (.A(net79));
 sg13g2_antennanp ANTENNA_858 (.A(net79));
 sg13g2_antennanp ANTENNA_859 (.A(net79));
 sg13g2_antennanp ANTENNA_860 (.A(net84));
 sg13g2_antennanp ANTENNA_861 (.A(net84));
 sg13g2_antennanp ANTENNA_862 (.A(net84));
 sg13g2_antennanp ANTENNA_863 (.A(net84));
 sg13g2_antennanp ANTENNA_864 (.A(net84));
 sg13g2_antennanp ANTENNA_865 (.A(net84));
 sg13g2_antennanp ANTENNA_866 (.A(net84));
 sg13g2_antennanp ANTENNA_867 (.A(net84));
 sg13g2_antennanp ANTENNA_868 (.A(net85));
 sg13g2_antennanp ANTENNA_869 (.A(net85));
 sg13g2_antennanp ANTENNA_870 (.A(net85));
 sg13g2_antennanp ANTENNA_871 (.A(net85));
 sg13g2_antennanp ANTENNA_872 (.A(net85));
 sg13g2_antennanp ANTENNA_873 (.A(net85));
 sg13g2_antennanp ANTENNA_874 (.A(net85));
 sg13g2_antennanp ANTENNA_875 (.A(net85));
 sg13g2_antennanp ANTENNA_876 (.A(net85));
 sg13g2_antennanp ANTENNA_877 (.A(net89));
 sg13g2_antennanp ANTENNA_878 (.A(net89));
 sg13g2_antennanp ANTENNA_879 (.A(net89));
 sg13g2_antennanp ANTENNA_880 (.A(net89));
 sg13g2_antennanp ANTENNA_881 (.A(net89));
 sg13g2_antennanp ANTENNA_882 (.A(net89));
 sg13g2_antennanp ANTENNA_883 (.A(net89));
 sg13g2_antennanp ANTENNA_884 (.A(net89));
 sg13g2_antennanp ANTENNA_885 (.A(net89));
 sg13g2_antennanp ANTENNA_886 (.A(net91));
 sg13g2_antennanp ANTENNA_887 (.A(net91));
 sg13g2_antennanp ANTENNA_888 (.A(net91));
 sg13g2_antennanp ANTENNA_889 (.A(net91));
 sg13g2_antennanp ANTENNA_890 (.A(net91));
 sg13g2_antennanp ANTENNA_891 (.A(net91));
 sg13g2_antennanp ANTENNA_892 (.A(net91));
 sg13g2_antennanp ANTENNA_893 (.A(net91));
 sg13g2_antennanp ANTENNA_894 (.A(net94));
 sg13g2_antennanp ANTENNA_895 (.A(net94));
 sg13g2_antennanp ANTENNA_896 (.A(net94));
 sg13g2_antennanp ANTENNA_897 (.A(net94));
 sg13g2_antennanp ANTENNA_898 (.A(net94));
 sg13g2_antennanp ANTENNA_899 (.A(net94));
 sg13g2_antennanp ANTENNA_900 (.A(net94));
 sg13g2_antennanp ANTENNA_901 (.A(net94));
 sg13g2_antennanp ANTENNA_902 (.A(net100));
 sg13g2_antennanp ANTENNA_903 (.A(net100));
 sg13g2_antennanp ANTENNA_904 (.A(net100));
 sg13g2_antennanp ANTENNA_905 (.A(net100));
 sg13g2_antennanp ANTENNA_906 (.A(net100));
 sg13g2_antennanp ANTENNA_907 (.A(net100));
 sg13g2_antennanp ANTENNA_908 (.A(net100));
 sg13g2_antennanp ANTENNA_909 (.A(net100));
 sg13g2_antennanp ANTENNA_910 (.A(net100));
 sg13g2_antennanp ANTENNA_911 (.A(net100));
 sg13g2_antennanp ANTENNA_912 (.A(net100));
 sg13g2_antennanp ANTENNA_913 (.A(net100));
 sg13g2_antennanp ANTENNA_914 (.A(net100));
 sg13g2_antennanp ANTENNA_915 (.A(net100));
 sg13g2_antennanp ANTENNA_916 (.A(net100));
 sg13g2_antennanp ANTENNA_917 (.A(net100));
 sg13g2_antennanp ANTENNA_918 (.A(net100));
 sg13g2_antennanp ANTENNA_919 (.A(net100));
 sg13g2_antennanp ANTENNA_920 (.A(net100));
 sg13g2_antennanp ANTENNA_921 (.A(net100));
 sg13g2_antennanp ANTENNA_922 (.A(net100));
 sg13g2_antennanp ANTENNA_923 (.A(net100));
 sg13g2_antennanp ANTENNA_924 (.A(net100));
 sg13g2_antennanp ANTENNA_925 (.A(net100));
 sg13g2_antennanp ANTENNA_926 (.A(net100));
 sg13g2_antennanp ANTENNA_927 (.A(net100));
 sg13g2_antennanp ANTENNA_928 (.A(net100));
 sg13g2_antennanp ANTENNA_929 (.A(net100));
 sg13g2_antennanp ANTENNA_930 (.A(net100));
 sg13g2_antennanp ANTENNA_931 (.A(net101));
 sg13g2_antennanp ANTENNA_932 (.A(net101));
 sg13g2_antennanp ANTENNA_933 (.A(net101));
 sg13g2_antennanp ANTENNA_934 (.A(net101));
 sg13g2_antennanp ANTENNA_935 (.A(net101));
 sg13g2_antennanp ANTENNA_936 (.A(net101));
 sg13g2_antennanp ANTENNA_937 (.A(net101));
 sg13g2_antennanp ANTENNA_938 (.A(net101));
 sg13g2_antennanp ANTENNA_939 (.A(net101));
 sg13g2_antennanp ANTENNA_940 (.A(net106));
 sg13g2_antennanp ANTENNA_941 (.A(net106));
 sg13g2_antennanp ANTENNA_942 (.A(net106));
 sg13g2_antennanp ANTENNA_943 (.A(net106));
 sg13g2_antennanp ANTENNA_944 (.A(net106));
 sg13g2_antennanp ANTENNA_945 (.A(net106));
 sg13g2_antennanp ANTENNA_946 (.A(net106));
 sg13g2_antennanp ANTENNA_947 (.A(net106));
 sg13g2_antennanp ANTENNA_948 (.A(net106));
 sg13g2_antennanp ANTENNA_949 (.A(net107));
 sg13g2_antennanp ANTENNA_950 (.A(net107));
 sg13g2_antennanp ANTENNA_951 (.A(net107));
 sg13g2_antennanp ANTENNA_952 (.A(net107));
 sg13g2_antennanp ANTENNA_953 (.A(net107));
 sg13g2_antennanp ANTENNA_954 (.A(net107));
 sg13g2_antennanp ANTENNA_955 (.A(net107));
 sg13g2_antennanp ANTENNA_956 (.A(net107));
 sg13g2_antennanp ANTENNA_957 (.A(net107));
 sg13g2_antennanp ANTENNA_958 (.A(net113));
 sg13g2_antennanp ANTENNA_959 (.A(net113));
 sg13g2_antennanp ANTENNA_960 (.A(net113));
 sg13g2_antennanp ANTENNA_961 (.A(net113));
 sg13g2_antennanp ANTENNA_962 (.A(net113));
 sg13g2_antennanp ANTENNA_963 (.A(net113));
 sg13g2_antennanp ANTENNA_964 (.A(net113));
 sg13g2_antennanp ANTENNA_965 (.A(net113));
 sg13g2_antennanp ANTENNA_966 (.A(net124));
 sg13g2_antennanp ANTENNA_967 (.A(net124));
 sg13g2_antennanp ANTENNA_968 (.A(net124));
 sg13g2_antennanp ANTENNA_969 (.A(net124));
 sg13g2_antennanp ANTENNA_970 (.A(net124));
 sg13g2_antennanp ANTENNA_971 (.A(net124));
 sg13g2_antennanp ANTENNA_972 (.A(net124));
 sg13g2_antennanp ANTENNA_973 (.A(net124));
 sg13g2_antennanp ANTENNA_974 (.A(net125));
 sg13g2_antennanp ANTENNA_975 (.A(net125));
 sg13g2_antennanp ANTENNA_976 (.A(net125));
 sg13g2_antennanp ANTENNA_977 (.A(net125));
 sg13g2_antennanp ANTENNA_978 (.A(net125));
 sg13g2_antennanp ANTENNA_979 (.A(net125));
 sg13g2_antennanp ANTENNA_980 (.A(net125));
 sg13g2_antennanp ANTENNA_981 (.A(net125));
 sg13g2_antennanp ANTENNA_982 (.A(net125));
 sg13g2_antennanp ANTENNA_983 (.A(net126));
 sg13g2_antennanp ANTENNA_984 (.A(net126));
 sg13g2_antennanp ANTENNA_985 (.A(net126));
 sg13g2_antennanp ANTENNA_986 (.A(net126));
 sg13g2_antennanp ANTENNA_987 (.A(net126));
 sg13g2_antennanp ANTENNA_988 (.A(net126));
 sg13g2_antennanp ANTENNA_989 (.A(net126));
 sg13g2_antennanp ANTENNA_990 (.A(net126));
 sg13g2_antennanp ANTENNA_991 (.A(net126));
 sg13g2_antennanp ANTENNA_992 (.A(net126));
 sg13g2_antennanp ANTENNA_993 (.A(net126));
 sg13g2_antennanp ANTENNA_994 (.A(net126));
 sg13g2_antennanp ANTENNA_995 (.A(net126));
 sg13g2_antennanp ANTENNA_996 (.A(net126));
 sg13g2_antennanp ANTENNA_997 (.A(net126));
 sg13g2_antennanp ANTENNA_998 (.A(net126));
 sg13g2_antennanp ANTENNA_999 (.A(net126));
 sg13g2_antennanp ANTENNA_1000 (.A(net126));
 sg13g2_antennanp ANTENNA_1001 (.A(net126));
 sg13g2_antennanp ANTENNA_1002 (.A(net126));
 sg13g2_antennanp ANTENNA_1003 (.A(net128));
 sg13g2_antennanp ANTENNA_1004 (.A(net128));
 sg13g2_antennanp ANTENNA_1005 (.A(net128));
 sg13g2_antennanp ANTENNA_1006 (.A(net128));
 sg13g2_antennanp ANTENNA_1007 (.A(net128));
 sg13g2_antennanp ANTENNA_1008 (.A(net128));
 sg13g2_antennanp ANTENNA_1009 (.A(net128));
 sg13g2_antennanp ANTENNA_1010 (.A(net128));
 sg13g2_antennanp ANTENNA_1011 (.A(net128));
 sg13g2_antennanp ANTENNA_1012 (.A(net129));
 sg13g2_antennanp ANTENNA_1013 (.A(net129));
 sg13g2_antennanp ANTENNA_1014 (.A(net129));
 sg13g2_antennanp ANTENNA_1015 (.A(net129));
 sg13g2_antennanp ANTENNA_1016 (.A(net129));
 sg13g2_antennanp ANTENNA_1017 (.A(net129));
 sg13g2_antennanp ANTENNA_1018 (.A(net129));
 sg13g2_antennanp ANTENNA_1019 (.A(net129));
 sg13g2_antennanp ANTENNA_1020 (.A(net129));
 sg13g2_antennanp ANTENNA_1021 (.A(net129));
 sg13g2_antennanp ANTENNA_1022 (.A(net129));
 sg13g2_antennanp ANTENNA_1023 (.A(net129));
 sg13g2_antennanp ANTENNA_1024 (.A(net129));
 sg13g2_antennanp ANTENNA_1025 (.A(net129));
 sg13g2_antennanp ANTENNA_1026 (.A(net129));
 sg13g2_antennanp ANTENNA_1027 (.A(net129));
 sg13g2_antennanp ANTENNA_1028 (.A(net134));
 sg13g2_antennanp ANTENNA_1029 (.A(net134));
 sg13g2_antennanp ANTENNA_1030 (.A(net134));
 sg13g2_antennanp ANTENNA_1031 (.A(net134));
 sg13g2_antennanp ANTENNA_1032 (.A(net134));
 sg13g2_antennanp ANTENNA_1033 (.A(net134));
 sg13g2_antennanp ANTENNA_1034 (.A(net134));
 sg13g2_antennanp ANTENNA_1035 (.A(net134));
 sg13g2_antennanp ANTENNA_1036 (.A(net134));
 sg13g2_antennanp ANTENNA_1037 (.A(net142));
 sg13g2_antennanp ANTENNA_1038 (.A(net142));
 sg13g2_antennanp ANTENNA_1039 (.A(net142));
 sg13g2_antennanp ANTENNA_1040 (.A(net142));
 sg13g2_antennanp ANTENNA_1041 (.A(net142));
 sg13g2_antennanp ANTENNA_1042 (.A(net142));
 sg13g2_antennanp ANTENNA_1043 (.A(net142));
 sg13g2_antennanp ANTENNA_1044 (.A(net142));
 sg13g2_antennanp ANTENNA_1045 (.A(net142));
 sg13g2_antennanp ANTENNA_1046 (.A(net144));
 sg13g2_antennanp ANTENNA_1047 (.A(net144));
 sg13g2_antennanp ANTENNA_1048 (.A(net144));
 sg13g2_antennanp ANTENNA_1049 (.A(net144));
 sg13g2_antennanp ANTENNA_1050 (.A(net144));
 sg13g2_antennanp ANTENNA_1051 (.A(net144));
 sg13g2_antennanp ANTENNA_1052 (.A(net144));
 sg13g2_antennanp ANTENNA_1053 (.A(net144));
 sg13g2_antennanp ANTENNA_1054 (.A(net149));
 sg13g2_antennanp ANTENNA_1055 (.A(net149));
 sg13g2_antennanp ANTENNA_1056 (.A(net149));
 sg13g2_antennanp ANTENNA_1057 (.A(net149));
 sg13g2_antennanp ANTENNA_1058 (.A(net149));
 sg13g2_antennanp ANTENNA_1059 (.A(net149));
 sg13g2_antennanp ANTENNA_1060 (.A(net149));
 sg13g2_antennanp ANTENNA_1061 (.A(net149));
 sg13g2_antennanp ANTENNA_1062 (.A(net153));
 sg13g2_antennanp ANTENNA_1063 (.A(net153));
 sg13g2_antennanp ANTENNA_1064 (.A(net153));
 sg13g2_antennanp ANTENNA_1065 (.A(net153));
 sg13g2_antennanp ANTENNA_1066 (.A(net153));
 sg13g2_antennanp ANTENNA_1067 (.A(net153));
 sg13g2_antennanp ANTENNA_1068 (.A(net153));
 sg13g2_antennanp ANTENNA_1069 (.A(net153));
 sg13g2_antennanp ANTENNA_1070 (.A(net153));
 sg13g2_antennanp ANTENNA_1071 (.A(net161));
 sg13g2_antennanp ANTENNA_1072 (.A(net161));
 sg13g2_antennanp ANTENNA_1073 (.A(net161));
 sg13g2_antennanp ANTENNA_1074 (.A(net161));
 sg13g2_antennanp ANTENNA_1075 (.A(net161));
 sg13g2_antennanp ANTENNA_1076 (.A(net161));
 sg13g2_antennanp ANTENNA_1077 (.A(net161));
 sg13g2_antennanp ANTENNA_1078 (.A(net161));
 sg13g2_antennanp ANTENNA_1079 (.A(net161));
 sg13g2_antennanp ANTENNA_1080 (.A(net164));
 sg13g2_antennanp ANTENNA_1081 (.A(net164));
 sg13g2_antennanp ANTENNA_1082 (.A(net164));
 sg13g2_antennanp ANTENNA_1083 (.A(net164));
 sg13g2_antennanp ANTENNA_1084 (.A(net164));
 sg13g2_antennanp ANTENNA_1085 (.A(net164));
 sg13g2_antennanp ANTENNA_1086 (.A(net164));
 sg13g2_antennanp ANTENNA_1087 (.A(net164));
 sg13g2_antennanp ANTENNA_1088 (.A(net164));
 sg13g2_antennanp ANTENNA_1089 (.A(net167));
 sg13g2_antennanp ANTENNA_1090 (.A(net167));
 sg13g2_antennanp ANTENNA_1091 (.A(net167));
 sg13g2_antennanp ANTENNA_1092 (.A(net167));
 sg13g2_antennanp ANTENNA_1093 (.A(net167));
 sg13g2_antennanp ANTENNA_1094 (.A(net167));
 sg13g2_antennanp ANTENNA_1095 (.A(net167));
 sg13g2_antennanp ANTENNA_1096 (.A(net167));
 sg13g2_antennanp ANTENNA_1097 (.A(net168));
 sg13g2_antennanp ANTENNA_1098 (.A(net168));
 sg13g2_antennanp ANTENNA_1099 (.A(net168));
 sg13g2_antennanp ANTENNA_1100 (.A(net168));
 sg13g2_antennanp ANTENNA_1101 (.A(net168));
 sg13g2_antennanp ANTENNA_1102 (.A(net168));
 sg13g2_antennanp ANTENNA_1103 (.A(net168));
 sg13g2_antennanp ANTENNA_1104 (.A(net168));
 sg13g2_antennanp ANTENNA_1105 (.A(net168));
 sg13g2_antennanp ANTENNA_1106 (.A(net171));
 sg13g2_antennanp ANTENNA_1107 (.A(net171));
 sg13g2_antennanp ANTENNA_1108 (.A(net171));
 sg13g2_antennanp ANTENNA_1109 (.A(net171));
 sg13g2_antennanp ANTENNA_1110 (.A(net171));
 sg13g2_antennanp ANTENNA_1111 (.A(net171));
 sg13g2_antennanp ANTENNA_1112 (.A(net171));
 sg13g2_antennanp ANTENNA_1113 (.A(net171));
 sg13g2_antennanp ANTENNA_1114 (.A(net171));
 sg13g2_antennanp ANTENNA_1115 (.A(net172));
 sg13g2_antennanp ANTENNA_1116 (.A(net172));
 sg13g2_antennanp ANTENNA_1117 (.A(net172));
 sg13g2_antennanp ANTENNA_1118 (.A(net172));
 sg13g2_antennanp ANTENNA_1119 (.A(net172));
 sg13g2_antennanp ANTENNA_1120 (.A(net172));
 sg13g2_antennanp ANTENNA_1121 (.A(net172));
 sg13g2_antennanp ANTENNA_1122 (.A(net172));
 sg13g2_antennanp ANTENNA_1123 (.A(net174));
 sg13g2_antennanp ANTENNA_1124 (.A(net174));
 sg13g2_antennanp ANTENNA_1125 (.A(net174));
 sg13g2_antennanp ANTENNA_1126 (.A(net174));
 sg13g2_antennanp ANTENNA_1127 (.A(net174));
 sg13g2_antennanp ANTENNA_1128 (.A(net174));
 sg13g2_antennanp ANTENNA_1129 (.A(net174));
 sg13g2_antennanp ANTENNA_1130 (.A(net174));
 sg13g2_antennanp ANTENNA_1131 (.A(net174));
 sg13g2_antennanp ANTENNA_1132 (.A(net182));
 sg13g2_antennanp ANTENNA_1133 (.A(net182));
 sg13g2_antennanp ANTENNA_1134 (.A(net182));
 sg13g2_antennanp ANTENNA_1135 (.A(net182));
 sg13g2_antennanp ANTENNA_1136 (.A(net182));
 sg13g2_antennanp ANTENNA_1137 (.A(net182));
 sg13g2_antennanp ANTENNA_1138 (.A(net182));
 sg13g2_antennanp ANTENNA_1139 (.A(net182));
 sg13g2_antennanp ANTENNA_1140 (.A(net185));
 sg13g2_antennanp ANTENNA_1141 (.A(net185));
 sg13g2_antennanp ANTENNA_1142 (.A(net185));
 sg13g2_antennanp ANTENNA_1143 (.A(net185));
 sg13g2_antennanp ANTENNA_1144 (.A(net185));
 sg13g2_antennanp ANTENNA_1145 (.A(net185));
 sg13g2_antennanp ANTENNA_1146 (.A(net185));
 sg13g2_antennanp ANTENNA_1147 (.A(net185));
 sg13g2_antennanp ANTENNA_1148 (.A(net185));
 sg13g2_antennanp ANTENNA_1149 (.A(net185));
 sg13g2_antennanp ANTENNA_1150 (.A(net185));
 sg13g2_antennanp ANTENNA_1151 (.A(net198));
 sg13g2_antennanp ANTENNA_1152 (.A(net198));
 sg13g2_antennanp ANTENNA_1153 (.A(net198));
 sg13g2_antennanp ANTENNA_1154 (.A(net198));
 sg13g2_antennanp ANTENNA_1155 (.A(net198));
 sg13g2_antennanp ANTENNA_1156 (.A(net198));
 sg13g2_antennanp ANTENNA_1157 (.A(net198));
 sg13g2_antennanp ANTENNA_1158 (.A(net198));
 sg13g2_antennanp ANTENNA_1159 (.A(net198));
 sg13g2_antennanp ANTENNA_1160 (.A(net198));
 sg13g2_antennanp ANTENNA_1161 (.A(net198));
 sg13g2_antennanp ANTENNA_1162 (.A(net198));
 sg13g2_antennanp ANTENNA_1163 (.A(net198));
 sg13g2_antennanp ANTENNA_1164 (.A(net198));
 sg13g2_antennanp ANTENNA_1165 (.A(net198));
 sg13g2_antennanp ANTENNA_1166 (.A(net198));
 sg13g2_antennanp ANTENNA_1167 (.A(net203));
 sg13g2_antennanp ANTENNA_1168 (.A(net203));
 sg13g2_antennanp ANTENNA_1169 (.A(net203));
 sg13g2_antennanp ANTENNA_1170 (.A(net203));
 sg13g2_antennanp ANTENNA_1171 (.A(net203));
 sg13g2_antennanp ANTENNA_1172 (.A(net203));
 sg13g2_antennanp ANTENNA_1173 (.A(net203));
 sg13g2_antennanp ANTENNA_1174 (.A(net203));
 sg13g2_antennanp ANTENNA_1175 (.A(net203));
 sg13g2_antennanp ANTENNA_1176 (.A(net203));
 sg13g2_antennanp ANTENNA_1177 (.A(net203));
 sg13g2_antennanp ANTENNA_1178 (.A(net203));
 sg13g2_antennanp ANTENNA_1179 (.A(net203));
 sg13g2_antennanp ANTENNA_1180 (.A(net203));
 sg13g2_antennanp ANTENNA_1181 (.A(net203));
 sg13g2_antennanp ANTENNA_1182 (.A(net203));
 sg13g2_antennanp ANTENNA_1183 (.A(net203));
 sg13g2_antennanp ANTENNA_1184 (.A(net203));
 sg13g2_antennanp ANTENNA_1185 (.A(net203));
 sg13g2_antennanp ANTENNA_1186 (.A(net203));
 sg13g2_antennanp ANTENNA_1187 (.A(net205));
 sg13g2_antennanp ANTENNA_1188 (.A(net205));
 sg13g2_antennanp ANTENNA_1189 (.A(net205));
 sg13g2_antennanp ANTENNA_1190 (.A(net205));
 sg13g2_antennanp ANTENNA_1191 (.A(net205));
 sg13g2_antennanp ANTENNA_1192 (.A(net205));
 sg13g2_antennanp ANTENNA_1193 (.A(net205));
 sg13g2_antennanp ANTENNA_1194 (.A(net205));
 sg13g2_antennanp ANTENNA_1195 (.A(net205));
 sg13g2_antennanp ANTENNA_1196 (.A(net210));
 sg13g2_antennanp ANTENNA_1197 (.A(net210));
 sg13g2_antennanp ANTENNA_1198 (.A(net210));
 sg13g2_antennanp ANTENNA_1199 (.A(net210));
 sg13g2_antennanp ANTENNA_1200 (.A(net210));
 sg13g2_antennanp ANTENNA_1201 (.A(net210));
 sg13g2_antennanp ANTENNA_1202 (.A(net210));
 sg13g2_antennanp ANTENNA_1203 (.A(net210));
 sg13g2_antennanp ANTENNA_1204 (.A(net210));
 sg13g2_antennanp ANTENNA_1205 (.A(clknet_level_2_1_38_clk));
 sg13g2_antennanp ANTENNA_1206 (.A(clknet_level_2_1_38_clk));
 sg13g2_antennanp ANTENNA_1207 (.A(clknet_level_2_1_38_clk));
 sg13g2_antennanp ANTENNA_1208 (.A(clknet_level_2_1_38_clk));
 sg13g2_antennanp ANTENNA_1209 (.A(clknet_level_2_1_38_clk));
 sg13g2_antennanp ANTENNA_1210 (.A(clknet_level_2_1_38_clk));
 sg13g2_antennanp ANTENNA_1211 (.A(clknet_level_2_1_38_clk));
 sg13g2_antennanp ANTENNA_1212 (.A(clknet_level_2_1_38_clk));
 sg13g2_antennanp ANTENNA_1213 (.A(_0003_));
 sg13g2_antennanp ANTENNA_1214 (.A(_0016_));
 sg13g2_antennanp ANTENNA_1215 (.A(_0018_));
 sg13g2_antennanp ANTENNA_1216 (.A(_0018_));
 sg13g2_antennanp ANTENNA_1217 (.A(_0021_));
 sg13g2_antennanp ANTENNA_1218 (.A(_0022_));
 sg13g2_antennanp ANTENNA_1219 (.A(_0023_));
 sg13g2_antennanp ANTENNA_1220 (.A(_0024_));
 sg13g2_antennanp ANTENNA_1221 (.A(_0025_));
 sg13g2_antennanp ANTENNA_1222 (.A(_0025_));
 sg13g2_antennanp ANTENNA_1223 (.A(_0027_));
 sg13g2_antennanp ANTENNA_1224 (.A(_0027_));
 sg13g2_antennanp ANTENNA_1225 (.A(_0028_));
 sg13g2_antennanp ANTENNA_1226 (.A(_0028_));
 sg13g2_antennanp ANTENNA_1227 (.A(_0038_));
 sg13g2_antennanp ANTENNA_1228 (.A(_0038_));
 sg13g2_antennanp ANTENNA_1229 (.A(_0038_));
 sg13g2_antennanp ANTENNA_1230 (.A(_0038_));
 sg13g2_antennanp ANTENNA_1231 (.A(_0038_));
 sg13g2_antennanp ANTENNA_1232 (.A(_0038_));
 sg13g2_antennanp ANTENNA_1233 (.A(_0038_));
 sg13g2_antennanp ANTENNA_1234 (.A(_0038_));
 sg13g2_antennanp ANTENNA_1235 (.A(_0038_));
 sg13g2_antennanp ANTENNA_1236 (.A(_0090_));
 sg13g2_antennanp ANTENNA_1237 (.A(_0090_));
 sg13g2_antennanp ANTENNA_1238 (.A(_0090_));
 sg13g2_antennanp ANTENNA_1239 (.A(_0100_));
 sg13g2_antennanp ANTENNA_1240 (.A(_0100_));
 sg13g2_antennanp ANTENNA_1241 (.A(_0100_));
 sg13g2_antennanp ANTENNA_1242 (.A(_0100_));
 sg13g2_antennanp ANTENNA_1243 (.A(_0100_));
 sg13g2_antennanp ANTENNA_1244 (.A(_0123_));
 sg13g2_antennanp ANTENNA_1245 (.A(_0123_));
 sg13g2_antennanp ANTENNA_1246 (.A(_0125_));
 sg13g2_antennanp ANTENNA_1247 (.A(_0125_));
 sg13g2_antennanp ANTENNA_1248 (.A(_0125_));
 sg13g2_antennanp ANTENNA_1249 (.A(_0150_));
 sg13g2_antennanp ANTENNA_1250 (.A(_0150_));
 sg13g2_antennanp ANTENNA_1251 (.A(_0150_));
 sg13g2_antennanp ANTENNA_1252 (.A(_0150_));
 sg13g2_antennanp ANTENNA_1253 (.A(_0150_));
 sg13g2_antennanp ANTENNA_1254 (.A(_0150_));
 sg13g2_antennanp ANTENNA_1255 (.A(_0150_));
 sg13g2_antennanp ANTENNA_1256 (.A(_0150_));
 sg13g2_antennanp ANTENNA_1257 (.A(_0150_));
 sg13g2_antennanp ANTENNA_1258 (.A(_0158_));
 sg13g2_antennanp ANTENNA_1259 (.A(_0165_));
 sg13g2_antennanp ANTENNA_1260 (.A(_0165_));
 sg13g2_antennanp ANTENNA_1261 (.A(_0165_));
 sg13g2_antennanp ANTENNA_1262 (.A(_0165_));
 sg13g2_antennanp ANTENNA_1263 (.A(_0167_));
 sg13g2_antennanp ANTENNA_1264 (.A(_0167_));
 sg13g2_antennanp ANTENNA_1265 (.A(_0167_));
 sg13g2_antennanp ANTENNA_1266 (.A(_0167_));
 sg13g2_antennanp ANTENNA_1267 (.A(_0167_));
 sg13g2_antennanp ANTENNA_1268 (.A(_0167_));
 sg13g2_antennanp ANTENNA_1269 (.A(_0167_));
 sg13g2_antennanp ANTENNA_1270 (.A(_0167_));
 sg13g2_antennanp ANTENNA_1271 (.A(_0168_));
 sg13g2_antennanp ANTENNA_1272 (.A(_0168_));
 sg13g2_antennanp ANTENNA_1273 (.A(_0168_));
 sg13g2_antennanp ANTENNA_1274 (.A(_0168_));
 sg13g2_antennanp ANTENNA_1275 (.A(_0168_));
 sg13g2_antennanp ANTENNA_1276 (.A(_0168_));
 sg13g2_antennanp ANTENNA_1277 (.A(_0189_));
 sg13g2_antennanp ANTENNA_1278 (.A(_0230_));
 sg13g2_antennanp ANTENNA_1279 (.A(_0260_));
 sg13g2_antennanp ANTENNA_1280 (.A(_0260_));
 sg13g2_antennanp ANTENNA_1281 (.A(_0260_));
 sg13g2_antennanp ANTENNA_1282 (.A(_0260_));
 sg13g2_antennanp ANTENNA_1283 (.A(_0269_));
 sg13g2_antennanp ANTENNA_1284 (.A(_0301_));
 sg13g2_antennanp ANTENNA_1285 (.A(_0345_));
 sg13g2_antennanp ANTENNA_1286 (.A(_0345_));
 sg13g2_antennanp ANTENNA_1287 (.A(_0345_));
 sg13g2_antennanp ANTENNA_1288 (.A(_0345_));
 sg13g2_antennanp ANTENNA_1289 (.A(_0346_));
 sg13g2_antennanp ANTENNA_1290 (.A(_0346_));
 sg13g2_antennanp ANTENNA_1291 (.A(_0346_));
 sg13g2_antennanp ANTENNA_1292 (.A(_0346_));
 sg13g2_antennanp ANTENNA_1293 (.A(_0360_));
 sg13g2_antennanp ANTENNA_1294 (.A(_0360_));
 sg13g2_antennanp ANTENNA_1295 (.A(_0360_));
 sg13g2_antennanp ANTENNA_1296 (.A(_0360_));
 sg13g2_antennanp ANTENNA_1297 (.A(_0360_));
 sg13g2_antennanp ANTENNA_1298 (.A(_0387_));
 sg13g2_antennanp ANTENNA_1299 (.A(_0387_));
 sg13g2_antennanp ANTENNA_1300 (.A(_0387_));
 sg13g2_antennanp ANTENNA_1301 (.A(_0387_));
 sg13g2_antennanp ANTENNA_1302 (.A(_0387_));
 sg13g2_antennanp ANTENNA_1303 (.A(_0387_));
 sg13g2_antennanp ANTENNA_1304 (.A(_0435_));
 sg13g2_antennanp ANTENNA_1305 (.A(_0435_));
 sg13g2_antennanp ANTENNA_1306 (.A(_0438_));
 sg13g2_antennanp ANTENNA_1307 (.A(_0438_));
 sg13g2_antennanp ANTENNA_1308 (.A(_0438_));
 sg13g2_antennanp ANTENNA_1309 (.A(_0438_));
 sg13g2_antennanp ANTENNA_1310 (.A(_0438_));
 sg13g2_antennanp ANTENNA_1311 (.A(_0438_));
 sg13g2_antennanp ANTENNA_1312 (.A(_0448_));
 sg13g2_antennanp ANTENNA_1313 (.A(_0477_));
 sg13g2_antennanp ANTENNA_1314 (.A(_0477_));
 sg13g2_antennanp ANTENNA_1315 (.A(_0477_));
 sg13g2_antennanp ANTENNA_1316 (.A(_0477_));
 sg13g2_antennanp ANTENNA_1317 (.A(_0477_));
 sg13g2_antennanp ANTENNA_1318 (.A(_0477_));
 sg13g2_antennanp ANTENNA_1319 (.A(_0477_));
 sg13g2_antennanp ANTENNA_1320 (.A(_0490_));
 sg13g2_antennanp ANTENNA_1321 (.A(_0490_));
 sg13g2_antennanp ANTENNA_1322 (.A(_0507_));
 sg13g2_antennanp ANTENNA_1323 (.A(_0507_));
 sg13g2_antennanp ANTENNA_1324 (.A(_0511_));
 sg13g2_antennanp ANTENNA_1325 (.A(_0511_));
 sg13g2_antennanp ANTENNA_1326 (.A(_0511_));
 sg13g2_antennanp ANTENNA_1327 (.A(_0521_));
 sg13g2_antennanp ANTENNA_1328 (.A(_0521_));
 sg13g2_antennanp ANTENNA_1329 (.A(_0521_));
 sg13g2_antennanp ANTENNA_1330 (.A(_0597_));
 sg13g2_antennanp ANTENNA_1331 (.A(_0597_));
 sg13g2_antennanp ANTENNA_1332 (.A(_0597_));
 sg13g2_antennanp ANTENNA_1333 (.A(_0597_));
 sg13g2_antennanp ANTENNA_1334 (.A(_0597_));
 sg13g2_antennanp ANTENNA_1335 (.A(_0598_));
 sg13g2_antennanp ANTENNA_1336 (.A(_0598_));
 sg13g2_antennanp ANTENNA_1337 (.A(_0598_));
 sg13g2_antennanp ANTENNA_1338 (.A(_0598_));
 sg13g2_antennanp ANTENNA_1339 (.A(_0598_));
 sg13g2_antennanp ANTENNA_1340 (.A(_0623_));
 sg13g2_antennanp ANTENNA_1341 (.A(_0780_));
 sg13g2_antennanp ANTENNA_1342 (.A(_0800_));
 sg13g2_antennanp ANTENNA_1343 (.A(_0824_));
 sg13g2_antennanp ANTENNA_1344 (.A(_0824_));
 sg13g2_antennanp ANTENNA_1345 (.A(_0824_));
 sg13g2_antennanp ANTENNA_1346 (.A(_0866_));
 sg13g2_antennanp ANTENNA_1347 (.A(_0866_));
 sg13g2_antennanp ANTENNA_1348 (.A(_0866_));
 sg13g2_antennanp ANTENNA_1349 (.A(_0878_));
 sg13g2_antennanp ANTENNA_1350 (.A(_0878_));
 sg13g2_antennanp ANTENNA_1351 (.A(_0878_));
 sg13g2_antennanp ANTENNA_1352 (.A(_0878_));
 sg13g2_antennanp ANTENNA_1353 (.A(_0878_));
 sg13g2_antennanp ANTENNA_1354 (.A(_0878_));
 sg13g2_antennanp ANTENNA_1355 (.A(_0878_));
 sg13g2_antennanp ANTENNA_1356 (.A(_0878_));
 sg13g2_antennanp ANTENNA_1357 (.A(_0878_));
 sg13g2_antennanp ANTENNA_1358 (.A(_1002_));
 sg13g2_antennanp ANTENNA_1359 (.A(_1002_));
 sg13g2_antennanp ANTENNA_1360 (.A(_1071_));
 sg13g2_antennanp ANTENNA_1361 (.A(_1071_));
 sg13g2_antennanp ANTENNA_1362 (.A(_1071_));
 sg13g2_antennanp ANTENNA_1363 (.A(_1085_));
 sg13g2_antennanp ANTENNA_1364 (.A(_1085_));
 sg13g2_antennanp ANTENNA_1365 (.A(_1085_));
 sg13g2_antennanp ANTENNA_1366 (.A(_1085_));
 sg13g2_antennanp ANTENNA_1367 (.A(_1085_));
 sg13g2_antennanp ANTENNA_1368 (.A(_1085_));
 sg13g2_antennanp ANTENNA_1369 (.A(_1151_));
 sg13g2_antennanp ANTENNA_1370 (.A(_1151_));
 sg13g2_antennanp ANTENNA_1371 (.A(_1151_));
 sg13g2_antennanp ANTENNA_1372 (.A(_1151_));
 sg13g2_antennanp ANTENNA_1373 (.A(_1151_));
 sg13g2_antennanp ANTENNA_1374 (.A(_1151_));
 sg13g2_antennanp ANTENNA_1375 (.A(_1162_));
 sg13g2_antennanp ANTENNA_1376 (.A(_1162_));
 sg13g2_antennanp ANTENNA_1377 (.A(_1162_));
 sg13g2_antennanp ANTENNA_1378 (.A(_1162_));
 sg13g2_antennanp ANTENNA_1379 (.A(_1162_));
 sg13g2_antennanp ANTENNA_1380 (.A(_1162_));
 sg13g2_antennanp ANTENNA_1381 (.A(_1162_));
 sg13g2_antennanp ANTENNA_1382 (.A(_1162_));
 sg13g2_antennanp ANTENNA_1383 (.A(_1225_));
 sg13g2_antennanp ANTENNA_1384 (.A(_1225_));
 sg13g2_antennanp ANTENNA_1385 (.A(_1292_));
 sg13g2_antennanp ANTENNA_1386 (.A(_1292_));
 sg13g2_antennanp ANTENNA_1387 (.A(_1326_));
 sg13g2_antennanp ANTENNA_1388 (.A(_1326_));
 sg13g2_antennanp ANTENNA_1389 (.A(_1326_));
 sg13g2_antennanp ANTENNA_1390 (.A(_1326_));
 sg13g2_antennanp ANTENNA_1391 (.A(_1326_));
 sg13g2_antennanp ANTENNA_1392 (.A(_1326_));
 sg13g2_antennanp ANTENNA_1393 (.A(_1326_));
 sg13g2_antennanp ANTENNA_1394 (.A(_1363_));
 sg13g2_antennanp ANTENNA_1395 (.A(_1411_));
 sg13g2_antennanp ANTENNA_1396 (.A(_1439_));
 sg13g2_antennanp ANTENNA_1397 (.A(_1470_));
 sg13g2_antennanp ANTENNA_1398 (.A(_1470_));
 sg13g2_antennanp ANTENNA_1399 (.A(_1519_));
 sg13g2_antennanp ANTENNA_1400 (.A(_1531_));
 sg13g2_antennanp ANTENNA_1401 (.A(_1531_));
 sg13g2_antennanp ANTENNA_1402 (.A(_1532_));
 sg13g2_antennanp ANTENNA_1403 (.A(_1532_));
 sg13g2_antennanp ANTENNA_1404 (.A(_1532_));
 sg13g2_antennanp ANTENNA_1405 (.A(_1544_));
 sg13g2_antennanp ANTENNA_1406 (.A(_1544_));
 sg13g2_antennanp ANTENNA_1407 (.A(_1544_));
 sg13g2_antennanp ANTENNA_1408 (.A(_1544_));
 sg13g2_antennanp ANTENNA_1409 (.A(_1544_));
 sg13g2_antennanp ANTENNA_1410 (.A(_1544_));
 sg13g2_antennanp ANTENNA_1411 (.A(_1544_));
 sg13g2_antennanp ANTENNA_1412 (.A(_1544_));
 sg13g2_antennanp ANTENNA_1413 (.A(_1553_));
 sg13g2_antennanp ANTENNA_1414 (.A(_1631_));
 sg13g2_antennanp ANTENNA_1415 (.A(_1631_));
 sg13g2_antennanp ANTENNA_1416 (.A(_1631_));
 sg13g2_antennanp ANTENNA_1417 (.A(_1631_));
 sg13g2_antennanp ANTENNA_1418 (.A(_1631_));
 sg13g2_antennanp ANTENNA_1419 (.A(_1631_));
 sg13g2_antennanp ANTENNA_1420 (.A(_1631_));
 sg13g2_antennanp ANTENNA_1421 (.A(_1631_));
 sg13g2_antennanp ANTENNA_1422 (.A(_1685_));
 sg13g2_antennanp ANTENNA_1423 (.A(_1685_));
 sg13g2_antennanp ANTENNA_1424 (.A(_1685_));
 sg13g2_antennanp ANTENNA_1425 (.A(_1685_));
 sg13g2_antennanp ANTENNA_1426 (.A(_1696_));
 sg13g2_antennanp ANTENNA_1427 (.A(_1696_));
 sg13g2_antennanp ANTENNA_1428 (.A(_1696_));
 sg13g2_antennanp ANTENNA_1429 (.A(_1696_));
 sg13g2_antennanp ANTENNA_1430 (.A(_1696_));
 sg13g2_antennanp ANTENNA_1431 (.A(_1696_));
 sg13g2_antennanp ANTENNA_1432 (.A(_1696_));
 sg13g2_antennanp ANTENNA_1433 (.A(_1696_));
 sg13g2_antennanp ANTENNA_1434 (.A(_1696_));
 sg13g2_antennanp ANTENNA_1435 (.A(_1696_));
 sg13g2_antennanp ANTENNA_1436 (.A(_1707_));
 sg13g2_antennanp ANTENNA_1437 (.A(_1707_));
 sg13g2_antennanp ANTENNA_1438 (.A(_1707_));
 sg13g2_antennanp ANTENNA_1439 (.A(_1707_));
 sg13g2_antennanp ANTENNA_1440 (.A(_1707_));
 sg13g2_antennanp ANTENNA_1441 (.A(_1716_));
 sg13g2_antennanp ANTENNA_1442 (.A(_1735_));
 sg13g2_antennanp ANTENNA_1443 (.A(_1735_));
 sg13g2_antennanp ANTENNA_1444 (.A(_1761_));
 sg13g2_antennanp ANTENNA_1445 (.A(_1761_));
 sg13g2_antennanp ANTENNA_1446 (.A(_2014_));
 sg13g2_antennanp ANTENNA_1447 (.A(_2014_));
 sg13g2_antennanp ANTENNA_1448 (.A(_2020_));
 sg13g2_antennanp ANTENNA_1449 (.A(_2020_));
 sg13g2_antennanp ANTENNA_1450 (.A(_2020_));
 sg13g2_antennanp ANTENNA_1451 (.A(_2020_));
 sg13g2_antennanp ANTENNA_1452 (.A(_2020_));
 sg13g2_antennanp ANTENNA_1453 (.A(_2020_));
 sg13g2_antennanp ANTENNA_1454 (.A(_2020_));
 sg13g2_antennanp ANTENNA_1455 (.A(_2020_));
 sg13g2_antennanp ANTENNA_1456 (.A(_2037_));
 sg13g2_antennanp ANTENNA_1457 (.A(_2053_));
 sg13g2_antennanp ANTENNA_1458 (.A(_2053_));
 sg13g2_antennanp ANTENNA_1459 (.A(_2053_));
 sg13g2_antennanp ANTENNA_1460 (.A(_2097_));
 sg13g2_antennanp ANTENNA_1461 (.A(_2097_));
 sg13g2_antennanp ANTENNA_1462 (.A(_2097_));
 sg13g2_antennanp ANTENNA_1463 (.A(_2097_));
 sg13g2_antennanp ANTENNA_1464 (.A(_2097_));
 sg13g2_antennanp ANTENNA_1465 (.A(_2110_));
 sg13g2_antennanp ANTENNA_1466 (.A(_2110_));
 sg13g2_antennanp ANTENNA_1467 (.A(_2112_));
 sg13g2_antennanp ANTENNA_1468 (.A(_2145_));
 sg13g2_antennanp ANTENNA_1469 (.A(_2171_));
 sg13g2_antennanp ANTENNA_1470 (.A(_2171_));
 sg13g2_antennanp ANTENNA_1471 (.A(_2171_));
 sg13g2_antennanp ANTENNA_1472 (.A(_2171_));
 sg13g2_antennanp ANTENNA_1473 (.A(_2171_));
 sg13g2_antennanp ANTENNA_1474 (.A(_2171_));
 sg13g2_antennanp ANTENNA_1475 (.A(_2171_));
 sg13g2_antennanp ANTENNA_1476 (.A(_2171_));
 sg13g2_antennanp ANTENNA_1477 (.A(_2171_));
 sg13g2_antennanp ANTENNA_1478 (.A(_2172_));
 sg13g2_antennanp ANTENNA_1479 (.A(_2172_));
 sg13g2_antennanp ANTENNA_1480 (.A(_2172_));
 sg13g2_antennanp ANTENNA_1481 (.A(_2172_));
 sg13g2_antennanp ANTENNA_1482 (.A(_2172_));
 sg13g2_antennanp ANTENNA_1483 (.A(_2172_));
 sg13g2_antennanp ANTENNA_1484 (.A(_2172_));
 sg13g2_antennanp ANTENNA_1485 (.A(_2172_));
 sg13g2_antennanp ANTENNA_1486 (.A(_2172_));
 sg13g2_antennanp ANTENNA_1487 (.A(_2172_));
 sg13g2_antennanp ANTENNA_1488 (.A(_2257_));
 sg13g2_antennanp ANTENNA_1489 (.A(_2257_));
 sg13g2_antennanp ANTENNA_1490 (.A(_2408_));
 sg13g2_antennanp ANTENNA_1491 (.A(_2408_));
 sg13g2_antennanp ANTENNA_1492 (.A(_2408_));
 sg13g2_antennanp ANTENNA_1493 (.A(_2430_));
 sg13g2_antennanp ANTENNA_1494 (.A(_2430_));
 sg13g2_antennanp ANTENNA_1495 (.A(_2430_));
 sg13g2_antennanp ANTENNA_1496 (.A(_2430_));
 sg13g2_antennanp ANTENNA_1497 (.A(_2430_));
 sg13g2_antennanp ANTENNA_1498 (.A(_2430_));
 sg13g2_antennanp ANTENNA_1499 (.A(_2444_));
 sg13g2_antennanp ANTENNA_1500 (.A(_2444_));
 sg13g2_antennanp ANTENNA_1501 (.A(_2444_));
 sg13g2_antennanp ANTENNA_1502 (.A(_2444_));
 sg13g2_antennanp ANTENNA_1503 (.A(_2444_));
 sg13g2_antennanp ANTENNA_1504 (.A(_2444_));
 sg13g2_antennanp ANTENNA_1505 (.A(_2444_));
 sg13g2_antennanp ANTENNA_1506 (.A(_2461_));
 sg13g2_antennanp ANTENNA_1507 (.A(_2461_));
 sg13g2_antennanp ANTENNA_1508 (.A(_2461_));
 sg13g2_antennanp ANTENNA_1509 (.A(_2461_));
 sg13g2_antennanp ANTENNA_1510 (.A(_2461_));
 sg13g2_antennanp ANTENNA_1511 (.A(_2467_));
 sg13g2_antennanp ANTENNA_1512 (.A(_2467_));
 sg13g2_antennanp ANTENNA_1513 (.A(_2467_));
 sg13g2_antennanp ANTENNA_1514 (.A(_2467_));
 sg13g2_antennanp ANTENNA_1515 (.A(_2467_));
 sg13g2_antennanp ANTENNA_1516 (.A(_2470_));
 sg13g2_antennanp ANTENNA_1517 (.A(_2470_));
 sg13g2_antennanp ANTENNA_1518 (.A(_2470_));
 sg13g2_antennanp ANTENNA_1519 (.A(_2470_));
 sg13g2_antennanp ANTENNA_1520 (.A(_2480_));
 sg13g2_antennanp ANTENNA_1521 (.A(_2480_));
 sg13g2_antennanp ANTENNA_1522 (.A(_2480_));
 sg13g2_antennanp ANTENNA_1523 (.A(_2480_));
 sg13g2_antennanp ANTENNA_1524 (.A(_2480_));
 sg13g2_antennanp ANTENNA_1525 (.A(_2482_));
 sg13g2_antennanp ANTENNA_1526 (.A(_2482_));
 sg13g2_antennanp ANTENNA_1527 (.A(_2482_));
 sg13g2_antennanp ANTENNA_1528 (.A(_2482_));
 sg13g2_antennanp ANTENNA_1529 (.A(_2482_));
 sg13g2_antennanp ANTENNA_1530 (.A(_2482_));
 sg13g2_antennanp ANTENNA_1531 (.A(_2482_));
 sg13g2_antennanp ANTENNA_1532 (.A(_2487_));
 sg13g2_antennanp ANTENNA_1533 (.A(_2487_));
 sg13g2_antennanp ANTENNA_1534 (.A(_2501_));
 sg13g2_antennanp ANTENNA_1535 (.A(_2501_));
 sg13g2_antennanp ANTENNA_1536 (.A(_2501_));
 sg13g2_antennanp ANTENNA_1537 (.A(_2520_));
 sg13g2_antennanp ANTENNA_1538 (.A(_2520_));
 sg13g2_antennanp ANTENNA_1539 (.A(_2520_));
 sg13g2_antennanp ANTENNA_1540 (.A(_2520_));
 sg13g2_antennanp ANTENNA_1541 (.A(_2520_));
 sg13g2_antennanp ANTENNA_1542 (.A(_2520_));
 sg13g2_antennanp ANTENNA_1543 (.A(_2530_));
 sg13g2_antennanp ANTENNA_1544 (.A(_2530_));
 sg13g2_antennanp ANTENNA_1545 (.A(_2530_));
 sg13g2_antennanp ANTENNA_1546 (.A(_2530_));
 sg13g2_antennanp ANTENNA_1547 (.A(_2532_));
 sg13g2_antennanp ANTENNA_1548 (.A(_2532_));
 sg13g2_antennanp ANTENNA_1549 (.A(_2532_));
 sg13g2_antennanp ANTENNA_1550 (.A(_2532_));
 sg13g2_antennanp ANTENNA_1551 (.A(_2532_));
 sg13g2_antennanp ANTENNA_1552 (.A(_2537_));
 sg13g2_antennanp ANTENNA_1553 (.A(_2537_));
 sg13g2_antennanp ANTENNA_1554 (.A(_2537_));
 sg13g2_antennanp ANTENNA_1555 (.A(_2537_));
 sg13g2_antennanp ANTENNA_1556 (.A(_2573_));
 sg13g2_antennanp ANTENNA_1557 (.A(_2573_));
 sg13g2_antennanp ANTENNA_1558 (.A(_2573_));
 sg13g2_antennanp ANTENNA_1559 (.A(_2573_));
 sg13g2_antennanp ANTENNA_1560 (.A(_2577_));
 sg13g2_antennanp ANTENNA_1561 (.A(_2577_));
 sg13g2_antennanp ANTENNA_1562 (.A(_2577_));
 sg13g2_antennanp ANTENNA_1563 (.A(_2577_));
 sg13g2_antennanp ANTENNA_1564 (.A(_2577_));
 sg13g2_antennanp ANTENNA_1565 (.A(_2577_));
 sg13g2_antennanp ANTENNA_1566 (.A(_2577_));
 sg13g2_antennanp ANTENNA_1567 (.A(_2577_));
 sg13g2_antennanp ANTENNA_1568 (.A(_2585_));
 sg13g2_antennanp ANTENNA_1569 (.A(_2585_));
 sg13g2_antennanp ANTENNA_1570 (.A(_2585_));
 sg13g2_antennanp ANTENNA_1571 (.A(_2588_));
 sg13g2_antennanp ANTENNA_1572 (.A(_2595_));
 sg13g2_antennanp ANTENNA_1573 (.A(_2595_));
 sg13g2_antennanp ANTENNA_1574 (.A(_2595_));
 sg13g2_antennanp ANTENNA_1575 (.A(_2600_));
 sg13g2_antennanp ANTENNA_1576 (.A(_2600_));
 sg13g2_antennanp ANTENNA_1577 (.A(_2600_));
 sg13g2_antennanp ANTENNA_1578 (.A(_2600_));
 sg13g2_antennanp ANTENNA_1579 (.A(_2601_));
 sg13g2_antennanp ANTENNA_1580 (.A(_2601_));
 sg13g2_antennanp ANTENNA_1581 (.A(_2601_));
 sg13g2_antennanp ANTENNA_1582 (.A(_2601_));
 sg13g2_antennanp ANTENNA_1583 (.A(_2607_));
 sg13g2_antennanp ANTENNA_1584 (.A(_2607_));
 sg13g2_antennanp ANTENNA_1585 (.A(_2615_));
 sg13g2_antennanp ANTENNA_1586 (.A(_2615_));
 sg13g2_antennanp ANTENNA_1587 (.A(_2615_));
 sg13g2_antennanp ANTENNA_1588 (.A(_2619_));
 sg13g2_antennanp ANTENNA_1589 (.A(_2619_));
 sg13g2_antennanp ANTENNA_1590 (.A(_2619_));
 sg13g2_antennanp ANTENNA_1591 (.A(_2619_));
 sg13g2_antennanp ANTENNA_1592 (.A(_2619_));
 sg13g2_antennanp ANTENNA_1593 (.A(_2619_));
 sg13g2_antennanp ANTENNA_1594 (.A(_2619_));
 sg13g2_antennanp ANTENNA_1595 (.A(_2619_));
 sg13g2_antennanp ANTENNA_1596 (.A(_2619_));
 sg13g2_antennanp ANTENNA_1597 (.A(_2622_));
 sg13g2_antennanp ANTENNA_1598 (.A(_2622_));
 sg13g2_antennanp ANTENNA_1599 (.A(_2622_));
 sg13g2_antennanp ANTENNA_1600 (.A(_2622_));
 sg13g2_antennanp ANTENNA_1601 (.A(_2622_));
 sg13g2_antennanp ANTENNA_1602 (.A(_2622_));
 sg13g2_antennanp ANTENNA_1603 (.A(_2625_));
 sg13g2_antennanp ANTENNA_1604 (.A(_2625_));
 sg13g2_antennanp ANTENNA_1605 (.A(_2625_));
 sg13g2_antennanp ANTENNA_1606 (.A(_2625_));
 sg13g2_antennanp ANTENNA_1607 (.A(_2659_));
 sg13g2_antennanp ANTENNA_1608 (.A(_2659_));
 sg13g2_antennanp ANTENNA_1609 (.A(_2659_));
 sg13g2_antennanp ANTENNA_1610 (.A(_2659_));
 sg13g2_antennanp ANTENNA_1611 (.A(_2659_));
 sg13g2_antennanp ANTENNA_1612 (.A(_2665_));
 sg13g2_antennanp ANTENNA_1613 (.A(_2665_));
 sg13g2_antennanp ANTENNA_1614 (.A(_2665_));
 sg13g2_antennanp ANTENNA_1615 (.A(_2665_));
 sg13g2_antennanp ANTENNA_1616 (.A(_2678_));
 sg13g2_antennanp ANTENNA_1617 (.A(_2678_));
 sg13g2_antennanp ANTENNA_1618 (.A(_2678_));
 sg13g2_antennanp ANTENNA_1619 (.A(_2678_));
 sg13g2_antennanp ANTENNA_1620 (.A(_2678_));
 sg13g2_antennanp ANTENNA_1621 (.A(_2678_));
 sg13g2_antennanp ANTENNA_1622 (.A(_2678_));
 sg13g2_antennanp ANTENNA_1623 (.A(_2681_));
 sg13g2_antennanp ANTENNA_1624 (.A(_2681_));
 sg13g2_antennanp ANTENNA_1625 (.A(_2681_));
 sg13g2_antennanp ANTENNA_1626 (.A(_2681_));
 sg13g2_antennanp ANTENNA_1627 (.A(_2732_));
 sg13g2_antennanp ANTENNA_1628 (.A(_2732_));
 sg13g2_antennanp ANTENNA_1629 (.A(_2732_));
 sg13g2_antennanp ANTENNA_1630 (.A(_2733_));
 sg13g2_antennanp ANTENNA_1631 (.A(_2733_));
 sg13g2_antennanp ANTENNA_1632 (.A(_2733_));
 sg13g2_antennanp ANTENNA_1633 (.A(_2733_));
 sg13g2_antennanp ANTENNA_1634 (.A(_2739_));
 sg13g2_antennanp ANTENNA_1635 (.A(_2739_));
 sg13g2_antennanp ANTENNA_1636 (.A(_2739_));
 sg13g2_antennanp ANTENNA_1637 (.A(_2739_));
 sg13g2_antennanp ANTENNA_1638 (.A(_2769_));
 sg13g2_antennanp ANTENNA_1639 (.A(_2769_));
 sg13g2_antennanp ANTENNA_1640 (.A(_2769_));
 sg13g2_antennanp ANTENNA_1641 (.A(_2769_));
 sg13g2_antennanp ANTENNA_1642 (.A(_2779_));
 sg13g2_antennanp ANTENNA_1643 (.A(_2779_));
 sg13g2_antennanp ANTENNA_1644 (.A(_2779_));
 sg13g2_antennanp ANTENNA_1645 (.A(_2779_));
 sg13g2_antennanp ANTENNA_1646 (.A(_2789_));
 sg13g2_antennanp ANTENNA_1647 (.A(_2789_));
 sg13g2_antennanp ANTENNA_1648 (.A(_2789_));
 sg13g2_antennanp ANTENNA_1649 (.A(_2789_));
 sg13g2_antennanp ANTENNA_1650 (.A(_2805_));
 sg13g2_antennanp ANTENNA_1651 (.A(_2805_));
 sg13g2_antennanp ANTENNA_1652 (.A(_2808_));
 sg13g2_antennanp ANTENNA_1653 (.A(_2808_));
 sg13g2_antennanp ANTENNA_1654 (.A(_2808_));
 sg13g2_antennanp ANTENNA_1655 (.A(_2808_));
 sg13g2_antennanp ANTENNA_1656 (.A(_2816_));
 sg13g2_antennanp ANTENNA_1657 (.A(_2816_));
 sg13g2_antennanp ANTENNA_1658 (.A(_2816_));
 sg13g2_antennanp ANTENNA_1659 (.A(_2816_));
 sg13g2_antennanp ANTENNA_1660 (.A(_2826_));
 sg13g2_antennanp ANTENNA_1661 (.A(_2826_));
 sg13g2_antennanp ANTENNA_1662 (.A(_2826_));
 sg13g2_antennanp ANTENNA_1663 (.A(_2826_));
 sg13g2_antennanp ANTENNA_1664 (.A(_2858_));
 sg13g2_antennanp ANTENNA_1665 (.A(_2858_));
 sg13g2_antennanp ANTENNA_1666 (.A(_2879_));
 sg13g2_antennanp ANTENNA_1667 (.A(_2879_));
 sg13g2_antennanp ANTENNA_1668 (.A(_2879_));
 sg13g2_antennanp ANTENNA_1669 (.A(_2879_));
 sg13g2_antennanp ANTENNA_1670 (.A(_2879_));
 sg13g2_antennanp ANTENNA_1671 (.A(_2879_));
 sg13g2_antennanp ANTENNA_1672 (.A(_2879_));
 sg13g2_antennanp ANTENNA_1673 (.A(_2879_));
 sg13g2_antennanp ANTENNA_1674 (.A(_2914_));
 sg13g2_antennanp ANTENNA_1675 (.A(_2914_));
 sg13g2_antennanp ANTENNA_1676 (.A(_2931_));
 sg13g2_antennanp ANTENNA_1677 (.A(_2931_));
 sg13g2_antennanp ANTENNA_1678 (.A(_2931_));
 sg13g2_antennanp ANTENNA_1679 (.A(_2931_));
 sg13g2_antennanp ANTENNA_1680 (.A(_2936_));
 sg13g2_antennanp ANTENNA_1681 (.A(_2936_));
 sg13g2_antennanp ANTENNA_1682 (.A(_2936_));
 sg13g2_antennanp ANTENNA_1683 (.A(_2957_));
 sg13g2_antennanp ANTENNA_1684 (.A(_2957_));
 sg13g2_antennanp ANTENNA_1685 (.A(_2957_));
 sg13g2_antennanp ANTENNA_1686 (.A(_2957_));
 sg13g2_antennanp ANTENNA_1687 (.A(_2967_));
 sg13g2_antennanp ANTENNA_1688 (.A(_2967_));
 sg13g2_antennanp ANTENNA_1689 (.A(_2967_));
 sg13g2_antennanp ANTENNA_1690 (.A(_2967_));
 sg13g2_antennanp ANTENNA_1691 (.A(_2967_));
 sg13g2_antennanp ANTENNA_1692 (.A(_2970_));
 sg13g2_antennanp ANTENNA_1693 (.A(_2970_));
 sg13g2_antennanp ANTENNA_1694 (.A(_2970_));
 sg13g2_antennanp ANTENNA_1695 (.A(_2970_));
 sg13g2_antennanp ANTENNA_1696 (.A(_2970_));
 sg13g2_antennanp ANTENNA_1697 (.A(_2970_));
 sg13g2_antennanp ANTENNA_1698 (.A(_2970_));
 sg13g2_antennanp ANTENNA_1699 (.A(_2974_));
 sg13g2_antennanp ANTENNA_1700 (.A(_2977_));
 sg13g2_antennanp ANTENNA_1701 (.A(_2977_));
 sg13g2_antennanp ANTENNA_1702 (.A(_2977_));
 sg13g2_antennanp ANTENNA_1703 (.A(_2977_));
 sg13g2_antennanp ANTENNA_1704 (.A(_2977_));
 sg13g2_antennanp ANTENNA_1705 (.A(_2986_));
 sg13g2_antennanp ANTENNA_1706 (.A(_2986_));
 sg13g2_antennanp ANTENNA_1707 (.A(_2986_));
 sg13g2_antennanp ANTENNA_1708 (.A(_2986_));
 sg13g2_antennanp ANTENNA_1709 (.A(_3018_));
 sg13g2_antennanp ANTENNA_1710 (.A(_3018_));
 sg13g2_antennanp ANTENNA_1711 (.A(_3018_));
 sg13g2_antennanp ANTENNA_1712 (.A(_3040_));
 sg13g2_antennanp ANTENNA_1713 (.A(_3040_));
 sg13g2_antennanp ANTENNA_1714 (.A(_3040_));
 sg13g2_antennanp ANTENNA_1715 (.A(clk));
 sg13g2_antennanp ANTENNA_1716 (.A(clk));
 sg13g2_antennanp ANTENNA_1717 (.A(net22));
 sg13g2_antennanp ANTENNA_1718 (.A(net22));
 sg13g2_antennanp ANTENNA_1719 (.A(net22));
 sg13g2_antennanp ANTENNA_1720 (.A(net22));
 sg13g2_antennanp ANTENNA_1721 (.A(net22));
 sg13g2_antennanp ANTENNA_1722 (.A(net22));
 sg13g2_antennanp ANTENNA_1723 (.A(net22));
 sg13g2_antennanp ANTENNA_1724 (.A(net22));
 sg13g2_antennanp ANTENNA_1725 (.A(net22));
 sg13g2_antennanp ANTENNA_1726 (.A(net23));
 sg13g2_antennanp ANTENNA_1727 (.A(net23));
 sg13g2_antennanp ANTENNA_1728 (.A(net23));
 sg13g2_antennanp ANTENNA_1729 (.A(net23));
 sg13g2_antennanp ANTENNA_1730 (.A(net23));
 sg13g2_antennanp ANTENNA_1731 (.A(net23));
 sg13g2_antennanp ANTENNA_1732 (.A(net23));
 sg13g2_antennanp ANTENNA_1733 (.A(net23));
 sg13g2_antennanp ANTENNA_1734 (.A(net29));
 sg13g2_antennanp ANTENNA_1735 (.A(net29));
 sg13g2_antennanp ANTENNA_1736 (.A(net29));
 sg13g2_antennanp ANTENNA_1737 (.A(net29));
 sg13g2_antennanp ANTENNA_1738 (.A(net29));
 sg13g2_antennanp ANTENNA_1739 (.A(net29));
 sg13g2_antennanp ANTENNA_1740 (.A(net29));
 sg13g2_antennanp ANTENNA_1741 (.A(net29));
 sg13g2_antennanp ANTENNA_1742 (.A(net29));
 sg13g2_antennanp ANTENNA_1743 (.A(net35));
 sg13g2_antennanp ANTENNA_1744 (.A(net35));
 sg13g2_antennanp ANTENNA_1745 (.A(net35));
 sg13g2_antennanp ANTENNA_1746 (.A(net35));
 sg13g2_antennanp ANTENNA_1747 (.A(net35));
 sg13g2_antennanp ANTENNA_1748 (.A(net35));
 sg13g2_antennanp ANTENNA_1749 (.A(net35));
 sg13g2_antennanp ANTENNA_1750 (.A(net35));
 sg13g2_antennanp ANTENNA_1751 (.A(net35));
 sg13g2_antennanp ANTENNA_1752 (.A(net40));
 sg13g2_antennanp ANTENNA_1753 (.A(net40));
 sg13g2_antennanp ANTENNA_1754 (.A(net40));
 sg13g2_antennanp ANTENNA_1755 (.A(net40));
 sg13g2_antennanp ANTENNA_1756 (.A(net40));
 sg13g2_antennanp ANTENNA_1757 (.A(net40));
 sg13g2_antennanp ANTENNA_1758 (.A(net40));
 sg13g2_antennanp ANTENNA_1759 (.A(net40));
 sg13g2_antennanp ANTENNA_1760 (.A(net40));
 sg13g2_antennanp ANTENNA_1761 (.A(net41));
 sg13g2_antennanp ANTENNA_1762 (.A(net41));
 sg13g2_antennanp ANTENNA_1763 (.A(net41));
 sg13g2_antennanp ANTENNA_1764 (.A(net41));
 sg13g2_antennanp ANTENNA_1765 (.A(net41));
 sg13g2_antennanp ANTENNA_1766 (.A(net41));
 sg13g2_antennanp ANTENNA_1767 (.A(net41));
 sg13g2_antennanp ANTENNA_1768 (.A(net41));
 sg13g2_antennanp ANTENNA_1769 (.A(net41));
 sg13g2_antennanp ANTENNA_1770 (.A(net46));
 sg13g2_antennanp ANTENNA_1771 (.A(net46));
 sg13g2_antennanp ANTENNA_1772 (.A(net46));
 sg13g2_antennanp ANTENNA_1773 (.A(net46));
 sg13g2_antennanp ANTENNA_1774 (.A(net46));
 sg13g2_antennanp ANTENNA_1775 (.A(net46));
 sg13g2_antennanp ANTENNA_1776 (.A(net46));
 sg13g2_antennanp ANTENNA_1777 (.A(net46));
 sg13g2_antennanp ANTENNA_1778 (.A(net46));
 sg13g2_antennanp ANTENNA_1779 (.A(net53));
 sg13g2_antennanp ANTENNA_1780 (.A(net53));
 sg13g2_antennanp ANTENNA_1781 (.A(net53));
 sg13g2_antennanp ANTENNA_1782 (.A(net53));
 sg13g2_antennanp ANTENNA_1783 (.A(net53));
 sg13g2_antennanp ANTENNA_1784 (.A(net53));
 sg13g2_antennanp ANTENNA_1785 (.A(net53));
 sg13g2_antennanp ANTENNA_1786 (.A(net53));
 sg13g2_antennanp ANTENNA_1787 (.A(net53));
 sg13g2_antennanp ANTENNA_1788 (.A(net59));
 sg13g2_antennanp ANTENNA_1789 (.A(net59));
 sg13g2_antennanp ANTENNA_1790 (.A(net59));
 sg13g2_antennanp ANTENNA_1791 (.A(net59));
 sg13g2_antennanp ANTENNA_1792 (.A(net59));
 sg13g2_antennanp ANTENNA_1793 (.A(net59));
 sg13g2_antennanp ANTENNA_1794 (.A(net59));
 sg13g2_antennanp ANTENNA_1795 (.A(net59));
 sg13g2_antennanp ANTENNA_1796 (.A(net59));
 sg13g2_antennanp ANTENNA_1797 (.A(net61));
 sg13g2_antennanp ANTENNA_1798 (.A(net61));
 sg13g2_antennanp ANTENNA_1799 (.A(net61));
 sg13g2_antennanp ANTENNA_1800 (.A(net61));
 sg13g2_antennanp ANTENNA_1801 (.A(net61));
 sg13g2_antennanp ANTENNA_1802 (.A(net61));
 sg13g2_antennanp ANTENNA_1803 (.A(net61));
 sg13g2_antennanp ANTENNA_1804 (.A(net61));
 sg13g2_antennanp ANTENNA_1805 (.A(net61));
 sg13g2_antennanp ANTENNA_1806 (.A(net61));
 sg13g2_antennanp ANTENNA_1807 (.A(net61));
 sg13g2_antennanp ANTENNA_1808 (.A(net61));
 sg13g2_antennanp ANTENNA_1809 (.A(net61));
 sg13g2_antennanp ANTENNA_1810 (.A(net61));
 sg13g2_antennanp ANTENNA_1811 (.A(net62));
 sg13g2_antennanp ANTENNA_1812 (.A(net62));
 sg13g2_antennanp ANTENNA_1813 (.A(net62));
 sg13g2_antennanp ANTENNA_1814 (.A(net62));
 sg13g2_antennanp ANTENNA_1815 (.A(net62));
 sg13g2_antennanp ANTENNA_1816 (.A(net62));
 sg13g2_antennanp ANTENNA_1817 (.A(net62));
 sg13g2_antennanp ANTENNA_1818 (.A(net62));
 sg13g2_antennanp ANTENNA_1819 (.A(net62));
 sg13g2_antennanp ANTENNA_1820 (.A(net64));
 sg13g2_antennanp ANTENNA_1821 (.A(net64));
 sg13g2_antennanp ANTENNA_1822 (.A(net64));
 sg13g2_antennanp ANTENNA_1823 (.A(net64));
 sg13g2_antennanp ANTENNA_1824 (.A(net64));
 sg13g2_antennanp ANTENNA_1825 (.A(net64));
 sg13g2_antennanp ANTENNA_1826 (.A(net64));
 sg13g2_antennanp ANTENNA_1827 (.A(net64));
 sg13g2_antennanp ANTENNA_1828 (.A(net70));
 sg13g2_antennanp ANTENNA_1829 (.A(net70));
 sg13g2_antennanp ANTENNA_1830 (.A(net70));
 sg13g2_antennanp ANTENNA_1831 (.A(net70));
 sg13g2_antennanp ANTENNA_1832 (.A(net70));
 sg13g2_antennanp ANTENNA_1833 (.A(net70));
 sg13g2_antennanp ANTENNA_1834 (.A(net70));
 sg13g2_antennanp ANTENNA_1835 (.A(net70));
 sg13g2_antennanp ANTENNA_1836 (.A(net70));
 sg13g2_antennanp ANTENNA_1837 (.A(net71));
 sg13g2_antennanp ANTENNA_1838 (.A(net71));
 sg13g2_antennanp ANTENNA_1839 (.A(net71));
 sg13g2_antennanp ANTENNA_1840 (.A(net71));
 sg13g2_antennanp ANTENNA_1841 (.A(net71));
 sg13g2_antennanp ANTENNA_1842 (.A(net71));
 sg13g2_antennanp ANTENNA_1843 (.A(net71));
 sg13g2_antennanp ANTENNA_1844 (.A(net71));
 sg13g2_antennanp ANTENNA_1845 (.A(net71));
 sg13g2_antennanp ANTENNA_1846 (.A(net71));
 sg13g2_antennanp ANTENNA_1847 (.A(net71));
 sg13g2_antennanp ANTENNA_1848 (.A(net71));
 sg13g2_antennanp ANTENNA_1849 (.A(net71));
 sg13g2_antennanp ANTENNA_1850 (.A(net71));
 sg13g2_antennanp ANTENNA_1851 (.A(net71));
 sg13g2_antennanp ANTENNA_1852 (.A(net71));
 sg13g2_antennanp ANTENNA_1853 (.A(net76));
 sg13g2_antennanp ANTENNA_1854 (.A(net76));
 sg13g2_antennanp ANTENNA_1855 (.A(net76));
 sg13g2_antennanp ANTENNA_1856 (.A(net76));
 sg13g2_antennanp ANTENNA_1857 (.A(net76));
 sg13g2_antennanp ANTENNA_1858 (.A(net76));
 sg13g2_antennanp ANTENNA_1859 (.A(net76));
 sg13g2_antennanp ANTENNA_1860 (.A(net76));
 sg13g2_antennanp ANTENNA_1861 (.A(net76));
 sg13g2_antennanp ANTENNA_1862 (.A(net78));
 sg13g2_antennanp ANTENNA_1863 (.A(net78));
 sg13g2_antennanp ANTENNA_1864 (.A(net78));
 sg13g2_antennanp ANTENNA_1865 (.A(net78));
 sg13g2_antennanp ANTENNA_1866 (.A(net78));
 sg13g2_antennanp ANTENNA_1867 (.A(net78));
 sg13g2_antennanp ANTENNA_1868 (.A(net78));
 sg13g2_antennanp ANTENNA_1869 (.A(net78));
 sg13g2_antennanp ANTENNA_1870 (.A(net78));
 sg13g2_antennanp ANTENNA_1871 (.A(net79));
 sg13g2_antennanp ANTENNA_1872 (.A(net79));
 sg13g2_antennanp ANTENNA_1873 (.A(net79));
 sg13g2_antennanp ANTENNA_1874 (.A(net79));
 sg13g2_antennanp ANTENNA_1875 (.A(net79));
 sg13g2_antennanp ANTENNA_1876 (.A(net79));
 sg13g2_antennanp ANTENNA_1877 (.A(net79));
 sg13g2_antennanp ANTENNA_1878 (.A(net79));
 sg13g2_antennanp ANTENNA_1879 (.A(net79));
 sg13g2_antennanp ANTENNA_1880 (.A(net79));
 sg13g2_antennanp ANTENNA_1881 (.A(net79));
 sg13g2_antennanp ANTENNA_1882 (.A(net79));
 sg13g2_antennanp ANTENNA_1883 (.A(net79));
 sg13g2_antennanp ANTENNA_1884 (.A(net79));
 sg13g2_antennanp ANTENNA_1885 (.A(net84));
 sg13g2_antennanp ANTENNA_1886 (.A(net84));
 sg13g2_antennanp ANTENNA_1887 (.A(net84));
 sg13g2_antennanp ANTENNA_1888 (.A(net84));
 sg13g2_antennanp ANTENNA_1889 (.A(net84));
 sg13g2_antennanp ANTENNA_1890 (.A(net84));
 sg13g2_antennanp ANTENNA_1891 (.A(net84));
 sg13g2_antennanp ANTENNA_1892 (.A(net84));
 sg13g2_antennanp ANTENNA_1893 (.A(net89));
 sg13g2_antennanp ANTENNA_1894 (.A(net89));
 sg13g2_antennanp ANTENNA_1895 (.A(net89));
 sg13g2_antennanp ANTENNA_1896 (.A(net89));
 sg13g2_antennanp ANTENNA_1897 (.A(net89));
 sg13g2_antennanp ANTENNA_1898 (.A(net89));
 sg13g2_antennanp ANTENNA_1899 (.A(net89));
 sg13g2_antennanp ANTENNA_1900 (.A(net89));
 sg13g2_antennanp ANTENNA_1901 (.A(net89));
 sg13g2_antennanp ANTENNA_1902 (.A(net91));
 sg13g2_antennanp ANTENNA_1903 (.A(net91));
 sg13g2_antennanp ANTENNA_1904 (.A(net91));
 sg13g2_antennanp ANTENNA_1905 (.A(net91));
 sg13g2_antennanp ANTENNA_1906 (.A(net91));
 sg13g2_antennanp ANTENNA_1907 (.A(net91));
 sg13g2_antennanp ANTENNA_1908 (.A(net91));
 sg13g2_antennanp ANTENNA_1909 (.A(net91));
 sg13g2_antennanp ANTENNA_1910 (.A(net94));
 sg13g2_antennanp ANTENNA_1911 (.A(net94));
 sg13g2_antennanp ANTENNA_1912 (.A(net94));
 sg13g2_antennanp ANTENNA_1913 (.A(net94));
 sg13g2_antennanp ANTENNA_1914 (.A(net94));
 sg13g2_antennanp ANTENNA_1915 (.A(net94));
 sg13g2_antennanp ANTENNA_1916 (.A(net94));
 sg13g2_antennanp ANTENNA_1917 (.A(net94));
 sg13g2_antennanp ANTENNA_1918 (.A(net100));
 sg13g2_antennanp ANTENNA_1919 (.A(net100));
 sg13g2_antennanp ANTENNA_1920 (.A(net100));
 sg13g2_antennanp ANTENNA_1921 (.A(net100));
 sg13g2_antennanp ANTENNA_1922 (.A(net100));
 sg13g2_antennanp ANTENNA_1923 (.A(net100));
 sg13g2_antennanp ANTENNA_1924 (.A(net100));
 sg13g2_antennanp ANTENNA_1925 (.A(net100));
 sg13g2_antennanp ANTENNA_1926 (.A(net100));
 sg13g2_antennanp ANTENNA_1927 (.A(net100));
 sg13g2_antennanp ANTENNA_1928 (.A(net100));
 sg13g2_antennanp ANTENNA_1929 (.A(net100));
 sg13g2_antennanp ANTENNA_1930 (.A(net100));
 sg13g2_antennanp ANTENNA_1931 (.A(net100));
 sg13g2_antennanp ANTENNA_1932 (.A(net100));
 sg13g2_antennanp ANTENNA_1933 (.A(net100));
 sg13g2_antennanp ANTENNA_1934 (.A(net100));
 sg13g2_antennanp ANTENNA_1935 (.A(net100));
 sg13g2_antennanp ANTENNA_1936 (.A(net101));
 sg13g2_antennanp ANTENNA_1937 (.A(net101));
 sg13g2_antennanp ANTENNA_1938 (.A(net101));
 sg13g2_antennanp ANTENNA_1939 (.A(net101));
 sg13g2_antennanp ANTENNA_1940 (.A(net101));
 sg13g2_antennanp ANTENNA_1941 (.A(net101));
 sg13g2_antennanp ANTENNA_1942 (.A(net101));
 sg13g2_antennanp ANTENNA_1943 (.A(net101));
 sg13g2_antennanp ANTENNA_1944 (.A(net101));
 sg13g2_antennanp ANTENNA_1945 (.A(net106));
 sg13g2_antennanp ANTENNA_1946 (.A(net106));
 sg13g2_antennanp ANTENNA_1947 (.A(net106));
 sg13g2_antennanp ANTENNA_1948 (.A(net106));
 sg13g2_antennanp ANTENNA_1949 (.A(net106));
 sg13g2_antennanp ANTENNA_1950 (.A(net106));
 sg13g2_antennanp ANTENNA_1951 (.A(net106));
 sg13g2_antennanp ANTENNA_1952 (.A(net106));
 sg13g2_antennanp ANTENNA_1953 (.A(net106));
 sg13g2_antennanp ANTENNA_1954 (.A(net107));
 sg13g2_antennanp ANTENNA_1955 (.A(net107));
 sg13g2_antennanp ANTENNA_1956 (.A(net107));
 sg13g2_antennanp ANTENNA_1957 (.A(net107));
 sg13g2_antennanp ANTENNA_1958 (.A(net107));
 sg13g2_antennanp ANTENNA_1959 (.A(net107));
 sg13g2_antennanp ANTENNA_1960 (.A(net107));
 sg13g2_antennanp ANTENNA_1961 (.A(net107));
 sg13g2_antennanp ANTENNA_1962 (.A(net107));
 sg13g2_antennanp ANTENNA_1963 (.A(net113));
 sg13g2_antennanp ANTENNA_1964 (.A(net113));
 sg13g2_antennanp ANTENNA_1965 (.A(net113));
 sg13g2_antennanp ANTENNA_1966 (.A(net113));
 sg13g2_antennanp ANTENNA_1967 (.A(net113));
 sg13g2_antennanp ANTENNA_1968 (.A(net113));
 sg13g2_antennanp ANTENNA_1969 (.A(net113));
 sg13g2_antennanp ANTENNA_1970 (.A(net113));
 sg13g2_antennanp ANTENNA_1971 (.A(net125));
 sg13g2_antennanp ANTENNA_1972 (.A(net125));
 sg13g2_antennanp ANTENNA_1973 (.A(net125));
 sg13g2_antennanp ANTENNA_1974 (.A(net125));
 sg13g2_antennanp ANTENNA_1975 (.A(net125));
 sg13g2_antennanp ANTENNA_1976 (.A(net125));
 sg13g2_antennanp ANTENNA_1977 (.A(net125));
 sg13g2_antennanp ANTENNA_1978 (.A(net125));
 sg13g2_antennanp ANTENNA_1979 (.A(net125));
 sg13g2_antennanp ANTENNA_1980 (.A(net128));
 sg13g2_antennanp ANTENNA_1981 (.A(net128));
 sg13g2_antennanp ANTENNA_1982 (.A(net128));
 sg13g2_antennanp ANTENNA_1983 (.A(net128));
 sg13g2_antennanp ANTENNA_1984 (.A(net128));
 sg13g2_antennanp ANTENNA_1985 (.A(net128));
 sg13g2_antennanp ANTENNA_1986 (.A(net128));
 sg13g2_antennanp ANTENNA_1987 (.A(net128));
 sg13g2_antennanp ANTENNA_1988 (.A(net128));
 sg13g2_antennanp ANTENNA_1989 (.A(net128));
 sg13g2_antennanp ANTENNA_1990 (.A(net128));
 sg13g2_antennanp ANTENNA_1991 (.A(net128));
 sg13g2_antennanp ANTENNA_1992 (.A(net128));
 sg13g2_antennanp ANTENNA_1993 (.A(net128));
 sg13g2_antennanp ANTENNA_1994 (.A(net128));
 sg13g2_antennanp ANTENNA_1995 (.A(net128));
 sg13g2_antennanp ANTENNA_1996 (.A(net128));
 sg13g2_antennanp ANTENNA_1997 (.A(net129));
 sg13g2_antennanp ANTENNA_1998 (.A(net129));
 sg13g2_antennanp ANTENNA_1999 (.A(net129));
 sg13g2_antennanp ANTENNA_2000 (.A(net129));
 sg13g2_antennanp ANTENNA_2001 (.A(net129));
 sg13g2_antennanp ANTENNA_2002 (.A(net129));
 sg13g2_antennanp ANTENNA_2003 (.A(net129));
 sg13g2_antennanp ANTENNA_2004 (.A(net129));
 sg13g2_antennanp ANTENNA_2005 (.A(net129));
 sg13g2_antennanp ANTENNA_2006 (.A(net134));
 sg13g2_antennanp ANTENNA_2007 (.A(net134));
 sg13g2_antennanp ANTENNA_2008 (.A(net134));
 sg13g2_antennanp ANTENNA_2009 (.A(net134));
 sg13g2_antennanp ANTENNA_2010 (.A(net134));
 sg13g2_antennanp ANTENNA_2011 (.A(net134));
 sg13g2_antennanp ANTENNA_2012 (.A(net134));
 sg13g2_antennanp ANTENNA_2013 (.A(net134));
 sg13g2_antennanp ANTENNA_2014 (.A(net134));
 sg13g2_antennanp ANTENNA_2015 (.A(net134));
 sg13g2_antennanp ANTENNA_2016 (.A(net134));
 sg13g2_antennanp ANTENNA_2017 (.A(net134));
 sg13g2_antennanp ANTENNA_2018 (.A(net134));
 sg13g2_antennanp ANTENNA_2019 (.A(net142));
 sg13g2_antennanp ANTENNA_2020 (.A(net142));
 sg13g2_antennanp ANTENNA_2021 (.A(net142));
 sg13g2_antennanp ANTENNA_2022 (.A(net142));
 sg13g2_antennanp ANTENNA_2023 (.A(net142));
 sg13g2_antennanp ANTENNA_2024 (.A(net142));
 sg13g2_antennanp ANTENNA_2025 (.A(net142));
 sg13g2_antennanp ANTENNA_2026 (.A(net142));
 sg13g2_antennanp ANTENNA_2027 (.A(net142));
 sg13g2_antennanp ANTENNA_2028 (.A(net144));
 sg13g2_antennanp ANTENNA_2029 (.A(net144));
 sg13g2_antennanp ANTENNA_2030 (.A(net144));
 sg13g2_antennanp ANTENNA_2031 (.A(net144));
 sg13g2_antennanp ANTENNA_2032 (.A(net144));
 sg13g2_antennanp ANTENNA_2033 (.A(net144));
 sg13g2_antennanp ANTENNA_2034 (.A(net144));
 sg13g2_antennanp ANTENNA_2035 (.A(net144));
 sg13g2_antennanp ANTENNA_2036 (.A(net153));
 sg13g2_antennanp ANTENNA_2037 (.A(net153));
 sg13g2_antennanp ANTENNA_2038 (.A(net153));
 sg13g2_antennanp ANTENNA_2039 (.A(net153));
 sg13g2_antennanp ANTENNA_2040 (.A(net153));
 sg13g2_antennanp ANTENNA_2041 (.A(net153));
 sg13g2_antennanp ANTENNA_2042 (.A(net153));
 sg13g2_antennanp ANTENNA_2043 (.A(net153));
 sg13g2_antennanp ANTENNA_2044 (.A(net153));
 sg13g2_antennanp ANTENNA_2045 (.A(net161));
 sg13g2_antennanp ANTENNA_2046 (.A(net161));
 sg13g2_antennanp ANTENNA_2047 (.A(net161));
 sg13g2_antennanp ANTENNA_2048 (.A(net161));
 sg13g2_antennanp ANTENNA_2049 (.A(net161));
 sg13g2_antennanp ANTENNA_2050 (.A(net161));
 sg13g2_antennanp ANTENNA_2051 (.A(net161));
 sg13g2_antennanp ANTENNA_2052 (.A(net161));
 sg13g2_antennanp ANTENNA_2053 (.A(net161));
 sg13g2_antennanp ANTENNA_2054 (.A(net164));
 sg13g2_antennanp ANTENNA_2055 (.A(net164));
 sg13g2_antennanp ANTENNA_2056 (.A(net164));
 sg13g2_antennanp ANTENNA_2057 (.A(net164));
 sg13g2_antennanp ANTENNA_2058 (.A(net164));
 sg13g2_antennanp ANTENNA_2059 (.A(net164));
 sg13g2_antennanp ANTENNA_2060 (.A(net164));
 sg13g2_antennanp ANTENNA_2061 (.A(net164));
 sg13g2_antennanp ANTENNA_2062 (.A(net164));
 sg13g2_antennanp ANTENNA_2063 (.A(net167));
 sg13g2_antennanp ANTENNA_2064 (.A(net167));
 sg13g2_antennanp ANTENNA_2065 (.A(net167));
 sg13g2_antennanp ANTENNA_2066 (.A(net167));
 sg13g2_antennanp ANTENNA_2067 (.A(net167));
 sg13g2_antennanp ANTENNA_2068 (.A(net167));
 sg13g2_antennanp ANTENNA_2069 (.A(net167));
 sg13g2_antennanp ANTENNA_2070 (.A(net167));
 sg13g2_antennanp ANTENNA_2071 (.A(net167));
 sg13g2_antennanp ANTENNA_2072 (.A(net171));
 sg13g2_antennanp ANTENNA_2073 (.A(net171));
 sg13g2_antennanp ANTENNA_2074 (.A(net171));
 sg13g2_antennanp ANTENNA_2075 (.A(net171));
 sg13g2_antennanp ANTENNA_2076 (.A(net171));
 sg13g2_antennanp ANTENNA_2077 (.A(net171));
 sg13g2_antennanp ANTENNA_2078 (.A(net171));
 sg13g2_antennanp ANTENNA_2079 (.A(net171));
 sg13g2_antennanp ANTENNA_2080 (.A(net171));
 sg13g2_antennanp ANTENNA_2081 (.A(net174));
 sg13g2_antennanp ANTENNA_2082 (.A(net174));
 sg13g2_antennanp ANTENNA_2083 (.A(net174));
 sg13g2_antennanp ANTENNA_2084 (.A(net174));
 sg13g2_antennanp ANTENNA_2085 (.A(net174));
 sg13g2_antennanp ANTENNA_2086 (.A(net174));
 sg13g2_antennanp ANTENNA_2087 (.A(net174));
 sg13g2_antennanp ANTENNA_2088 (.A(net174));
 sg13g2_antennanp ANTENNA_2089 (.A(net174));
 sg13g2_antennanp ANTENNA_2090 (.A(net182));
 sg13g2_antennanp ANTENNA_2091 (.A(net182));
 sg13g2_antennanp ANTENNA_2092 (.A(net182));
 sg13g2_antennanp ANTENNA_2093 (.A(net182));
 sg13g2_antennanp ANTENNA_2094 (.A(net182));
 sg13g2_antennanp ANTENNA_2095 (.A(net182));
 sg13g2_antennanp ANTENNA_2096 (.A(net182));
 sg13g2_antennanp ANTENNA_2097 (.A(net182));
 sg13g2_antennanp ANTENNA_2098 (.A(net185));
 sg13g2_antennanp ANTENNA_2099 (.A(net185));
 sg13g2_antennanp ANTENNA_2100 (.A(net185));
 sg13g2_antennanp ANTENNA_2101 (.A(net185));
 sg13g2_antennanp ANTENNA_2102 (.A(net185));
 sg13g2_antennanp ANTENNA_2103 (.A(net185));
 sg13g2_antennanp ANTENNA_2104 (.A(net185));
 sg13g2_antennanp ANTENNA_2105 (.A(net185));
 sg13g2_antennanp ANTENNA_2106 (.A(net185));
 sg13g2_antennanp ANTENNA_2107 (.A(net198));
 sg13g2_antennanp ANTENNA_2108 (.A(net198));
 sg13g2_antennanp ANTENNA_2109 (.A(net198));
 sg13g2_antennanp ANTENNA_2110 (.A(net198));
 sg13g2_antennanp ANTENNA_2111 (.A(net198));
 sg13g2_antennanp ANTENNA_2112 (.A(net198));
 sg13g2_antennanp ANTENNA_2113 (.A(net198));
 sg13g2_antennanp ANTENNA_2114 (.A(net198));
 sg13g2_antennanp ANTENNA_2115 (.A(net210));
 sg13g2_antennanp ANTENNA_2116 (.A(net210));
 sg13g2_antennanp ANTENNA_2117 (.A(net210));
 sg13g2_antennanp ANTENNA_2118 (.A(net210));
 sg13g2_antennanp ANTENNA_2119 (.A(net210));
 sg13g2_antennanp ANTENNA_2120 (.A(net210));
 sg13g2_antennanp ANTENNA_2121 (.A(net210));
 sg13g2_antennanp ANTENNA_2122 (.A(net210));
 sg13g2_antennanp ANTENNA_2123 (.A(net210));
 sg13g2_antennanp ANTENNA_2124 (.A(_0003_));
 sg13g2_antennanp ANTENNA_2125 (.A(_0016_));
 sg13g2_antennanp ANTENNA_2126 (.A(_0016_));
 sg13g2_antennanp ANTENNA_2127 (.A(_0018_));
 sg13g2_antennanp ANTENNA_2128 (.A(_0018_));
 sg13g2_antennanp ANTENNA_2129 (.A(_0021_));
 sg13g2_antennanp ANTENNA_2130 (.A(_0022_));
 sg13g2_antennanp ANTENNA_2131 (.A(_0023_));
 sg13g2_antennanp ANTENNA_2132 (.A(_0024_));
 sg13g2_antennanp ANTENNA_2133 (.A(_0025_));
 sg13g2_antennanp ANTENNA_2134 (.A(_0025_));
 sg13g2_antennanp ANTENNA_2135 (.A(_0027_));
 sg13g2_antennanp ANTENNA_2136 (.A(_0027_));
 sg13g2_antennanp ANTENNA_2137 (.A(_0028_));
 sg13g2_antennanp ANTENNA_2138 (.A(_0028_));
 sg13g2_antennanp ANTENNA_2139 (.A(_0038_));
 sg13g2_antennanp ANTENNA_2140 (.A(_0038_));
 sg13g2_antennanp ANTENNA_2141 (.A(_0038_));
 sg13g2_antennanp ANTENNA_2142 (.A(_0038_));
 sg13g2_antennanp ANTENNA_2143 (.A(_0038_));
 sg13g2_antennanp ANTENNA_2144 (.A(_0038_));
 sg13g2_antennanp ANTENNA_2145 (.A(_0038_));
 sg13g2_antennanp ANTENNA_2146 (.A(_0038_));
 sg13g2_antennanp ANTENNA_2147 (.A(_0038_));
 sg13g2_antennanp ANTENNA_2148 (.A(_0123_));
 sg13g2_antennanp ANTENNA_2149 (.A(_0123_));
 sg13g2_antennanp ANTENNA_2150 (.A(_0125_));
 sg13g2_antennanp ANTENNA_2151 (.A(_0125_));
 sg13g2_antennanp ANTENNA_2152 (.A(_0125_));
 sg13g2_antennanp ANTENNA_2153 (.A(_0150_));
 sg13g2_antennanp ANTENNA_2154 (.A(_0150_));
 sg13g2_antennanp ANTENNA_2155 (.A(_0150_));
 sg13g2_antennanp ANTENNA_2156 (.A(_0150_));
 sg13g2_antennanp ANTENNA_2157 (.A(_0150_));
 sg13g2_antennanp ANTENNA_2158 (.A(_0158_));
 sg13g2_antennanp ANTENNA_2159 (.A(_0165_));
 sg13g2_antennanp ANTENNA_2160 (.A(_0165_));
 sg13g2_antennanp ANTENNA_2161 (.A(_0165_));
 sg13g2_antennanp ANTENNA_2162 (.A(_0165_));
 sg13g2_antennanp ANTENNA_2163 (.A(_0167_));
 sg13g2_antennanp ANTENNA_2164 (.A(_0167_));
 sg13g2_antennanp ANTENNA_2165 (.A(_0167_));
 sg13g2_antennanp ANTENNA_2166 (.A(_0167_));
 sg13g2_antennanp ANTENNA_2167 (.A(_0167_));
 sg13g2_antennanp ANTENNA_2168 (.A(_0167_));
 sg13g2_antennanp ANTENNA_2169 (.A(_0167_));
 sg13g2_antennanp ANTENNA_2170 (.A(_0167_));
 sg13g2_antennanp ANTENNA_2171 (.A(_0168_));
 sg13g2_antennanp ANTENNA_2172 (.A(_0168_));
 sg13g2_antennanp ANTENNA_2173 (.A(_0168_));
 sg13g2_antennanp ANTENNA_2174 (.A(_0168_));
 sg13g2_antennanp ANTENNA_2175 (.A(_0168_));
 sg13g2_antennanp ANTENNA_2176 (.A(_0168_));
 sg13g2_antennanp ANTENNA_2177 (.A(_0189_));
 sg13g2_antennanp ANTENNA_2178 (.A(_0230_));
 sg13g2_antennanp ANTENNA_2179 (.A(_0230_));
 sg13g2_antennanp ANTENNA_2180 (.A(_0260_));
 sg13g2_antennanp ANTENNA_2181 (.A(_0260_));
 sg13g2_antennanp ANTENNA_2182 (.A(_0260_));
 sg13g2_antennanp ANTENNA_2183 (.A(_0260_));
 sg13g2_antennanp ANTENNA_2184 (.A(_0269_));
 sg13g2_antennanp ANTENNA_2185 (.A(_0301_));
 sg13g2_antennanp ANTENNA_2186 (.A(_0345_));
 sg13g2_antennanp ANTENNA_2187 (.A(_0345_));
 sg13g2_antennanp ANTENNA_2188 (.A(_0345_));
 sg13g2_antennanp ANTENNA_2189 (.A(_0345_));
 sg13g2_antennanp ANTENNA_2190 (.A(_0346_));
 sg13g2_antennanp ANTENNA_2191 (.A(_0346_));
 sg13g2_antennanp ANTENNA_2192 (.A(_0346_));
 sg13g2_antennanp ANTENNA_2193 (.A(_0346_));
 sg13g2_antennanp ANTENNA_2194 (.A(_0360_));
 sg13g2_antennanp ANTENNA_2195 (.A(_0360_));
 sg13g2_antennanp ANTENNA_2196 (.A(_0360_));
 sg13g2_antennanp ANTENNA_2197 (.A(_0360_));
 sg13g2_antennanp ANTENNA_2198 (.A(_0360_));
 sg13g2_antennanp ANTENNA_2199 (.A(_0387_));
 sg13g2_antennanp ANTENNA_2200 (.A(_0387_));
 sg13g2_antennanp ANTENNA_2201 (.A(_0387_));
 sg13g2_antennanp ANTENNA_2202 (.A(_0387_));
 sg13g2_antennanp ANTENNA_2203 (.A(_0387_));
 sg13g2_antennanp ANTENNA_2204 (.A(_0387_));
 sg13g2_antennanp ANTENNA_2205 (.A(_0435_));
 sg13g2_antennanp ANTENNA_2206 (.A(_0435_));
 sg13g2_antennanp ANTENNA_2207 (.A(_0438_));
 sg13g2_antennanp ANTENNA_2208 (.A(_0438_));
 sg13g2_antennanp ANTENNA_2209 (.A(_0438_));
 sg13g2_antennanp ANTENNA_2210 (.A(_0438_));
 sg13g2_antennanp ANTENNA_2211 (.A(_0438_));
 sg13g2_antennanp ANTENNA_2212 (.A(_0438_));
 sg13g2_antennanp ANTENNA_2213 (.A(_0448_));
 sg13g2_antennanp ANTENNA_2214 (.A(_0477_));
 sg13g2_antennanp ANTENNA_2215 (.A(_0477_));
 sg13g2_antennanp ANTENNA_2216 (.A(_0477_));
 sg13g2_antennanp ANTENNA_2217 (.A(_0477_));
 sg13g2_antennanp ANTENNA_2218 (.A(_0477_));
 sg13g2_antennanp ANTENNA_2219 (.A(_0477_));
 sg13g2_antennanp ANTENNA_2220 (.A(_0477_));
 sg13g2_antennanp ANTENNA_2221 (.A(_0507_));
 sg13g2_antennanp ANTENNA_2222 (.A(_0507_));
 sg13g2_antennanp ANTENNA_2223 (.A(_0511_));
 sg13g2_antennanp ANTENNA_2224 (.A(_0511_));
 sg13g2_antennanp ANTENNA_2225 (.A(_0511_));
 sg13g2_antennanp ANTENNA_2226 (.A(_0521_));
 sg13g2_antennanp ANTENNA_2227 (.A(_0521_));
 sg13g2_antennanp ANTENNA_2228 (.A(_0521_));
 sg13g2_antennanp ANTENNA_2229 (.A(_0597_));
 sg13g2_antennanp ANTENNA_2230 (.A(_0597_));
 sg13g2_antennanp ANTENNA_2231 (.A(_0597_));
 sg13g2_antennanp ANTENNA_2232 (.A(_0597_));
 sg13g2_antennanp ANTENNA_2233 (.A(_0597_));
 sg13g2_antennanp ANTENNA_2234 (.A(_0598_));
 sg13g2_antennanp ANTENNA_2235 (.A(_0598_));
 sg13g2_antennanp ANTENNA_2236 (.A(_0598_));
 sg13g2_antennanp ANTENNA_2237 (.A(_0598_));
 sg13g2_antennanp ANTENNA_2238 (.A(_0598_));
 sg13g2_antennanp ANTENNA_2239 (.A(_0623_));
 sg13g2_antennanp ANTENNA_2240 (.A(_0780_));
 sg13g2_antennanp ANTENNA_2241 (.A(_0800_));
 sg13g2_antennanp ANTENNA_2242 (.A(_0866_));
 sg13g2_antennanp ANTENNA_2243 (.A(_0866_));
 sg13g2_antennanp ANTENNA_2244 (.A(_0866_));
 sg13g2_antennanp ANTENNA_2245 (.A(_0878_));
 sg13g2_antennanp ANTENNA_2246 (.A(_0878_));
 sg13g2_antennanp ANTENNA_2247 (.A(_0878_));
 sg13g2_antennanp ANTENNA_2248 (.A(_0878_));
 sg13g2_antennanp ANTENNA_2249 (.A(_0878_));
 sg13g2_antennanp ANTENNA_2250 (.A(_0878_));
 sg13g2_antennanp ANTENNA_2251 (.A(_0878_));
 sg13g2_antennanp ANTENNA_2252 (.A(_0878_));
 sg13g2_antennanp ANTENNA_2253 (.A(_0878_));
 sg13g2_antennanp ANTENNA_2254 (.A(_1002_));
 sg13g2_antennanp ANTENNA_2255 (.A(_1002_));
 sg13g2_antennanp ANTENNA_2256 (.A(_1071_));
 sg13g2_antennanp ANTENNA_2257 (.A(_1071_));
 sg13g2_antennanp ANTENNA_2258 (.A(_1071_));
 sg13g2_antennanp ANTENNA_2259 (.A(_1085_));
 sg13g2_antennanp ANTENNA_2260 (.A(_1085_));
 sg13g2_antennanp ANTENNA_2261 (.A(_1085_));
 sg13g2_antennanp ANTENNA_2262 (.A(_1085_));
 sg13g2_antennanp ANTENNA_2263 (.A(_1085_));
 sg13g2_antennanp ANTENNA_2264 (.A(_1085_));
 sg13g2_antennanp ANTENNA_2265 (.A(_1225_));
 sg13g2_antennanp ANTENNA_2266 (.A(_1225_));
 sg13g2_antennanp ANTENNA_2267 (.A(_1292_));
 sg13g2_antennanp ANTENNA_2268 (.A(_1292_));
 sg13g2_antennanp ANTENNA_2269 (.A(_1326_));
 sg13g2_antennanp ANTENNA_2270 (.A(_1326_));
 sg13g2_antennanp ANTENNA_2271 (.A(_1326_));
 sg13g2_antennanp ANTENNA_2272 (.A(_1326_));
 sg13g2_antennanp ANTENNA_2273 (.A(_1326_));
 sg13g2_antennanp ANTENNA_2274 (.A(_1326_));
 sg13g2_antennanp ANTENNA_2275 (.A(_1326_));
 sg13g2_antennanp ANTENNA_2276 (.A(_1326_));
 sg13g2_antennanp ANTENNA_2277 (.A(_1326_));
 sg13g2_antennanp ANTENNA_2278 (.A(_1363_));
 sg13g2_antennanp ANTENNA_2279 (.A(_1411_));
 sg13g2_antennanp ANTENNA_2280 (.A(_1439_));
 sg13g2_antennanp ANTENNA_2281 (.A(_1439_));
 sg13g2_antennanp ANTENNA_2282 (.A(_1470_));
 sg13g2_antennanp ANTENNA_2283 (.A(_1470_));
 sg13g2_antennanp ANTENNA_2284 (.A(_1519_));
 sg13g2_antennanp ANTENNA_2285 (.A(_1531_));
 sg13g2_antennanp ANTENNA_2286 (.A(_1531_));
 sg13g2_antennanp ANTENNA_2287 (.A(_1532_));
 sg13g2_antennanp ANTENNA_2288 (.A(_1532_));
 sg13g2_antennanp ANTENNA_2289 (.A(_1532_));
 sg13g2_antennanp ANTENNA_2290 (.A(_1544_));
 sg13g2_antennanp ANTENNA_2291 (.A(_1544_));
 sg13g2_antennanp ANTENNA_2292 (.A(_1544_));
 sg13g2_antennanp ANTENNA_2293 (.A(_1544_));
 sg13g2_antennanp ANTENNA_2294 (.A(_1544_));
 sg13g2_antennanp ANTENNA_2295 (.A(_1553_));
 sg13g2_antennanp ANTENNA_2296 (.A(_1631_));
 sg13g2_antennanp ANTENNA_2297 (.A(_1631_));
 sg13g2_antennanp ANTENNA_2298 (.A(_1631_));
 sg13g2_antennanp ANTENNA_2299 (.A(_1685_));
 sg13g2_antennanp ANTENNA_2300 (.A(_1685_));
 sg13g2_antennanp ANTENNA_2301 (.A(_1685_));
 sg13g2_antennanp ANTENNA_2302 (.A(_1685_));
 sg13g2_antennanp ANTENNA_2303 (.A(_1696_));
 sg13g2_antennanp ANTENNA_2304 (.A(_1696_));
 sg13g2_antennanp ANTENNA_2305 (.A(_1696_));
 sg13g2_antennanp ANTENNA_2306 (.A(_1696_));
 sg13g2_antennanp ANTENNA_2307 (.A(_1696_));
 sg13g2_antennanp ANTENNA_2308 (.A(_1696_));
 sg13g2_antennanp ANTENNA_2309 (.A(_1696_));
 sg13g2_antennanp ANTENNA_2310 (.A(_1696_));
 sg13g2_antennanp ANTENNA_2311 (.A(_1696_));
 sg13g2_antennanp ANTENNA_2312 (.A(_1696_));
 sg13g2_antennanp ANTENNA_2313 (.A(_1707_));
 sg13g2_antennanp ANTENNA_2314 (.A(_1707_));
 sg13g2_antennanp ANTENNA_2315 (.A(_1707_));
 sg13g2_antennanp ANTENNA_2316 (.A(_1707_));
 sg13g2_antennanp ANTENNA_2317 (.A(_1707_));
 sg13g2_antennanp ANTENNA_2318 (.A(_1716_));
 sg13g2_antennanp ANTENNA_2319 (.A(_1735_));
 sg13g2_antennanp ANTENNA_2320 (.A(_1735_));
 sg13g2_antennanp ANTENNA_2321 (.A(_1761_));
 sg13g2_antennanp ANTENNA_2322 (.A(_2014_));
 sg13g2_antennanp ANTENNA_2323 (.A(_2014_));
 sg13g2_antennanp ANTENNA_2324 (.A(_2020_));
 sg13g2_antennanp ANTENNA_2325 (.A(_2020_));
 sg13g2_antennanp ANTENNA_2326 (.A(_2020_));
 sg13g2_antennanp ANTENNA_2327 (.A(_2020_));
 sg13g2_antennanp ANTENNA_2328 (.A(_2020_));
 sg13g2_antennanp ANTENNA_2329 (.A(_2020_));
 sg13g2_antennanp ANTENNA_2330 (.A(_2020_));
 sg13g2_antennanp ANTENNA_2331 (.A(_2020_));
 sg13g2_antennanp ANTENNA_2332 (.A(_2020_));
 sg13g2_antennanp ANTENNA_2333 (.A(_2020_));
 sg13g2_antennanp ANTENNA_2334 (.A(_2020_));
 sg13g2_antennanp ANTENNA_2335 (.A(_2020_));
 sg13g2_antennanp ANTENNA_2336 (.A(_2020_));
 sg13g2_antennanp ANTENNA_2337 (.A(_2037_));
 sg13g2_antennanp ANTENNA_2338 (.A(_2097_));
 sg13g2_antennanp ANTENNA_2339 (.A(_2097_));
 sg13g2_antennanp ANTENNA_2340 (.A(_2097_));
 sg13g2_antennanp ANTENNA_2341 (.A(_2097_));
 sg13g2_antennanp ANTENNA_2342 (.A(_2097_));
 sg13g2_antennanp ANTENNA_2343 (.A(_2110_));
 sg13g2_antennanp ANTENNA_2344 (.A(_2110_));
 sg13g2_antennanp ANTENNA_2345 (.A(_2112_));
 sg13g2_antennanp ANTENNA_2346 (.A(_2145_));
 sg13g2_antennanp ANTENNA_2347 (.A(_2171_));
 sg13g2_antennanp ANTENNA_2348 (.A(_2171_));
 sg13g2_antennanp ANTENNA_2349 (.A(_2171_));
 sg13g2_antennanp ANTENNA_2350 (.A(_2171_));
 sg13g2_antennanp ANTENNA_2351 (.A(_2171_));
 sg13g2_antennanp ANTENNA_2352 (.A(_2171_));
 sg13g2_antennanp ANTENNA_2353 (.A(_2171_));
 sg13g2_antennanp ANTENNA_2354 (.A(_2171_));
 sg13g2_antennanp ANTENNA_2355 (.A(_2171_));
 sg13g2_antennanp ANTENNA_2356 (.A(_2172_));
 sg13g2_antennanp ANTENNA_2357 (.A(_2172_));
 sg13g2_antennanp ANTENNA_2358 (.A(_2172_));
 sg13g2_antennanp ANTENNA_2359 (.A(_2172_));
 sg13g2_antennanp ANTENNA_2360 (.A(_2172_));
 sg13g2_antennanp ANTENNA_2361 (.A(_2172_));
 sg13g2_antennanp ANTENNA_2362 (.A(_2172_));
 sg13g2_antennanp ANTENNA_2363 (.A(_2172_));
 sg13g2_antennanp ANTENNA_2364 (.A(_2172_));
 sg13g2_antennanp ANTENNA_2365 (.A(_2172_));
 sg13g2_antennanp ANTENNA_2366 (.A(_2257_));
 sg13g2_antennanp ANTENNA_2367 (.A(_2257_));
 sg13g2_antennanp ANTENNA_2368 (.A(_2408_));
 sg13g2_antennanp ANTENNA_2369 (.A(_2408_));
 sg13g2_antennanp ANTENNA_2370 (.A(_2408_));
 sg13g2_antennanp ANTENNA_2371 (.A(_2430_));
 sg13g2_antennanp ANTENNA_2372 (.A(_2430_));
 sg13g2_antennanp ANTENNA_2373 (.A(_2430_));
 sg13g2_antennanp ANTENNA_2374 (.A(_2430_));
 sg13g2_antennanp ANTENNA_2375 (.A(_2430_));
 sg13g2_antennanp ANTENNA_2376 (.A(_2430_));
 sg13g2_antennanp ANTENNA_2377 (.A(_2461_));
 sg13g2_antennanp ANTENNA_2378 (.A(_2461_));
 sg13g2_antennanp ANTENNA_2379 (.A(_2461_));
 sg13g2_antennanp ANTENNA_2380 (.A(_2461_));
 sg13g2_antennanp ANTENNA_2381 (.A(_2461_));
 sg13g2_antennanp ANTENNA_2382 (.A(_2467_));
 sg13g2_antennanp ANTENNA_2383 (.A(_2467_));
 sg13g2_antennanp ANTENNA_2384 (.A(_2467_));
 sg13g2_antennanp ANTENNA_2385 (.A(_2467_));
 sg13g2_antennanp ANTENNA_2386 (.A(_2467_));
 sg13g2_antennanp ANTENNA_2387 (.A(_2470_));
 sg13g2_antennanp ANTENNA_2388 (.A(_2470_));
 sg13g2_antennanp ANTENNA_2389 (.A(_2470_));
 sg13g2_antennanp ANTENNA_2390 (.A(_2470_));
 sg13g2_antennanp ANTENNA_2391 (.A(_2480_));
 sg13g2_antennanp ANTENNA_2392 (.A(_2480_));
 sg13g2_antennanp ANTENNA_2393 (.A(_2480_));
 sg13g2_antennanp ANTENNA_2394 (.A(_2480_));
 sg13g2_antennanp ANTENNA_2395 (.A(_2482_));
 sg13g2_antennanp ANTENNA_2396 (.A(_2482_));
 sg13g2_antennanp ANTENNA_2397 (.A(_2482_));
 sg13g2_antennanp ANTENNA_2398 (.A(_2482_));
 sg13g2_antennanp ANTENNA_2399 (.A(_2482_));
 sg13g2_antennanp ANTENNA_2400 (.A(_2482_));
 sg13g2_antennanp ANTENNA_2401 (.A(_2482_));
 sg13g2_antennanp ANTENNA_2402 (.A(_2482_));
 sg13g2_antennanp ANTENNA_2403 (.A(_2487_));
 sg13g2_antennanp ANTENNA_2404 (.A(_2487_));
 sg13g2_antennanp ANTENNA_2405 (.A(_2501_));
 sg13g2_antennanp ANTENNA_2406 (.A(_2501_));
 sg13g2_antennanp ANTENNA_2407 (.A(_2501_));
 sg13g2_antennanp ANTENNA_2408 (.A(_2501_));
 sg13g2_antennanp ANTENNA_2409 (.A(_2501_));
 sg13g2_antennanp ANTENNA_2410 (.A(_2501_));
 sg13g2_antennanp ANTENNA_2411 (.A(_2520_));
 sg13g2_antennanp ANTENNA_2412 (.A(_2520_));
 sg13g2_antennanp ANTENNA_2413 (.A(_2520_));
 sg13g2_antennanp ANTENNA_2414 (.A(_2520_));
 sg13g2_antennanp ANTENNA_2415 (.A(_2530_));
 sg13g2_antennanp ANTENNA_2416 (.A(_2530_));
 sg13g2_antennanp ANTENNA_2417 (.A(_2530_));
 sg13g2_antennanp ANTENNA_2418 (.A(_2530_));
 sg13g2_antennanp ANTENNA_2419 (.A(_2532_));
 sg13g2_antennanp ANTENNA_2420 (.A(_2532_));
 sg13g2_antennanp ANTENNA_2421 (.A(_2532_));
 sg13g2_antennanp ANTENNA_2422 (.A(_2532_));
 sg13g2_antennanp ANTENNA_2423 (.A(_2532_));
 sg13g2_antennanp ANTENNA_2424 (.A(_2532_));
 sg13g2_antennanp ANTENNA_2425 (.A(_2532_));
 sg13g2_antennanp ANTENNA_2426 (.A(_2532_));
 sg13g2_antennanp ANTENNA_2427 (.A(_2532_));
 sg13g2_antennanp ANTENNA_2428 (.A(_2532_));
 sg13g2_antennanp ANTENNA_2429 (.A(_2537_));
 sg13g2_antennanp ANTENNA_2430 (.A(_2537_));
 sg13g2_antennanp ANTENNA_2431 (.A(_2537_));
 sg13g2_antennanp ANTENNA_2432 (.A(_2537_));
 sg13g2_antennanp ANTENNA_2433 (.A(_2573_));
 sg13g2_antennanp ANTENNA_2434 (.A(_2573_));
 sg13g2_antennanp ANTENNA_2435 (.A(_2573_));
 sg13g2_antennanp ANTENNA_2436 (.A(_2573_));
 sg13g2_antennanp ANTENNA_2437 (.A(_2577_));
 sg13g2_antennanp ANTENNA_2438 (.A(_2577_));
 sg13g2_antennanp ANTENNA_2439 (.A(_2577_));
 sg13g2_antennanp ANTENNA_2440 (.A(_2577_));
 sg13g2_antennanp ANTENNA_2441 (.A(_2577_));
 sg13g2_antennanp ANTENNA_2442 (.A(_2577_));
 sg13g2_antennanp ANTENNA_2443 (.A(_2577_));
 sg13g2_antennanp ANTENNA_2444 (.A(_2577_));
 sg13g2_antennanp ANTENNA_2445 (.A(_2585_));
 sg13g2_antennanp ANTENNA_2446 (.A(_2585_));
 sg13g2_antennanp ANTENNA_2447 (.A(_2585_));
 sg13g2_antennanp ANTENNA_2448 (.A(_2588_));
 sg13g2_antennanp ANTENNA_2449 (.A(_2595_));
 sg13g2_antennanp ANTENNA_2450 (.A(_2595_));
 sg13g2_antennanp ANTENNA_2451 (.A(_2595_));
 sg13g2_antennanp ANTENNA_2452 (.A(_2595_));
 sg13g2_antennanp ANTENNA_2453 (.A(_2595_));
 sg13g2_antennanp ANTENNA_2454 (.A(_2595_));
 sg13g2_antennanp ANTENNA_2455 (.A(_2600_));
 sg13g2_antennanp ANTENNA_2456 (.A(_2600_));
 sg13g2_antennanp ANTENNA_2457 (.A(_2600_));
 sg13g2_antennanp ANTENNA_2458 (.A(_2600_));
 sg13g2_antennanp ANTENNA_2459 (.A(_2601_));
 sg13g2_antennanp ANTENNA_2460 (.A(_2601_));
 sg13g2_antennanp ANTENNA_2461 (.A(_2601_));
 sg13g2_antennanp ANTENNA_2462 (.A(_2601_));
 sg13g2_antennanp ANTENNA_2463 (.A(_2607_));
 sg13g2_antennanp ANTENNA_2464 (.A(_2607_));
 sg13g2_antennanp ANTENNA_2465 (.A(_2615_));
 sg13g2_antennanp ANTENNA_2466 (.A(_2615_));
 sg13g2_antennanp ANTENNA_2467 (.A(_2615_));
 sg13g2_antennanp ANTENNA_2468 (.A(_2619_));
 sg13g2_antennanp ANTENNA_2469 (.A(_2619_));
 sg13g2_antennanp ANTENNA_2470 (.A(_2619_));
 sg13g2_antennanp ANTENNA_2471 (.A(_2619_));
 sg13g2_antennanp ANTENNA_2472 (.A(_2619_));
 sg13g2_antennanp ANTENNA_2473 (.A(_2619_));
 sg13g2_antennanp ANTENNA_2474 (.A(_2622_));
 sg13g2_antennanp ANTENNA_2475 (.A(_2622_));
 sg13g2_antennanp ANTENNA_2476 (.A(_2622_));
 sg13g2_antennanp ANTENNA_2477 (.A(_2622_));
 sg13g2_antennanp ANTENNA_2478 (.A(_2622_));
 sg13g2_antennanp ANTENNA_2479 (.A(_2622_));
 sg13g2_antennanp ANTENNA_2480 (.A(_2625_));
 sg13g2_antennanp ANTENNA_2481 (.A(_2625_));
 sg13g2_antennanp ANTENNA_2482 (.A(_2625_));
 sg13g2_antennanp ANTENNA_2483 (.A(_2625_));
 sg13g2_antennanp ANTENNA_2484 (.A(_2659_));
 sg13g2_antennanp ANTENNA_2485 (.A(_2659_));
 sg13g2_antennanp ANTENNA_2486 (.A(_2659_));
 sg13g2_antennanp ANTENNA_2487 (.A(_2659_));
 sg13g2_antennanp ANTENNA_2488 (.A(_2659_));
 sg13g2_antennanp ANTENNA_2489 (.A(_2665_));
 sg13g2_antennanp ANTENNA_2490 (.A(_2665_));
 sg13g2_antennanp ANTENNA_2491 (.A(_2665_));
 sg13g2_antennanp ANTENNA_2492 (.A(_2678_));
 sg13g2_antennanp ANTENNA_2493 (.A(_2678_));
 sg13g2_antennanp ANTENNA_2494 (.A(_2678_));
 sg13g2_antennanp ANTENNA_2495 (.A(_2678_));
 sg13g2_antennanp ANTENNA_2496 (.A(_2678_));
 sg13g2_antennanp ANTENNA_2497 (.A(_2678_));
 sg13g2_antennanp ANTENNA_2498 (.A(_2678_));
 sg13g2_antennanp ANTENNA_2499 (.A(_2732_));
 sg13g2_antennanp ANTENNA_2500 (.A(_2732_));
 sg13g2_antennanp ANTENNA_2501 (.A(_2732_));
 sg13g2_antennanp ANTENNA_2502 (.A(_2733_));
 sg13g2_antennanp ANTENNA_2503 (.A(_2733_));
 sg13g2_antennanp ANTENNA_2504 (.A(_2733_));
 sg13g2_antennanp ANTENNA_2505 (.A(_2733_));
 sg13g2_antennanp ANTENNA_2506 (.A(_2739_));
 sg13g2_antennanp ANTENNA_2507 (.A(_2739_));
 sg13g2_antennanp ANTENNA_2508 (.A(_2739_));
 sg13g2_antennanp ANTENNA_2509 (.A(_2739_));
 sg13g2_antennanp ANTENNA_2510 (.A(_2769_));
 sg13g2_antennanp ANTENNA_2511 (.A(_2769_));
 sg13g2_antennanp ANTENNA_2512 (.A(_2769_));
 sg13g2_antennanp ANTENNA_2513 (.A(_2769_));
 sg13g2_antennanp ANTENNA_2514 (.A(_2779_));
 sg13g2_antennanp ANTENNA_2515 (.A(_2779_));
 sg13g2_antennanp ANTENNA_2516 (.A(_2779_));
 sg13g2_antennanp ANTENNA_2517 (.A(_2779_));
 sg13g2_antennanp ANTENNA_2518 (.A(_2789_));
 sg13g2_antennanp ANTENNA_2519 (.A(_2789_));
 sg13g2_antennanp ANTENNA_2520 (.A(_2789_));
 sg13g2_antennanp ANTENNA_2521 (.A(_2789_));
 sg13g2_antennanp ANTENNA_2522 (.A(_2805_));
 sg13g2_antennanp ANTENNA_2523 (.A(_2805_));
 sg13g2_antennanp ANTENNA_2524 (.A(_2808_));
 sg13g2_antennanp ANTENNA_2525 (.A(_2808_));
 sg13g2_antennanp ANTENNA_2526 (.A(_2808_));
 sg13g2_antennanp ANTENNA_2527 (.A(_2808_));
 sg13g2_antennanp ANTENNA_2528 (.A(_2816_));
 sg13g2_antennanp ANTENNA_2529 (.A(_2816_));
 sg13g2_antennanp ANTENNA_2530 (.A(_2816_));
 sg13g2_antennanp ANTENNA_2531 (.A(_2816_));
 sg13g2_antennanp ANTENNA_2532 (.A(_2826_));
 sg13g2_antennanp ANTENNA_2533 (.A(_2826_));
 sg13g2_antennanp ANTENNA_2534 (.A(_2826_));
 sg13g2_antennanp ANTENNA_2535 (.A(_2826_));
 sg13g2_antennanp ANTENNA_2536 (.A(_2858_));
 sg13g2_antennanp ANTENNA_2537 (.A(_2858_));
 sg13g2_antennanp ANTENNA_2538 (.A(_2879_));
 sg13g2_antennanp ANTENNA_2539 (.A(_2879_));
 sg13g2_antennanp ANTENNA_2540 (.A(_2879_));
 sg13g2_antennanp ANTENNA_2541 (.A(_2879_));
 sg13g2_antennanp ANTENNA_2542 (.A(_2879_));
 sg13g2_antennanp ANTENNA_2543 (.A(_2879_));
 sg13g2_antennanp ANTENNA_2544 (.A(_2879_));
 sg13g2_antennanp ANTENNA_2545 (.A(_2879_));
 sg13g2_antennanp ANTENNA_2546 (.A(_2914_));
 sg13g2_antennanp ANTENNA_2547 (.A(_2931_));
 sg13g2_antennanp ANTENNA_2548 (.A(_2931_));
 sg13g2_antennanp ANTENNA_2549 (.A(_2931_));
 sg13g2_antennanp ANTENNA_2550 (.A(_2931_));
 sg13g2_antennanp ANTENNA_2551 (.A(_2936_));
 sg13g2_antennanp ANTENNA_2552 (.A(_2936_));
 sg13g2_antennanp ANTENNA_2553 (.A(_2936_));
 sg13g2_antennanp ANTENNA_2554 (.A(_2957_));
 sg13g2_antennanp ANTENNA_2555 (.A(_2957_));
 sg13g2_antennanp ANTENNA_2556 (.A(_2957_));
 sg13g2_antennanp ANTENNA_2557 (.A(_2957_));
 sg13g2_antennanp ANTENNA_2558 (.A(_2967_));
 sg13g2_antennanp ANTENNA_2559 (.A(_2967_));
 sg13g2_antennanp ANTENNA_2560 (.A(_2967_));
 sg13g2_antennanp ANTENNA_2561 (.A(_2967_));
 sg13g2_antennanp ANTENNA_2562 (.A(_2967_));
 sg13g2_antennanp ANTENNA_2563 (.A(_2967_));
 sg13g2_antennanp ANTENNA_2564 (.A(_2967_));
 sg13g2_antennanp ANTENNA_2565 (.A(_2967_));
 sg13g2_antennanp ANTENNA_2566 (.A(_2967_));
 sg13g2_antennanp ANTENNA_2567 (.A(_2967_));
 sg13g2_antennanp ANTENNA_2568 (.A(_2967_));
 sg13g2_antennanp ANTENNA_2569 (.A(_2967_));
 sg13g2_antennanp ANTENNA_2570 (.A(_2967_));
 sg13g2_antennanp ANTENNA_2571 (.A(_2970_));
 sg13g2_antennanp ANTENNA_2572 (.A(_2970_));
 sg13g2_antennanp ANTENNA_2573 (.A(_2970_));
 sg13g2_antennanp ANTENNA_2574 (.A(_2970_));
 sg13g2_antennanp ANTENNA_2575 (.A(_2974_));
 sg13g2_antennanp ANTENNA_2576 (.A(_2974_));
 sg13g2_antennanp ANTENNA_2577 (.A(_2977_));
 sg13g2_antennanp ANTENNA_2578 (.A(_2977_));
 sg13g2_antennanp ANTENNA_2579 (.A(_2977_));
 sg13g2_antennanp ANTENNA_2580 (.A(_2977_));
 sg13g2_antennanp ANTENNA_2581 (.A(_2977_));
 sg13g2_antennanp ANTENNA_2582 (.A(_2986_));
 sg13g2_antennanp ANTENNA_2583 (.A(_2986_));
 sg13g2_antennanp ANTENNA_2584 (.A(_2986_));
 sg13g2_antennanp ANTENNA_2585 (.A(_2986_));
 sg13g2_antennanp ANTENNA_2586 (.A(_3018_));
 sg13g2_antennanp ANTENNA_2587 (.A(_3018_));
 sg13g2_antennanp ANTENNA_2588 (.A(_3018_));
 sg13g2_antennanp ANTENNA_2589 (.A(_3040_));
 sg13g2_antennanp ANTENNA_2590 (.A(_3040_));
 sg13g2_antennanp ANTENNA_2591 (.A(_3040_));
 sg13g2_antennanp ANTENNA_2592 (.A(clk));
 sg13g2_antennanp ANTENNA_2593 (.A(clk));
 sg13g2_antennanp ANTENNA_2594 (.A(net22));
 sg13g2_antennanp ANTENNA_2595 (.A(net22));
 sg13g2_antennanp ANTENNA_2596 (.A(net22));
 sg13g2_antennanp ANTENNA_2597 (.A(net22));
 sg13g2_antennanp ANTENNA_2598 (.A(net22));
 sg13g2_antennanp ANTENNA_2599 (.A(net22));
 sg13g2_antennanp ANTENNA_2600 (.A(net22));
 sg13g2_antennanp ANTENNA_2601 (.A(net22));
 sg13g2_antennanp ANTENNA_2602 (.A(net22));
 sg13g2_antennanp ANTENNA_2603 (.A(net23));
 sg13g2_antennanp ANTENNA_2604 (.A(net23));
 sg13g2_antennanp ANTENNA_2605 (.A(net23));
 sg13g2_antennanp ANTENNA_2606 (.A(net23));
 sg13g2_antennanp ANTENNA_2607 (.A(net23));
 sg13g2_antennanp ANTENNA_2608 (.A(net23));
 sg13g2_antennanp ANTENNA_2609 (.A(net23));
 sg13g2_antennanp ANTENNA_2610 (.A(net23));
 sg13g2_antennanp ANTENNA_2611 (.A(net29));
 sg13g2_antennanp ANTENNA_2612 (.A(net29));
 sg13g2_antennanp ANTENNA_2613 (.A(net29));
 sg13g2_antennanp ANTENNA_2614 (.A(net29));
 sg13g2_antennanp ANTENNA_2615 (.A(net29));
 sg13g2_antennanp ANTENNA_2616 (.A(net29));
 sg13g2_antennanp ANTENNA_2617 (.A(net29));
 sg13g2_antennanp ANTENNA_2618 (.A(net29));
 sg13g2_antennanp ANTENNA_2619 (.A(net29));
 sg13g2_antennanp ANTENNA_2620 (.A(net35));
 sg13g2_antennanp ANTENNA_2621 (.A(net35));
 sg13g2_antennanp ANTENNA_2622 (.A(net35));
 sg13g2_antennanp ANTENNA_2623 (.A(net35));
 sg13g2_antennanp ANTENNA_2624 (.A(net35));
 sg13g2_antennanp ANTENNA_2625 (.A(net35));
 sg13g2_antennanp ANTENNA_2626 (.A(net35));
 sg13g2_antennanp ANTENNA_2627 (.A(net35));
 sg13g2_antennanp ANTENNA_2628 (.A(net35));
 sg13g2_antennanp ANTENNA_2629 (.A(net40));
 sg13g2_antennanp ANTENNA_2630 (.A(net40));
 sg13g2_antennanp ANTENNA_2631 (.A(net40));
 sg13g2_antennanp ANTENNA_2632 (.A(net40));
 sg13g2_antennanp ANTENNA_2633 (.A(net40));
 sg13g2_antennanp ANTENNA_2634 (.A(net40));
 sg13g2_antennanp ANTENNA_2635 (.A(net40));
 sg13g2_antennanp ANTENNA_2636 (.A(net40));
 sg13g2_antennanp ANTENNA_2637 (.A(net40));
 sg13g2_antennanp ANTENNA_2638 (.A(net46));
 sg13g2_antennanp ANTENNA_2639 (.A(net46));
 sg13g2_antennanp ANTENNA_2640 (.A(net46));
 sg13g2_antennanp ANTENNA_2641 (.A(net46));
 sg13g2_antennanp ANTENNA_2642 (.A(net46));
 sg13g2_antennanp ANTENNA_2643 (.A(net46));
 sg13g2_antennanp ANTENNA_2644 (.A(net46));
 sg13g2_antennanp ANTENNA_2645 (.A(net46));
 sg13g2_antennanp ANTENNA_2646 (.A(net46));
 sg13g2_antennanp ANTENNA_2647 (.A(net53));
 sg13g2_antennanp ANTENNA_2648 (.A(net53));
 sg13g2_antennanp ANTENNA_2649 (.A(net53));
 sg13g2_antennanp ANTENNA_2650 (.A(net53));
 sg13g2_antennanp ANTENNA_2651 (.A(net53));
 sg13g2_antennanp ANTENNA_2652 (.A(net53));
 sg13g2_antennanp ANTENNA_2653 (.A(net53));
 sg13g2_antennanp ANTENNA_2654 (.A(net53));
 sg13g2_antennanp ANTENNA_2655 (.A(net53));
 sg13g2_antennanp ANTENNA_2656 (.A(net59));
 sg13g2_antennanp ANTENNA_2657 (.A(net59));
 sg13g2_antennanp ANTENNA_2658 (.A(net59));
 sg13g2_antennanp ANTENNA_2659 (.A(net59));
 sg13g2_antennanp ANTENNA_2660 (.A(net59));
 sg13g2_antennanp ANTENNA_2661 (.A(net59));
 sg13g2_antennanp ANTENNA_2662 (.A(net59));
 sg13g2_antennanp ANTENNA_2663 (.A(net59));
 sg13g2_antennanp ANTENNA_2664 (.A(net59));
 sg13g2_antennanp ANTENNA_2665 (.A(net61));
 sg13g2_antennanp ANTENNA_2666 (.A(net61));
 sg13g2_antennanp ANTENNA_2667 (.A(net61));
 sg13g2_antennanp ANTENNA_2668 (.A(net61));
 sg13g2_antennanp ANTENNA_2669 (.A(net61));
 sg13g2_antennanp ANTENNA_2670 (.A(net61));
 sg13g2_antennanp ANTENNA_2671 (.A(net61));
 sg13g2_antennanp ANTENNA_2672 (.A(net61));
 sg13g2_antennanp ANTENNA_2673 (.A(net61));
 sg13g2_antennanp ANTENNA_2674 (.A(net62));
 sg13g2_antennanp ANTENNA_2675 (.A(net62));
 sg13g2_antennanp ANTENNA_2676 (.A(net62));
 sg13g2_antennanp ANTENNA_2677 (.A(net62));
 sg13g2_antennanp ANTENNA_2678 (.A(net62));
 sg13g2_antennanp ANTENNA_2679 (.A(net62));
 sg13g2_antennanp ANTENNA_2680 (.A(net62));
 sg13g2_antennanp ANTENNA_2681 (.A(net62));
 sg13g2_antennanp ANTENNA_2682 (.A(net62));
 sg13g2_antennanp ANTENNA_2683 (.A(net64));
 sg13g2_antennanp ANTENNA_2684 (.A(net64));
 sg13g2_antennanp ANTENNA_2685 (.A(net64));
 sg13g2_antennanp ANTENNA_2686 (.A(net64));
 sg13g2_antennanp ANTENNA_2687 (.A(net64));
 sg13g2_antennanp ANTENNA_2688 (.A(net64));
 sg13g2_antennanp ANTENNA_2689 (.A(net64));
 sg13g2_antennanp ANTENNA_2690 (.A(net64));
 sg13g2_antennanp ANTENNA_2691 (.A(net70));
 sg13g2_antennanp ANTENNA_2692 (.A(net70));
 sg13g2_antennanp ANTENNA_2693 (.A(net70));
 sg13g2_antennanp ANTENNA_2694 (.A(net70));
 sg13g2_antennanp ANTENNA_2695 (.A(net70));
 sg13g2_antennanp ANTENNA_2696 (.A(net70));
 sg13g2_antennanp ANTENNA_2697 (.A(net70));
 sg13g2_antennanp ANTENNA_2698 (.A(net70));
 sg13g2_antennanp ANTENNA_2699 (.A(net71));
 sg13g2_antennanp ANTENNA_2700 (.A(net71));
 sg13g2_antennanp ANTENNA_2701 (.A(net71));
 sg13g2_antennanp ANTENNA_2702 (.A(net71));
 sg13g2_antennanp ANTENNA_2703 (.A(net71));
 sg13g2_antennanp ANTENNA_2704 (.A(net71));
 sg13g2_antennanp ANTENNA_2705 (.A(net71));
 sg13g2_antennanp ANTENNA_2706 (.A(net71));
 sg13g2_antennanp ANTENNA_2707 (.A(net71));
 sg13g2_antennanp ANTENNA_2708 (.A(net71));
 sg13g2_antennanp ANTENNA_2709 (.A(net71));
 sg13g2_antennanp ANTENNA_2710 (.A(net71));
 sg13g2_antennanp ANTENNA_2711 (.A(net71));
 sg13g2_antennanp ANTENNA_2712 (.A(net71));
 sg13g2_antennanp ANTENNA_2713 (.A(net71));
 sg13g2_antennanp ANTENNA_2714 (.A(net71));
 sg13g2_antennanp ANTENNA_2715 (.A(net76));
 sg13g2_antennanp ANTENNA_2716 (.A(net76));
 sg13g2_antennanp ANTENNA_2717 (.A(net76));
 sg13g2_antennanp ANTENNA_2718 (.A(net76));
 sg13g2_antennanp ANTENNA_2719 (.A(net76));
 sg13g2_antennanp ANTENNA_2720 (.A(net76));
 sg13g2_antennanp ANTENNA_2721 (.A(net76));
 sg13g2_antennanp ANTENNA_2722 (.A(net76));
 sg13g2_antennanp ANTENNA_2723 (.A(net76));
 sg13g2_antennanp ANTENNA_2724 (.A(net78));
 sg13g2_antennanp ANTENNA_2725 (.A(net78));
 sg13g2_antennanp ANTENNA_2726 (.A(net78));
 sg13g2_antennanp ANTENNA_2727 (.A(net78));
 sg13g2_antennanp ANTENNA_2728 (.A(net78));
 sg13g2_antennanp ANTENNA_2729 (.A(net78));
 sg13g2_antennanp ANTENNA_2730 (.A(net78));
 sg13g2_antennanp ANTENNA_2731 (.A(net78));
 sg13g2_antennanp ANTENNA_2732 (.A(net78));
 sg13g2_antennanp ANTENNA_2733 (.A(net79));
 sg13g2_antennanp ANTENNA_2734 (.A(net79));
 sg13g2_antennanp ANTENNA_2735 (.A(net79));
 sg13g2_antennanp ANTENNA_2736 (.A(net79));
 sg13g2_antennanp ANTENNA_2737 (.A(net79));
 sg13g2_antennanp ANTENNA_2738 (.A(net79));
 sg13g2_antennanp ANTENNA_2739 (.A(net79));
 sg13g2_antennanp ANTENNA_2740 (.A(net79));
 sg13g2_antennanp ANTENNA_2741 (.A(net79));
 sg13g2_antennanp ANTENNA_2742 (.A(net84));
 sg13g2_antennanp ANTENNA_2743 (.A(net84));
 sg13g2_antennanp ANTENNA_2744 (.A(net84));
 sg13g2_antennanp ANTENNA_2745 (.A(net84));
 sg13g2_antennanp ANTENNA_2746 (.A(net84));
 sg13g2_antennanp ANTENNA_2747 (.A(net84));
 sg13g2_antennanp ANTENNA_2748 (.A(net84));
 sg13g2_antennanp ANTENNA_2749 (.A(net84));
 sg13g2_antennanp ANTENNA_2750 (.A(net89));
 sg13g2_antennanp ANTENNA_2751 (.A(net89));
 sg13g2_antennanp ANTENNA_2752 (.A(net89));
 sg13g2_antennanp ANTENNA_2753 (.A(net89));
 sg13g2_antennanp ANTENNA_2754 (.A(net89));
 sg13g2_antennanp ANTENNA_2755 (.A(net89));
 sg13g2_antennanp ANTENNA_2756 (.A(net89));
 sg13g2_antennanp ANTENNA_2757 (.A(net89));
 sg13g2_antennanp ANTENNA_2758 (.A(net89));
 sg13g2_antennanp ANTENNA_2759 (.A(net91));
 sg13g2_antennanp ANTENNA_2760 (.A(net91));
 sg13g2_antennanp ANTENNA_2761 (.A(net91));
 sg13g2_antennanp ANTENNA_2762 (.A(net91));
 sg13g2_antennanp ANTENNA_2763 (.A(net91));
 sg13g2_antennanp ANTENNA_2764 (.A(net91));
 sg13g2_antennanp ANTENNA_2765 (.A(net91));
 sg13g2_antennanp ANTENNA_2766 (.A(net91));
 sg13g2_antennanp ANTENNA_2767 (.A(net91));
 sg13g2_antennanp ANTENNA_2768 (.A(net91));
 sg13g2_antennanp ANTENNA_2769 (.A(net91));
 sg13g2_antennanp ANTENNA_2770 (.A(net91));
 sg13g2_antennanp ANTENNA_2771 (.A(net91));
 sg13g2_antennanp ANTENNA_2772 (.A(net91));
 sg13g2_antennanp ANTENNA_2773 (.A(net91));
 sg13g2_antennanp ANTENNA_2774 (.A(net91));
 sg13g2_antennanp ANTENNA_2775 (.A(net94));
 sg13g2_antennanp ANTENNA_2776 (.A(net94));
 sg13g2_antennanp ANTENNA_2777 (.A(net94));
 sg13g2_antennanp ANTENNA_2778 (.A(net94));
 sg13g2_antennanp ANTENNA_2779 (.A(net94));
 sg13g2_antennanp ANTENNA_2780 (.A(net94));
 sg13g2_antennanp ANTENNA_2781 (.A(net94));
 sg13g2_antennanp ANTENNA_2782 (.A(net94));
 sg13g2_antennanp ANTENNA_2783 (.A(net100));
 sg13g2_antennanp ANTENNA_2784 (.A(net100));
 sg13g2_antennanp ANTENNA_2785 (.A(net100));
 sg13g2_antennanp ANTENNA_2786 (.A(net100));
 sg13g2_antennanp ANTENNA_2787 (.A(net100));
 sg13g2_antennanp ANTENNA_2788 (.A(net100));
 sg13g2_antennanp ANTENNA_2789 (.A(net100));
 sg13g2_antennanp ANTENNA_2790 (.A(net100));
 sg13g2_antennanp ANTENNA_2791 (.A(net100));
 sg13g2_antennanp ANTENNA_2792 (.A(net106));
 sg13g2_antennanp ANTENNA_2793 (.A(net106));
 sg13g2_antennanp ANTENNA_2794 (.A(net106));
 sg13g2_antennanp ANTENNA_2795 (.A(net106));
 sg13g2_antennanp ANTENNA_2796 (.A(net106));
 sg13g2_antennanp ANTENNA_2797 (.A(net106));
 sg13g2_antennanp ANTENNA_2798 (.A(net106));
 sg13g2_antennanp ANTENNA_2799 (.A(net106));
 sg13g2_antennanp ANTENNA_2800 (.A(net106));
 sg13g2_antennanp ANTENNA_2801 (.A(net107));
 sg13g2_antennanp ANTENNA_2802 (.A(net107));
 sg13g2_antennanp ANTENNA_2803 (.A(net107));
 sg13g2_antennanp ANTENNA_2804 (.A(net107));
 sg13g2_antennanp ANTENNA_2805 (.A(net107));
 sg13g2_antennanp ANTENNA_2806 (.A(net107));
 sg13g2_antennanp ANTENNA_2807 (.A(net107));
 sg13g2_antennanp ANTENNA_2808 (.A(net107));
 sg13g2_antennanp ANTENNA_2809 (.A(net107));
 sg13g2_antennanp ANTENNA_2810 (.A(net113));
 sg13g2_antennanp ANTENNA_2811 (.A(net113));
 sg13g2_antennanp ANTENNA_2812 (.A(net113));
 sg13g2_antennanp ANTENNA_2813 (.A(net113));
 sg13g2_antennanp ANTENNA_2814 (.A(net113));
 sg13g2_antennanp ANTENNA_2815 (.A(net113));
 sg13g2_antennanp ANTENNA_2816 (.A(net113));
 sg13g2_antennanp ANTENNA_2817 (.A(net113));
 sg13g2_antennanp ANTENNA_2818 (.A(net125));
 sg13g2_antennanp ANTENNA_2819 (.A(net125));
 sg13g2_antennanp ANTENNA_2820 (.A(net125));
 sg13g2_antennanp ANTENNA_2821 (.A(net125));
 sg13g2_antennanp ANTENNA_2822 (.A(net125));
 sg13g2_antennanp ANTENNA_2823 (.A(net125));
 sg13g2_antennanp ANTENNA_2824 (.A(net125));
 sg13g2_antennanp ANTENNA_2825 (.A(net125));
 sg13g2_antennanp ANTENNA_2826 (.A(net125));
 sg13g2_antennanp ANTENNA_2827 (.A(net128));
 sg13g2_antennanp ANTENNA_2828 (.A(net128));
 sg13g2_antennanp ANTENNA_2829 (.A(net128));
 sg13g2_antennanp ANTENNA_2830 (.A(net128));
 sg13g2_antennanp ANTENNA_2831 (.A(net128));
 sg13g2_antennanp ANTENNA_2832 (.A(net128));
 sg13g2_antennanp ANTENNA_2833 (.A(net128));
 sg13g2_antennanp ANTENNA_2834 (.A(net128));
 sg13g2_antennanp ANTENNA_2835 (.A(net129));
 sg13g2_antennanp ANTENNA_2836 (.A(net129));
 sg13g2_antennanp ANTENNA_2837 (.A(net129));
 sg13g2_antennanp ANTENNA_2838 (.A(net129));
 sg13g2_antennanp ANTENNA_2839 (.A(net129));
 sg13g2_antennanp ANTENNA_2840 (.A(net129));
 sg13g2_antennanp ANTENNA_2841 (.A(net129));
 sg13g2_antennanp ANTENNA_2842 (.A(net129));
 sg13g2_antennanp ANTENNA_2843 (.A(net129));
 sg13g2_antennanp ANTENNA_2844 (.A(net144));
 sg13g2_antennanp ANTENNA_2845 (.A(net144));
 sg13g2_antennanp ANTENNA_2846 (.A(net144));
 sg13g2_antennanp ANTENNA_2847 (.A(net144));
 sg13g2_antennanp ANTENNA_2848 (.A(net144));
 sg13g2_antennanp ANTENNA_2849 (.A(net144));
 sg13g2_antennanp ANTENNA_2850 (.A(net144));
 sg13g2_antennanp ANTENNA_2851 (.A(net144));
 sg13g2_antennanp ANTENNA_2852 (.A(net144));
 sg13g2_antennanp ANTENNA_2853 (.A(net153));
 sg13g2_antennanp ANTENNA_2854 (.A(net153));
 sg13g2_antennanp ANTENNA_2855 (.A(net153));
 sg13g2_antennanp ANTENNA_2856 (.A(net153));
 sg13g2_antennanp ANTENNA_2857 (.A(net153));
 sg13g2_antennanp ANTENNA_2858 (.A(net153));
 sg13g2_antennanp ANTENNA_2859 (.A(net153));
 sg13g2_antennanp ANTENNA_2860 (.A(net153));
 sg13g2_antennanp ANTENNA_2861 (.A(net153));
 sg13g2_antennanp ANTENNA_2862 (.A(net161));
 sg13g2_antennanp ANTENNA_2863 (.A(net161));
 sg13g2_antennanp ANTENNA_2864 (.A(net161));
 sg13g2_antennanp ANTENNA_2865 (.A(net161));
 sg13g2_antennanp ANTENNA_2866 (.A(net161));
 sg13g2_antennanp ANTENNA_2867 (.A(net161));
 sg13g2_antennanp ANTENNA_2868 (.A(net161));
 sg13g2_antennanp ANTENNA_2869 (.A(net161));
 sg13g2_antennanp ANTENNA_2870 (.A(net161));
 sg13g2_antennanp ANTENNA_2871 (.A(net164));
 sg13g2_antennanp ANTENNA_2872 (.A(net164));
 sg13g2_antennanp ANTENNA_2873 (.A(net164));
 sg13g2_antennanp ANTENNA_2874 (.A(net164));
 sg13g2_antennanp ANTENNA_2875 (.A(net164));
 sg13g2_antennanp ANTENNA_2876 (.A(net164));
 sg13g2_antennanp ANTENNA_2877 (.A(net164));
 sg13g2_antennanp ANTENNA_2878 (.A(net164));
 sg13g2_antennanp ANTENNA_2879 (.A(net164));
 sg13g2_antennanp ANTENNA_2880 (.A(net167));
 sg13g2_antennanp ANTENNA_2881 (.A(net167));
 sg13g2_antennanp ANTENNA_2882 (.A(net167));
 sg13g2_antennanp ANTENNA_2883 (.A(net167));
 sg13g2_antennanp ANTENNA_2884 (.A(net167));
 sg13g2_antennanp ANTENNA_2885 (.A(net167));
 sg13g2_antennanp ANTENNA_2886 (.A(net167));
 sg13g2_antennanp ANTENNA_2887 (.A(net167));
 sg13g2_antennanp ANTENNA_2888 (.A(net167));
 sg13g2_antennanp ANTENNA_2889 (.A(net174));
 sg13g2_antennanp ANTENNA_2890 (.A(net174));
 sg13g2_antennanp ANTENNA_2891 (.A(net174));
 sg13g2_antennanp ANTENNA_2892 (.A(net174));
 sg13g2_antennanp ANTENNA_2893 (.A(net174));
 sg13g2_antennanp ANTENNA_2894 (.A(net174));
 sg13g2_antennanp ANTENNA_2895 (.A(net174));
 sg13g2_antennanp ANTENNA_2896 (.A(net174));
 sg13g2_antennanp ANTENNA_2897 (.A(net174));
 sg13g2_antennanp ANTENNA_2898 (.A(net182));
 sg13g2_antennanp ANTENNA_2899 (.A(net182));
 sg13g2_antennanp ANTENNA_2900 (.A(net182));
 sg13g2_antennanp ANTENNA_2901 (.A(net182));
 sg13g2_antennanp ANTENNA_2902 (.A(net182));
 sg13g2_antennanp ANTENNA_2903 (.A(net182));
 sg13g2_antennanp ANTENNA_2904 (.A(net182));
 sg13g2_antennanp ANTENNA_2905 (.A(net182));
 sg13g2_antennanp ANTENNA_2906 (.A(net185));
 sg13g2_antennanp ANTENNA_2907 (.A(net185));
 sg13g2_antennanp ANTENNA_2908 (.A(net185));
 sg13g2_antennanp ANTENNA_2909 (.A(net185));
 sg13g2_antennanp ANTENNA_2910 (.A(net185));
 sg13g2_antennanp ANTENNA_2911 (.A(net185));
 sg13g2_antennanp ANTENNA_2912 (.A(net185));
 sg13g2_antennanp ANTENNA_2913 (.A(net185));
 sg13g2_antennanp ANTENNA_2914 (.A(net185));
 sg13g2_antennanp ANTENNA_2915 (.A(net210));
 sg13g2_antennanp ANTENNA_2916 (.A(net210));
 sg13g2_antennanp ANTENNA_2917 (.A(net210));
 sg13g2_antennanp ANTENNA_2918 (.A(net210));
 sg13g2_antennanp ANTENNA_2919 (.A(net210));
 sg13g2_antennanp ANTENNA_2920 (.A(net210));
 sg13g2_antennanp ANTENNA_2921 (.A(net210));
 sg13g2_antennanp ANTENNA_2922 (.A(net210));
 sg13g2_antennanp ANTENNA_2923 (.A(net210));
 sg13g2_antennanp ANTENNA_2924 (.A(_0003_));
 sg13g2_antennanp ANTENNA_2925 (.A(_0016_));
 sg13g2_antennanp ANTENNA_2926 (.A(_0016_));
 sg13g2_antennanp ANTENNA_2927 (.A(_0018_));
 sg13g2_antennanp ANTENNA_2928 (.A(_0018_));
 sg13g2_antennanp ANTENNA_2929 (.A(_0021_));
 sg13g2_antennanp ANTENNA_2930 (.A(_0022_));
 sg13g2_antennanp ANTENNA_2931 (.A(_0023_));
 sg13g2_antennanp ANTENNA_2932 (.A(_0024_));
 sg13g2_antennanp ANTENNA_2933 (.A(_0025_));
 sg13g2_antennanp ANTENNA_2934 (.A(_0025_));
 sg13g2_antennanp ANTENNA_2935 (.A(_0027_));
 sg13g2_antennanp ANTENNA_2936 (.A(_0027_));
 sg13g2_antennanp ANTENNA_2937 (.A(_0028_));
 sg13g2_antennanp ANTENNA_2938 (.A(_0028_));
 sg13g2_antennanp ANTENNA_2939 (.A(_0038_));
 sg13g2_antennanp ANTENNA_2940 (.A(_0038_));
 sg13g2_antennanp ANTENNA_2941 (.A(_0038_));
 sg13g2_antennanp ANTENNA_2942 (.A(_0038_));
 sg13g2_antennanp ANTENNA_2943 (.A(_0038_));
 sg13g2_antennanp ANTENNA_2944 (.A(_0038_));
 sg13g2_antennanp ANTENNA_2945 (.A(_0038_));
 sg13g2_antennanp ANTENNA_2946 (.A(_0038_));
 sg13g2_antennanp ANTENNA_2947 (.A(_0038_));
 sg13g2_antennanp ANTENNA_2948 (.A(_0123_));
 sg13g2_antennanp ANTENNA_2949 (.A(_0123_));
 sg13g2_antennanp ANTENNA_2950 (.A(_0125_));
 sg13g2_antennanp ANTENNA_2951 (.A(_0125_));
 sg13g2_antennanp ANTENNA_2952 (.A(_0125_));
 sg13g2_antennanp ANTENNA_2953 (.A(_0150_));
 sg13g2_antennanp ANTENNA_2954 (.A(_0150_));
 sg13g2_antennanp ANTENNA_2955 (.A(_0150_));
 sg13g2_antennanp ANTENNA_2956 (.A(_0150_));
 sg13g2_antennanp ANTENNA_2957 (.A(_0150_));
 sg13g2_antennanp ANTENNA_2958 (.A(_0150_));
 sg13g2_antennanp ANTENNA_2959 (.A(_0158_));
 sg13g2_antennanp ANTENNA_2960 (.A(_0165_));
 sg13g2_antennanp ANTENNA_2961 (.A(_0165_));
 sg13g2_antennanp ANTENNA_2962 (.A(_0165_));
 sg13g2_antennanp ANTENNA_2963 (.A(_0165_));
 sg13g2_antennanp ANTENNA_2964 (.A(_0167_));
 sg13g2_antennanp ANTENNA_2965 (.A(_0167_));
 sg13g2_antennanp ANTENNA_2966 (.A(_0167_));
 sg13g2_antennanp ANTENNA_2967 (.A(_0167_));
 sg13g2_antennanp ANTENNA_2968 (.A(_0167_));
 sg13g2_antennanp ANTENNA_2969 (.A(_0167_));
 sg13g2_antennanp ANTENNA_2970 (.A(_0167_));
 sg13g2_antennanp ANTENNA_2971 (.A(_0167_));
 sg13g2_antennanp ANTENNA_2972 (.A(_0168_));
 sg13g2_antennanp ANTENNA_2973 (.A(_0168_));
 sg13g2_antennanp ANTENNA_2974 (.A(_0168_));
 sg13g2_antennanp ANTENNA_2975 (.A(_0168_));
 sg13g2_antennanp ANTENNA_2976 (.A(_0168_));
 sg13g2_antennanp ANTENNA_2977 (.A(_0168_));
 sg13g2_antennanp ANTENNA_2978 (.A(_0189_));
 sg13g2_antennanp ANTENNA_2979 (.A(_0230_));
 sg13g2_antennanp ANTENNA_2980 (.A(_0230_));
 sg13g2_antennanp ANTENNA_2981 (.A(_0260_));
 sg13g2_antennanp ANTENNA_2982 (.A(_0260_));
 sg13g2_antennanp ANTENNA_2983 (.A(_0260_));
 sg13g2_antennanp ANTENNA_2984 (.A(_0260_));
 sg13g2_antennanp ANTENNA_2985 (.A(_0269_));
 sg13g2_antennanp ANTENNA_2986 (.A(_0301_));
 sg13g2_antennanp ANTENNA_2987 (.A(_0345_));
 sg13g2_antennanp ANTENNA_2988 (.A(_0345_));
 sg13g2_antennanp ANTENNA_2989 (.A(_0345_));
 sg13g2_antennanp ANTENNA_2990 (.A(_0345_));
 sg13g2_antennanp ANTENNA_2991 (.A(_0346_));
 sg13g2_antennanp ANTENNA_2992 (.A(_0346_));
 sg13g2_antennanp ANTENNA_2993 (.A(_0346_));
 sg13g2_antennanp ANTENNA_2994 (.A(_0346_));
 sg13g2_antennanp ANTENNA_2995 (.A(_0360_));
 sg13g2_antennanp ANTENNA_2996 (.A(_0360_));
 sg13g2_antennanp ANTENNA_2997 (.A(_0360_));
 sg13g2_antennanp ANTENNA_2998 (.A(_0360_));
 sg13g2_antennanp ANTENNA_2999 (.A(_0360_));
 sg13g2_antennanp ANTENNA_3000 (.A(_0387_));
 sg13g2_antennanp ANTENNA_3001 (.A(_0387_));
 sg13g2_antennanp ANTENNA_3002 (.A(_0387_));
 sg13g2_antennanp ANTENNA_3003 (.A(_0387_));
 sg13g2_antennanp ANTENNA_3004 (.A(_0387_));
 sg13g2_antennanp ANTENNA_3005 (.A(_0387_));
 sg13g2_antennanp ANTENNA_3006 (.A(_0435_));
 sg13g2_antennanp ANTENNA_3007 (.A(_0435_));
 sg13g2_antennanp ANTENNA_3008 (.A(_0438_));
 sg13g2_antennanp ANTENNA_3009 (.A(_0438_));
 sg13g2_antennanp ANTENNA_3010 (.A(_0438_));
 sg13g2_antennanp ANTENNA_3011 (.A(_0438_));
 sg13g2_antennanp ANTENNA_3012 (.A(_0438_));
 sg13g2_antennanp ANTENNA_3013 (.A(_0438_));
 sg13g2_antennanp ANTENNA_3014 (.A(_0448_));
 sg13g2_antennanp ANTENNA_3015 (.A(_0490_));
 sg13g2_antennanp ANTENNA_3016 (.A(_0490_));
 sg13g2_antennanp ANTENNA_3017 (.A(_0507_));
 sg13g2_antennanp ANTENNA_3018 (.A(_0507_));
 sg13g2_antennanp ANTENNA_3019 (.A(_0511_));
 sg13g2_antennanp ANTENNA_3020 (.A(_0511_));
 sg13g2_antennanp ANTENNA_3021 (.A(_0511_));
 sg13g2_antennanp ANTENNA_3022 (.A(_0521_));
 sg13g2_antennanp ANTENNA_3023 (.A(_0521_));
 sg13g2_antennanp ANTENNA_3024 (.A(_0521_));
 sg13g2_antennanp ANTENNA_3025 (.A(_0597_));
 sg13g2_antennanp ANTENNA_3026 (.A(_0597_));
 sg13g2_antennanp ANTENNA_3027 (.A(_0597_));
 sg13g2_antennanp ANTENNA_3028 (.A(_0597_));
 sg13g2_antennanp ANTENNA_3029 (.A(_0597_));
 sg13g2_antennanp ANTENNA_3030 (.A(_0598_));
 sg13g2_antennanp ANTENNA_3031 (.A(_0598_));
 sg13g2_antennanp ANTENNA_3032 (.A(_0598_));
 sg13g2_antennanp ANTENNA_3033 (.A(_0598_));
 sg13g2_antennanp ANTENNA_3034 (.A(_0598_));
 sg13g2_antennanp ANTENNA_3035 (.A(_0623_));
 sg13g2_antennanp ANTENNA_3036 (.A(_0780_));
 sg13g2_antennanp ANTENNA_3037 (.A(_0800_));
 sg13g2_antennanp ANTENNA_3038 (.A(_0866_));
 sg13g2_antennanp ANTENNA_3039 (.A(_0866_));
 sg13g2_antennanp ANTENNA_3040 (.A(_0866_));
 sg13g2_antennanp ANTENNA_3041 (.A(_0878_));
 sg13g2_antennanp ANTENNA_3042 (.A(_0878_));
 sg13g2_antennanp ANTENNA_3043 (.A(_0878_));
 sg13g2_antennanp ANTENNA_3044 (.A(_0878_));
 sg13g2_antennanp ANTENNA_3045 (.A(_0878_));
 sg13g2_antennanp ANTENNA_3046 (.A(_0878_));
 sg13g2_antennanp ANTENNA_3047 (.A(_0878_));
 sg13g2_antennanp ANTENNA_3048 (.A(_0878_));
 sg13g2_antennanp ANTENNA_3049 (.A(_0878_));
 sg13g2_antennanp ANTENNA_3050 (.A(_1002_));
 sg13g2_antennanp ANTENNA_3051 (.A(_1002_));
 sg13g2_antennanp ANTENNA_3052 (.A(_1071_));
 sg13g2_antennanp ANTENNA_3053 (.A(_1071_));
 sg13g2_antennanp ANTENNA_3054 (.A(_1071_));
 sg13g2_antennanp ANTENNA_3055 (.A(_1085_));
 sg13g2_antennanp ANTENNA_3056 (.A(_1085_));
 sg13g2_antennanp ANTENNA_3057 (.A(_1085_));
 sg13g2_antennanp ANTENNA_3058 (.A(_1085_));
 sg13g2_antennanp ANTENNA_3059 (.A(_1085_));
 sg13g2_antennanp ANTENNA_3060 (.A(_1085_));
 sg13g2_antennanp ANTENNA_3061 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3062 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3063 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3064 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3065 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3066 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3067 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3068 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3069 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3070 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3071 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3072 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3073 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3074 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3075 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3076 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3077 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3078 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3079 (.A(_1225_));
 sg13g2_antennanp ANTENNA_3080 (.A(_1225_));
 sg13g2_antennanp ANTENNA_3081 (.A(_1292_));
 sg13g2_antennanp ANTENNA_3082 (.A(_1292_));
 sg13g2_antennanp ANTENNA_3083 (.A(_1326_));
 sg13g2_antennanp ANTENNA_3084 (.A(_1326_));
 sg13g2_antennanp ANTENNA_3085 (.A(_1326_));
 sg13g2_antennanp ANTENNA_3086 (.A(_1326_));
 sg13g2_antennanp ANTENNA_3087 (.A(_1326_));
 sg13g2_antennanp ANTENNA_3088 (.A(_1326_));
 sg13g2_antennanp ANTENNA_3089 (.A(_1326_));
 sg13g2_antennanp ANTENNA_3090 (.A(_1326_));
 sg13g2_antennanp ANTENNA_3091 (.A(_1326_));
 sg13g2_antennanp ANTENNA_3092 (.A(_1363_));
 sg13g2_antennanp ANTENNA_3093 (.A(_1363_));
 sg13g2_antennanp ANTENNA_3094 (.A(_1411_));
 sg13g2_antennanp ANTENNA_3095 (.A(_1439_));
 sg13g2_antennanp ANTENNA_3096 (.A(_1470_));
 sg13g2_antennanp ANTENNA_3097 (.A(_1470_));
 sg13g2_antennanp ANTENNA_3098 (.A(_1519_));
 sg13g2_antennanp ANTENNA_3099 (.A(_1531_));
 sg13g2_antennanp ANTENNA_3100 (.A(_1531_));
 sg13g2_antennanp ANTENNA_3101 (.A(_1532_));
 sg13g2_antennanp ANTENNA_3102 (.A(_1532_));
 sg13g2_antennanp ANTENNA_3103 (.A(_1532_));
 sg13g2_antennanp ANTENNA_3104 (.A(_1544_));
 sg13g2_antennanp ANTENNA_3105 (.A(_1544_));
 sg13g2_antennanp ANTENNA_3106 (.A(_1544_));
 sg13g2_antennanp ANTENNA_3107 (.A(_1544_));
 sg13g2_antennanp ANTENNA_3108 (.A(_1544_));
 sg13g2_antennanp ANTENNA_3109 (.A(_1553_));
 sg13g2_antennanp ANTENNA_3110 (.A(_1631_));
 sg13g2_antennanp ANTENNA_3111 (.A(_1631_));
 sg13g2_antennanp ANTENNA_3112 (.A(_1631_));
 sg13g2_antennanp ANTENNA_3113 (.A(_1685_));
 sg13g2_antennanp ANTENNA_3114 (.A(_1685_));
 sg13g2_antennanp ANTENNA_3115 (.A(_1685_));
 sg13g2_antennanp ANTENNA_3116 (.A(_1685_));
 sg13g2_antennanp ANTENNA_3117 (.A(_1696_));
 sg13g2_antennanp ANTENNA_3118 (.A(_1696_));
 sg13g2_antennanp ANTENNA_3119 (.A(_1696_));
 sg13g2_antennanp ANTENNA_3120 (.A(_1696_));
 sg13g2_antennanp ANTENNA_3121 (.A(_1696_));
 sg13g2_antennanp ANTENNA_3122 (.A(_1696_));
 sg13g2_antennanp ANTENNA_3123 (.A(_1696_));
 sg13g2_antennanp ANTENNA_3124 (.A(_1696_));
 sg13g2_antennanp ANTENNA_3125 (.A(_1696_));
 sg13g2_antennanp ANTENNA_3126 (.A(_1696_));
 sg13g2_antennanp ANTENNA_3127 (.A(_1707_));
 sg13g2_antennanp ANTENNA_3128 (.A(_1707_));
 sg13g2_antennanp ANTENNA_3129 (.A(_1707_));
 sg13g2_antennanp ANTENNA_3130 (.A(_1716_));
 sg13g2_antennanp ANTENNA_3131 (.A(_1735_));
 sg13g2_antennanp ANTENNA_3132 (.A(_1761_));
 sg13g2_antennanp ANTENNA_3133 (.A(_2014_));
 sg13g2_antennanp ANTENNA_3134 (.A(_2014_));
 sg13g2_antennanp ANTENNA_3135 (.A(_2037_));
 sg13g2_antennanp ANTENNA_3136 (.A(_2053_));
 sg13g2_antennanp ANTENNA_3137 (.A(_2053_));
 sg13g2_antennanp ANTENNA_3138 (.A(_2053_));
 sg13g2_antennanp ANTENNA_3139 (.A(_2097_));
 sg13g2_antennanp ANTENNA_3140 (.A(_2097_));
 sg13g2_antennanp ANTENNA_3141 (.A(_2097_));
 sg13g2_antennanp ANTENNA_3142 (.A(_2097_));
 sg13g2_antennanp ANTENNA_3143 (.A(_2097_));
 sg13g2_antennanp ANTENNA_3144 (.A(_2110_));
 sg13g2_antennanp ANTENNA_3145 (.A(_2110_));
 sg13g2_antennanp ANTENNA_3146 (.A(_2112_));
 sg13g2_antennanp ANTENNA_3147 (.A(_2145_));
 sg13g2_antennanp ANTENNA_3148 (.A(_2171_));
 sg13g2_antennanp ANTENNA_3149 (.A(_2171_));
 sg13g2_antennanp ANTENNA_3150 (.A(_2171_));
 sg13g2_antennanp ANTENNA_3151 (.A(_2171_));
 sg13g2_antennanp ANTENNA_3152 (.A(_2171_));
 sg13g2_antennanp ANTENNA_3153 (.A(_2171_));
 sg13g2_antennanp ANTENNA_3154 (.A(_2171_));
 sg13g2_antennanp ANTENNA_3155 (.A(_2171_));
 sg13g2_antennanp ANTENNA_3156 (.A(_2171_));
 sg13g2_antennanp ANTENNA_3157 (.A(_2172_));
 sg13g2_antennanp ANTENNA_3158 (.A(_2172_));
 sg13g2_antennanp ANTENNA_3159 (.A(_2172_));
 sg13g2_antennanp ANTENNA_3160 (.A(_2172_));
 sg13g2_antennanp ANTENNA_3161 (.A(_2172_));
 sg13g2_antennanp ANTENNA_3162 (.A(_2172_));
 sg13g2_antennanp ANTENNA_3163 (.A(_2172_));
 sg13g2_antennanp ANTENNA_3164 (.A(_2172_));
 sg13g2_antennanp ANTENNA_3165 (.A(_2172_));
 sg13g2_antennanp ANTENNA_3166 (.A(_2172_));
 sg13g2_antennanp ANTENNA_3167 (.A(_2257_));
 sg13g2_antennanp ANTENNA_3168 (.A(_2257_));
 sg13g2_antennanp ANTENNA_3169 (.A(_2430_));
 sg13g2_antennanp ANTENNA_3170 (.A(_2430_));
 sg13g2_antennanp ANTENNA_3171 (.A(_2430_));
 sg13g2_antennanp ANTENNA_3172 (.A(_2430_));
 sg13g2_antennanp ANTENNA_3173 (.A(_2430_));
 sg13g2_antennanp ANTENNA_3174 (.A(_2430_));
 sg13g2_antennanp ANTENNA_3175 (.A(_2467_));
 sg13g2_antennanp ANTENNA_3176 (.A(_2467_));
 sg13g2_antennanp ANTENNA_3177 (.A(_2467_));
 sg13g2_antennanp ANTENNA_3178 (.A(_2467_));
 sg13g2_antennanp ANTENNA_3179 (.A(_2467_));
 sg13g2_antennanp ANTENNA_3180 (.A(_2470_));
 sg13g2_antennanp ANTENNA_3181 (.A(_2470_));
 sg13g2_antennanp ANTENNA_3182 (.A(_2470_));
 sg13g2_antennanp ANTENNA_3183 (.A(_2470_));
 sg13g2_antennanp ANTENNA_3184 (.A(_2480_));
 sg13g2_antennanp ANTENNA_3185 (.A(_2480_));
 sg13g2_antennanp ANTENNA_3186 (.A(_2480_));
 sg13g2_antennanp ANTENNA_3187 (.A(_2480_));
 sg13g2_antennanp ANTENNA_3188 (.A(_2480_));
 sg13g2_antennanp ANTENNA_3189 (.A(_2480_));
 sg13g2_antennanp ANTENNA_3190 (.A(_2480_));
 sg13g2_antennanp ANTENNA_3191 (.A(_2480_));
 sg13g2_antennanp ANTENNA_3192 (.A(_2482_));
 sg13g2_antennanp ANTENNA_3193 (.A(_2482_));
 sg13g2_antennanp ANTENNA_3194 (.A(_2482_));
 sg13g2_antennanp ANTENNA_3195 (.A(_2482_));
 sg13g2_antennanp ANTENNA_3196 (.A(_2482_));
 sg13g2_antennanp ANTENNA_3197 (.A(_2482_));
 sg13g2_antennanp ANTENNA_3198 (.A(_2482_));
 sg13g2_antennanp ANTENNA_3199 (.A(_2487_));
 sg13g2_antennanp ANTENNA_3200 (.A(_2487_));
 sg13g2_antennanp ANTENNA_3201 (.A(_2501_));
 sg13g2_antennanp ANTENNA_3202 (.A(_2501_));
 sg13g2_antennanp ANTENNA_3203 (.A(_2501_));
 sg13g2_antennanp ANTENNA_3204 (.A(_2501_));
 sg13g2_antennanp ANTENNA_3205 (.A(_2501_));
 sg13g2_antennanp ANTENNA_3206 (.A(_2501_));
 sg13g2_antennanp ANTENNA_3207 (.A(_2520_));
 sg13g2_antennanp ANTENNA_3208 (.A(_2520_));
 sg13g2_antennanp ANTENNA_3209 (.A(_2520_));
 sg13g2_antennanp ANTENNA_3210 (.A(_2520_));
 sg13g2_antennanp ANTENNA_3211 (.A(_2520_));
 sg13g2_antennanp ANTENNA_3212 (.A(_2520_));
 sg13g2_antennanp ANTENNA_3213 (.A(_2530_));
 sg13g2_antennanp ANTENNA_3214 (.A(_2530_));
 sg13g2_antennanp ANTENNA_3215 (.A(_2530_));
 sg13g2_antennanp ANTENNA_3216 (.A(_2530_));
 sg13g2_antennanp ANTENNA_3217 (.A(_2537_));
 sg13g2_antennanp ANTENNA_3218 (.A(_2537_));
 sg13g2_antennanp ANTENNA_3219 (.A(_2537_));
 sg13g2_antennanp ANTENNA_3220 (.A(_2537_));
 sg13g2_antennanp ANTENNA_3221 (.A(_2573_));
 sg13g2_antennanp ANTENNA_3222 (.A(_2573_));
 sg13g2_antennanp ANTENNA_3223 (.A(_2573_));
 sg13g2_antennanp ANTENNA_3224 (.A(_2573_));
 sg13g2_antennanp ANTENNA_3225 (.A(_2577_));
 sg13g2_antennanp ANTENNA_3226 (.A(_2577_));
 sg13g2_antennanp ANTENNA_3227 (.A(_2577_));
 sg13g2_antennanp ANTENNA_3228 (.A(_2577_));
 sg13g2_antennanp ANTENNA_3229 (.A(_2577_));
 sg13g2_antennanp ANTENNA_3230 (.A(_2577_));
 sg13g2_antennanp ANTENNA_3231 (.A(_2577_));
 sg13g2_antennanp ANTENNA_3232 (.A(_2577_));
 sg13g2_antennanp ANTENNA_3233 (.A(_2585_));
 sg13g2_antennanp ANTENNA_3234 (.A(_2585_));
 sg13g2_antennanp ANTENNA_3235 (.A(_2585_));
 sg13g2_antennanp ANTENNA_3236 (.A(_2585_));
 sg13g2_antennanp ANTENNA_3237 (.A(_2588_));
 sg13g2_antennanp ANTENNA_3238 (.A(_2595_));
 sg13g2_antennanp ANTENNA_3239 (.A(_2595_));
 sg13g2_antennanp ANTENNA_3240 (.A(_2595_));
 sg13g2_antennanp ANTENNA_3241 (.A(_2595_));
 sg13g2_antennanp ANTENNA_3242 (.A(_2600_));
 sg13g2_antennanp ANTENNA_3243 (.A(_2600_));
 sg13g2_antennanp ANTENNA_3244 (.A(_2600_));
 sg13g2_antennanp ANTENNA_3245 (.A(_2600_));
 sg13g2_antennanp ANTENNA_3246 (.A(_2607_));
 sg13g2_antennanp ANTENNA_3247 (.A(_2607_));
 sg13g2_antennanp ANTENNA_3248 (.A(_2615_));
 sg13g2_antennanp ANTENNA_3249 (.A(_2615_));
 sg13g2_antennanp ANTENNA_3250 (.A(_2615_));
 sg13g2_antennanp ANTENNA_3251 (.A(_2619_));
 sg13g2_antennanp ANTENNA_3252 (.A(_2619_));
 sg13g2_antennanp ANTENNA_3253 (.A(_2619_));
 sg13g2_antennanp ANTENNA_3254 (.A(_2619_));
 sg13g2_antennanp ANTENNA_3255 (.A(_2619_));
 sg13g2_antennanp ANTENNA_3256 (.A(_2619_));
 sg13g2_antennanp ANTENNA_3257 (.A(_2622_));
 sg13g2_antennanp ANTENNA_3258 (.A(_2622_));
 sg13g2_antennanp ANTENNA_3259 (.A(_2622_));
 sg13g2_antennanp ANTENNA_3260 (.A(_2622_));
 sg13g2_antennanp ANTENNA_3261 (.A(_2622_));
 sg13g2_antennanp ANTENNA_3262 (.A(_2622_));
 sg13g2_antennanp ANTENNA_3263 (.A(_2625_));
 sg13g2_antennanp ANTENNA_3264 (.A(_2625_));
 sg13g2_antennanp ANTENNA_3265 (.A(_2625_));
 sg13g2_antennanp ANTENNA_3266 (.A(_2625_));
 sg13g2_antennanp ANTENNA_3267 (.A(_2659_));
 sg13g2_antennanp ANTENNA_3268 (.A(_2659_));
 sg13g2_antennanp ANTENNA_3269 (.A(_2659_));
 sg13g2_antennanp ANTENNA_3270 (.A(_2659_));
 sg13g2_antennanp ANTENNA_3271 (.A(_2659_));
 sg13g2_antennanp ANTENNA_3272 (.A(_2665_));
 sg13g2_antennanp ANTENNA_3273 (.A(_2665_));
 sg13g2_antennanp ANTENNA_3274 (.A(_2665_));
 sg13g2_antennanp ANTENNA_3275 (.A(_2665_));
 sg13g2_antennanp ANTENNA_3276 (.A(_2678_));
 sg13g2_antennanp ANTENNA_3277 (.A(_2678_));
 sg13g2_antennanp ANTENNA_3278 (.A(_2678_));
 sg13g2_antennanp ANTENNA_3279 (.A(_2678_));
 sg13g2_antennanp ANTENNA_3280 (.A(_2678_));
 sg13g2_antennanp ANTENNA_3281 (.A(_2678_));
 sg13g2_antennanp ANTENNA_3282 (.A(_2678_));
 sg13g2_antennanp ANTENNA_3283 (.A(_2732_));
 sg13g2_antennanp ANTENNA_3284 (.A(_2732_));
 sg13g2_antennanp ANTENNA_3285 (.A(_2732_));
 sg13g2_antennanp ANTENNA_3286 (.A(_2733_));
 sg13g2_antennanp ANTENNA_3287 (.A(_2733_));
 sg13g2_antennanp ANTENNA_3288 (.A(_2733_));
 sg13g2_antennanp ANTENNA_3289 (.A(_2733_));
 sg13g2_antennanp ANTENNA_3290 (.A(_2739_));
 sg13g2_antennanp ANTENNA_3291 (.A(_2739_));
 sg13g2_antennanp ANTENNA_3292 (.A(_2739_));
 sg13g2_antennanp ANTENNA_3293 (.A(_2739_));
 sg13g2_antennanp ANTENNA_3294 (.A(_2769_));
 sg13g2_antennanp ANTENNA_3295 (.A(_2769_));
 sg13g2_antennanp ANTENNA_3296 (.A(_2769_));
 sg13g2_antennanp ANTENNA_3297 (.A(_2769_));
 sg13g2_antennanp ANTENNA_3298 (.A(_2789_));
 sg13g2_antennanp ANTENNA_3299 (.A(_2789_));
 sg13g2_antennanp ANTENNA_3300 (.A(_2789_));
 sg13g2_antennanp ANTENNA_3301 (.A(_2789_));
 sg13g2_antennanp ANTENNA_3302 (.A(_2805_));
 sg13g2_antennanp ANTENNA_3303 (.A(_2805_));
 sg13g2_antennanp ANTENNA_3304 (.A(_2808_));
 sg13g2_antennanp ANTENNA_3305 (.A(_2808_));
 sg13g2_antennanp ANTENNA_3306 (.A(_2808_));
 sg13g2_antennanp ANTENNA_3307 (.A(_2808_));
 sg13g2_antennanp ANTENNA_3308 (.A(_2826_));
 sg13g2_antennanp ANTENNA_3309 (.A(_2826_));
 sg13g2_antennanp ANTENNA_3310 (.A(_2826_));
 sg13g2_antennanp ANTENNA_3311 (.A(_2826_));
 sg13g2_antennanp ANTENNA_3312 (.A(_2858_));
 sg13g2_antennanp ANTENNA_3313 (.A(_2858_));
 sg13g2_antennanp ANTENNA_3314 (.A(_2879_));
 sg13g2_antennanp ANTENNA_3315 (.A(_2879_));
 sg13g2_antennanp ANTENNA_3316 (.A(_2879_));
 sg13g2_antennanp ANTENNA_3317 (.A(_2879_));
 sg13g2_antennanp ANTENNA_3318 (.A(_2879_));
 sg13g2_antennanp ANTENNA_3319 (.A(_2879_));
 sg13g2_antennanp ANTENNA_3320 (.A(_2879_));
 sg13g2_antennanp ANTENNA_3321 (.A(_2879_));
 sg13g2_antennanp ANTENNA_3322 (.A(_2914_));
 sg13g2_antennanp ANTENNA_3323 (.A(_2931_));
 sg13g2_antennanp ANTENNA_3324 (.A(_2931_));
 sg13g2_antennanp ANTENNA_3325 (.A(_2931_));
 sg13g2_antennanp ANTENNA_3326 (.A(_2931_));
 sg13g2_antennanp ANTENNA_3327 (.A(_2936_));
 sg13g2_antennanp ANTENNA_3328 (.A(_2936_));
 sg13g2_antennanp ANTENNA_3329 (.A(_2936_));
 sg13g2_antennanp ANTENNA_3330 (.A(_2957_));
 sg13g2_antennanp ANTENNA_3331 (.A(_2957_));
 sg13g2_antennanp ANTENNA_3332 (.A(_2957_));
 sg13g2_antennanp ANTENNA_3333 (.A(_2957_));
 sg13g2_antennanp ANTENNA_3334 (.A(_2970_));
 sg13g2_antennanp ANTENNA_3335 (.A(_2970_));
 sg13g2_antennanp ANTENNA_3336 (.A(_2970_));
 sg13g2_antennanp ANTENNA_3337 (.A(_2970_));
 sg13g2_antennanp ANTENNA_3338 (.A(_2974_));
 sg13g2_antennanp ANTENNA_3339 (.A(_2974_));
 sg13g2_antennanp ANTENNA_3340 (.A(_2977_));
 sg13g2_antennanp ANTENNA_3341 (.A(_2977_));
 sg13g2_antennanp ANTENNA_3342 (.A(_2977_));
 sg13g2_antennanp ANTENNA_3343 (.A(_2977_));
 sg13g2_antennanp ANTENNA_3344 (.A(_2977_));
 sg13g2_antennanp ANTENNA_3345 (.A(_2986_));
 sg13g2_antennanp ANTENNA_3346 (.A(_2986_));
 sg13g2_antennanp ANTENNA_3347 (.A(_2986_));
 sg13g2_antennanp ANTENNA_3348 (.A(_2986_));
 sg13g2_antennanp ANTENNA_3349 (.A(_3018_));
 sg13g2_antennanp ANTENNA_3350 (.A(_3018_));
 sg13g2_antennanp ANTENNA_3351 (.A(_3018_));
 sg13g2_antennanp ANTENNA_3352 (.A(clk));
 sg13g2_antennanp ANTENNA_3353 (.A(clk));
 sg13g2_antennanp ANTENNA_3354 (.A(net22));
 sg13g2_antennanp ANTENNA_3355 (.A(net22));
 sg13g2_antennanp ANTENNA_3356 (.A(net22));
 sg13g2_antennanp ANTENNA_3357 (.A(net22));
 sg13g2_antennanp ANTENNA_3358 (.A(net22));
 sg13g2_antennanp ANTENNA_3359 (.A(net22));
 sg13g2_antennanp ANTENNA_3360 (.A(net22));
 sg13g2_antennanp ANTENNA_3361 (.A(net22));
 sg13g2_antennanp ANTENNA_3362 (.A(net22));
 sg13g2_antennanp ANTENNA_3363 (.A(net23));
 sg13g2_antennanp ANTENNA_3364 (.A(net23));
 sg13g2_antennanp ANTENNA_3365 (.A(net23));
 sg13g2_antennanp ANTENNA_3366 (.A(net23));
 sg13g2_antennanp ANTENNA_3367 (.A(net23));
 sg13g2_antennanp ANTENNA_3368 (.A(net23));
 sg13g2_antennanp ANTENNA_3369 (.A(net23));
 sg13g2_antennanp ANTENNA_3370 (.A(net23));
 sg13g2_antennanp ANTENNA_3371 (.A(net29));
 sg13g2_antennanp ANTENNA_3372 (.A(net29));
 sg13g2_antennanp ANTENNA_3373 (.A(net29));
 sg13g2_antennanp ANTENNA_3374 (.A(net29));
 sg13g2_antennanp ANTENNA_3375 (.A(net29));
 sg13g2_antennanp ANTENNA_3376 (.A(net29));
 sg13g2_antennanp ANTENNA_3377 (.A(net29));
 sg13g2_antennanp ANTENNA_3378 (.A(net29));
 sg13g2_antennanp ANTENNA_3379 (.A(net29));
 sg13g2_antennanp ANTENNA_3380 (.A(net35));
 sg13g2_antennanp ANTENNA_3381 (.A(net35));
 sg13g2_antennanp ANTENNA_3382 (.A(net35));
 sg13g2_antennanp ANTENNA_3383 (.A(net35));
 sg13g2_antennanp ANTENNA_3384 (.A(net35));
 sg13g2_antennanp ANTENNA_3385 (.A(net35));
 sg13g2_antennanp ANTENNA_3386 (.A(net35));
 sg13g2_antennanp ANTENNA_3387 (.A(net35));
 sg13g2_antennanp ANTENNA_3388 (.A(net35));
 sg13g2_antennanp ANTENNA_3389 (.A(net46));
 sg13g2_antennanp ANTENNA_3390 (.A(net46));
 sg13g2_antennanp ANTENNA_3391 (.A(net46));
 sg13g2_antennanp ANTENNA_3392 (.A(net46));
 sg13g2_antennanp ANTENNA_3393 (.A(net46));
 sg13g2_antennanp ANTENNA_3394 (.A(net46));
 sg13g2_antennanp ANTENNA_3395 (.A(net46));
 sg13g2_antennanp ANTENNA_3396 (.A(net46));
 sg13g2_antennanp ANTENNA_3397 (.A(net53));
 sg13g2_antennanp ANTENNA_3398 (.A(net53));
 sg13g2_antennanp ANTENNA_3399 (.A(net53));
 sg13g2_antennanp ANTENNA_3400 (.A(net53));
 sg13g2_antennanp ANTENNA_3401 (.A(net53));
 sg13g2_antennanp ANTENNA_3402 (.A(net53));
 sg13g2_antennanp ANTENNA_3403 (.A(net53));
 sg13g2_antennanp ANTENNA_3404 (.A(net53));
 sg13g2_antennanp ANTENNA_3405 (.A(net59));
 sg13g2_antennanp ANTENNA_3406 (.A(net59));
 sg13g2_antennanp ANTENNA_3407 (.A(net59));
 sg13g2_antennanp ANTENNA_3408 (.A(net59));
 sg13g2_antennanp ANTENNA_3409 (.A(net59));
 sg13g2_antennanp ANTENNA_3410 (.A(net59));
 sg13g2_antennanp ANTENNA_3411 (.A(net59));
 sg13g2_antennanp ANTENNA_3412 (.A(net59));
 sg13g2_antennanp ANTENNA_3413 (.A(net59));
 sg13g2_antennanp ANTENNA_3414 (.A(net61));
 sg13g2_antennanp ANTENNA_3415 (.A(net61));
 sg13g2_antennanp ANTENNA_3416 (.A(net61));
 sg13g2_antennanp ANTENNA_3417 (.A(net61));
 sg13g2_antennanp ANTENNA_3418 (.A(net61));
 sg13g2_antennanp ANTENNA_3419 (.A(net61));
 sg13g2_antennanp ANTENNA_3420 (.A(net61));
 sg13g2_antennanp ANTENNA_3421 (.A(net61));
 sg13g2_antennanp ANTENNA_3422 (.A(net61));
 sg13g2_antennanp ANTENNA_3423 (.A(net62));
 sg13g2_antennanp ANTENNA_3424 (.A(net62));
 sg13g2_antennanp ANTENNA_3425 (.A(net62));
 sg13g2_antennanp ANTENNA_3426 (.A(net62));
 sg13g2_antennanp ANTENNA_3427 (.A(net62));
 sg13g2_antennanp ANTENNA_3428 (.A(net62));
 sg13g2_antennanp ANTENNA_3429 (.A(net62));
 sg13g2_antennanp ANTENNA_3430 (.A(net62));
 sg13g2_antennanp ANTENNA_3431 (.A(net62));
 sg13g2_antennanp ANTENNA_3432 (.A(net64));
 sg13g2_antennanp ANTENNA_3433 (.A(net64));
 sg13g2_antennanp ANTENNA_3434 (.A(net64));
 sg13g2_antennanp ANTENNA_3435 (.A(net64));
 sg13g2_antennanp ANTENNA_3436 (.A(net64));
 sg13g2_antennanp ANTENNA_3437 (.A(net64));
 sg13g2_antennanp ANTENNA_3438 (.A(net64));
 sg13g2_antennanp ANTENNA_3439 (.A(net64));
 sg13g2_antennanp ANTENNA_3440 (.A(net70));
 sg13g2_antennanp ANTENNA_3441 (.A(net70));
 sg13g2_antennanp ANTENNA_3442 (.A(net70));
 sg13g2_antennanp ANTENNA_3443 (.A(net70));
 sg13g2_antennanp ANTENNA_3444 (.A(net70));
 sg13g2_antennanp ANTENNA_3445 (.A(net70));
 sg13g2_antennanp ANTENNA_3446 (.A(net70));
 sg13g2_antennanp ANTENNA_3447 (.A(net70));
 sg13g2_antennanp ANTENNA_3448 (.A(net71));
 sg13g2_antennanp ANTENNA_3449 (.A(net71));
 sg13g2_antennanp ANTENNA_3450 (.A(net71));
 sg13g2_antennanp ANTENNA_3451 (.A(net71));
 sg13g2_antennanp ANTENNA_3452 (.A(net71));
 sg13g2_antennanp ANTENNA_3453 (.A(net71));
 sg13g2_antennanp ANTENNA_3454 (.A(net71));
 sg13g2_antennanp ANTENNA_3455 (.A(net71));
 sg13g2_antennanp ANTENNA_3456 (.A(net71));
 sg13g2_antennanp ANTENNA_3457 (.A(net71));
 sg13g2_antennanp ANTENNA_3458 (.A(net71));
 sg13g2_antennanp ANTENNA_3459 (.A(net71));
 sg13g2_antennanp ANTENNA_3460 (.A(net71));
 sg13g2_antennanp ANTENNA_3461 (.A(net71));
 sg13g2_antennanp ANTENNA_3462 (.A(net71));
 sg13g2_antennanp ANTENNA_3463 (.A(net71));
 sg13g2_antennanp ANTENNA_3464 (.A(net76));
 sg13g2_antennanp ANTENNA_3465 (.A(net76));
 sg13g2_antennanp ANTENNA_3466 (.A(net76));
 sg13g2_antennanp ANTENNA_3467 (.A(net76));
 sg13g2_antennanp ANTENNA_3468 (.A(net76));
 sg13g2_antennanp ANTENNA_3469 (.A(net76));
 sg13g2_antennanp ANTENNA_3470 (.A(net76));
 sg13g2_antennanp ANTENNA_3471 (.A(net76));
 sg13g2_antennanp ANTENNA_3472 (.A(net76));
 sg13g2_antennanp ANTENNA_3473 (.A(net78));
 sg13g2_antennanp ANTENNA_3474 (.A(net78));
 sg13g2_antennanp ANTENNA_3475 (.A(net78));
 sg13g2_antennanp ANTENNA_3476 (.A(net78));
 sg13g2_antennanp ANTENNA_3477 (.A(net78));
 sg13g2_antennanp ANTENNA_3478 (.A(net78));
 sg13g2_antennanp ANTENNA_3479 (.A(net78));
 sg13g2_antennanp ANTENNA_3480 (.A(net78));
 sg13g2_antennanp ANTENNA_3481 (.A(net78));
 sg13g2_antennanp ANTENNA_3482 (.A(net79));
 sg13g2_antennanp ANTENNA_3483 (.A(net79));
 sg13g2_antennanp ANTENNA_3484 (.A(net79));
 sg13g2_antennanp ANTENNA_3485 (.A(net79));
 sg13g2_antennanp ANTENNA_3486 (.A(net79));
 sg13g2_antennanp ANTENNA_3487 (.A(net79));
 sg13g2_antennanp ANTENNA_3488 (.A(net79));
 sg13g2_antennanp ANTENNA_3489 (.A(net79));
 sg13g2_antennanp ANTENNA_3490 (.A(net79));
 sg13g2_antennanp ANTENNA_3491 (.A(net84));
 sg13g2_antennanp ANTENNA_3492 (.A(net84));
 sg13g2_antennanp ANTENNA_3493 (.A(net84));
 sg13g2_antennanp ANTENNA_3494 (.A(net84));
 sg13g2_antennanp ANTENNA_3495 (.A(net84));
 sg13g2_antennanp ANTENNA_3496 (.A(net84));
 sg13g2_antennanp ANTENNA_3497 (.A(net84));
 sg13g2_antennanp ANTENNA_3498 (.A(net84));
 sg13g2_antennanp ANTENNA_3499 (.A(net89));
 sg13g2_antennanp ANTENNA_3500 (.A(net89));
 sg13g2_antennanp ANTENNA_3501 (.A(net89));
 sg13g2_antennanp ANTENNA_3502 (.A(net89));
 sg13g2_antennanp ANTENNA_3503 (.A(net89));
 sg13g2_antennanp ANTENNA_3504 (.A(net89));
 sg13g2_antennanp ANTENNA_3505 (.A(net89));
 sg13g2_antennanp ANTENNA_3506 (.A(net89));
 sg13g2_antennanp ANTENNA_3507 (.A(net89));
 sg13g2_antennanp ANTENNA_3508 (.A(net91));
 sg13g2_antennanp ANTENNA_3509 (.A(net91));
 sg13g2_antennanp ANTENNA_3510 (.A(net91));
 sg13g2_antennanp ANTENNA_3511 (.A(net91));
 sg13g2_antennanp ANTENNA_3512 (.A(net91));
 sg13g2_antennanp ANTENNA_3513 (.A(net91));
 sg13g2_antennanp ANTENNA_3514 (.A(net91));
 sg13g2_antennanp ANTENNA_3515 (.A(net91));
 sg13g2_antennanp ANTENNA_3516 (.A(net94));
 sg13g2_antennanp ANTENNA_3517 (.A(net94));
 sg13g2_antennanp ANTENNA_3518 (.A(net94));
 sg13g2_antennanp ANTENNA_3519 (.A(net94));
 sg13g2_antennanp ANTENNA_3520 (.A(net94));
 sg13g2_antennanp ANTENNA_3521 (.A(net94));
 sg13g2_antennanp ANTENNA_3522 (.A(net94));
 sg13g2_antennanp ANTENNA_3523 (.A(net94));
 sg13g2_antennanp ANTENNA_3524 (.A(net100));
 sg13g2_antennanp ANTENNA_3525 (.A(net100));
 sg13g2_antennanp ANTENNA_3526 (.A(net100));
 sg13g2_antennanp ANTENNA_3527 (.A(net100));
 sg13g2_antennanp ANTENNA_3528 (.A(net100));
 sg13g2_antennanp ANTENNA_3529 (.A(net100));
 sg13g2_antennanp ANTENNA_3530 (.A(net100));
 sg13g2_antennanp ANTENNA_3531 (.A(net100));
 sg13g2_antennanp ANTENNA_3532 (.A(net100));
 sg13g2_antennanp ANTENNA_3533 (.A(net106));
 sg13g2_antennanp ANTENNA_3534 (.A(net106));
 sg13g2_antennanp ANTENNA_3535 (.A(net106));
 sg13g2_antennanp ANTENNA_3536 (.A(net106));
 sg13g2_antennanp ANTENNA_3537 (.A(net106));
 sg13g2_antennanp ANTENNA_3538 (.A(net106));
 sg13g2_antennanp ANTENNA_3539 (.A(net106));
 sg13g2_antennanp ANTENNA_3540 (.A(net106));
 sg13g2_antennanp ANTENNA_3541 (.A(net106));
 sg13g2_antennanp ANTENNA_3542 (.A(net107));
 sg13g2_antennanp ANTENNA_3543 (.A(net107));
 sg13g2_antennanp ANTENNA_3544 (.A(net107));
 sg13g2_antennanp ANTENNA_3545 (.A(net107));
 sg13g2_antennanp ANTENNA_3546 (.A(net107));
 sg13g2_antennanp ANTENNA_3547 (.A(net107));
 sg13g2_antennanp ANTENNA_3548 (.A(net107));
 sg13g2_antennanp ANTENNA_3549 (.A(net107));
 sg13g2_antennanp ANTENNA_3550 (.A(net107));
 sg13g2_antennanp ANTENNA_3551 (.A(net113));
 sg13g2_antennanp ANTENNA_3552 (.A(net113));
 sg13g2_antennanp ANTENNA_3553 (.A(net113));
 sg13g2_antennanp ANTENNA_3554 (.A(net113));
 sg13g2_antennanp ANTENNA_3555 (.A(net113));
 sg13g2_antennanp ANTENNA_3556 (.A(net113));
 sg13g2_antennanp ANTENNA_3557 (.A(net113));
 sg13g2_antennanp ANTENNA_3558 (.A(net113));
 sg13g2_antennanp ANTENNA_3559 (.A(net125));
 sg13g2_antennanp ANTENNA_3560 (.A(net125));
 sg13g2_antennanp ANTENNA_3561 (.A(net125));
 sg13g2_antennanp ANTENNA_3562 (.A(net125));
 sg13g2_antennanp ANTENNA_3563 (.A(net125));
 sg13g2_antennanp ANTENNA_3564 (.A(net125));
 sg13g2_antennanp ANTENNA_3565 (.A(net125));
 sg13g2_antennanp ANTENNA_3566 (.A(net125));
 sg13g2_antennanp ANTENNA_3567 (.A(net125));
 sg13g2_antennanp ANTENNA_3568 (.A(net128));
 sg13g2_antennanp ANTENNA_3569 (.A(net128));
 sg13g2_antennanp ANTENNA_3570 (.A(net128));
 sg13g2_antennanp ANTENNA_3571 (.A(net128));
 sg13g2_antennanp ANTENNA_3572 (.A(net128));
 sg13g2_antennanp ANTENNA_3573 (.A(net128));
 sg13g2_antennanp ANTENNA_3574 (.A(net128));
 sg13g2_antennanp ANTENNA_3575 (.A(net128));
 sg13g2_antennanp ANTENNA_3576 (.A(net129));
 sg13g2_antennanp ANTENNA_3577 (.A(net129));
 sg13g2_antennanp ANTENNA_3578 (.A(net129));
 sg13g2_antennanp ANTENNA_3579 (.A(net129));
 sg13g2_antennanp ANTENNA_3580 (.A(net129));
 sg13g2_antennanp ANTENNA_3581 (.A(net129));
 sg13g2_antennanp ANTENNA_3582 (.A(net129));
 sg13g2_antennanp ANTENNA_3583 (.A(net129));
 sg13g2_antennanp ANTENNA_3584 (.A(net129));
 sg13g2_antennanp ANTENNA_3585 (.A(net129));
 sg13g2_antennanp ANTENNA_3586 (.A(net129));
 sg13g2_antennanp ANTENNA_3587 (.A(net129));
 sg13g2_antennanp ANTENNA_3588 (.A(net129));
 sg13g2_antennanp ANTENNA_3589 (.A(net129));
 sg13g2_antennanp ANTENNA_3590 (.A(net129));
 sg13g2_antennanp ANTENNA_3591 (.A(net129));
 sg13g2_antennanp ANTENNA_3592 (.A(net142));
 sg13g2_antennanp ANTENNA_3593 (.A(net142));
 sg13g2_antennanp ANTENNA_3594 (.A(net142));
 sg13g2_antennanp ANTENNA_3595 (.A(net142));
 sg13g2_antennanp ANTENNA_3596 (.A(net142));
 sg13g2_antennanp ANTENNA_3597 (.A(net142));
 sg13g2_antennanp ANTENNA_3598 (.A(net142));
 sg13g2_antennanp ANTENNA_3599 (.A(net142));
 sg13g2_antennanp ANTENNA_3600 (.A(net142));
 sg13g2_antennanp ANTENNA_3601 (.A(net144));
 sg13g2_antennanp ANTENNA_3602 (.A(net144));
 sg13g2_antennanp ANTENNA_3603 (.A(net144));
 sg13g2_antennanp ANTENNA_3604 (.A(net144));
 sg13g2_antennanp ANTENNA_3605 (.A(net144));
 sg13g2_antennanp ANTENNA_3606 (.A(net144));
 sg13g2_antennanp ANTENNA_3607 (.A(net144));
 sg13g2_antennanp ANTENNA_3608 (.A(net144));
 sg13g2_antennanp ANTENNA_3609 (.A(net144));
 sg13g2_antennanp ANTENNA_3610 (.A(net153));
 sg13g2_antennanp ANTENNA_3611 (.A(net153));
 sg13g2_antennanp ANTENNA_3612 (.A(net153));
 sg13g2_antennanp ANTENNA_3613 (.A(net153));
 sg13g2_antennanp ANTENNA_3614 (.A(net153));
 sg13g2_antennanp ANTENNA_3615 (.A(net153));
 sg13g2_antennanp ANTENNA_3616 (.A(net153));
 sg13g2_antennanp ANTENNA_3617 (.A(net153));
 sg13g2_antennanp ANTENNA_3618 (.A(net153));
 sg13g2_antennanp ANTENNA_3619 (.A(net161));
 sg13g2_antennanp ANTENNA_3620 (.A(net161));
 sg13g2_antennanp ANTENNA_3621 (.A(net161));
 sg13g2_antennanp ANTENNA_3622 (.A(net161));
 sg13g2_antennanp ANTENNA_3623 (.A(net161));
 sg13g2_antennanp ANTENNA_3624 (.A(net161));
 sg13g2_antennanp ANTENNA_3625 (.A(net161));
 sg13g2_antennanp ANTENNA_3626 (.A(net161));
 sg13g2_antennanp ANTENNA_3627 (.A(net161));
 sg13g2_antennanp ANTENNA_3628 (.A(net164));
 sg13g2_antennanp ANTENNA_3629 (.A(net164));
 sg13g2_antennanp ANTENNA_3630 (.A(net164));
 sg13g2_antennanp ANTENNA_3631 (.A(net164));
 sg13g2_antennanp ANTENNA_3632 (.A(net164));
 sg13g2_antennanp ANTENNA_3633 (.A(net164));
 sg13g2_antennanp ANTENNA_3634 (.A(net164));
 sg13g2_antennanp ANTENNA_3635 (.A(net164));
 sg13g2_antennanp ANTENNA_3636 (.A(net164));
 sg13g2_antennanp ANTENNA_3637 (.A(net167));
 sg13g2_antennanp ANTENNA_3638 (.A(net167));
 sg13g2_antennanp ANTENNA_3639 (.A(net167));
 sg13g2_antennanp ANTENNA_3640 (.A(net167));
 sg13g2_antennanp ANTENNA_3641 (.A(net167));
 sg13g2_antennanp ANTENNA_3642 (.A(net167));
 sg13g2_antennanp ANTENNA_3643 (.A(net167));
 sg13g2_antennanp ANTENNA_3644 (.A(net167));
 sg13g2_antennanp ANTENNA_3645 (.A(net167));
 sg13g2_antennanp ANTENNA_3646 (.A(net174));
 sg13g2_antennanp ANTENNA_3647 (.A(net174));
 sg13g2_antennanp ANTENNA_3648 (.A(net174));
 sg13g2_antennanp ANTENNA_3649 (.A(net174));
 sg13g2_antennanp ANTENNA_3650 (.A(net174));
 sg13g2_antennanp ANTENNA_3651 (.A(net174));
 sg13g2_antennanp ANTENNA_3652 (.A(net174));
 sg13g2_antennanp ANTENNA_3653 (.A(net174));
 sg13g2_antennanp ANTENNA_3654 (.A(net174));
 sg13g2_antennanp ANTENNA_3655 (.A(net182));
 sg13g2_antennanp ANTENNA_3656 (.A(net182));
 sg13g2_antennanp ANTENNA_3657 (.A(net182));
 sg13g2_antennanp ANTENNA_3658 (.A(net182));
 sg13g2_antennanp ANTENNA_3659 (.A(net182));
 sg13g2_antennanp ANTENNA_3660 (.A(net182));
 sg13g2_antennanp ANTENNA_3661 (.A(net182));
 sg13g2_antennanp ANTENNA_3662 (.A(net182));
 sg13g2_antennanp ANTENNA_3663 (.A(net185));
 sg13g2_antennanp ANTENNA_3664 (.A(net185));
 sg13g2_antennanp ANTENNA_3665 (.A(net185));
 sg13g2_antennanp ANTENNA_3666 (.A(net185));
 sg13g2_antennanp ANTENNA_3667 (.A(net185));
 sg13g2_antennanp ANTENNA_3668 (.A(net185));
 sg13g2_antennanp ANTENNA_3669 (.A(net185));
 sg13g2_antennanp ANTENNA_3670 (.A(net185));
 sg13g2_antennanp ANTENNA_3671 (.A(net185));
 sg13g2_antennanp ANTENNA_3672 (.A(net210));
 sg13g2_antennanp ANTENNA_3673 (.A(net210));
 sg13g2_antennanp ANTENNA_3674 (.A(net210));
 sg13g2_antennanp ANTENNA_3675 (.A(net210));
 sg13g2_antennanp ANTENNA_3676 (.A(net210));
 sg13g2_antennanp ANTENNA_3677 (.A(net210));
 sg13g2_antennanp ANTENNA_3678 (.A(net210));
 sg13g2_antennanp ANTENNA_3679 (.A(net210));
 sg13g2_antennanp ANTENNA_3680 (.A(net210));
 sg13g2_antennanp ANTENNA_3681 (.A(_0003_));
 sg13g2_antennanp ANTENNA_3682 (.A(_0016_));
 sg13g2_antennanp ANTENNA_3683 (.A(_0016_));
 sg13g2_antennanp ANTENNA_3684 (.A(_0018_));
 sg13g2_antennanp ANTENNA_3685 (.A(_0018_));
 sg13g2_antennanp ANTENNA_3686 (.A(_0021_));
 sg13g2_antennanp ANTENNA_3687 (.A(_0022_));
 sg13g2_antennanp ANTENNA_3688 (.A(_0023_));
 sg13g2_antennanp ANTENNA_3689 (.A(_0024_));
 sg13g2_antennanp ANTENNA_3690 (.A(_0025_));
 sg13g2_antennanp ANTENNA_3691 (.A(_0025_));
 sg13g2_antennanp ANTENNA_3692 (.A(_0027_));
 sg13g2_antennanp ANTENNA_3693 (.A(_0027_));
 sg13g2_antennanp ANTENNA_3694 (.A(_0028_));
 sg13g2_antennanp ANTENNA_3695 (.A(_0028_));
 sg13g2_antennanp ANTENNA_3696 (.A(_0038_));
 sg13g2_antennanp ANTENNA_3697 (.A(_0038_));
 sg13g2_antennanp ANTENNA_3698 (.A(_0038_));
 sg13g2_antennanp ANTENNA_3699 (.A(_0038_));
 sg13g2_antennanp ANTENNA_3700 (.A(_0038_));
 sg13g2_antennanp ANTENNA_3701 (.A(_0038_));
 sg13g2_antennanp ANTENNA_3702 (.A(_0038_));
 sg13g2_antennanp ANTENNA_3703 (.A(_0038_));
 sg13g2_antennanp ANTENNA_3704 (.A(_0038_));
 sg13g2_antennanp ANTENNA_3705 (.A(_0123_));
 sg13g2_antennanp ANTENNA_3706 (.A(_0123_));
 sg13g2_antennanp ANTENNA_3707 (.A(_0125_));
 sg13g2_antennanp ANTENNA_3708 (.A(_0125_));
 sg13g2_antennanp ANTENNA_3709 (.A(_0125_));
 sg13g2_antennanp ANTENNA_3710 (.A(_0150_));
 sg13g2_antennanp ANTENNA_3711 (.A(_0150_));
 sg13g2_antennanp ANTENNA_3712 (.A(_0150_));
 sg13g2_antennanp ANTENNA_3713 (.A(_0150_));
 sg13g2_antennanp ANTENNA_3714 (.A(_0150_));
 sg13g2_antennanp ANTENNA_3715 (.A(_0150_));
 sg13g2_antennanp ANTENNA_3716 (.A(_0150_));
 sg13g2_antennanp ANTENNA_3717 (.A(_0150_));
 sg13g2_antennanp ANTENNA_3718 (.A(_0150_));
 sg13g2_antennanp ANTENNA_3719 (.A(_0150_));
 sg13g2_antennanp ANTENNA_3720 (.A(_0158_));
 sg13g2_antennanp ANTENNA_3721 (.A(_0165_));
 sg13g2_antennanp ANTENNA_3722 (.A(_0165_));
 sg13g2_antennanp ANTENNA_3723 (.A(_0165_));
 sg13g2_antennanp ANTENNA_3724 (.A(_0165_));
 sg13g2_antennanp ANTENNA_3725 (.A(_0167_));
 sg13g2_antennanp ANTENNA_3726 (.A(_0167_));
 sg13g2_antennanp ANTENNA_3727 (.A(_0167_));
 sg13g2_antennanp ANTENNA_3728 (.A(_0167_));
 sg13g2_antennanp ANTENNA_3729 (.A(_0167_));
 sg13g2_antennanp ANTENNA_3730 (.A(_0167_));
 sg13g2_antennanp ANTENNA_3731 (.A(_0167_));
 sg13g2_antennanp ANTENNA_3732 (.A(_0167_));
 sg13g2_antennanp ANTENNA_3733 (.A(_0168_));
 sg13g2_antennanp ANTENNA_3734 (.A(_0168_));
 sg13g2_antennanp ANTENNA_3735 (.A(_0168_));
 sg13g2_antennanp ANTENNA_3736 (.A(_0168_));
 sg13g2_antennanp ANTENNA_3737 (.A(_0168_));
 sg13g2_antennanp ANTENNA_3738 (.A(_0168_));
 sg13g2_antennanp ANTENNA_3739 (.A(_0189_));
 sg13g2_antennanp ANTENNA_3740 (.A(_0230_));
 sg13g2_antennanp ANTENNA_3741 (.A(_0260_));
 sg13g2_antennanp ANTENNA_3742 (.A(_0260_));
 sg13g2_antennanp ANTENNA_3743 (.A(_0260_));
 sg13g2_antennanp ANTENNA_3744 (.A(_0260_));
 sg13g2_antennanp ANTENNA_3745 (.A(_0269_));
 sg13g2_antennanp ANTENNA_3746 (.A(_0301_));
 sg13g2_antennanp ANTENNA_3747 (.A(_0345_));
 sg13g2_antennanp ANTENNA_3748 (.A(_0345_));
 sg13g2_antennanp ANTENNA_3749 (.A(_0345_));
 sg13g2_antennanp ANTENNA_3750 (.A(_0345_));
 sg13g2_antennanp ANTENNA_3751 (.A(_0346_));
 sg13g2_antennanp ANTENNA_3752 (.A(_0346_));
 sg13g2_antennanp ANTENNA_3753 (.A(_0346_));
 sg13g2_antennanp ANTENNA_3754 (.A(_0346_));
 sg13g2_antennanp ANTENNA_3755 (.A(_0346_));
 sg13g2_antennanp ANTENNA_3756 (.A(_0346_));
 sg13g2_antennanp ANTENNA_3757 (.A(_0346_));
 sg13g2_antennanp ANTENNA_3758 (.A(_0346_));
 sg13g2_antennanp ANTENNA_3759 (.A(_0360_));
 sg13g2_antennanp ANTENNA_3760 (.A(_0360_));
 sg13g2_antennanp ANTENNA_3761 (.A(_0360_));
 sg13g2_antennanp ANTENNA_3762 (.A(_0360_));
 sg13g2_antennanp ANTENNA_3763 (.A(_0360_));
 sg13g2_antennanp ANTENNA_3764 (.A(_0387_));
 sg13g2_antennanp ANTENNA_3765 (.A(_0387_));
 sg13g2_antennanp ANTENNA_3766 (.A(_0387_));
 sg13g2_antennanp ANTENNA_3767 (.A(_0387_));
 sg13g2_antennanp ANTENNA_3768 (.A(_0387_));
 sg13g2_antennanp ANTENNA_3769 (.A(_0387_));
 sg13g2_antennanp ANTENNA_3770 (.A(_0435_));
 sg13g2_antennanp ANTENNA_3771 (.A(_0435_));
 sg13g2_antennanp ANTENNA_3772 (.A(_0448_));
 sg13g2_antennanp ANTENNA_3773 (.A(_0490_));
 sg13g2_antennanp ANTENNA_3774 (.A(_0490_));
 sg13g2_antennanp ANTENNA_3775 (.A(_0507_));
 sg13g2_antennanp ANTENNA_3776 (.A(_0507_));
 sg13g2_antennanp ANTENNA_3777 (.A(_0511_));
 sg13g2_antennanp ANTENNA_3778 (.A(_0511_));
 sg13g2_antennanp ANTENNA_3779 (.A(_0511_));
 sg13g2_antennanp ANTENNA_3780 (.A(_0521_));
 sg13g2_antennanp ANTENNA_3781 (.A(_0521_));
 sg13g2_antennanp ANTENNA_3782 (.A(_0521_));
 sg13g2_antennanp ANTENNA_3783 (.A(_0597_));
 sg13g2_antennanp ANTENNA_3784 (.A(_0597_));
 sg13g2_antennanp ANTENNA_3785 (.A(_0597_));
 sg13g2_antennanp ANTENNA_3786 (.A(_0597_));
 sg13g2_antennanp ANTENNA_3787 (.A(_0598_));
 sg13g2_antennanp ANTENNA_3788 (.A(_0598_));
 sg13g2_antennanp ANTENNA_3789 (.A(_0598_));
 sg13g2_antennanp ANTENNA_3790 (.A(_0598_));
 sg13g2_antennanp ANTENNA_3791 (.A(_0598_));
 sg13g2_antennanp ANTENNA_3792 (.A(_0623_));
 sg13g2_antennanp ANTENNA_3793 (.A(_0780_));
 sg13g2_antennanp ANTENNA_3794 (.A(_0800_));
 sg13g2_antennanp ANTENNA_3795 (.A(_0866_));
 sg13g2_antennanp ANTENNA_3796 (.A(_0866_));
 sg13g2_antennanp ANTENNA_3797 (.A(_0866_));
 sg13g2_antennanp ANTENNA_3798 (.A(_0878_));
 sg13g2_antennanp ANTENNA_3799 (.A(_0878_));
 sg13g2_antennanp ANTENNA_3800 (.A(_0878_));
 sg13g2_antennanp ANTENNA_3801 (.A(_0878_));
 sg13g2_antennanp ANTENNA_3802 (.A(_0878_));
 sg13g2_antennanp ANTENNA_3803 (.A(_0878_));
 sg13g2_antennanp ANTENNA_3804 (.A(_0878_));
 sg13g2_antennanp ANTENNA_3805 (.A(_0878_));
 sg13g2_antennanp ANTENNA_3806 (.A(_0878_));
 sg13g2_antennanp ANTENNA_3807 (.A(_1002_));
 sg13g2_antennanp ANTENNA_3808 (.A(_1002_));
 sg13g2_antennanp ANTENNA_3809 (.A(_1071_));
 sg13g2_antennanp ANTENNA_3810 (.A(_1071_));
 sg13g2_antennanp ANTENNA_3811 (.A(_1071_));
 sg13g2_antennanp ANTENNA_3812 (.A(_1085_));
 sg13g2_antennanp ANTENNA_3813 (.A(_1085_));
 sg13g2_antennanp ANTENNA_3814 (.A(_1085_));
 sg13g2_antennanp ANTENNA_3815 (.A(_1085_));
 sg13g2_antennanp ANTENNA_3816 (.A(_1085_));
 sg13g2_antennanp ANTENNA_3817 (.A(_1085_));
 sg13g2_antennanp ANTENNA_3818 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3819 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3820 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3821 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3822 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3823 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3824 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3825 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3826 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3827 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3828 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3829 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3830 (.A(_1162_));
 sg13g2_antennanp ANTENNA_3831 (.A(_1225_));
 sg13g2_antennanp ANTENNA_3832 (.A(_1225_));
 sg13g2_antennanp ANTENNA_3833 (.A(_1292_));
 sg13g2_antennanp ANTENNA_3834 (.A(_1292_));
 sg13g2_antennanp ANTENNA_3835 (.A(_1326_));
 sg13g2_antennanp ANTENNA_3836 (.A(_1326_));
 sg13g2_antennanp ANTENNA_3837 (.A(_1326_));
 sg13g2_antennanp ANTENNA_3838 (.A(_1326_));
 sg13g2_antennanp ANTENNA_3839 (.A(_1326_));
 sg13g2_antennanp ANTENNA_3840 (.A(_1326_));
 sg13g2_antennanp ANTENNA_3841 (.A(_1326_));
 sg13g2_antennanp ANTENNA_3842 (.A(_1326_));
 sg13g2_antennanp ANTENNA_3843 (.A(_1326_));
 sg13g2_antennanp ANTENNA_3844 (.A(_1363_));
 sg13g2_antennanp ANTENNA_3845 (.A(_1411_));
 sg13g2_antennanp ANTENNA_3846 (.A(_1439_));
 sg13g2_antennanp ANTENNA_3847 (.A(_1470_));
 sg13g2_antennanp ANTENNA_3848 (.A(_1470_));
 sg13g2_antennanp ANTENNA_3849 (.A(_1519_));
 sg13g2_antennanp ANTENNA_3850 (.A(_1531_));
 sg13g2_antennanp ANTENNA_3851 (.A(_1531_));
 sg13g2_antennanp ANTENNA_3852 (.A(_1532_));
 sg13g2_antennanp ANTENNA_3853 (.A(_1532_));
 sg13g2_antennanp ANTENNA_3854 (.A(_1532_));
 sg13g2_antennanp ANTENNA_3855 (.A(_1544_));
 sg13g2_antennanp ANTENNA_3856 (.A(_1544_));
 sg13g2_antennanp ANTENNA_3857 (.A(_1544_));
 sg13g2_antennanp ANTENNA_3858 (.A(_1544_));
 sg13g2_antennanp ANTENNA_3859 (.A(_1544_));
 sg13g2_antennanp ANTENNA_3860 (.A(_1553_));
 sg13g2_antennanp ANTENNA_3861 (.A(_1631_));
 sg13g2_antennanp ANTENNA_3862 (.A(_1631_));
 sg13g2_antennanp ANTENNA_3863 (.A(_1631_));
 sg13g2_antennanp ANTENNA_3864 (.A(_1685_));
 sg13g2_antennanp ANTENNA_3865 (.A(_1685_));
 sg13g2_antennanp ANTENNA_3866 (.A(_1685_));
 sg13g2_antennanp ANTENNA_3867 (.A(_1685_));
 sg13g2_antennanp ANTENNA_3868 (.A(_1696_));
 sg13g2_antennanp ANTENNA_3869 (.A(_1696_));
 sg13g2_antennanp ANTENNA_3870 (.A(_1696_));
 sg13g2_antennanp ANTENNA_3871 (.A(_1696_));
 sg13g2_antennanp ANTENNA_3872 (.A(_1696_));
 sg13g2_antennanp ANTENNA_3873 (.A(_1696_));
 sg13g2_antennanp ANTENNA_3874 (.A(_1696_));
 sg13g2_antennanp ANTENNA_3875 (.A(_1696_));
 sg13g2_antennanp ANTENNA_3876 (.A(_1696_));
 sg13g2_antennanp ANTENNA_3877 (.A(_1696_));
 sg13g2_antennanp ANTENNA_3878 (.A(_1707_));
 sg13g2_antennanp ANTENNA_3879 (.A(_1707_));
 sg13g2_antennanp ANTENNA_3880 (.A(_1707_));
 sg13g2_antennanp ANTENNA_3881 (.A(_1707_));
 sg13g2_antennanp ANTENNA_3882 (.A(_1707_));
 sg13g2_antennanp ANTENNA_3883 (.A(_1707_));
 sg13g2_antennanp ANTENNA_3884 (.A(_1707_));
 sg13g2_antennanp ANTENNA_3885 (.A(_1707_));
 sg13g2_antennanp ANTENNA_3886 (.A(_1716_));
 sg13g2_antennanp ANTENNA_3887 (.A(_1735_));
 sg13g2_antennanp ANTENNA_3888 (.A(_1761_));
 sg13g2_antennanp ANTENNA_3889 (.A(_2014_));
 sg13g2_antennanp ANTENNA_3890 (.A(_2014_));
 sg13g2_antennanp ANTENNA_3891 (.A(_2020_));
 sg13g2_antennanp ANTENNA_3892 (.A(_2020_));
 sg13g2_antennanp ANTENNA_3893 (.A(_2020_));
 sg13g2_antennanp ANTENNA_3894 (.A(_2020_));
 sg13g2_antennanp ANTENNA_3895 (.A(_2020_));
 sg13g2_antennanp ANTENNA_3896 (.A(_2020_));
 sg13g2_antennanp ANTENNA_3897 (.A(_2020_));
 sg13g2_antennanp ANTENNA_3898 (.A(_2020_));
 sg13g2_antennanp ANTENNA_3899 (.A(_2020_));
 sg13g2_antennanp ANTENNA_3900 (.A(_2020_));
 sg13g2_antennanp ANTENNA_3901 (.A(_2020_));
 sg13g2_antennanp ANTENNA_3902 (.A(_2020_));
 sg13g2_antennanp ANTENNA_3903 (.A(_2020_));
 sg13g2_antennanp ANTENNA_3904 (.A(_2037_));
 sg13g2_antennanp ANTENNA_3905 (.A(_2053_));
 sg13g2_antennanp ANTENNA_3906 (.A(_2053_));
 sg13g2_antennanp ANTENNA_3907 (.A(_2053_));
 sg13g2_antennanp ANTENNA_3908 (.A(_2097_));
 sg13g2_antennanp ANTENNA_3909 (.A(_2097_));
 sg13g2_antennanp ANTENNA_3910 (.A(_2097_));
 sg13g2_antennanp ANTENNA_3911 (.A(_2097_));
 sg13g2_antennanp ANTENNA_3912 (.A(_2097_));
 sg13g2_antennanp ANTENNA_3913 (.A(_2110_));
 sg13g2_antennanp ANTENNA_3914 (.A(_2110_));
 sg13g2_antennanp ANTENNA_3915 (.A(_2112_));
 sg13g2_antennanp ANTENNA_3916 (.A(_2145_));
 sg13g2_antennanp ANTENNA_3917 (.A(_2171_));
 sg13g2_antennanp ANTENNA_3918 (.A(_2171_));
 sg13g2_antennanp ANTENNA_3919 (.A(_2171_));
 sg13g2_antennanp ANTENNA_3920 (.A(_2171_));
 sg13g2_antennanp ANTENNA_3921 (.A(_2171_));
 sg13g2_antennanp ANTENNA_3922 (.A(_2171_));
 sg13g2_antennanp ANTENNA_3923 (.A(_2171_));
 sg13g2_antennanp ANTENNA_3924 (.A(_2171_));
 sg13g2_antennanp ANTENNA_3925 (.A(_2171_));
 sg13g2_antennanp ANTENNA_3926 (.A(_2172_));
 sg13g2_antennanp ANTENNA_3927 (.A(_2172_));
 sg13g2_antennanp ANTENNA_3928 (.A(_2172_));
 sg13g2_antennanp ANTENNA_3929 (.A(_2172_));
 sg13g2_antennanp ANTENNA_3930 (.A(_2172_));
 sg13g2_antennanp ANTENNA_3931 (.A(_2172_));
 sg13g2_antennanp ANTENNA_3932 (.A(_2172_));
 sg13g2_antennanp ANTENNA_3933 (.A(_2172_));
 sg13g2_antennanp ANTENNA_3934 (.A(_2172_));
 sg13g2_antennanp ANTENNA_3935 (.A(_2172_));
 sg13g2_antennanp ANTENNA_3936 (.A(_2257_));
 sg13g2_antennanp ANTENNA_3937 (.A(_2257_));
 sg13g2_antennanp ANTENNA_3938 (.A(_2430_));
 sg13g2_antennanp ANTENNA_3939 (.A(_2430_));
 sg13g2_antennanp ANTENNA_3940 (.A(_2430_));
 sg13g2_antennanp ANTENNA_3941 (.A(_2430_));
 sg13g2_antennanp ANTENNA_3942 (.A(_2430_));
 sg13g2_antennanp ANTENNA_3943 (.A(_2430_));
 sg13g2_antennanp ANTENNA_3944 (.A(_2467_));
 sg13g2_antennanp ANTENNA_3945 (.A(_2467_));
 sg13g2_antennanp ANTENNA_3946 (.A(_2467_));
 sg13g2_antennanp ANTENNA_3947 (.A(_2467_));
 sg13g2_antennanp ANTENNA_3948 (.A(_2467_));
 sg13g2_antennanp ANTENNA_3949 (.A(_2470_));
 sg13g2_antennanp ANTENNA_3950 (.A(_2470_));
 sg13g2_antennanp ANTENNA_3951 (.A(_2470_));
 sg13g2_antennanp ANTENNA_3952 (.A(_2470_));
 sg13g2_antennanp ANTENNA_3953 (.A(_2480_));
 sg13g2_antennanp ANTENNA_3954 (.A(_2480_));
 sg13g2_antennanp ANTENNA_3955 (.A(_2480_));
 sg13g2_antennanp ANTENNA_3956 (.A(_2480_));
 sg13g2_antennanp ANTENNA_3957 (.A(_2480_));
 sg13g2_antennanp ANTENNA_3958 (.A(_2480_));
 sg13g2_antennanp ANTENNA_3959 (.A(_2480_));
 sg13g2_antennanp ANTENNA_3960 (.A(_2480_));
 sg13g2_antennanp ANTENNA_3961 (.A(_2482_));
 sg13g2_antennanp ANTENNA_3962 (.A(_2482_));
 sg13g2_antennanp ANTENNA_3963 (.A(_2482_));
 sg13g2_antennanp ANTENNA_3964 (.A(_2482_));
 sg13g2_antennanp ANTENNA_3965 (.A(_2482_));
 sg13g2_antennanp ANTENNA_3966 (.A(_2482_));
 sg13g2_antennanp ANTENNA_3967 (.A(_2482_));
 sg13g2_antennanp ANTENNA_3968 (.A(_2482_));
 sg13g2_antennanp ANTENNA_3969 (.A(_2487_));
 sg13g2_antennanp ANTENNA_3970 (.A(_2487_));
 sg13g2_antennanp ANTENNA_3971 (.A(_2501_));
 sg13g2_antennanp ANTENNA_3972 (.A(_2501_));
 sg13g2_antennanp ANTENNA_3973 (.A(_2501_));
 sg13g2_antennanp ANTENNA_3974 (.A(_2501_));
 sg13g2_antennanp ANTENNA_3975 (.A(_2520_));
 sg13g2_antennanp ANTENNA_3976 (.A(_2520_));
 sg13g2_antennanp ANTENNA_3977 (.A(_2520_));
 sg13g2_antennanp ANTENNA_3978 (.A(_2520_));
 sg13g2_antennanp ANTENNA_3979 (.A(_2520_));
 sg13g2_antennanp ANTENNA_3980 (.A(_2520_));
 sg13g2_antennanp ANTENNA_3981 (.A(_2530_));
 sg13g2_antennanp ANTENNA_3982 (.A(_2530_));
 sg13g2_antennanp ANTENNA_3983 (.A(_2530_));
 sg13g2_antennanp ANTENNA_3984 (.A(_2530_));
 sg13g2_antennanp ANTENNA_3985 (.A(_2537_));
 sg13g2_antennanp ANTENNA_3986 (.A(_2537_));
 sg13g2_antennanp ANTENNA_3987 (.A(_2537_));
 sg13g2_antennanp ANTENNA_3988 (.A(_2537_));
 sg13g2_antennanp ANTENNA_3989 (.A(_2573_));
 sg13g2_antennanp ANTENNA_3990 (.A(_2573_));
 sg13g2_antennanp ANTENNA_3991 (.A(_2573_));
 sg13g2_antennanp ANTENNA_3992 (.A(_2573_));
 sg13g2_antennanp ANTENNA_3993 (.A(_2577_));
 sg13g2_antennanp ANTENNA_3994 (.A(_2577_));
 sg13g2_antennanp ANTENNA_3995 (.A(_2577_));
 sg13g2_antennanp ANTENNA_3996 (.A(_2577_));
 sg13g2_antennanp ANTENNA_3997 (.A(_2577_));
 sg13g2_antennanp ANTENNA_3998 (.A(_2577_));
 sg13g2_antennanp ANTENNA_3999 (.A(_2577_));
 sg13g2_antennanp ANTENNA_4000 (.A(_2577_));
 sg13g2_antennanp ANTENNA_4001 (.A(_2585_));
 sg13g2_antennanp ANTENNA_4002 (.A(_2585_));
 sg13g2_antennanp ANTENNA_4003 (.A(_2585_));
 sg13g2_antennanp ANTENNA_4004 (.A(_2585_));
 sg13g2_antennanp ANTENNA_4005 (.A(_2588_));
 sg13g2_antennanp ANTENNA_4006 (.A(_2600_));
 sg13g2_antennanp ANTENNA_4007 (.A(_2600_));
 sg13g2_antennanp ANTENNA_4008 (.A(_2600_));
 sg13g2_antennanp ANTENNA_4009 (.A(_2600_));
 sg13g2_antennanp ANTENNA_4010 (.A(_2607_));
 sg13g2_antennanp ANTENNA_4011 (.A(_2607_));
 sg13g2_antennanp ANTENNA_4012 (.A(_2615_));
 sg13g2_antennanp ANTENNA_4013 (.A(_2615_));
 sg13g2_antennanp ANTENNA_4014 (.A(_2615_));
 sg13g2_antennanp ANTENNA_4015 (.A(_2622_));
 sg13g2_antennanp ANTENNA_4016 (.A(_2622_));
 sg13g2_antennanp ANTENNA_4017 (.A(_2622_));
 sg13g2_antennanp ANTENNA_4018 (.A(_2622_));
 sg13g2_antennanp ANTENNA_4019 (.A(_2622_));
 sg13g2_antennanp ANTENNA_4020 (.A(_2622_));
 sg13g2_antennanp ANTENNA_4021 (.A(_2625_));
 sg13g2_antennanp ANTENNA_4022 (.A(_2625_));
 sg13g2_antennanp ANTENNA_4023 (.A(_2625_));
 sg13g2_antennanp ANTENNA_4024 (.A(_2625_));
 sg13g2_antennanp ANTENNA_4025 (.A(_2625_));
 sg13g2_antennanp ANTENNA_4026 (.A(_2659_));
 sg13g2_antennanp ANTENNA_4027 (.A(_2659_));
 sg13g2_antennanp ANTENNA_4028 (.A(_2659_));
 sg13g2_antennanp ANTENNA_4029 (.A(_2659_));
 sg13g2_antennanp ANTENNA_4030 (.A(_2659_));
 sg13g2_antennanp ANTENNA_4031 (.A(_2665_));
 sg13g2_antennanp ANTENNA_4032 (.A(_2665_));
 sg13g2_antennanp ANTENNA_4033 (.A(_2665_));
 sg13g2_antennanp ANTENNA_4034 (.A(_2665_));
 sg13g2_antennanp ANTENNA_4035 (.A(_2678_));
 sg13g2_antennanp ANTENNA_4036 (.A(_2678_));
 sg13g2_antennanp ANTENNA_4037 (.A(_2678_));
 sg13g2_antennanp ANTENNA_4038 (.A(_2678_));
 sg13g2_antennanp ANTENNA_4039 (.A(_2678_));
 sg13g2_antennanp ANTENNA_4040 (.A(_2678_));
 sg13g2_antennanp ANTENNA_4041 (.A(_2732_));
 sg13g2_antennanp ANTENNA_4042 (.A(_2732_));
 sg13g2_antennanp ANTENNA_4043 (.A(_2732_));
 sg13g2_antennanp ANTENNA_4044 (.A(_2733_));
 sg13g2_antennanp ANTENNA_4045 (.A(_2733_));
 sg13g2_antennanp ANTENNA_4046 (.A(_2733_));
 sg13g2_antennanp ANTENNA_4047 (.A(_2733_));
 sg13g2_antennanp ANTENNA_4048 (.A(_2739_));
 sg13g2_antennanp ANTENNA_4049 (.A(_2739_));
 sg13g2_antennanp ANTENNA_4050 (.A(_2739_));
 sg13g2_antennanp ANTENNA_4051 (.A(_2739_));
 sg13g2_antennanp ANTENNA_4052 (.A(_2739_));
 sg13g2_antennanp ANTENNA_4053 (.A(_2769_));
 sg13g2_antennanp ANTENNA_4054 (.A(_2769_));
 sg13g2_antennanp ANTENNA_4055 (.A(_2769_));
 sg13g2_antennanp ANTENNA_4056 (.A(_2769_));
 sg13g2_antennanp ANTENNA_4057 (.A(_2789_));
 sg13g2_antennanp ANTENNA_4058 (.A(_2789_));
 sg13g2_antennanp ANTENNA_4059 (.A(_2789_));
 sg13g2_antennanp ANTENNA_4060 (.A(_2789_));
 sg13g2_antennanp ANTENNA_4061 (.A(_2805_));
 sg13g2_antennanp ANTENNA_4062 (.A(_2805_));
 sg13g2_antennanp ANTENNA_4063 (.A(_2808_));
 sg13g2_antennanp ANTENNA_4064 (.A(_2808_));
 sg13g2_antennanp ANTENNA_4065 (.A(_2808_));
 sg13g2_antennanp ANTENNA_4066 (.A(_2808_));
 sg13g2_antennanp ANTENNA_4067 (.A(_2816_));
 sg13g2_antennanp ANTENNA_4068 (.A(_2816_));
 sg13g2_antennanp ANTENNA_4069 (.A(_2816_));
 sg13g2_antennanp ANTENNA_4070 (.A(_2816_));
 sg13g2_antennanp ANTENNA_4071 (.A(_2826_));
 sg13g2_antennanp ANTENNA_4072 (.A(_2826_));
 sg13g2_antennanp ANTENNA_4073 (.A(_2826_));
 sg13g2_antennanp ANTENNA_4074 (.A(_2826_));
 sg13g2_antennanp ANTENNA_4075 (.A(_2858_));
 sg13g2_antennanp ANTENNA_4076 (.A(_2858_));
 sg13g2_antennanp ANTENNA_4077 (.A(_2879_));
 sg13g2_antennanp ANTENNA_4078 (.A(_2879_));
 sg13g2_antennanp ANTENNA_4079 (.A(_2879_));
 sg13g2_antennanp ANTENNA_4080 (.A(_2879_));
 sg13g2_antennanp ANTENNA_4081 (.A(_2879_));
 sg13g2_antennanp ANTENNA_4082 (.A(_2879_));
 sg13g2_antennanp ANTENNA_4083 (.A(_2879_));
 sg13g2_antennanp ANTENNA_4084 (.A(_2879_));
 sg13g2_antennanp ANTENNA_4085 (.A(_2914_));
 sg13g2_antennanp ANTENNA_4086 (.A(_2931_));
 sg13g2_antennanp ANTENNA_4087 (.A(_2931_));
 sg13g2_antennanp ANTENNA_4088 (.A(_2931_));
 sg13g2_antennanp ANTENNA_4089 (.A(_2936_));
 sg13g2_antennanp ANTENNA_4090 (.A(_2936_));
 sg13g2_antennanp ANTENNA_4091 (.A(_2936_));
 sg13g2_antennanp ANTENNA_4092 (.A(_2970_));
 sg13g2_antennanp ANTENNA_4093 (.A(_2970_));
 sg13g2_antennanp ANTENNA_4094 (.A(_2970_));
 sg13g2_antennanp ANTENNA_4095 (.A(_2970_));
 sg13g2_antennanp ANTENNA_4096 (.A(_2974_));
 sg13g2_antennanp ANTENNA_4097 (.A(_2974_));
 sg13g2_antennanp ANTENNA_4098 (.A(_2986_));
 sg13g2_antennanp ANTENNA_4099 (.A(_2986_));
 sg13g2_antennanp ANTENNA_4100 (.A(_2986_));
 sg13g2_antennanp ANTENNA_4101 (.A(_2986_));
 sg13g2_antennanp ANTENNA_4102 (.A(_3018_));
 sg13g2_antennanp ANTENNA_4103 (.A(_3018_));
 sg13g2_antennanp ANTENNA_4104 (.A(_3018_));
 sg13g2_antennanp ANTENNA_4105 (.A(clk));
 sg13g2_antennanp ANTENNA_4106 (.A(clk));
 sg13g2_antennanp ANTENNA_4107 (.A(net22));
 sg13g2_antennanp ANTENNA_4108 (.A(net22));
 sg13g2_antennanp ANTENNA_4109 (.A(net22));
 sg13g2_antennanp ANTENNA_4110 (.A(net22));
 sg13g2_antennanp ANTENNA_4111 (.A(net22));
 sg13g2_antennanp ANTENNA_4112 (.A(net22));
 sg13g2_antennanp ANTENNA_4113 (.A(net22));
 sg13g2_antennanp ANTENNA_4114 (.A(net22));
 sg13g2_antennanp ANTENNA_4115 (.A(net22));
 sg13g2_antennanp ANTENNA_4116 (.A(net23));
 sg13g2_antennanp ANTENNA_4117 (.A(net23));
 sg13g2_antennanp ANTENNA_4118 (.A(net23));
 sg13g2_antennanp ANTENNA_4119 (.A(net23));
 sg13g2_antennanp ANTENNA_4120 (.A(net23));
 sg13g2_antennanp ANTENNA_4121 (.A(net23));
 sg13g2_antennanp ANTENNA_4122 (.A(net23));
 sg13g2_antennanp ANTENNA_4123 (.A(net23));
 sg13g2_antennanp ANTENNA_4124 (.A(net29));
 sg13g2_antennanp ANTENNA_4125 (.A(net29));
 sg13g2_antennanp ANTENNA_4126 (.A(net29));
 sg13g2_antennanp ANTENNA_4127 (.A(net29));
 sg13g2_antennanp ANTENNA_4128 (.A(net29));
 sg13g2_antennanp ANTENNA_4129 (.A(net29));
 sg13g2_antennanp ANTENNA_4130 (.A(net29));
 sg13g2_antennanp ANTENNA_4131 (.A(net29));
 sg13g2_antennanp ANTENNA_4132 (.A(net29));
 sg13g2_antennanp ANTENNA_4133 (.A(net35));
 sg13g2_antennanp ANTENNA_4134 (.A(net35));
 sg13g2_antennanp ANTENNA_4135 (.A(net35));
 sg13g2_antennanp ANTENNA_4136 (.A(net35));
 sg13g2_antennanp ANTENNA_4137 (.A(net35));
 sg13g2_antennanp ANTENNA_4138 (.A(net35));
 sg13g2_antennanp ANTENNA_4139 (.A(net35));
 sg13g2_antennanp ANTENNA_4140 (.A(net35));
 sg13g2_antennanp ANTENNA_4141 (.A(net35));
 sg13g2_antennanp ANTENNA_4142 (.A(net46));
 sg13g2_antennanp ANTENNA_4143 (.A(net46));
 sg13g2_antennanp ANTENNA_4144 (.A(net46));
 sg13g2_antennanp ANTENNA_4145 (.A(net46));
 sg13g2_antennanp ANTENNA_4146 (.A(net46));
 sg13g2_antennanp ANTENNA_4147 (.A(net46));
 sg13g2_antennanp ANTENNA_4148 (.A(net46));
 sg13g2_antennanp ANTENNA_4149 (.A(net46));
 sg13g2_antennanp ANTENNA_4150 (.A(net53));
 sg13g2_antennanp ANTENNA_4151 (.A(net53));
 sg13g2_antennanp ANTENNA_4152 (.A(net53));
 sg13g2_antennanp ANTENNA_4153 (.A(net53));
 sg13g2_antennanp ANTENNA_4154 (.A(net53));
 sg13g2_antennanp ANTENNA_4155 (.A(net53));
 sg13g2_antennanp ANTENNA_4156 (.A(net53));
 sg13g2_antennanp ANTENNA_4157 (.A(net53));
 sg13g2_antennanp ANTENNA_4158 (.A(net59));
 sg13g2_antennanp ANTENNA_4159 (.A(net59));
 sg13g2_antennanp ANTENNA_4160 (.A(net59));
 sg13g2_antennanp ANTENNA_4161 (.A(net59));
 sg13g2_antennanp ANTENNA_4162 (.A(net59));
 sg13g2_antennanp ANTENNA_4163 (.A(net59));
 sg13g2_antennanp ANTENNA_4164 (.A(net59));
 sg13g2_antennanp ANTENNA_4165 (.A(net59));
 sg13g2_antennanp ANTENNA_4166 (.A(net59));
 sg13g2_antennanp ANTENNA_4167 (.A(net59));
 sg13g2_antennanp ANTENNA_4168 (.A(net59));
 sg13g2_antennanp ANTENNA_4169 (.A(net59));
 sg13g2_antennanp ANTENNA_4170 (.A(net59));
 sg13g2_antennanp ANTENNA_4171 (.A(net59));
 sg13g2_antennanp ANTENNA_4172 (.A(net59));
 sg13g2_antennanp ANTENNA_4173 (.A(net61));
 sg13g2_antennanp ANTENNA_4174 (.A(net61));
 sg13g2_antennanp ANTENNA_4175 (.A(net61));
 sg13g2_antennanp ANTENNA_4176 (.A(net61));
 sg13g2_antennanp ANTENNA_4177 (.A(net61));
 sg13g2_antennanp ANTENNA_4178 (.A(net61));
 sg13g2_antennanp ANTENNA_4179 (.A(net61));
 sg13g2_antennanp ANTENNA_4180 (.A(net61));
 sg13g2_antennanp ANTENNA_4181 (.A(net61));
 sg13g2_antennanp ANTENNA_4182 (.A(net70));
 sg13g2_antennanp ANTENNA_4183 (.A(net70));
 sg13g2_antennanp ANTENNA_4184 (.A(net70));
 sg13g2_antennanp ANTENNA_4185 (.A(net70));
 sg13g2_antennanp ANTENNA_4186 (.A(net70));
 sg13g2_antennanp ANTENNA_4187 (.A(net70));
 sg13g2_antennanp ANTENNA_4188 (.A(net70));
 sg13g2_antennanp ANTENNA_4189 (.A(net70));
 sg13g2_antennanp ANTENNA_4190 (.A(net71));
 sg13g2_antennanp ANTENNA_4191 (.A(net71));
 sg13g2_antennanp ANTENNA_4192 (.A(net71));
 sg13g2_antennanp ANTENNA_4193 (.A(net71));
 sg13g2_antennanp ANTENNA_4194 (.A(net71));
 sg13g2_antennanp ANTENNA_4195 (.A(net71));
 sg13g2_antennanp ANTENNA_4196 (.A(net71));
 sg13g2_antennanp ANTENNA_4197 (.A(net71));
 sg13g2_antennanp ANTENNA_4198 (.A(net71));
 sg13g2_antennanp ANTENNA_4199 (.A(net71));
 sg13g2_antennanp ANTENNA_4200 (.A(net71));
 sg13g2_antennanp ANTENNA_4201 (.A(net71));
 sg13g2_antennanp ANTENNA_4202 (.A(net71));
 sg13g2_antennanp ANTENNA_4203 (.A(net71));
 sg13g2_antennanp ANTENNA_4204 (.A(net71));
 sg13g2_antennanp ANTENNA_4205 (.A(net71));
 sg13g2_antennanp ANTENNA_4206 (.A(net76));
 sg13g2_antennanp ANTENNA_4207 (.A(net76));
 sg13g2_antennanp ANTENNA_4208 (.A(net76));
 sg13g2_antennanp ANTENNA_4209 (.A(net76));
 sg13g2_antennanp ANTENNA_4210 (.A(net76));
 sg13g2_antennanp ANTENNA_4211 (.A(net76));
 sg13g2_antennanp ANTENNA_4212 (.A(net76));
 sg13g2_antennanp ANTENNA_4213 (.A(net76));
 sg13g2_antennanp ANTENNA_4214 (.A(net76));
 sg13g2_antennanp ANTENNA_4215 (.A(net78));
 sg13g2_antennanp ANTENNA_4216 (.A(net78));
 sg13g2_antennanp ANTENNA_4217 (.A(net78));
 sg13g2_antennanp ANTENNA_4218 (.A(net78));
 sg13g2_antennanp ANTENNA_4219 (.A(net78));
 sg13g2_antennanp ANTENNA_4220 (.A(net78));
 sg13g2_antennanp ANTENNA_4221 (.A(net78));
 sg13g2_antennanp ANTENNA_4222 (.A(net78));
 sg13g2_antennanp ANTENNA_4223 (.A(net78));
 sg13g2_antennanp ANTENNA_4224 (.A(net84));
 sg13g2_antennanp ANTENNA_4225 (.A(net84));
 sg13g2_antennanp ANTENNA_4226 (.A(net84));
 sg13g2_antennanp ANTENNA_4227 (.A(net84));
 sg13g2_antennanp ANTENNA_4228 (.A(net84));
 sg13g2_antennanp ANTENNA_4229 (.A(net84));
 sg13g2_antennanp ANTENNA_4230 (.A(net84));
 sg13g2_antennanp ANTENNA_4231 (.A(net84));
 sg13g2_antennanp ANTENNA_4232 (.A(net89));
 sg13g2_antennanp ANTENNA_4233 (.A(net89));
 sg13g2_antennanp ANTENNA_4234 (.A(net89));
 sg13g2_antennanp ANTENNA_4235 (.A(net89));
 sg13g2_antennanp ANTENNA_4236 (.A(net89));
 sg13g2_antennanp ANTENNA_4237 (.A(net89));
 sg13g2_antennanp ANTENNA_4238 (.A(net89));
 sg13g2_antennanp ANTENNA_4239 (.A(net89));
 sg13g2_antennanp ANTENNA_4240 (.A(net89));
 sg13g2_antennanp ANTENNA_4241 (.A(net91));
 sg13g2_antennanp ANTENNA_4242 (.A(net91));
 sg13g2_antennanp ANTENNA_4243 (.A(net91));
 sg13g2_antennanp ANTENNA_4244 (.A(net91));
 sg13g2_antennanp ANTENNA_4245 (.A(net91));
 sg13g2_antennanp ANTENNA_4246 (.A(net91));
 sg13g2_antennanp ANTENNA_4247 (.A(net91));
 sg13g2_antennanp ANTENNA_4248 (.A(net91));
 sg13g2_antennanp ANTENNA_4249 (.A(net94));
 sg13g2_antennanp ANTENNA_4250 (.A(net94));
 sg13g2_antennanp ANTENNA_4251 (.A(net94));
 sg13g2_antennanp ANTENNA_4252 (.A(net94));
 sg13g2_antennanp ANTENNA_4253 (.A(net94));
 sg13g2_antennanp ANTENNA_4254 (.A(net94));
 sg13g2_antennanp ANTENNA_4255 (.A(net94));
 sg13g2_antennanp ANTENNA_4256 (.A(net94));
 sg13g2_antennanp ANTENNA_4257 (.A(net100));
 sg13g2_antennanp ANTENNA_4258 (.A(net100));
 sg13g2_antennanp ANTENNA_4259 (.A(net100));
 sg13g2_antennanp ANTENNA_4260 (.A(net100));
 sg13g2_antennanp ANTENNA_4261 (.A(net100));
 sg13g2_antennanp ANTENNA_4262 (.A(net100));
 sg13g2_antennanp ANTENNA_4263 (.A(net100));
 sg13g2_antennanp ANTENNA_4264 (.A(net100));
 sg13g2_antennanp ANTENNA_4265 (.A(net100));
 sg13g2_antennanp ANTENNA_4266 (.A(net106));
 sg13g2_antennanp ANTENNA_4267 (.A(net106));
 sg13g2_antennanp ANTENNA_4268 (.A(net106));
 sg13g2_antennanp ANTENNA_4269 (.A(net106));
 sg13g2_antennanp ANTENNA_4270 (.A(net106));
 sg13g2_antennanp ANTENNA_4271 (.A(net106));
 sg13g2_antennanp ANTENNA_4272 (.A(net106));
 sg13g2_antennanp ANTENNA_4273 (.A(net106));
 sg13g2_antennanp ANTENNA_4274 (.A(net106));
 sg13g2_antennanp ANTENNA_4275 (.A(net107));
 sg13g2_antennanp ANTENNA_4276 (.A(net107));
 sg13g2_antennanp ANTENNA_4277 (.A(net107));
 sg13g2_antennanp ANTENNA_4278 (.A(net107));
 sg13g2_antennanp ANTENNA_4279 (.A(net107));
 sg13g2_antennanp ANTENNA_4280 (.A(net107));
 sg13g2_antennanp ANTENNA_4281 (.A(net107));
 sg13g2_antennanp ANTENNA_4282 (.A(net107));
 sg13g2_antennanp ANTENNA_4283 (.A(net107));
 sg13g2_antennanp ANTENNA_4284 (.A(net113));
 sg13g2_antennanp ANTENNA_4285 (.A(net113));
 sg13g2_antennanp ANTENNA_4286 (.A(net113));
 sg13g2_antennanp ANTENNA_4287 (.A(net113));
 sg13g2_antennanp ANTENNA_4288 (.A(net113));
 sg13g2_antennanp ANTENNA_4289 (.A(net113));
 sg13g2_antennanp ANTENNA_4290 (.A(net113));
 sg13g2_antennanp ANTENNA_4291 (.A(net113));
 sg13g2_antennanp ANTENNA_4292 (.A(net125));
 sg13g2_antennanp ANTENNA_4293 (.A(net125));
 sg13g2_antennanp ANTENNA_4294 (.A(net125));
 sg13g2_antennanp ANTENNA_4295 (.A(net125));
 sg13g2_antennanp ANTENNA_4296 (.A(net125));
 sg13g2_antennanp ANTENNA_4297 (.A(net125));
 sg13g2_antennanp ANTENNA_4298 (.A(net125));
 sg13g2_antennanp ANTENNA_4299 (.A(net125));
 sg13g2_antennanp ANTENNA_4300 (.A(net125));
 sg13g2_antennanp ANTENNA_4301 (.A(net128));
 sg13g2_antennanp ANTENNA_4302 (.A(net128));
 sg13g2_antennanp ANTENNA_4303 (.A(net128));
 sg13g2_antennanp ANTENNA_4304 (.A(net128));
 sg13g2_antennanp ANTENNA_4305 (.A(net128));
 sg13g2_antennanp ANTENNA_4306 (.A(net128));
 sg13g2_antennanp ANTENNA_4307 (.A(net128));
 sg13g2_antennanp ANTENNA_4308 (.A(net128));
 sg13g2_antennanp ANTENNA_4309 (.A(net129));
 sg13g2_antennanp ANTENNA_4310 (.A(net129));
 sg13g2_antennanp ANTENNA_4311 (.A(net129));
 sg13g2_antennanp ANTENNA_4312 (.A(net129));
 sg13g2_antennanp ANTENNA_4313 (.A(net129));
 sg13g2_antennanp ANTENNA_4314 (.A(net129));
 sg13g2_antennanp ANTENNA_4315 (.A(net129));
 sg13g2_antennanp ANTENNA_4316 (.A(net129));
 sg13g2_antennanp ANTENNA_4317 (.A(net129));
 sg13g2_antennanp ANTENNA_4318 (.A(net142));
 sg13g2_antennanp ANTENNA_4319 (.A(net142));
 sg13g2_antennanp ANTENNA_4320 (.A(net142));
 sg13g2_antennanp ANTENNA_4321 (.A(net142));
 sg13g2_antennanp ANTENNA_4322 (.A(net142));
 sg13g2_antennanp ANTENNA_4323 (.A(net142));
 sg13g2_antennanp ANTENNA_4324 (.A(net142));
 sg13g2_antennanp ANTENNA_4325 (.A(net142));
 sg13g2_antennanp ANTENNA_4326 (.A(net142));
 sg13g2_antennanp ANTENNA_4327 (.A(net144));
 sg13g2_antennanp ANTENNA_4328 (.A(net144));
 sg13g2_antennanp ANTENNA_4329 (.A(net144));
 sg13g2_antennanp ANTENNA_4330 (.A(net144));
 sg13g2_antennanp ANTENNA_4331 (.A(net144));
 sg13g2_antennanp ANTENNA_4332 (.A(net144));
 sg13g2_antennanp ANTENNA_4333 (.A(net144));
 sg13g2_antennanp ANTENNA_4334 (.A(net144));
 sg13g2_antennanp ANTENNA_4335 (.A(net144));
 sg13g2_antennanp ANTENNA_4336 (.A(net153));
 sg13g2_antennanp ANTENNA_4337 (.A(net153));
 sg13g2_antennanp ANTENNA_4338 (.A(net153));
 sg13g2_antennanp ANTENNA_4339 (.A(net153));
 sg13g2_antennanp ANTENNA_4340 (.A(net153));
 sg13g2_antennanp ANTENNA_4341 (.A(net153));
 sg13g2_antennanp ANTENNA_4342 (.A(net153));
 sg13g2_antennanp ANTENNA_4343 (.A(net153));
 sg13g2_antennanp ANTENNA_4344 (.A(net153));
 sg13g2_antennanp ANTENNA_4345 (.A(net153));
 sg13g2_antennanp ANTENNA_4346 (.A(net153));
 sg13g2_antennanp ANTENNA_4347 (.A(net153));
 sg13g2_antennanp ANTENNA_4348 (.A(net153));
 sg13g2_antennanp ANTENNA_4349 (.A(net153));
 sg13g2_antennanp ANTENNA_4350 (.A(net153));
 sg13g2_antennanp ANTENNA_4351 (.A(net153));
 sg13g2_antennanp ANTENNA_4352 (.A(net153));
 sg13g2_antennanp ANTENNA_4353 (.A(net153));
 sg13g2_antennanp ANTENNA_4354 (.A(net164));
 sg13g2_antennanp ANTENNA_4355 (.A(net164));
 sg13g2_antennanp ANTENNA_4356 (.A(net164));
 sg13g2_antennanp ANTENNA_4357 (.A(net164));
 sg13g2_antennanp ANTENNA_4358 (.A(net164));
 sg13g2_antennanp ANTENNA_4359 (.A(net164));
 sg13g2_antennanp ANTENNA_4360 (.A(net164));
 sg13g2_antennanp ANTENNA_4361 (.A(net164));
 sg13g2_antennanp ANTENNA_4362 (.A(net164));
 sg13g2_antennanp ANTENNA_4363 (.A(net167));
 sg13g2_antennanp ANTENNA_4364 (.A(net167));
 sg13g2_antennanp ANTENNA_4365 (.A(net167));
 sg13g2_antennanp ANTENNA_4366 (.A(net167));
 sg13g2_antennanp ANTENNA_4367 (.A(net167));
 sg13g2_antennanp ANTENNA_4368 (.A(net167));
 sg13g2_antennanp ANTENNA_4369 (.A(net167));
 sg13g2_antennanp ANTENNA_4370 (.A(net167));
 sg13g2_antennanp ANTENNA_4371 (.A(net167));
 sg13g2_antennanp ANTENNA_4372 (.A(net182));
 sg13g2_antennanp ANTENNA_4373 (.A(net182));
 sg13g2_antennanp ANTENNA_4374 (.A(net182));
 sg13g2_antennanp ANTENNA_4375 (.A(net182));
 sg13g2_antennanp ANTENNA_4376 (.A(net182));
 sg13g2_antennanp ANTENNA_4377 (.A(net182));
 sg13g2_antennanp ANTENNA_4378 (.A(net182));
 sg13g2_antennanp ANTENNA_4379 (.A(net182));
 sg13g2_antennanp ANTENNA_4380 (.A(net185));
 sg13g2_antennanp ANTENNA_4381 (.A(net185));
 sg13g2_antennanp ANTENNA_4382 (.A(net185));
 sg13g2_antennanp ANTENNA_4383 (.A(net185));
 sg13g2_antennanp ANTENNA_4384 (.A(net185));
 sg13g2_antennanp ANTENNA_4385 (.A(net185));
 sg13g2_antennanp ANTENNA_4386 (.A(net185));
 sg13g2_antennanp ANTENNA_4387 (.A(net185));
 sg13g2_antennanp ANTENNA_4388 (.A(net185));
 sg13g2_antennanp ANTENNA_4389 (.A(net185));
 sg13g2_antennanp ANTENNA_4390 (.A(net185));
 sg13g2_antennanp ANTENNA_4391 (.A(net185));
 sg13g2_antennanp ANTENNA_4392 (.A(net198));
 sg13g2_antennanp ANTENNA_4393 (.A(net198));
 sg13g2_antennanp ANTENNA_4394 (.A(net198));
 sg13g2_antennanp ANTENNA_4395 (.A(net198));
 sg13g2_antennanp ANTENNA_4396 (.A(net198));
 sg13g2_antennanp ANTENNA_4397 (.A(net198));
 sg13g2_antennanp ANTENNA_4398 (.A(net198));
 sg13g2_antennanp ANTENNA_4399 (.A(net198));
 sg13g2_antennanp ANTENNA_4400 (.A(net210));
 sg13g2_antennanp ANTENNA_4401 (.A(net210));
 sg13g2_antennanp ANTENNA_4402 (.A(net210));
 sg13g2_antennanp ANTENNA_4403 (.A(net210));
 sg13g2_antennanp ANTENNA_4404 (.A(net210));
 sg13g2_antennanp ANTENNA_4405 (.A(net210));
 sg13g2_antennanp ANTENNA_4406 (.A(net210));
 sg13g2_antennanp ANTENNA_4407 (.A(net210));
 sg13g2_antennanp ANTENNA_4408 (.A(net210));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_4 FILLER_0_630 ();
 sg13g2_fill_2 FILLER_0_634 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_decap_8 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_0_868 ();
 sg13g2_decap_8 FILLER_0_875 ();
 sg13g2_decap_8 FILLER_0_882 ();
 sg13g2_decap_8 FILLER_0_889 ();
 sg13g2_decap_8 FILLER_0_896 ();
 sg13g2_decap_8 FILLER_0_903 ();
 sg13g2_decap_8 FILLER_0_910 ();
 sg13g2_decap_8 FILLER_0_917 ();
 sg13g2_decap_8 FILLER_0_924 ();
 sg13g2_decap_8 FILLER_0_931 ();
 sg13g2_decap_8 FILLER_0_938 ();
 sg13g2_decap_8 FILLER_0_945 ();
 sg13g2_decap_8 FILLER_0_952 ();
 sg13g2_decap_8 FILLER_0_959 ();
 sg13g2_decap_8 FILLER_0_966 ();
 sg13g2_decap_8 FILLER_0_973 ();
 sg13g2_decap_8 FILLER_0_980 ();
 sg13g2_decap_8 FILLER_0_987 ();
 sg13g2_decap_8 FILLER_0_994 ();
 sg13g2_decap_8 FILLER_0_1001 ();
 sg13g2_decap_8 FILLER_0_1008 ();
 sg13g2_decap_8 FILLER_0_1015 ();
 sg13g2_decap_8 FILLER_0_1022 ();
 sg13g2_decap_8 FILLER_0_1029 ();
 sg13g2_decap_8 FILLER_0_1036 ();
 sg13g2_decap_8 FILLER_0_1043 ();
 sg13g2_decap_8 FILLER_0_1050 ();
 sg13g2_decap_8 FILLER_0_1057 ();
 sg13g2_decap_8 FILLER_0_1064 ();
 sg13g2_decap_8 FILLER_0_1071 ();
 sg13g2_decap_8 FILLER_0_1078 ();
 sg13g2_decap_8 FILLER_0_1085 ();
 sg13g2_decap_8 FILLER_0_1092 ();
 sg13g2_decap_8 FILLER_0_1099 ();
 sg13g2_decap_8 FILLER_0_1106 ();
 sg13g2_decap_8 FILLER_0_1113 ();
 sg13g2_decap_8 FILLER_0_1120 ();
 sg13g2_decap_8 FILLER_0_1127 ();
 sg13g2_decap_8 FILLER_0_1134 ();
 sg13g2_decap_8 FILLER_0_1141 ();
 sg13g2_decap_8 FILLER_0_1148 ();
 sg13g2_decap_8 FILLER_0_1155 ();
 sg13g2_decap_8 FILLER_0_1162 ();
 sg13g2_decap_8 FILLER_0_1169 ();
 sg13g2_decap_8 FILLER_0_1176 ();
 sg13g2_decap_8 FILLER_0_1183 ();
 sg13g2_decap_8 FILLER_0_1190 ();
 sg13g2_decap_8 FILLER_0_1197 ();
 sg13g2_decap_8 FILLER_0_1204 ();
 sg13g2_decap_8 FILLER_0_1211 ();
 sg13g2_decap_8 FILLER_0_1218 ();
 sg13g2_decap_8 FILLER_0_1225 ();
 sg13g2_decap_8 FILLER_0_1232 ();
 sg13g2_decap_8 FILLER_0_1239 ();
 sg13g2_decap_8 FILLER_0_1246 ();
 sg13g2_decap_8 FILLER_0_1253 ();
 sg13g2_decap_8 FILLER_0_1260 ();
 sg13g2_decap_8 FILLER_0_1267 ();
 sg13g2_decap_8 FILLER_0_1274 ();
 sg13g2_decap_8 FILLER_0_1281 ();
 sg13g2_decap_8 FILLER_0_1288 ();
 sg13g2_decap_8 FILLER_0_1295 ();
 sg13g2_decap_8 FILLER_0_1302 ();
 sg13g2_decap_8 FILLER_0_1309 ();
 sg13g2_decap_8 FILLER_0_1316 ();
 sg13g2_decap_8 FILLER_0_1323 ();
 sg13g2_decap_8 FILLER_0_1330 ();
 sg13g2_decap_8 FILLER_0_1337 ();
 sg13g2_decap_8 FILLER_0_1344 ();
 sg13g2_decap_8 FILLER_0_1351 ();
 sg13g2_decap_8 FILLER_0_1358 ();
 sg13g2_decap_8 FILLER_0_1365 ();
 sg13g2_decap_8 FILLER_0_1372 ();
 sg13g2_decap_8 FILLER_0_1379 ();
 sg13g2_decap_8 FILLER_0_1386 ();
 sg13g2_decap_8 FILLER_0_1393 ();
 sg13g2_decap_8 FILLER_0_1400 ();
 sg13g2_decap_8 FILLER_0_1407 ();
 sg13g2_decap_8 FILLER_0_1414 ();
 sg13g2_decap_8 FILLER_0_1421 ();
 sg13g2_decap_8 FILLER_0_1428 ();
 sg13g2_decap_8 FILLER_0_1435 ();
 sg13g2_decap_8 FILLER_0_1442 ();
 sg13g2_decap_8 FILLER_0_1449 ();
 sg13g2_decap_8 FILLER_0_1456 ();
 sg13g2_decap_8 FILLER_0_1463 ();
 sg13g2_decap_8 FILLER_0_1470 ();
 sg13g2_decap_8 FILLER_0_1477 ();
 sg13g2_decap_8 FILLER_0_1484 ();
 sg13g2_decap_8 FILLER_0_1491 ();
 sg13g2_decap_8 FILLER_0_1498 ();
 sg13g2_decap_8 FILLER_0_1505 ();
 sg13g2_decap_8 FILLER_0_1512 ();
 sg13g2_decap_8 FILLER_0_1519 ();
 sg13g2_decap_8 FILLER_0_1526 ();
 sg13g2_decap_8 FILLER_0_1533 ();
 sg13g2_decap_8 FILLER_0_1540 ();
 sg13g2_decap_8 FILLER_0_1547 ();
 sg13g2_decap_8 FILLER_0_1554 ();
 sg13g2_decap_8 FILLER_0_1561 ();
 sg13g2_decap_8 FILLER_0_1568 ();
 sg13g2_decap_8 FILLER_0_1575 ();
 sg13g2_decap_8 FILLER_0_1582 ();
 sg13g2_decap_8 FILLER_0_1589 ();
 sg13g2_decap_8 FILLER_0_1596 ();
 sg13g2_decap_8 FILLER_0_1603 ();
 sg13g2_decap_8 FILLER_0_1610 ();
 sg13g2_decap_8 FILLER_0_1617 ();
 sg13g2_decap_8 FILLER_0_1624 ();
 sg13g2_decap_8 FILLER_0_1631 ();
 sg13g2_decap_8 FILLER_0_1638 ();
 sg13g2_decap_8 FILLER_0_1645 ();
 sg13g2_decap_8 FILLER_0_1652 ();
 sg13g2_decap_8 FILLER_0_1659 ();
 sg13g2_decap_8 FILLER_0_1666 ();
 sg13g2_decap_8 FILLER_0_1673 ();
 sg13g2_decap_8 FILLER_0_1680 ();
 sg13g2_decap_8 FILLER_0_1687 ();
 sg13g2_decap_8 FILLER_0_1694 ();
 sg13g2_decap_8 FILLER_0_1701 ();
 sg13g2_decap_8 FILLER_0_1708 ();
 sg13g2_decap_8 FILLER_0_1715 ();
 sg13g2_decap_8 FILLER_0_1722 ();
 sg13g2_decap_8 FILLER_0_1729 ();
 sg13g2_decap_8 FILLER_0_1736 ();
 sg13g2_decap_8 FILLER_0_1743 ();
 sg13g2_decap_8 FILLER_0_1750 ();
 sg13g2_decap_8 FILLER_0_1757 ();
 sg13g2_decap_8 FILLER_0_1764 ();
 sg13g2_decap_8 FILLER_0_1771 ();
 sg13g2_decap_8 FILLER_0_1778 ();
 sg13g2_decap_8 FILLER_0_1785 ();
 sg13g2_decap_8 FILLER_0_1792 ();
 sg13g2_decap_8 FILLER_0_1799 ();
 sg13g2_decap_8 FILLER_0_1806 ();
 sg13g2_decap_8 FILLER_0_1813 ();
 sg13g2_decap_8 FILLER_0_1820 ();
 sg13g2_decap_8 FILLER_0_1827 ();
 sg13g2_decap_8 FILLER_0_1834 ();
 sg13g2_decap_8 FILLER_0_1841 ();
 sg13g2_decap_8 FILLER_0_1848 ();
 sg13g2_decap_8 FILLER_0_1855 ();
 sg13g2_decap_8 FILLER_0_1862 ();
 sg13g2_decap_8 FILLER_0_1869 ();
 sg13g2_decap_8 FILLER_0_1876 ();
 sg13g2_decap_8 FILLER_0_1883 ();
 sg13g2_decap_8 FILLER_0_1890 ();
 sg13g2_decap_8 FILLER_0_1897 ();
 sg13g2_decap_8 FILLER_0_1904 ();
 sg13g2_decap_8 FILLER_0_1911 ();
 sg13g2_decap_8 FILLER_0_1918 ();
 sg13g2_decap_8 FILLER_0_1925 ();
 sg13g2_decap_8 FILLER_0_1932 ();
 sg13g2_decap_8 FILLER_0_1939 ();
 sg13g2_decap_8 FILLER_0_1946 ();
 sg13g2_decap_8 FILLER_0_1953 ();
 sg13g2_decap_8 FILLER_0_1960 ();
 sg13g2_decap_8 FILLER_0_1967 ();
 sg13g2_decap_8 FILLER_0_1974 ();
 sg13g2_decap_8 FILLER_0_1981 ();
 sg13g2_decap_8 FILLER_0_1988 ();
 sg13g2_decap_8 FILLER_0_1995 ();
 sg13g2_decap_8 FILLER_0_2002 ();
 sg13g2_decap_8 FILLER_0_2009 ();
 sg13g2_decap_8 FILLER_0_2016 ();
 sg13g2_decap_8 FILLER_0_2023 ();
 sg13g2_decap_8 FILLER_0_2030 ();
 sg13g2_decap_8 FILLER_0_2037 ();
 sg13g2_decap_8 FILLER_0_2044 ();
 sg13g2_decap_8 FILLER_0_2051 ();
 sg13g2_decap_8 FILLER_0_2058 ();
 sg13g2_decap_8 FILLER_0_2065 ();
 sg13g2_decap_8 FILLER_0_2072 ();
 sg13g2_decap_8 FILLER_0_2079 ();
 sg13g2_decap_8 FILLER_0_2086 ();
 sg13g2_decap_8 FILLER_0_2093 ();
 sg13g2_decap_8 FILLER_0_2100 ();
 sg13g2_decap_8 FILLER_0_2107 ();
 sg13g2_decap_8 FILLER_0_2114 ();
 sg13g2_decap_8 FILLER_0_2121 ();
 sg13g2_decap_8 FILLER_0_2128 ();
 sg13g2_decap_8 FILLER_0_2135 ();
 sg13g2_decap_8 FILLER_0_2142 ();
 sg13g2_decap_8 FILLER_0_2149 ();
 sg13g2_decap_8 FILLER_0_2156 ();
 sg13g2_decap_8 FILLER_0_2163 ();
 sg13g2_decap_8 FILLER_0_2170 ();
 sg13g2_decap_8 FILLER_0_2177 ();
 sg13g2_decap_8 FILLER_0_2184 ();
 sg13g2_decap_8 FILLER_0_2191 ();
 sg13g2_decap_8 FILLER_0_2198 ();
 sg13g2_decap_8 FILLER_0_2205 ();
 sg13g2_decap_8 FILLER_0_2212 ();
 sg13g2_decap_8 FILLER_0_2219 ();
 sg13g2_decap_8 FILLER_0_2226 ();
 sg13g2_decap_8 FILLER_0_2233 ();
 sg13g2_decap_8 FILLER_0_2240 ();
 sg13g2_decap_8 FILLER_0_2247 ();
 sg13g2_decap_8 FILLER_0_2254 ();
 sg13g2_decap_8 FILLER_0_2261 ();
 sg13g2_decap_8 FILLER_0_2268 ();
 sg13g2_decap_8 FILLER_0_2275 ();
 sg13g2_decap_8 FILLER_0_2282 ();
 sg13g2_decap_8 FILLER_0_2289 ();
 sg13g2_decap_8 FILLER_0_2296 ();
 sg13g2_decap_8 FILLER_0_2303 ();
 sg13g2_decap_8 FILLER_0_2310 ();
 sg13g2_decap_8 FILLER_0_2317 ();
 sg13g2_decap_8 FILLER_0_2324 ();
 sg13g2_decap_8 FILLER_0_2331 ();
 sg13g2_decap_8 FILLER_0_2338 ();
 sg13g2_decap_8 FILLER_0_2345 ();
 sg13g2_decap_8 FILLER_0_2352 ();
 sg13g2_decap_8 FILLER_0_2359 ();
 sg13g2_decap_8 FILLER_0_2366 ();
 sg13g2_decap_8 FILLER_0_2373 ();
 sg13g2_decap_8 FILLER_0_2380 ();
 sg13g2_decap_8 FILLER_0_2387 ();
 sg13g2_decap_8 FILLER_0_2394 ();
 sg13g2_decap_8 FILLER_0_2401 ();
 sg13g2_decap_8 FILLER_0_2408 ();
 sg13g2_decap_8 FILLER_0_2415 ();
 sg13g2_decap_8 FILLER_0_2422 ();
 sg13g2_decap_8 FILLER_0_2429 ();
 sg13g2_decap_8 FILLER_0_2436 ();
 sg13g2_decap_8 FILLER_0_2443 ();
 sg13g2_decap_8 FILLER_0_2450 ();
 sg13g2_decap_8 FILLER_0_2457 ();
 sg13g2_decap_8 FILLER_0_2464 ();
 sg13g2_decap_8 FILLER_0_2471 ();
 sg13g2_decap_8 FILLER_0_2478 ();
 sg13g2_decap_8 FILLER_0_2485 ();
 sg13g2_decap_8 FILLER_0_2492 ();
 sg13g2_decap_8 FILLER_0_2499 ();
 sg13g2_decap_8 FILLER_0_2506 ();
 sg13g2_decap_8 FILLER_0_2513 ();
 sg13g2_decap_8 FILLER_0_2520 ();
 sg13g2_decap_8 FILLER_0_2527 ();
 sg13g2_decap_8 FILLER_0_2534 ();
 sg13g2_decap_8 FILLER_0_2541 ();
 sg13g2_decap_8 FILLER_0_2548 ();
 sg13g2_decap_8 FILLER_0_2555 ();
 sg13g2_decap_8 FILLER_0_2562 ();
 sg13g2_decap_8 FILLER_0_2569 ();
 sg13g2_decap_8 FILLER_0_2576 ();
 sg13g2_decap_8 FILLER_0_2583 ();
 sg13g2_decap_8 FILLER_0_2590 ();
 sg13g2_decap_8 FILLER_0_2597 ();
 sg13g2_decap_8 FILLER_0_2604 ();
 sg13g2_decap_8 FILLER_0_2611 ();
 sg13g2_decap_8 FILLER_0_2618 ();
 sg13g2_decap_8 FILLER_0_2625 ();
 sg13g2_decap_8 FILLER_0_2632 ();
 sg13g2_decap_8 FILLER_0_2639 ();
 sg13g2_decap_8 FILLER_0_2646 ();
 sg13g2_decap_8 FILLER_0_2653 ();
 sg13g2_decap_8 FILLER_0_2660 ();
 sg13g2_fill_2 FILLER_0_2667 ();
 sg13g2_fill_1 FILLER_0_2669 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_fill_1 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_424 ();
 sg13g2_decap_8 FILLER_1_431 ();
 sg13g2_decap_8 FILLER_1_438 ();
 sg13g2_decap_8 FILLER_1_445 ();
 sg13g2_decap_8 FILLER_1_452 ();
 sg13g2_decap_8 FILLER_1_459 ();
 sg13g2_fill_2 FILLER_1_466 ();
 sg13g2_decap_8 FILLER_1_472 ();
 sg13g2_decap_8 FILLER_1_479 ();
 sg13g2_decap_8 FILLER_1_486 ();
 sg13g2_decap_4 FILLER_1_493 ();
 sg13g2_fill_1 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_502 ();
 sg13g2_decap_8 FILLER_1_509 ();
 sg13g2_decap_8 FILLER_1_516 ();
 sg13g2_decap_8 FILLER_1_523 ();
 sg13g2_decap_4 FILLER_1_530 ();
 sg13g2_fill_1 FILLER_1_534 ();
 sg13g2_decap_8 FILLER_1_538 ();
 sg13g2_decap_8 FILLER_1_545 ();
 sg13g2_decap_8 FILLER_1_552 ();
 sg13g2_decap_8 FILLER_1_559 ();
 sg13g2_decap_8 FILLER_1_566 ();
 sg13g2_decap_8 FILLER_1_573 ();
 sg13g2_decap_8 FILLER_1_580 ();
 sg13g2_fill_1 FILLER_1_587 ();
 sg13g2_decap_8 FILLER_1_592 ();
 sg13g2_decap_8 FILLER_1_599 ();
 sg13g2_decap_8 FILLER_1_606 ();
 sg13g2_decap_8 FILLER_1_613 ();
 sg13g2_decap_8 FILLER_1_620 ();
 sg13g2_decap_8 FILLER_1_646 ();
 sg13g2_decap_8 FILLER_1_653 ();
 sg13g2_fill_2 FILLER_1_660 ();
 sg13g2_decap_8 FILLER_1_671 ();
 sg13g2_decap_8 FILLER_1_678 ();
 sg13g2_decap_8 FILLER_1_685 ();
 sg13g2_decap_8 FILLER_1_692 ();
 sg13g2_decap_8 FILLER_1_699 ();
 sg13g2_fill_2 FILLER_1_706 ();
 sg13g2_fill_1 FILLER_1_708 ();
 sg13g2_decap_8 FILLER_1_712 ();
 sg13g2_decap_8 FILLER_1_719 ();
 sg13g2_decap_8 FILLER_1_726 ();
 sg13g2_decap_8 FILLER_1_733 ();
 sg13g2_decap_8 FILLER_1_740 ();
 sg13g2_decap_8 FILLER_1_747 ();
 sg13g2_decap_8 FILLER_1_754 ();
 sg13g2_decap_8 FILLER_1_761 ();
 sg13g2_decap_8 FILLER_1_768 ();
 sg13g2_decap_8 FILLER_1_775 ();
 sg13g2_decap_8 FILLER_1_782 ();
 sg13g2_decap_8 FILLER_1_789 ();
 sg13g2_decap_8 FILLER_1_796 ();
 sg13g2_decap_8 FILLER_1_803 ();
 sg13g2_decap_8 FILLER_1_810 ();
 sg13g2_decap_8 FILLER_1_817 ();
 sg13g2_decap_8 FILLER_1_824 ();
 sg13g2_decap_8 FILLER_1_831 ();
 sg13g2_decap_8 FILLER_1_838 ();
 sg13g2_decap_4 FILLER_1_845 ();
 sg13g2_fill_2 FILLER_1_849 ();
 sg13g2_decap_8 FILLER_1_859 ();
 sg13g2_decap_8 FILLER_1_866 ();
 sg13g2_decap_8 FILLER_1_873 ();
 sg13g2_decap_8 FILLER_1_880 ();
 sg13g2_decap_8 FILLER_1_887 ();
 sg13g2_decap_8 FILLER_1_894 ();
 sg13g2_decap_8 FILLER_1_901 ();
 sg13g2_decap_8 FILLER_1_908 ();
 sg13g2_decap_8 FILLER_1_915 ();
 sg13g2_decap_8 FILLER_1_922 ();
 sg13g2_decap_8 FILLER_1_929 ();
 sg13g2_decap_8 FILLER_1_936 ();
 sg13g2_decap_8 FILLER_1_943 ();
 sg13g2_decap_8 FILLER_1_950 ();
 sg13g2_decap_8 FILLER_1_957 ();
 sg13g2_decap_8 FILLER_1_964 ();
 sg13g2_decap_8 FILLER_1_971 ();
 sg13g2_decap_8 FILLER_1_978 ();
 sg13g2_decap_8 FILLER_1_985 ();
 sg13g2_decap_8 FILLER_1_992 ();
 sg13g2_decap_8 FILLER_1_999 ();
 sg13g2_decap_8 FILLER_1_1006 ();
 sg13g2_decap_8 FILLER_1_1013 ();
 sg13g2_decap_4 FILLER_1_1020 ();
 sg13g2_fill_1 FILLER_1_1024 ();
 sg13g2_decap_8 FILLER_1_1028 ();
 sg13g2_decap_8 FILLER_1_1035 ();
 sg13g2_decap_8 FILLER_1_1042 ();
 sg13g2_decap_8 FILLER_1_1049 ();
 sg13g2_decap_8 FILLER_1_1056 ();
 sg13g2_decap_8 FILLER_1_1063 ();
 sg13g2_decap_8 FILLER_1_1070 ();
 sg13g2_decap_8 FILLER_1_1077 ();
 sg13g2_decap_8 FILLER_1_1084 ();
 sg13g2_decap_4 FILLER_1_1091 ();
 sg13g2_decap_8 FILLER_1_1106 ();
 sg13g2_decap_8 FILLER_1_1113 ();
 sg13g2_decap_8 FILLER_1_1120 ();
 sg13g2_decap_8 FILLER_1_1127 ();
 sg13g2_decap_8 FILLER_1_1134 ();
 sg13g2_decap_8 FILLER_1_1141 ();
 sg13g2_decap_8 FILLER_1_1148 ();
 sg13g2_decap_8 FILLER_1_1155 ();
 sg13g2_decap_8 FILLER_1_1162 ();
 sg13g2_decap_8 FILLER_1_1169 ();
 sg13g2_decap_8 FILLER_1_1176 ();
 sg13g2_decap_8 FILLER_1_1183 ();
 sg13g2_fill_2 FILLER_1_1190 ();
 sg13g2_fill_1 FILLER_1_1207 ();
 sg13g2_fill_2 FILLER_1_1223 ();
 sg13g2_decap_8 FILLER_1_1237 ();
 sg13g2_decap_8 FILLER_1_1244 ();
 sg13g2_decap_8 FILLER_1_1251 ();
 sg13g2_decap_8 FILLER_1_1258 ();
 sg13g2_fill_1 FILLER_1_1265 ();
 sg13g2_decap_8 FILLER_1_1269 ();
 sg13g2_decap_8 FILLER_1_1276 ();
 sg13g2_decap_8 FILLER_1_1283 ();
 sg13g2_decap_8 FILLER_1_1290 ();
 sg13g2_decap_8 FILLER_1_1297 ();
 sg13g2_decap_8 FILLER_1_1304 ();
 sg13g2_decap_8 FILLER_1_1311 ();
 sg13g2_decap_8 FILLER_1_1318 ();
 sg13g2_decap_8 FILLER_1_1325 ();
 sg13g2_decap_8 FILLER_1_1332 ();
 sg13g2_decap_8 FILLER_1_1339 ();
 sg13g2_decap_8 FILLER_1_1346 ();
 sg13g2_decap_8 FILLER_1_1353 ();
 sg13g2_decap_8 FILLER_1_1360 ();
 sg13g2_decap_8 FILLER_1_1367 ();
 sg13g2_decap_8 FILLER_1_1374 ();
 sg13g2_decap_8 FILLER_1_1381 ();
 sg13g2_decap_8 FILLER_1_1388 ();
 sg13g2_decap_8 FILLER_1_1395 ();
 sg13g2_decap_8 FILLER_1_1402 ();
 sg13g2_decap_8 FILLER_1_1409 ();
 sg13g2_decap_8 FILLER_1_1416 ();
 sg13g2_decap_8 FILLER_1_1423 ();
 sg13g2_decap_8 FILLER_1_1430 ();
 sg13g2_decap_8 FILLER_1_1437 ();
 sg13g2_decap_8 FILLER_1_1444 ();
 sg13g2_decap_8 FILLER_1_1451 ();
 sg13g2_decap_8 FILLER_1_1458 ();
 sg13g2_decap_8 FILLER_1_1465 ();
 sg13g2_decap_8 FILLER_1_1472 ();
 sg13g2_decap_8 FILLER_1_1479 ();
 sg13g2_decap_8 FILLER_1_1486 ();
 sg13g2_decap_8 FILLER_1_1493 ();
 sg13g2_decap_8 FILLER_1_1500 ();
 sg13g2_decap_4 FILLER_1_1507 ();
 sg13g2_decap_8 FILLER_1_1526 ();
 sg13g2_decap_8 FILLER_1_1533 ();
 sg13g2_decap_8 FILLER_1_1540 ();
 sg13g2_decap_8 FILLER_1_1547 ();
 sg13g2_fill_2 FILLER_1_1554 ();
 sg13g2_fill_1 FILLER_1_1556 ();
 sg13g2_decap_8 FILLER_1_1564 ();
 sg13g2_decap_8 FILLER_1_1571 ();
 sg13g2_decap_8 FILLER_1_1578 ();
 sg13g2_decap_8 FILLER_1_1585 ();
 sg13g2_decap_8 FILLER_1_1592 ();
 sg13g2_decap_8 FILLER_1_1599 ();
 sg13g2_decap_8 FILLER_1_1606 ();
 sg13g2_decap_8 FILLER_1_1613 ();
 sg13g2_decap_8 FILLER_1_1620 ();
 sg13g2_decap_8 FILLER_1_1627 ();
 sg13g2_decap_8 FILLER_1_1634 ();
 sg13g2_decap_8 FILLER_1_1641 ();
 sg13g2_decap_8 FILLER_1_1648 ();
 sg13g2_decap_8 FILLER_1_1655 ();
 sg13g2_decap_8 FILLER_1_1662 ();
 sg13g2_decap_8 FILLER_1_1669 ();
 sg13g2_decap_8 FILLER_1_1676 ();
 sg13g2_decap_8 FILLER_1_1683 ();
 sg13g2_decap_8 FILLER_1_1690 ();
 sg13g2_decap_8 FILLER_1_1697 ();
 sg13g2_decap_8 FILLER_1_1704 ();
 sg13g2_decap_8 FILLER_1_1711 ();
 sg13g2_decap_8 FILLER_1_1718 ();
 sg13g2_decap_8 FILLER_1_1725 ();
 sg13g2_decap_8 FILLER_1_1732 ();
 sg13g2_decap_8 FILLER_1_1739 ();
 sg13g2_decap_8 FILLER_1_1746 ();
 sg13g2_decap_8 FILLER_1_1753 ();
 sg13g2_decap_8 FILLER_1_1760 ();
 sg13g2_decap_8 FILLER_1_1767 ();
 sg13g2_decap_8 FILLER_1_1774 ();
 sg13g2_decap_8 FILLER_1_1781 ();
 sg13g2_decap_8 FILLER_1_1788 ();
 sg13g2_decap_8 FILLER_1_1795 ();
 sg13g2_decap_8 FILLER_1_1802 ();
 sg13g2_decap_8 FILLER_1_1809 ();
 sg13g2_decap_8 FILLER_1_1816 ();
 sg13g2_decap_8 FILLER_1_1823 ();
 sg13g2_decap_8 FILLER_1_1830 ();
 sg13g2_decap_8 FILLER_1_1837 ();
 sg13g2_decap_8 FILLER_1_1844 ();
 sg13g2_decap_8 FILLER_1_1851 ();
 sg13g2_decap_8 FILLER_1_1858 ();
 sg13g2_decap_8 FILLER_1_1865 ();
 sg13g2_decap_8 FILLER_1_1872 ();
 sg13g2_decap_8 FILLER_1_1879 ();
 sg13g2_decap_8 FILLER_1_1886 ();
 sg13g2_decap_8 FILLER_1_1893 ();
 sg13g2_decap_8 FILLER_1_1900 ();
 sg13g2_decap_8 FILLER_1_1907 ();
 sg13g2_decap_8 FILLER_1_1914 ();
 sg13g2_decap_8 FILLER_1_1921 ();
 sg13g2_decap_8 FILLER_1_1928 ();
 sg13g2_decap_8 FILLER_1_1935 ();
 sg13g2_decap_8 FILLER_1_1942 ();
 sg13g2_decap_8 FILLER_1_1949 ();
 sg13g2_decap_8 FILLER_1_1956 ();
 sg13g2_decap_8 FILLER_1_1963 ();
 sg13g2_decap_8 FILLER_1_1970 ();
 sg13g2_decap_8 FILLER_1_1977 ();
 sg13g2_decap_8 FILLER_1_1984 ();
 sg13g2_decap_8 FILLER_1_1991 ();
 sg13g2_decap_8 FILLER_1_1998 ();
 sg13g2_decap_8 FILLER_1_2005 ();
 sg13g2_decap_8 FILLER_1_2012 ();
 sg13g2_decap_8 FILLER_1_2019 ();
 sg13g2_decap_8 FILLER_1_2026 ();
 sg13g2_decap_8 FILLER_1_2033 ();
 sg13g2_decap_8 FILLER_1_2040 ();
 sg13g2_decap_8 FILLER_1_2047 ();
 sg13g2_decap_8 FILLER_1_2054 ();
 sg13g2_decap_8 FILLER_1_2061 ();
 sg13g2_decap_8 FILLER_1_2068 ();
 sg13g2_decap_8 FILLER_1_2075 ();
 sg13g2_decap_8 FILLER_1_2082 ();
 sg13g2_decap_8 FILLER_1_2089 ();
 sg13g2_decap_8 FILLER_1_2096 ();
 sg13g2_decap_8 FILLER_1_2103 ();
 sg13g2_decap_8 FILLER_1_2110 ();
 sg13g2_decap_8 FILLER_1_2117 ();
 sg13g2_decap_8 FILLER_1_2124 ();
 sg13g2_decap_8 FILLER_1_2131 ();
 sg13g2_decap_8 FILLER_1_2138 ();
 sg13g2_decap_8 FILLER_1_2145 ();
 sg13g2_decap_8 FILLER_1_2152 ();
 sg13g2_decap_8 FILLER_1_2159 ();
 sg13g2_decap_8 FILLER_1_2166 ();
 sg13g2_decap_8 FILLER_1_2173 ();
 sg13g2_decap_8 FILLER_1_2180 ();
 sg13g2_decap_8 FILLER_1_2187 ();
 sg13g2_decap_8 FILLER_1_2194 ();
 sg13g2_decap_8 FILLER_1_2201 ();
 sg13g2_decap_8 FILLER_1_2208 ();
 sg13g2_decap_8 FILLER_1_2215 ();
 sg13g2_decap_8 FILLER_1_2222 ();
 sg13g2_decap_8 FILLER_1_2229 ();
 sg13g2_decap_8 FILLER_1_2236 ();
 sg13g2_decap_8 FILLER_1_2243 ();
 sg13g2_decap_8 FILLER_1_2250 ();
 sg13g2_decap_8 FILLER_1_2257 ();
 sg13g2_decap_8 FILLER_1_2264 ();
 sg13g2_decap_8 FILLER_1_2271 ();
 sg13g2_decap_8 FILLER_1_2278 ();
 sg13g2_decap_8 FILLER_1_2285 ();
 sg13g2_decap_8 FILLER_1_2292 ();
 sg13g2_decap_8 FILLER_1_2299 ();
 sg13g2_decap_8 FILLER_1_2306 ();
 sg13g2_decap_8 FILLER_1_2313 ();
 sg13g2_decap_8 FILLER_1_2320 ();
 sg13g2_decap_8 FILLER_1_2327 ();
 sg13g2_decap_8 FILLER_1_2334 ();
 sg13g2_decap_8 FILLER_1_2341 ();
 sg13g2_decap_8 FILLER_1_2348 ();
 sg13g2_decap_8 FILLER_1_2355 ();
 sg13g2_decap_8 FILLER_1_2362 ();
 sg13g2_decap_8 FILLER_1_2369 ();
 sg13g2_decap_8 FILLER_1_2376 ();
 sg13g2_decap_8 FILLER_1_2383 ();
 sg13g2_decap_8 FILLER_1_2390 ();
 sg13g2_decap_8 FILLER_1_2397 ();
 sg13g2_decap_8 FILLER_1_2404 ();
 sg13g2_decap_8 FILLER_1_2411 ();
 sg13g2_decap_8 FILLER_1_2418 ();
 sg13g2_decap_8 FILLER_1_2425 ();
 sg13g2_decap_8 FILLER_1_2432 ();
 sg13g2_decap_8 FILLER_1_2439 ();
 sg13g2_decap_8 FILLER_1_2446 ();
 sg13g2_decap_8 FILLER_1_2453 ();
 sg13g2_decap_8 FILLER_1_2460 ();
 sg13g2_decap_8 FILLER_1_2467 ();
 sg13g2_decap_8 FILLER_1_2474 ();
 sg13g2_decap_8 FILLER_1_2481 ();
 sg13g2_decap_8 FILLER_1_2488 ();
 sg13g2_decap_8 FILLER_1_2495 ();
 sg13g2_decap_8 FILLER_1_2502 ();
 sg13g2_decap_8 FILLER_1_2509 ();
 sg13g2_decap_8 FILLER_1_2516 ();
 sg13g2_decap_8 FILLER_1_2523 ();
 sg13g2_decap_8 FILLER_1_2530 ();
 sg13g2_decap_8 FILLER_1_2537 ();
 sg13g2_decap_8 FILLER_1_2544 ();
 sg13g2_decap_8 FILLER_1_2551 ();
 sg13g2_decap_8 FILLER_1_2558 ();
 sg13g2_decap_8 FILLER_1_2565 ();
 sg13g2_decap_8 FILLER_1_2572 ();
 sg13g2_decap_8 FILLER_1_2579 ();
 sg13g2_decap_8 FILLER_1_2586 ();
 sg13g2_decap_8 FILLER_1_2593 ();
 sg13g2_decap_8 FILLER_1_2600 ();
 sg13g2_decap_8 FILLER_1_2607 ();
 sg13g2_decap_8 FILLER_1_2614 ();
 sg13g2_decap_8 FILLER_1_2621 ();
 sg13g2_decap_8 FILLER_1_2628 ();
 sg13g2_decap_8 FILLER_1_2635 ();
 sg13g2_decap_8 FILLER_1_2642 ();
 sg13g2_decap_8 FILLER_1_2649 ();
 sg13g2_decap_8 FILLER_1_2656 ();
 sg13g2_decap_8 FILLER_1_2663 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_4 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_4 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_296 ();
 sg13g2_decap_8 FILLER_2_303 ();
 sg13g2_decap_8 FILLER_2_310 ();
 sg13g2_decap_8 FILLER_2_317 ();
 sg13g2_decap_8 FILLER_2_324 ();
 sg13g2_decap_8 FILLER_2_331 ();
 sg13g2_decap_8 FILLER_2_338 ();
 sg13g2_decap_8 FILLER_2_345 ();
 sg13g2_decap_8 FILLER_2_352 ();
 sg13g2_decap_8 FILLER_2_359 ();
 sg13g2_decap_8 FILLER_2_366 ();
 sg13g2_decap_8 FILLER_2_373 ();
 sg13g2_decap_8 FILLER_2_380 ();
 sg13g2_decap_8 FILLER_2_387 ();
 sg13g2_fill_2 FILLER_2_394 ();
 sg13g2_fill_1 FILLER_2_396 ();
 sg13g2_fill_2 FILLER_2_400 ();
 sg13g2_fill_1 FILLER_2_402 ();
 sg13g2_decap_4 FILLER_2_409 ();
 sg13g2_fill_2 FILLER_2_413 ();
 sg13g2_fill_1 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_433 ();
 sg13g2_decap_8 FILLER_2_440 ();
 sg13g2_decap_8 FILLER_2_447 ();
 sg13g2_decap_8 FILLER_2_454 ();
 sg13g2_fill_2 FILLER_2_461 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_fill_2 FILLER_2_511 ();
 sg13g2_fill_1 FILLER_2_513 ();
 sg13g2_decap_8 FILLER_2_517 ();
 sg13g2_decap_8 FILLER_2_524 ();
 sg13g2_decap_4 FILLER_2_531 ();
 sg13g2_decap_8 FILLER_2_540 ();
 sg13g2_decap_8 FILLER_2_547 ();
 sg13g2_decap_8 FILLER_2_554 ();
 sg13g2_decap_8 FILLER_2_561 ();
 sg13g2_decap_8 FILLER_2_568 ();
 sg13g2_decap_8 FILLER_2_575 ();
 sg13g2_decap_4 FILLER_2_582 ();
 sg13g2_fill_1 FILLER_2_586 ();
 sg13g2_decap_8 FILLER_2_591 ();
 sg13g2_decap_4 FILLER_2_598 ();
 sg13g2_fill_2 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_608 ();
 sg13g2_decap_8 FILLER_2_615 ();
 sg13g2_decap_8 FILLER_2_622 ();
 sg13g2_decap_8 FILLER_2_629 ();
 sg13g2_decap_8 FILLER_2_636 ();
 sg13g2_decap_8 FILLER_2_643 ();
 sg13g2_decap_4 FILLER_2_650 ();
 sg13g2_fill_2 FILLER_2_654 ();
 sg13g2_fill_2 FILLER_2_660 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_fill_2 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_696 ();
 sg13g2_fill_2 FILLER_2_703 ();
 sg13g2_fill_1 FILLER_2_705 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_4 FILLER_2_742 ();
 sg13g2_fill_1 FILLER_2_746 ();
 sg13g2_decap_8 FILLER_2_750 ();
 sg13g2_decap_8 FILLER_2_757 ();
 sg13g2_decap_8 FILLER_2_764 ();
 sg13g2_decap_8 FILLER_2_771 ();
 sg13g2_decap_8 FILLER_2_778 ();
 sg13g2_fill_1 FILLER_2_785 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_fill_1 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_820 ();
 sg13g2_decap_8 FILLER_2_827 ();
 sg13g2_fill_2 FILLER_2_834 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_fill_2 FILLER_2_854 ();
 sg13g2_decap_8 FILLER_2_860 ();
 sg13g2_decap_8 FILLER_2_867 ();
 sg13g2_decap_8 FILLER_2_874 ();
 sg13g2_decap_8 FILLER_2_881 ();
 sg13g2_decap_8 FILLER_2_888 ();
 sg13g2_decap_8 FILLER_2_895 ();
 sg13g2_fill_1 FILLER_2_902 ();
 sg13g2_decap_8 FILLER_2_915 ();
 sg13g2_decap_8 FILLER_2_922 ();
 sg13g2_decap_8 FILLER_2_929 ();
 sg13g2_decap_4 FILLER_2_936 ();
 sg13g2_fill_1 FILLER_2_940 ();
 sg13g2_decap_4 FILLER_2_965 ();
 sg13g2_decap_8 FILLER_2_984 ();
 sg13g2_decap_8 FILLER_2_991 ();
 sg13g2_decap_8 FILLER_2_998 ();
 sg13g2_decap_8 FILLER_2_1005 ();
 sg13g2_decap_8 FILLER_2_1012 ();
 sg13g2_decap_4 FILLER_2_1019 ();
 sg13g2_fill_2 FILLER_2_1023 ();
 sg13g2_decap_8 FILLER_2_1030 ();
 sg13g2_decap_4 FILLER_2_1037 ();
 sg13g2_fill_2 FILLER_2_1057 ();
 sg13g2_fill_2 FILLER_2_1063 ();
 sg13g2_decap_8 FILLER_2_1068 ();
 sg13g2_decap_8 FILLER_2_1075 ();
 sg13g2_decap_8 FILLER_2_1082 ();
 sg13g2_decap_8 FILLER_2_1089 ();
 sg13g2_decap_8 FILLER_2_1096 ();
 sg13g2_decap_8 FILLER_2_1103 ();
 sg13g2_decap_8 FILLER_2_1110 ();
 sg13g2_decap_8 FILLER_2_1117 ();
 sg13g2_decap_8 FILLER_2_1124 ();
 sg13g2_decap_8 FILLER_2_1131 ();
 sg13g2_fill_1 FILLER_2_1138 ();
 sg13g2_decap_8 FILLER_2_1147 ();
 sg13g2_decap_8 FILLER_2_1154 ();
 sg13g2_decap_8 FILLER_2_1161 ();
 sg13g2_decap_8 FILLER_2_1168 ();
 sg13g2_decap_4 FILLER_2_1175 ();
 sg13g2_fill_1 FILLER_2_1179 ();
 sg13g2_decap_8 FILLER_2_1188 ();
 sg13g2_decap_8 FILLER_2_1195 ();
 sg13g2_fill_2 FILLER_2_1202 ();
 sg13g2_decap_8 FILLER_2_1208 ();
 sg13g2_fill_2 FILLER_2_1215 ();
 sg13g2_decap_4 FILLER_2_1221 ();
 sg13g2_decap_8 FILLER_2_1229 ();
 sg13g2_decap_8 FILLER_2_1236 ();
 sg13g2_decap_4 FILLER_2_1243 ();
 sg13g2_fill_2 FILLER_2_1247 ();
 sg13g2_fill_2 FILLER_2_1264 ();
 sg13g2_decap_8 FILLER_2_1276 ();
 sg13g2_decap_4 FILLER_2_1283 ();
 sg13g2_fill_1 FILLER_2_1287 ();
 sg13g2_decap_8 FILLER_2_1294 ();
 sg13g2_decap_8 FILLER_2_1301 ();
 sg13g2_decap_8 FILLER_2_1308 ();
 sg13g2_decap_8 FILLER_2_1315 ();
 sg13g2_decap_8 FILLER_2_1322 ();
 sg13g2_fill_2 FILLER_2_1329 ();
 sg13g2_decap_4 FILLER_2_1335 ();
 sg13g2_fill_1 FILLER_2_1339 ();
 sg13g2_decap_8 FILLER_2_1345 ();
 sg13g2_decap_8 FILLER_2_1352 ();
 sg13g2_decap_8 FILLER_2_1359 ();
 sg13g2_decap_4 FILLER_2_1366 ();
 sg13g2_fill_2 FILLER_2_1376 ();
 sg13g2_decap_8 FILLER_2_1391 ();
 sg13g2_decap_8 FILLER_2_1398 ();
 sg13g2_decap_8 FILLER_2_1405 ();
 sg13g2_decap_8 FILLER_2_1412 ();
 sg13g2_decap_8 FILLER_2_1419 ();
 sg13g2_decap_8 FILLER_2_1426 ();
 sg13g2_fill_2 FILLER_2_1433 ();
 sg13g2_decap_8 FILLER_2_1441 ();
 sg13g2_decap_4 FILLER_2_1448 ();
 sg13g2_fill_1 FILLER_2_1452 ();
 sg13g2_decap_8 FILLER_2_1457 ();
 sg13g2_decap_8 FILLER_2_1464 ();
 sg13g2_decap_8 FILLER_2_1471 ();
 sg13g2_decap_8 FILLER_2_1478 ();
 sg13g2_decap_8 FILLER_2_1485 ();
 sg13g2_decap_8 FILLER_2_1492 ();
 sg13g2_decap_8 FILLER_2_1499 ();
 sg13g2_decap_4 FILLER_2_1506 ();
 sg13g2_fill_1 FILLER_2_1510 ();
 sg13g2_fill_2 FILLER_2_1519 ();
 sg13g2_decap_8 FILLER_2_1525 ();
 sg13g2_decap_8 FILLER_2_1532 ();
 sg13g2_decap_8 FILLER_2_1539 ();
 sg13g2_decap_4 FILLER_2_1552 ();
 sg13g2_fill_1 FILLER_2_1556 ();
 sg13g2_decap_8 FILLER_2_1567 ();
 sg13g2_decap_8 FILLER_2_1574 ();
 sg13g2_decap_8 FILLER_2_1581 ();
 sg13g2_decap_8 FILLER_2_1588 ();
 sg13g2_decap_8 FILLER_2_1595 ();
 sg13g2_decap_8 FILLER_2_1602 ();
 sg13g2_decap_8 FILLER_2_1609 ();
 sg13g2_decap_8 FILLER_2_1616 ();
 sg13g2_decap_4 FILLER_2_1623 ();
 sg13g2_decap_4 FILLER_2_1635 ();
 sg13g2_fill_1 FILLER_2_1639 ();
 sg13g2_decap_8 FILLER_2_1653 ();
 sg13g2_decap_8 FILLER_2_1660 ();
 sg13g2_decap_8 FILLER_2_1667 ();
 sg13g2_fill_1 FILLER_2_1674 ();
 sg13g2_decap_8 FILLER_2_1679 ();
 sg13g2_decap_8 FILLER_2_1686 ();
 sg13g2_fill_2 FILLER_2_1693 ();
 sg13g2_decap_8 FILLER_2_1699 ();
 sg13g2_decap_8 FILLER_2_1714 ();
 sg13g2_decap_8 FILLER_2_1734 ();
 sg13g2_decap_8 FILLER_2_1741 ();
 sg13g2_decap_8 FILLER_2_1748 ();
 sg13g2_decap_8 FILLER_2_1755 ();
 sg13g2_decap_8 FILLER_2_1762 ();
 sg13g2_decap_8 FILLER_2_1769 ();
 sg13g2_decap_8 FILLER_2_1776 ();
 sg13g2_decap_8 FILLER_2_1783 ();
 sg13g2_decap_8 FILLER_2_1790 ();
 sg13g2_decap_8 FILLER_2_1797 ();
 sg13g2_decap_8 FILLER_2_1804 ();
 sg13g2_decap_8 FILLER_2_1811 ();
 sg13g2_decap_8 FILLER_2_1818 ();
 sg13g2_decap_8 FILLER_2_1825 ();
 sg13g2_decap_8 FILLER_2_1832 ();
 sg13g2_decap_8 FILLER_2_1839 ();
 sg13g2_decap_8 FILLER_2_1846 ();
 sg13g2_decap_8 FILLER_2_1853 ();
 sg13g2_decap_8 FILLER_2_1860 ();
 sg13g2_decap_8 FILLER_2_1867 ();
 sg13g2_decap_8 FILLER_2_1874 ();
 sg13g2_decap_8 FILLER_2_1881 ();
 sg13g2_decap_8 FILLER_2_1888 ();
 sg13g2_decap_8 FILLER_2_1895 ();
 sg13g2_decap_8 FILLER_2_1902 ();
 sg13g2_decap_8 FILLER_2_1909 ();
 sg13g2_decap_8 FILLER_2_1916 ();
 sg13g2_decap_8 FILLER_2_1923 ();
 sg13g2_decap_8 FILLER_2_1930 ();
 sg13g2_decap_8 FILLER_2_1937 ();
 sg13g2_decap_8 FILLER_2_1944 ();
 sg13g2_decap_8 FILLER_2_1951 ();
 sg13g2_decap_8 FILLER_2_1958 ();
 sg13g2_decap_8 FILLER_2_1965 ();
 sg13g2_decap_8 FILLER_2_1972 ();
 sg13g2_decap_8 FILLER_2_1979 ();
 sg13g2_decap_8 FILLER_2_1986 ();
 sg13g2_decap_8 FILLER_2_1993 ();
 sg13g2_decap_8 FILLER_2_2000 ();
 sg13g2_decap_8 FILLER_2_2007 ();
 sg13g2_decap_8 FILLER_2_2014 ();
 sg13g2_decap_8 FILLER_2_2021 ();
 sg13g2_decap_8 FILLER_2_2028 ();
 sg13g2_decap_8 FILLER_2_2035 ();
 sg13g2_decap_8 FILLER_2_2042 ();
 sg13g2_decap_8 FILLER_2_2049 ();
 sg13g2_decap_8 FILLER_2_2056 ();
 sg13g2_decap_8 FILLER_2_2063 ();
 sg13g2_decap_8 FILLER_2_2070 ();
 sg13g2_decap_8 FILLER_2_2077 ();
 sg13g2_decap_8 FILLER_2_2084 ();
 sg13g2_decap_8 FILLER_2_2091 ();
 sg13g2_decap_8 FILLER_2_2098 ();
 sg13g2_decap_8 FILLER_2_2105 ();
 sg13g2_decap_8 FILLER_2_2112 ();
 sg13g2_decap_8 FILLER_2_2119 ();
 sg13g2_decap_8 FILLER_2_2126 ();
 sg13g2_decap_8 FILLER_2_2133 ();
 sg13g2_decap_8 FILLER_2_2140 ();
 sg13g2_decap_8 FILLER_2_2147 ();
 sg13g2_decap_8 FILLER_2_2154 ();
 sg13g2_decap_8 FILLER_2_2161 ();
 sg13g2_decap_8 FILLER_2_2168 ();
 sg13g2_decap_8 FILLER_2_2175 ();
 sg13g2_decap_8 FILLER_2_2182 ();
 sg13g2_decap_8 FILLER_2_2189 ();
 sg13g2_decap_8 FILLER_2_2196 ();
 sg13g2_decap_8 FILLER_2_2203 ();
 sg13g2_decap_8 FILLER_2_2210 ();
 sg13g2_decap_8 FILLER_2_2217 ();
 sg13g2_decap_8 FILLER_2_2224 ();
 sg13g2_decap_8 FILLER_2_2231 ();
 sg13g2_decap_8 FILLER_2_2238 ();
 sg13g2_decap_8 FILLER_2_2245 ();
 sg13g2_decap_8 FILLER_2_2252 ();
 sg13g2_decap_8 FILLER_2_2259 ();
 sg13g2_decap_8 FILLER_2_2266 ();
 sg13g2_decap_8 FILLER_2_2273 ();
 sg13g2_decap_8 FILLER_2_2280 ();
 sg13g2_decap_8 FILLER_2_2287 ();
 sg13g2_decap_8 FILLER_2_2294 ();
 sg13g2_decap_8 FILLER_2_2301 ();
 sg13g2_decap_8 FILLER_2_2308 ();
 sg13g2_decap_8 FILLER_2_2315 ();
 sg13g2_decap_8 FILLER_2_2322 ();
 sg13g2_decap_8 FILLER_2_2329 ();
 sg13g2_decap_8 FILLER_2_2336 ();
 sg13g2_decap_8 FILLER_2_2343 ();
 sg13g2_decap_8 FILLER_2_2350 ();
 sg13g2_decap_8 FILLER_2_2357 ();
 sg13g2_decap_8 FILLER_2_2364 ();
 sg13g2_decap_8 FILLER_2_2371 ();
 sg13g2_decap_8 FILLER_2_2378 ();
 sg13g2_decap_8 FILLER_2_2385 ();
 sg13g2_decap_8 FILLER_2_2392 ();
 sg13g2_decap_8 FILLER_2_2399 ();
 sg13g2_decap_8 FILLER_2_2406 ();
 sg13g2_decap_8 FILLER_2_2413 ();
 sg13g2_decap_8 FILLER_2_2420 ();
 sg13g2_decap_8 FILLER_2_2427 ();
 sg13g2_decap_8 FILLER_2_2434 ();
 sg13g2_decap_8 FILLER_2_2441 ();
 sg13g2_decap_8 FILLER_2_2448 ();
 sg13g2_decap_8 FILLER_2_2455 ();
 sg13g2_decap_8 FILLER_2_2462 ();
 sg13g2_decap_8 FILLER_2_2469 ();
 sg13g2_decap_8 FILLER_2_2476 ();
 sg13g2_decap_8 FILLER_2_2483 ();
 sg13g2_decap_8 FILLER_2_2490 ();
 sg13g2_decap_8 FILLER_2_2497 ();
 sg13g2_decap_8 FILLER_2_2504 ();
 sg13g2_decap_8 FILLER_2_2511 ();
 sg13g2_decap_8 FILLER_2_2518 ();
 sg13g2_decap_8 FILLER_2_2525 ();
 sg13g2_decap_8 FILLER_2_2532 ();
 sg13g2_decap_8 FILLER_2_2539 ();
 sg13g2_decap_8 FILLER_2_2546 ();
 sg13g2_decap_8 FILLER_2_2553 ();
 sg13g2_decap_8 FILLER_2_2560 ();
 sg13g2_decap_8 FILLER_2_2567 ();
 sg13g2_decap_8 FILLER_2_2574 ();
 sg13g2_decap_8 FILLER_2_2581 ();
 sg13g2_decap_8 FILLER_2_2588 ();
 sg13g2_decap_8 FILLER_2_2595 ();
 sg13g2_decap_8 FILLER_2_2602 ();
 sg13g2_decap_8 FILLER_2_2609 ();
 sg13g2_decap_8 FILLER_2_2616 ();
 sg13g2_decap_8 FILLER_2_2623 ();
 sg13g2_decap_8 FILLER_2_2630 ();
 sg13g2_decap_8 FILLER_2_2637 ();
 sg13g2_decap_8 FILLER_2_2644 ();
 sg13g2_decap_8 FILLER_2_2651 ();
 sg13g2_decap_8 FILLER_2_2658 ();
 sg13g2_decap_4 FILLER_2_2665 ();
 sg13g2_fill_1 FILLER_2_2669 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_4 FILLER_3_189 ();
 sg13g2_fill_1 FILLER_3_193 ();
 sg13g2_fill_2 FILLER_3_220 ();
 sg13g2_fill_1 FILLER_3_222 ();
 sg13g2_decap_8 FILLER_3_228 ();
 sg13g2_decap_8 FILLER_3_235 ();
 sg13g2_decap_8 FILLER_3_242 ();
 sg13g2_fill_1 FILLER_3_249 ();
 sg13g2_decap_8 FILLER_3_254 ();
 sg13g2_decap_4 FILLER_3_261 ();
 sg13g2_fill_2 FILLER_3_265 ();
 sg13g2_decap_4 FILLER_3_272 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_4 FILLER_3_287 ();
 sg13g2_fill_1 FILLER_3_291 ();
 sg13g2_decap_8 FILLER_3_318 ();
 sg13g2_decap_8 FILLER_3_325 ();
 sg13g2_decap_8 FILLER_3_332 ();
 sg13g2_decap_8 FILLER_3_339 ();
 sg13g2_decap_8 FILLER_3_346 ();
 sg13g2_decap_8 FILLER_3_353 ();
 sg13g2_decap_8 FILLER_3_360 ();
 sg13g2_decap_8 FILLER_3_367 ();
 sg13g2_decap_8 FILLER_3_374 ();
 sg13g2_decap_8 FILLER_3_381 ();
 sg13g2_decap_8 FILLER_3_388 ();
 sg13g2_fill_2 FILLER_3_395 ();
 sg13g2_fill_2 FILLER_3_401 ();
 sg13g2_fill_2 FILLER_3_440 ();
 sg13g2_fill_1 FILLER_3_442 ();
 sg13g2_decap_8 FILLER_3_447 ();
 sg13g2_decap_4 FILLER_3_454 ();
 sg13g2_fill_1 FILLER_3_458 ();
 sg13g2_decap_8 FILLER_3_468 ();
 sg13g2_decap_8 FILLER_3_475 ();
 sg13g2_decap_8 FILLER_3_482 ();
 sg13g2_decap_4 FILLER_3_489 ();
 sg13g2_fill_2 FILLER_3_493 ();
 sg13g2_decap_8 FILLER_3_499 ();
 sg13g2_decap_4 FILLER_3_506 ();
 sg13g2_fill_1 FILLER_3_510 ();
 sg13g2_fill_1 FILLER_3_534 ();
 sg13g2_fill_1 FILLER_3_538 ();
 sg13g2_decap_8 FILLER_3_547 ();
 sg13g2_decap_4 FILLER_3_554 ();
 sg13g2_fill_2 FILLER_3_558 ();
 sg13g2_decap_4 FILLER_3_568 ();
 sg13g2_decap_8 FILLER_3_576 ();
 sg13g2_fill_2 FILLER_3_583 ();
 sg13g2_decap_4 FILLER_3_593 ();
 sg13g2_decap_4 FILLER_3_612 ();
 sg13g2_decap_8 FILLER_3_619 ();
 sg13g2_decap_8 FILLER_3_626 ();
 sg13g2_decap_8 FILLER_3_633 ();
 sg13g2_decap_8 FILLER_3_640 ();
 sg13g2_decap_8 FILLER_3_647 ();
 sg13g2_decap_8 FILLER_3_654 ();
 sg13g2_fill_1 FILLER_3_661 ();
 sg13g2_decap_8 FILLER_3_667 ();
 sg13g2_decap_8 FILLER_3_674 ();
 sg13g2_fill_2 FILLER_3_681 ();
 sg13g2_fill_1 FILLER_3_683 ();
 sg13g2_decap_4 FILLER_3_693 ();
 sg13g2_fill_1 FILLER_3_697 ();
 sg13g2_fill_1 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_719 ();
 sg13g2_decap_8 FILLER_3_726 ();
 sg13g2_fill_2 FILLER_3_733 ();
 sg13g2_fill_1 FILLER_3_735 ();
 sg13g2_fill_2 FILLER_3_741 ();
 sg13g2_fill_1 FILLER_3_743 ();
 sg13g2_decap_8 FILLER_3_758 ();
 sg13g2_decap_8 FILLER_3_765 ();
 sg13g2_decap_8 FILLER_3_772 ();
 sg13g2_fill_2 FILLER_3_779 ();
 sg13g2_decap_8 FILLER_3_790 ();
 sg13g2_fill_2 FILLER_3_816 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_4 FILLER_3_833 ();
 sg13g2_fill_2 FILLER_3_837 ();
 sg13g2_decap_8 FILLER_3_843 ();
 sg13g2_decap_8 FILLER_3_850 ();
 sg13g2_decap_8 FILLER_3_857 ();
 sg13g2_decap_4 FILLER_3_864 ();
 sg13g2_fill_1 FILLER_3_868 ();
 sg13g2_decap_8 FILLER_3_873 ();
 sg13g2_decap_8 FILLER_3_880 ();
 sg13g2_decap_4 FILLER_3_887 ();
 sg13g2_fill_2 FILLER_3_901 ();
 sg13g2_decap_8 FILLER_3_918 ();
 sg13g2_decap_8 FILLER_3_925 ();
 sg13g2_decap_8 FILLER_3_932 ();
 sg13g2_decap_4 FILLER_3_939 ();
 sg13g2_fill_1 FILLER_3_943 ();
 sg13g2_fill_1 FILLER_3_952 ();
 sg13g2_decap_4 FILLER_3_963 ();
 sg13g2_fill_2 FILLER_3_967 ();
 sg13g2_decap_8 FILLER_3_980 ();
 sg13g2_decap_8 FILLER_3_987 ();
 sg13g2_decap_8 FILLER_3_994 ();
 sg13g2_fill_1 FILLER_3_1001 ();
 sg13g2_decap_8 FILLER_3_1010 ();
 sg13g2_decap_8 FILLER_3_1017 ();
 sg13g2_decap_8 FILLER_3_1024 ();
 sg13g2_decap_8 FILLER_3_1031 ();
 sg13g2_decap_4 FILLER_3_1038 ();
 sg13g2_fill_1 FILLER_3_1042 ();
 sg13g2_fill_1 FILLER_3_1055 ();
 sg13g2_decap_8 FILLER_3_1069 ();
 sg13g2_fill_1 FILLER_3_1076 ();
 sg13g2_fill_2 FILLER_3_1081 ();
 sg13g2_fill_1 FILLER_3_1083 ();
 sg13g2_fill_2 FILLER_3_1099 ();
 sg13g2_decap_8 FILLER_3_1105 ();
 sg13g2_decap_8 FILLER_3_1112 ();
 sg13g2_decap_8 FILLER_3_1119 ();
 sg13g2_decap_8 FILLER_3_1126 ();
 sg13g2_decap_8 FILLER_3_1133 ();
 sg13g2_fill_1 FILLER_3_1140 ();
 sg13g2_decap_8 FILLER_3_1145 ();
 sg13g2_decap_8 FILLER_3_1152 ();
 sg13g2_decap_8 FILLER_3_1159 ();
 sg13g2_decap_8 FILLER_3_1166 ();
 sg13g2_decap_8 FILLER_3_1173 ();
 sg13g2_decap_8 FILLER_3_1180 ();
 sg13g2_decap_8 FILLER_3_1187 ();
 sg13g2_fill_1 FILLER_3_1194 ();
 sg13g2_fill_2 FILLER_3_1210 ();
 sg13g2_decap_8 FILLER_3_1224 ();
 sg13g2_decap_8 FILLER_3_1231 ();
 sg13g2_decap_8 FILLER_3_1238 ();
 sg13g2_decap_8 FILLER_3_1245 ();
 sg13g2_fill_1 FILLER_3_1252 ();
 sg13g2_fill_1 FILLER_3_1260 ();
 sg13g2_decap_4 FILLER_3_1278 ();
 sg13g2_fill_2 FILLER_3_1286 ();
 sg13g2_decap_8 FILLER_3_1301 ();
 sg13g2_decap_8 FILLER_3_1308 ();
 sg13g2_fill_2 FILLER_3_1315 ();
 sg13g2_decap_8 FILLER_3_1352 ();
 sg13g2_decap_8 FILLER_3_1359 ();
 sg13g2_fill_1 FILLER_3_1366 ();
 sg13g2_decap_8 FILLER_3_1383 ();
 sg13g2_decap_8 FILLER_3_1390 ();
 sg13g2_decap_8 FILLER_3_1397 ();
 sg13g2_decap_4 FILLER_3_1404 ();
 sg13g2_fill_2 FILLER_3_1408 ();
 sg13g2_decap_8 FILLER_3_1416 ();
 sg13g2_decap_4 FILLER_3_1423 ();
 sg13g2_decap_4 FILLER_3_1431 ();
 sg13g2_fill_2 FILLER_3_1439 ();
 sg13g2_decap_4 FILLER_3_1446 ();
 sg13g2_fill_1 FILLER_3_1450 ();
 sg13g2_decap_8 FILLER_3_1464 ();
 sg13g2_decap_8 FILLER_3_1471 ();
 sg13g2_decap_8 FILLER_3_1478 ();
 sg13g2_decap_8 FILLER_3_1485 ();
 sg13g2_decap_8 FILLER_3_1492 ();
 sg13g2_decap_8 FILLER_3_1499 ();
 sg13g2_decap_8 FILLER_3_1506 ();
 sg13g2_decap_8 FILLER_3_1513 ();
 sg13g2_decap_8 FILLER_3_1520 ();
 sg13g2_decap_8 FILLER_3_1527 ();
 sg13g2_decap_4 FILLER_3_1534 ();
 sg13g2_fill_2 FILLER_3_1538 ();
 sg13g2_decap_8 FILLER_3_1557 ();
 sg13g2_decap_8 FILLER_3_1564 ();
 sg13g2_decap_8 FILLER_3_1571 ();
 sg13g2_decap_8 FILLER_3_1578 ();
 sg13g2_decap_8 FILLER_3_1585 ();
 sg13g2_fill_2 FILLER_3_1617 ();
 sg13g2_fill_1 FILLER_3_1619 ();
 sg13g2_decap_8 FILLER_3_1624 ();
 sg13g2_decap_8 FILLER_3_1631 ();
 sg13g2_decap_8 FILLER_3_1638 ();
 sg13g2_decap_8 FILLER_3_1645 ();
 sg13g2_decap_8 FILLER_3_1652 ();
 sg13g2_decap_8 FILLER_3_1659 ();
 sg13g2_decap_8 FILLER_3_1666 ();
 sg13g2_decap_8 FILLER_3_1673 ();
 sg13g2_decap_8 FILLER_3_1680 ();
 sg13g2_decap_8 FILLER_3_1687 ();
 sg13g2_fill_1 FILLER_3_1694 ();
 sg13g2_decap_8 FILLER_3_1703 ();
 sg13g2_decap_8 FILLER_3_1710 ();
 sg13g2_decap_8 FILLER_3_1717 ();
 sg13g2_decap_8 FILLER_3_1724 ();
 sg13g2_decap_8 FILLER_3_1731 ();
 sg13g2_decap_8 FILLER_3_1738 ();
 sg13g2_decap_8 FILLER_3_1745 ();
 sg13g2_fill_2 FILLER_3_1752 ();
 sg13g2_decap_8 FILLER_3_1767 ();
 sg13g2_decap_8 FILLER_3_1774 ();
 sg13g2_decap_8 FILLER_3_1781 ();
 sg13g2_decap_8 FILLER_3_1788 ();
 sg13g2_decap_8 FILLER_3_1795 ();
 sg13g2_decap_8 FILLER_3_1802 ();
 sg13g2_decap_8 FILLER_3_1809 ();
 sg13g2_decap_8 FILLER_3_1816 ();
 sg13g2_decap_8 FILLER_3_1823 ();
 sg13g2_decap_8 FILLER_3_1830 ();
 sg13g2_decap_8 FILLER_3_1837 ();
 sg13g2_decap_8 FILLER_3_1844 ();
 sg13g2_decap_8 FILLER_3_1851 ();
 sg13g2_decap_8 FILLER_3_1858 ();
 sg13g2_decap_8 FILLER_3_1865 ();
 sg13g2_decap_8 FILLER_3_1872 ();
 sg13g2_decap_8 FILLER_3_1879 ();
 sg13g2_decap_8 FILLER_3_1886 ();
 sg13g2_decap_8 FILLER_3_1893 ();
 sg13g2_decap_8 FILLER_3_1900 ();
 sg13g2_decap_8 FILLER_3_1907 ();
 sg13g2_decap_8 FILLER_3_1914 ();
 sg13g2_decap_8 FILLER_3_1921 ();
 sg13g2_decap_8 FILLER_3_1928 ();
 sg13g2_decap_8 FILLER_3_1935 ();
 sg13g2_decap_8 FILLER_3_1942 ();
 sg13g2_decap_8 FILLER_3_1949 ();
 sg13g2_decap_8 FILLER_3_1956 ();
 sg13g2_decap_8 FILLER_3_1963 ();
 sg13g2_decap_8 FILLER_3_1970 ();
 sg13g2_decap_8 FILLER_3_1977 ();
 sg13g2_decap_8 FILLER_3_1984 ();
 sg13g2_decap_8 FILLER_3_1991 ();
 sg13g2_decap_8 FILLER_3_1998 ();
 sg13g2_decap_8 FILLER_3_2005 ();
 sg13g2_decap_8 FILLER_3_2012 ();
 sg13g2_decap_8 FILLER_3_2019 ();
 sg13g2_decap_8 FILLER_3_2026 ();
 sg13g2_decap_8 FILLER_3_2033 ();
 sg13g2_decap_8 FILLER_3_2040 ();
 sg13g2_decap_8 FILLER_3_2047 ();
 sg13g2_decap_8 FILLER_3_2054 ();
 sg13g2_decap_8 FILLER_3_2061 ();
 sg13g2_decap_8 FILLER_3_2068 ();
 sg13g2_decap_8 FILLER_3_2075 ();
 sg13g2_decap_8 FILLER_3_2082 ();
 sg13g2_decap_8 FILLER_3_2089 ();
 sg13g2_decap_8 FILLER_3_2096 ();
 sg13g2_decap_8 FILLER_3_2103 ();
 sg13g2_decap_8 FILLER_3_2110 ();
 sg13g2_decap_8 FILLER_3_2117 ();
 sg13g2_decap_8 FILLER_3_2124 ();
 sg13g2_decap_8 FILLER_3_2131 ();
 sg13g2_decap_8 FILLER_3_2138 ();
 sg13g2_decap_8 FILLER_3_2145 ();
 sg13g2_decap_8 FILLER_3_2152 ();
 sg13g2_decap_8 FILLER_3_2159 ();
 sg13g2_decap_8 FILLER_3_2166 ();
 sg13g2_decap_8 FILLER_3_2173 ();
 sg13g2_decap_8 FILLER_3_2180 ();
 sg13g2_decap_8 FILLER_3_2187 ();
 sg13g2_decap_8 FILLER_3_2194 ();
 sg13g2_decap_8 FILLER_3_2201 ();
 sg13g2_decap_8 FILLER_3_2208 ();
 sg13g2_decap_8 FILLER_3_2215 ();
 sg13g2_decap_8 FILLER_3_2222 ();
 sg13g2_decap_8 FILLER_3_2229 ();
 sg13g2_decap_8 FILLER_3_2236 ();
 sg13g2_decap_8 FILLER_3_2243 ();
 sg13g2_decap_8 FILLER_3_2250 ();
 sg13g2_decap_8 FILLER_3_2257 ();
 sg13g2_decap_8 FILLER_3_2264 ();
 sg13g2_decap_8 FILLER_3_2271 ();
 sg13g2_decap_8 FILLER_3_2278 ();
 sg13g2_decap_8 FILLER_3_2285 ();
 sg13g2_decap_8 FILLER_3_2292 ();
 sg13g2_decap_8 FILLER_3_2299 ();
 sg13g2_decap_8 FILLER_3_2306 ();
 sg13g2_decap_8 FILLER_3_2313 ();
 sg13g2_decap_8 FILLER_3_2320 ();
 sg13g2_decap_8 FILLER_3_2327 ();
 sg13g2_decap_8 FILLER_3_2334 ();
 sg13g2_decap_8 FILLER_3_2341 ();
 sg13g2_decap_8 FILLER_3_2348 ();
 sg13g2_decap_8 FILLER_3_2355 ();
 sg13g2_decap_8 FILLER_3_2362 ();
 sg13g2_decap_8 FILLER_3_2369 ();
 sg13g2_decap_8 FILLER_3_2376 ();
 sg13g2_decap_8 FILLER_3_2383 ();
 sg13g2_decap_8 FILLER_3_2390 ();
 sg13g2_decap_8 FILLER_3_2397 ();
 sg13g2_decap_8 FILLER_3_2404 ();
 sg13g2_decap_8 FILLER_3_2411 ();
 sg13g2_decap_8 FILLER_3_2418 ();
 sg13g2_decap_8 FILLER_3_2425 ();
 sg13g2_decap_8 FILLER_3_2432 ();
 sg13g2_decap_8 FILLER_3_2439 ();
 sg13g2_decap_8 FILLER_3_2446 ();
 sg13g2_decap_8 FILLER_3_2453 ();
 sg13g2_decap_8 FILLER_3_2460 ();
 sg13g2_decap_8 FILLER_3_2467 ();
 sg13g2_decap_8 FILLER_3_2474 ();
 sg13g2_decap_8 FILLER_3_2481 ();
 sg13g2_decap_8 FILLER_3_2488 ();
 sg13g2_decap_8 FILLER_3_2495 ();
 sg13g2_decap_8 FILLER_3_2502 ();
 sg13g2_decap_8 FILLER_3_2509 ();
 sg13g2_decap_8 FILLER_3_2516 ();
 sg13g2_decap_8 FILLER_3_2523 ();
 sg13g2_decap_8 FILLER_3_2530 ();
 sg13g2_decap_8 FILLER_3_2537 ();
 sg13g2_decap_8 FILLER_3_2544 ();
 sg13g2_decap_8 FILLER_3_2551 ();
 sg13g2_decap_8 FILLER_3_2558 ();
 sg13g2_decap_8 FILLER_3_2565 ();
 sg13g2_decap_8 FILLER_3_2572 ();
 sg13g2_decap_8 FILLER_3_2579 ();
 sg13g2_decap_8 FILLER_3_2586 ();
 sg13g2_decap_8 FILLER_3_2593 ();
 sg13g2_decap_8 FILLER_3_2600 ();
 sg13g2_decap_8 FILLER_3_2607 ();
 sg13g2_decap_8 FILLER_3_2614 ();
 sg13g2_decap_8 FILLER_3_2621 ();
 sg13g2_decap_8 FILLER_3_2628 ();
 sg13g2_decap_8 FILLER_3_2635 ();
 sg13g2_decap_8 FILLER_3_2642 ();
 sg13g2_decap_8 FILLER_3_2649 ();
 sg13g2_decap_8 FILLER_3_2656 ();
 sg13g2_decap_8 FILLER_3_2663 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_4 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_204 ();
 sg13g2_decap_8 FILLER_4_211 ();
 sg13g2_decap_8 FILLER_4_218 ();
 sg13g2_decap_8 FILLER_4_229 ();
 sg13g2_decap_8 FILLER_4_236 ();
 sg13g2_decap_8 FILLER_4_243 ();
 sg13g2_decap_8 FILLER_4_250 ();
 sg13g2_decap_8 FILLER_4_257 ();
 sg13g2_decap_8 FILLER_4_264 ();
 sg13g2_decap_8 FILLER_4_271 ();
 sg13g2_decap_8 FILLER_4_278 ();
 sg13g2_decap_8 FILLER_4_285 ();
 sg13g2_decap_8 FILLER_4_292 ();
 sg13g2_decap_8 FILLER_4_303 ();
 sg13g2_decap_8 FILLER_4_310 ();
 sg13g2_decap_8 FILLER_4_317 ();
 sg13g2_decap_8 FILLER_4_324 ();
 sg13g2_decap_8 FILLER_4_331 ();
 sg13g2_decap_8 FILLER_4_338 ();
 sg13g2_decap_8 FILLER_4_345 ();
 sg13g2_decap_8 FILLER_4_352 ();
 sg13g2_decap_8 FILLER_4_359 ();
 sg13g2_decap_8 FILLER_4_366 ();
 sg13g2_decap_8 FILLER_4_373 ();
 sg13g2_decap_8 FILLER_4_380 ();
 sg13g2_decap_8 FILLER_4_387 ();
 sg13g2_decap_8 FILLER_4_394 ();
 sg13g2_decap_8 FILLER_4_401 ();
 sg13g2_decap_8 FILLER_4_408 ();
 sg13g2_decap_4 FILLER_4_415 ();
 sg13g2_decap_8 FILLER_4_433 ();
 sg13g2_fill_2 FILLER_4_440 ();
 sg13g2_decap_8 FILLER_4_447 ();
 sg13g2_decap_8 FILLER_4_454 ();
 sg13g2_decap_8 FILLER_4_461 ();
 sg13g2_decap_8 FILLER_4_468 ();
 sg13g2_decap_8 FILLER_4_475 ();
 sg13g2_decap_8 FILLER_4_482 ();
 sg13g2_decap_8 FILLER_4_489 ();
 sg13g2_fill_2 FILLER_4_496 ();
 sg13g2_fill_1 FILLER_4_498 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_fill_2 FILLER_4_511 ();
 sg13g2_fill_1 FILLER_4_513 ();
 sg13g2_decap_8 FILLER_4_517 ();
 sg13g2_decap_8 FILLER_4_524 ();
 sg13g2_decap_8 FILLER_4_531 ();
 sg13g2_decap_8 FILLER_4_538 ();
 sg13g2_decap_8 FILLER_4_545 ();
 sg13g2_decap_8 FILLER_4_552 ();
 sg13g2_decap_8 FILLER_4_559 ();
 sg13g2_decap_8 FILLER_4_566 ();
 sg13g2_decap_8 FILLER_4_573 ();
 sg13g2_decap_4 FILLER_4_580 ();
 sg13g2_fill_1 FILLER_4_584 ();
 sg13g2_decap_4 FILLER_4_610 ();
 sg13g2_fill_2 FILLER_4_614 ();
 sg13g2_decap_8 FILLER_4_621 ();
 sg13g2_decap_8 FILLER_4_628 ();
 sg13g2_decap_4 FILLER_4_635 ();
 sg13g2_fill_2 FILLER_4_639 ();
 sg13g2_decap_8 FILLER_4_645 ();
 sg13g2_decap_8 FILLER_4_652 ();
 sg13g2_decap_8 FILLER_4_659 ();
 sg13g2_decap_8 FILLER_4_666 ();
 sg13g2_decap_8 FILLER_4_673 ();
 sg13g2_decap_4 FILLER_4_680 ();
 sg13g2_decap_8 FILLER_4_687 ();
 sg13g2_decap_8 FILLER_4_694 ();
 sg13g2_decap_4 FILLER_4_701 ();
 sg13g2_fill_1 FILLER_4_705 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_4 FILLER_4_742 ();
 sg13g2_fill_1 FILLER_4_746 ();
 sg13g2_decap_8 FILLER_4_750 ();
 sg13g2_decap_8 FILLER_4_757 ();
 sg13g2_decap_8 FILLER_4_764 ();
 sg13g2_decap_8 FILLER_4_771 ();
 sg13g2_fill_2 FILLER_4_778 ();
 sg13g2_fill_1 FILLER_4_780 ();
 sg13g2_decap_8 FILLER_4_786 ();
 sg13g2_decap_8 FILLER_4_793 ();
 sg13g2_decap_8 FILLER_4_800 ();
 sg13g2_fill_1 FILLER_4_807 ();
 sg13g2_decap_8 FILLER_4_813 ();
 sg13g2_decap_8 FILLER_4_820 ();
 sg13g2_decap_8 FILLER_4_827 ();
 sg13g2_decap_8 FILLER_4_834 ();
 sg13g2_decap_8 FILLER_4_841 ();
 sg13g2_decap_8 FILLER_4_848 ();
 sg13g2_decap_8 FILLER_4_855 ();
 sg13g2_decap_4 FILLER_4_862 ();
 sg13g2_decap_8 FILLER_4_878 ();
 sg13g2_decap_8 FILLER_4_885 ();
 sg13g2_decap_4 FILLER_4_892 ();
 sg13g2_fill_1 FILLER_4_896 ();
 sg13g2_decap_8 FILLER_4_913 ();
 sg13g2_decap_8 FILLER_4_920 ();
 sg13g2_decap_8 FILLER_4_927 ();
 sg13g2_decap_8 FILLER_4_934 ();
 sg13g2_decap_8 FILLER_4_941 ();
 sg13g2_decap_8 FILLER_4_948 ();
 sg13g2_decap_8 FILLER_4_955 ();
 sg13g2_decap_8 FILLER_4_962 ();
 sg13g2_decap_8 FILLER_4_969 ();
 sg13g2_decap_8 FILLER_4_976 ();
 sg13g2_decap_8 FILLER_4_983 ();
 sg13g2_decap_8 FILLER_4_990 ();
 sg13g2_decap_8 FILLER_4_997 ();
 sg13g2_decap_4 FILLER_4_1004 ();
 sg13g2_fill_1 FILLER_4_1008 ();
 sg13g2_decap_8 FILLER_4_1014 ();
 sg13g2_decap_8 FILLER_4_1021 ();
 sg13g2_decap_8 FILLER_4_1028 ();
 sg13g2_decap_8 FILLER_4_1035 ();
 sg13g2_decap_8 FILLER_4_1042 ();
 sg13g2_fill_2 FILLER_4_1049 ();
 sg13g2_fill_1 FILLER_4_1051 ();
 sg13g2_decap_8 FILLER_4_1056 ();
 sg13g2_decap_8 FILLER_4_1063 ();
 sg13g2_decap_8 FILLER_4_1070 ();
 sg13g2_decap_8 FILLER_4_1077 ();
 sg13g2_fill_2 FILLER_4_1094 ();
 sg13g2_fill_1 FILLER_4_1096 ();
 sg13g2_decap_8 FILLER_4_1112 ();
 sg13g2_decap_8 FILLER_4_1119 ();
 sg13g2_decap_8 FILLER_4_1126 ();
 sg13g2_decap_8 FILLER_4_1133 ();
 sg13g2_decap_8 FILLER_4_1140 ();
 sg13g2_decap_8 FILLER_4_1147 ();
 sg13g2_decap_8 FILLER_4_1154 ();
 sg13g2_decap_8 FILLER_4_1161 ();
 sg13g2_fill_2 FILLER_4_1168 ();
 sg13g2_fill_1 FILLER_4_1170 ();
 sg13g2_decap_8 FILLER_4_1176 ();
 sg13g2_fill_2 FILLER_4_1183 ();
 sg13g2_decap_8 FILLER_4_1189 ();
 sg13g2_decap_8 FILLER_4_1196 ();
 sg13g2_decap_4 FILLER_4_1203 ();
 sg13g2_fill_2 FILLER_4_1207 ();
 sg13g2_fill_1 FILLER_4_1220 ();
 sg13g2_decap_8 FILLER_4_1236 ();
 sg13g2_decap_8 FILLER_4_1243 ();
 sg13g2_decap_8 FILLER_4_1250 ();
 sg13g2_decap_8 FILLER_4_1257 ();
 sg13g2_decap_8 FILLER_4_1264 ();
 sg13g2_decap_8 FILLER_4_1271 ();
 sg13g2_decap_8 FILLER_4_1278 ();
 sg13g2_decap_4 FILLER_4_1285 ();
 sg13g2_fill_2 FILLER_4_1289 ();
 sg13g2_decap_8 FILLER_4_1296 ();
 sg13g2_decap_8 FILLER_4_1303 ();
 sg13g2_fill_2 FILLER_4_1310 ();
 sg13g2_fill_1 FILLER_4_1312 ();
 sg13g2_decap_8 FILLER_4_1318 ();
 sg13g2_decap_8 FILLER_4_1325 ();
 sg13g2_decap_8 FILLER_4_1332 ();
 sg13g2_decap_8 FILLER_4_1339 ();
 sg13g2_decap_8 FILLER_4_1346 ();
 sg13g2_decap_8 FILLER_4_1353 ();
 sg13g2_fill_2 FILLER_4_1360 ();
 sg13g2_fill_2 FILLER_4_1367 ();
 sg13g2_fill_1 FILLER_4_1369 ();
 sg13g2_decap_8 FILLER_4_1373 ();
 sg13g2_decap_8 FILLER_4_1380 ();
 sg13g2_decap_8 FILLER_4_1387 ();
 sg13g2_decap_8 FILLER_4_1394 ();
 sg13g2_decap_8 FILLER_4_1401 ();
 sg13g2_decap_8 FILLER_4_1408 ();
 sg13g2_decap_8 FILLER_4_1415 ();
 sg13g2_decap_8 FILLER_4_1422 ();
 sg13g2_decap_8 FILLER_4_1429 ();
 sg13g2_fill_1 FILLER_4_1436 ();
 sg13g2_decap_8 FILLER_4_1442 ();
 sg13g2_decap_8 FILLER_4_1449 ();
 sg13g2_decap_8 FILLER_4_1456 ();
 sg13g2_decap_8 FILLER_4_1463 ();
 sg13g2_decap_8 FILLER_4_1470 ();
 sg13g2_decap_8 FILLER_4_1477 ();
 sg13g2_decap_8 FILLER_4_1484 ();
 sg13g2_decap_8 FILLER_4_1491 ();
 sg13g2_decap_8 FILLER_4_1498 ();
 sg13g2_decap_8 FILLER_4_1505 ();
 sg13g2_fill_2 FILLER_4_1512 ();
 sg13g2_decap_8 FILLER_4_1525 ();
 sg13g2_decap_8 FILLER_4_1532 ();
 sg13g2_decap_4 FILLER_4_1539 ();
 sg13g2_decap_8 FILLER_4_1551 ();
 sg13g2_fill_1 FILLER_4_1558 ();
 sg13g2_decap_8 FILLER_4_1564 ();
 sg13g2_decap_8 FILLER_4_1571 ();
 sg13g2_decap_8 FILLER_4_1578 ();
 sg13g2_decap_8 FILLER_4_1585 ();
 sg13g2_decap_8 FILLER_4_1597 ();
 sg13g2_decap_8 FILLER_4_1604 ();
 sg13g2_decap_8 FILLER_4_1611 ();
 sg13g2_decap_8 FILLER_4_1618 ();
 sg13g2_decap_8 FILLER_4_1625 ();
 sg13g2_decap_8 FILLER_4_1632 ();
 sg13g2_decap_8 FILLER_4_1639 ();
 sg13g2_decap_8 FILLER_4_1646 ();
 sg13g2_decap_8 FILLER_4_1653 ();
 sg13g2_decap_8 FILLER_4_1660 ();
 sg13g2_decap_8 FILLER_4_1667 ();
 sg13g2_decap_8 FILLER_4_1674 ();
 sg13g2_decap_8 FILLER_4_1681 ();
 sg13g2_decap_8 FILLER_4_1688 ();
 sg13g2_decap_8 FILLER_4_1695 ();
 sg13g2_decap_8 FILLER_4_1702 ();
 sg13g2_decap_8 FILLER_4_1709 ();
 sg13g2_decap_8 FILLER_4_1716 ();
 sg13g2_decap_8 FILLER_4_1723 ();
 sg13g2_decap_8 FILLER_4_1730 ();
 sg13g2_decap_8 FILLER_4_1737 ();
 sg13g2_decap_8 FILLER_4_1744 ();
 sg13g2_decap_8 FILLER_4_1751 ();
 sg13g2_fill_1 FILLER_4_1758 ();
 sg13g2_decap_8 FILLER_4_1767 ();
 sg13g2_decap_8 FILLER_4_1774 ();
 sg13g2_decap_8 FILLER_4_1781 ();
 sg13g2_decap_8 FILLER_4_1788 ();
 sg13g2_decap_8 FILLER_4_1795 ();
 sg13g2_decap_8 FILLER_4_1802 ();
 sg13g2_decap_8 FILLER_4_1809 ();
 sg13g2_decap_8 FILLER_4_1816 ();
 sg13g2_decap_8 FILLER_4_1823 ();
 sg13g2_decap_8 FILLER_4_1830 ();
 sg13g2_decap_8 FILLER_4_1837 ();
 sg13g2_decap_8 FILLER_4_1844 ();
 sg13g2_decap_8 FILLER_4_1851 ();
 sg13g2_decap_8 FILLER_4_1858 ();
 sg13g2_decap_8 FILLER_4_1865 ();
 sg13g2_decap_8 FILLER_4_1872 ();
 sg13g2_decap_8 FILLER_4_1879 ();
 sg13g2_decap_8 FILLER_4_1886 ();
 sg13g2_decap_8 FILLER_4_1893 ();
 sg13g2_decap_8 FILLER_4_1900 ();
 sg13g2_decap_8 FILLER_4_1907 ();
 sg13g2_decap_8 FILLER_4_1914 ();
 sg13g2_decap_8 FILLER_4_1921 ();
 sg13g2_decap_8 FILLER_4_1928 ();
 sg13g2_decap_8 FILLER_4_1935 ();
 sg13g2_decap_8 FILLER_4_1942 ();
 sg13g2_decap_8 FILLER_4_1949 ();
 sg13g2_decap_8 FILLER_4_1956 ();
 sg13g2_decap_8 FILLER_4_1963 ();
 sg13g2_decap_8 FILLER_4_1970 ();
 sg13g2_decap_8 FILLER_4_1977 ();
 sg13g2_decap_8 FILLER_4_1984 ();
 sg13g2_decap_8 FILLER_4_1991 ();
 sg13g2_decap_8 FILLER_4_1998 ();
 sg13g2_decap_8 FILLER_4_2005 ();
 sg13g2_decap_8 FILLER_4_2012 ();
 sg13g2_decap_8 FILLER_4_2019 ();
 sg13g2_decap_8 FILLER_4_2026 ();
 sg13g2_decap_8 FILLER_4_2033 ();
 sg13g2_decap_8 FILLER_4_2040 ();
 sg13g2_decap_8 FILLER_4_2047 ();
 sg13g2_decap_8 FILLER_4_2054 ();
 sg13g2_decap_8 FILLER_4_2061 ();
 sg13g2_decap_8 FILLER_4_2068 ();
 sg13g2_decap_8 FILLER_4_2075 ();
 sg13g2_decap_8 FILLER_4_2082 ();
 sg13g2_decap_8 FILLER_4_2089 ();
 sg13g2_decap_8 FILLER_4_2096 ();
 sg13g2_decap_8 FILLER_4_2103 ();
 sg13g2_decap_8 FILLER_4_2110 ();
 sg13g2_decap_8 FILLER_4_2117 ();
 sg13g2_decap_8 FILLER_4_2124 ();
 sg13g2_decap_8 FILLER_4_2131 ();
 sg13g2_decap_8 FILLER_4_2138 ();
 sg13g2_decap_8 FILLER_4_2145 ();
 sg13g2_decap_8 FILLER_4_2152 ();
 sg13g2_decap_8 FILLER_4_2159 ();
 sg13g2_decap_8 FILLER_4_2166 ();
 sg13g2_decap_8 FILLER_4_2173 ();
 sg13g2_decap_8 FILLER_4_2180 ();
 sg13g2_decap_8 FILLER_4_2187 ();
 sg13g2_decap_8 FILLER_4_2194 ();
 sg13g2_decap_8 FILLER_4_2201 ();
 sg13g2_decap_8 FILLER_4_2208 ();
 sg13g2_decap_8 FILLER_4_2215 ();
 sg13g2_decap_8 FILLER_4_2222 ();
 sg13g2_decap_8 FILLER_4_2229 ();
 sg13g2_decap_8 FILLER_4_2236 ();
 sg13g2_decap_8 FILLER_4_2243 ();
 sg13g2_decap_8 FILLER_4_2250 ();
 sg13g2_decap_8 FILLER_4_2257 ();
 sg13g2_decap_8 FILLER_4_2264 ();
 sg13g2_decap_8 FILLER_4_2271 ();
 sg13g2_decap_8 FILLER_4_2278 ();
 sg13g2_decap_8 FILLER_4_2285 ();
 sg13g2_decap_8 FILLER_4_2292 ();
 sg13g2_decap_8 FILLER_4_2299 ();
 sg13g2_decap_8 FILLER_4_2306 ();
 sg13g2_decap_8 FILLER_4_2313 ();
 sg13g2_decap_8 FILLER_4_2320 ();
 sg13g2_decap_8 FILLER_4_2327 ();
 sg13g2_decap_8 FILLER_4_2334 ();
 sg13g2_decap_8 FILLER_4_2341 ();
 sg13g2_decap_8 FILLER_4_2348 ();
 sg13g2_decap_8 FILLER_4_2355 ();
 sg13g2_decap_8 FILLER_4_2362 ();
 sg13g2_decap_8 FILLER_4_2369 ();
 sg13g2_decap_8 FILLER_4_2376 ();
 sg13g2_decap_8 FILLER_4_2383 ();
 sg13g2_decap_8 FILLER_4_2390 ();
 sg13g2_decap_8 FILLER_4_2397 ();
 sg13g2_decap_8 FILLER_4_2404 ();
 sg13g2_decap_8 FILLER_4_2411 ();
 sg13g2_decap_8 FILLER_4_2418 ();
 sg13g2_decap_8 FILLER_4_2425 ();
 sg13g2_decap_8 FILLER_4_2432 ();
 sg13g2_decap_8 FILLER_4_2439 ();
 sg13g2_decap_8 FILLER_4_2446 ();
 sg13g2_decap_8 FILLER_4_2453 ();
 sg13g2_decap_8 FILLER_4_2460 ();
 sg13g2_decap_8 FILLER_4_2467 ();
 sg13g2_decap_8 FILLER_4_2474 ();
 sg13g2_decap_8 FILLER_4_2481 ();
 sg13g2_decap_8 FILLER_4_2488 ();
 sg13g2_decap_8 FILLER_4_2495 ();
 sg13g2_decap_8 FILLER_4_2502 ();
 sg13g2_decap_8 FILLER_4_2509 ();
 sg13g2_decap_8 FILLER_4_2516 ();
 sg13g2_decap_8 FILLER_4_2523 ();
 sg13g2_decap_8 FILLER_4_2530 ();
 sg13g2_decap_8 FILLER_4_2537 ();
 sg13g2_decap_8 FILLER_4_2544 ();
 sg13g2_decap_8 FILLER_4_2551 ();
 sg13g2_decap_8 FILLER_4_2558 ();
 sg13g2_decap_8 FILLER_4_2565 ();
 sg13g2_decap_8 FILLER_4_2572 ();
 sg13g2_decap_8 FILLER_4_2579 ();
 sg13g2_decap_8 FILLER_4_2586 ();
 sg13g2_decap_8 FILLER_4_2593 ();
 sg13g2_decap_8 FILLER_4_2600 ();
 sg13g2_decap_8 FILLER_4_2607 ();
 sg13g2_decap_8 FILLER_4_2614 ();
 sg13g2_decap_8 FILLER_4_2621 ();
 sg13g2_decap_8 FILLER_4_2628 ();
 sg13g2_decap_8 FILLER_4_2635 ();
 sg13g2_decap_8 FILLER_4_2642 ();
 sg13g2_decap_8 FILLER_4_2649 ();
 sg13g2_decap_8 FILLER_4_2656 ();
 sg13g2_decap_8 FILLER_4_2663 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_4 FILLER_5_224 ();
 sg13g2_fill_2 FILLER_5_228 ();
 sg13g2_decap_8 FILLER_5_234 ();
 sg13g2_decap_8 FILLER_5_241 ();
 sg13g2_decap_8 FILLER_5_248 ();
 sg13g2_decap_8 FILLER_5_255 ();
 sg13g2_fill_2 FILLER_5_262 ();
 sg13g2_decap_4 FILLER_5_269 ();
 sg13g2_fill_1 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_284 ();
 sg13g2_decap_8 FILLER_5_291 ();
 sg13g2_decap_4 FILLER_5_298 ();
 sg13g2_fill_2 FILLER_5_302 ();
 sg13g2_decap_8 FILLER_5_307 ();
 sg13g2_decap_8 FILLER_5_314 ();
 sg13g2_decap_8 FILLER_5_321 ();
 sg13g2_decap_8 FILLER_5_328 ();
 sg13g2_decap_8 FILLER_5_335 ();
 sg13g2_decap_8 FILLER_5_342 ();
 sg13g2_decap_8 FILLER_5_349 ();
 sg13g2_decap_8 FILLER_5_356 ();
 sg13g2_decap_8 FILLER_5_363 ();
 sg13g2_decap_8 FILLER_5_370 ();
 sg13g2_decap_8 FILLER_5_377 ();
 sg13g2_decap_8 FILLER_5_384 ();
 sg13g2_decap_8 FILLER_5_391 ();
 sg13g2_decap_8 FILLER_5_398 ();
 sg13g2_decap_4 FILLER_5_405 ();
 sg13g2_fill_1 FILLER_5_409 ();
 sg13g2_decap_8 FILLER_5_433 ();
 sg13g2_decap_8 FILLER_5_440 ();
 sg13g2_decap_8 FILLER_5_447 ();
 sg13g2_decap_8 FILLER_5_454 ();
 sg13g2_decap_8 FILLER_5_461 ();
 sg13g2_decap_8 FILLER_5_468 ();
 sg13g2_decap_4 FILLER_5_475 ();
 sg13g2_fill_1 FILLER_5_479 ();
 sg13g2_decap_8 FILLER_5_496 ();
 sg13g2_decap_8 FILLER_5_503 ();
 sg13g2_decap_8 FILLER_5_510 ();
 sg13g2_decap_8 FILLER_5_517 ();
 sg13g2_decap_8 FILLER_5_524 ();
 sg13g2_decap_8 FILLER_5_531 ();
 sg13g2_decap_8 FILLER_5_538 ();
 sg13g2_decap_8 FILLER_5_545 ();
 sg13g2_decap_8 FILLER_5_552 ();
 sg13g2_decap_8 FILLER_5_559 ();
 sg13g2_decap_8 FILLER_5_566 ();
 sg13g2_decap_8 FILLER_5_573 ();
 sg13g2_decap_8 FILLER_5_580 ();
 sg13g2_decap_8 FILLER_5_587 ();
 sg13g2_decap_8 FILLER_5_594 ();
 sg13g2_decap_8 FILLER_5_601 ();
 sg13g2_fill_1 FILLER_5_612 ();
 sg13g2_decap_8 FILLER_5_617 ();
 sg13g2_decap_8 FILLER_5_624 ();
 sg13g2_decap_8 FILLER_5_631 ();
 sg13g2_decap_8 FILLER_5_638 ();
 sg13g2_fill_2 FILLER_5_645 ();
 sg13g2_fill_1 FILLER_5_647 ();
 sg13g2_decap_8 FILLER_5_653 ();
 sg13g2_decap_8 FILLER_5_660 ();
 sg13g2_decap_8 FILLER_5_667 ();
 sg13g2_decap_8 FILLER_5_674 ();
 sg13g2_decap_8 FILLER_5_681 ();
 sg13g2_decap_8 FILLER_5_688 ();
 sg13g2_decap_8 FILLER_5_695 ();
 sg13g2_decap_8 FILLER_5_702 ();
 sg13g2_decap_8 FILLER_5_709 ();
 sg13g2_decap_8 FILLER_5_716 ();
 sg13g2_decap_8 FILLER_5_723 ();
 sg13g2_decap_8 FILLER_5_730 ();
 sg13g2_decap_8 FILLER_5_737 ();
 sg13g2_decap_8 FILLER_5_744 ();
 sg13g2_decap_8 FILLER_5_751 ();
 sg13g2_decap_8 FILLER_5_758 ();
 sg13g2_decap_8 FILLER_5_765 ();
 sg13g2_decap_8 FILLER_5_772 ();
 sg13g2_decap_8 FILLER_5_779 ();
 sg13g2_decap_8 FILLER_5_786 ();
 sg13g2_decap_8 FILLER_5_793 ();
 sg13g2_decap_4 FILLER_5_800 ();
 sg13g2_fill_1 FILLER_5_804 ();
 sg13g2_decap_8 FILLER_5_820 ();
 sg13g2_decap_8 FILLER_5_827 ();
 sg13g2_decap_8 FILLER_5_834 ();
 sg13g2_decap_8 FILLER_5_841 ();
 sg13g2_decap_8 FILLER_5_848 ();
 sg13g2_decap_8 FILLER_5_855 ();
 sg13g2_fill_1 FILLER_5_862 ();
 sg13g2_decap_8 FILLER_5_871 ();
 sg13g2_decap_8 FILLER_5_878 ();
 sg13g2_decap_8 FILLER_5_885 ();
 sg13g2_decap_8 FILLER_5_892 ();
 sg13g2_decap_8 FILLER_5_899 ();
 sg13g2_decap_8 FILLER_5_918 ();
 sg13g2_decap_8 FILLER_5_925 ();
 sg13g2_fill_1 FILLER_5_932 ();
 sg13g2_decap_8 FILLER_5_948 ();
 sg13g2_decap_8 FILLER_5_955 ();
 sg13g2_decap_8 FILLER_5_962 ();
 sg13g2_decap_8 FILLER_5_969 ();
 sg13g2_decap_8 FILLER_5_976 ();
 sg13g2_decap_8 FILLER_5_983 ();
 sg13g2_decap_8 FILLER_5_990 ();
 sg13g2_decap_8 FILLER_5_997 ();
 sg13g2_decap_8 FILLER_5_1004 ();
 sg13g2_decap_8 FILLER_5_1011 ();
 sg13g2_decap_8 FILLER_5_1018 ();
 sg13g2_fill_2 FILLER_5_1025 ();
 sg13g2_decap_8 FILLER_5_1031 ();
 sg13g2_decap_8 FILLER_5_1038 ();
 sg13g2_decap_8 FILLER_5_1045 ();
 sg13g2_decap_8 FILLER_5_1052 ();
 sg13g2_decap_8 FILLER_5_1059 ();
 sg13g2_decap_8 FILLER_5_1066 ();
 sg13g2_decap_8 FILLER_5_1073 ();
 sg13g2_decap_4 FILLER_5_1080 ();
 sg13g2_fill_1 FILLER_5_1084 ();
 sg13g2_decap_8 FILLER_5_1108 ();
 sg13g2_decap_8 FILLER_5_1115 ();
 sg13g2_fill_2 FILLER_5_1122 ();
 sg13g2_fill_1 FILLER_5_1124 ();
 sg13g2_fill_2 FILLER_5_1140 ();
 sg13g2_decap_8 FILLER_5_1146 ();
 sg13g2_decap_8 FILLER_5_1153 ();
 sg13g2_decap_8 FILLER_5_1160 ();
 sg13g2_decap_8 FILLER_5_1167 ();
 sg13g2_fill_2 FILLER_5_1174 ();
 sg13g2_decap_8 FILLER_5_1181 ();
 sg13g2_decap_8 FILLER_5_1188 ();
 sg13g2_decap_8 FILLER_5_1195 ();
 sg13g2_decap_8 FILLER_5_1202 ();
 sg13g2_fill_2 FILLER_5_1209 ();
 sg13g2_fill_1 FILLER_5_1211 ();
 sg13g2_fill_2 FILLER_5_1221 ();
 sg13g2_fill_1 FILLER_5_1223 ();
 sg13g2_decap_8 FILLER_5_1228 ();
 sg13g2_decap_8 FILLER_5_1235 ();
 sg13g2_decap_4 FILLER_5_1242 ();
 sg13g2_fill_2 FILLER_5_1246 ();
 sg13g2_decap_8 FILLER_5_1264 ();
 sg13g2_decap_8 FILLER_5_1271 ();
 sg13g2_decap_8 FILLER_5_1278 ();
 sg13g2_decap_8 FILLER_5_1285 ();
 sg13g2_decap_8 FILLER_5_1292 ();
 sg13g2_decap_8 FILLER_5_1299 ();
 sg13g2_decap_8 FILLER_5_1306 ();
 sg13g2_decap_8 FILLER_5_1313 ();
 sg13g2_decap_8 FILLER_5_1320 ();
 sg13g2_decap_8 FILLER_5_1327 ();
 sg13g2_decap_8 FILLER_5_1334 ();
 sg13g2_decap_8 FILLER_5_1341 ();
 sg13g2_fill_2 FILLER_5_1348 ();
 sg13g2_fill_1 FILLER_5_1350 ();
 sg13g2_decap_8 FILLER_5_1355 ();
 sg13g2_decap_4 FILLER_5_1362 ();
 sg13g2_fill_1 FILLER_5_1366 ();
 sg13g2_decap_8 FILLER_5_1371 ();
 sg13g2_decap_8 FILLER_5_1378 ();
 sg13g2_decap_4 FILLER_5_1385 ();
 sg13g2_fill_1 FILLER_5_1389 ();
 sg13g2_decap_8 FILLER_5_1405 ();
 sg13g2_decap_8 FILLER_5_1412 ();
 sg13g2_decap_8 FILLER_5_1419 ();
 sg13g2_decap_8 FILLER_5_1426 ();
 sg13g2_decap_8 FILLER_5_1433 ();
 sg13g2_decap_8 FILLER_5_1440 ();
 sg13g2_decap_8 FILLER_5_1447 ();
 sg13g2_decap_8 FILLER_5_1454 ();
 sg13g2_decap_8 FILLER_5_1461 ();
 sg13g2_decap_8 FILLER_5_1468 ();
 sg13g2_decap_8 FILLER_5_1475 ();
 sg13g2_decap_8 FILLER_5_1482 ();
 sg13g2_decap_8 FILLER_5_1489 ();
 sg13g2_decap_8 FILLER_5_1496 ();
 sg13g2_decap_8 FILLER_5_1503 ();
 sg13g2_decap_4 FILLER_5_1510 ();
 sg13g2_decap_8 FILLER_5_1522 ();
 sg13g2_decap_8 FILLER_5_1529 ();
 sg13g2_decap_8 FILLER_5_1536 ();
 sg13g2_fill_2 FILLER_5_1543 ();
 sg13g2_fill_1 FILLER_5_1545 ();
 sg13g2_fill_2 FILLER_5_1554 ();
 sg13g2_decap_8 FILLER_5_1570 ();
 sg13g2_decap_8 FILLER_5_1577 ();
 sg13g2_decap_8 FILLER_5_1584 ();
 sg13g2_decap_8 FILLER_5_1591 ();
 sg13g2_decap_8 FILLER_5_1598 ();
 sg13g2_decap_8 FILLER_5_1605 ();
 sg13g2_decap_8 FILLER_5_1612 ();
 sg13g2_fill_2 FILLER_5_1619 ();
 sg13g2_fill_2 FILLER_5_1629 ();
 sg13g2_decap_8 FILLER_5_1635 ();
 sg13g2_decap_8 FILLER_5_1642 ();
 sg13g2_decap_8 FILLER_5_1649 ();
 sg13g2_decap_8 FILLER_5_1656 ();
 sg13g2_decap_8 FILLER_5_1663 ();
 sg13g2_fill_2 FILLER_5_1670 ();
 sg13g2_fill_1 FILLER_5_1672 ();
 sg13g2_decap_8 FILLER_5_1686 ();
 sg13g2_decap_8 FILLER_5_1693 ();
 sg13g2_decap_8 FILLER_5_1700 ();
 sg13g2_decap_8 FILLER_5_1707 ();
 sg13g2_decap_8 FILLER_5_1714 ();
 sg13g2_decap_8 FILLER_5_1721 ();
 sg13g2_decap_8 FILLER_5_1728 ();
 sg13g2_decap_8 FILLER_5_1735 ();
 sg13g2_decap_8 FILLER_5_1742 ();
 sg13g2_decap_8 FILLER_5_1749 ();
 sg13g2_decap_8 FILLER_5_1756 ();
 sg13g2_decap_8 FILLER_5_1763 ();
 sg13g2_decap_8 FILLER_5_1770 ();
 sg13g2_decap_8 FILLER_5_1777 ();
 sg13g2_decap_8 FILLER_5_1784 ();
 sg13g2_decap_8 FILLER_5_1791 ();
 sg13g2_decap_8 FILLER_5_1798 ();
 sg13g2_decap_8 FILLER_5_1805 ();
 sg13g2_decap_8 FILLER_5_1812 ();
 sg13g2_decap_8 FILLER_5_1819 ();
 sg13g2_decap_8 FILLER_5_1826 ();
 sg13g2_decap_8 FILLER_5_1833 ();
 sg13g2_decap_8 FILLER_5_1840 ();
 sg13g2_decap_8 FILLER_5_1847 ();
 sg13g2_decap_8 FILLER_5_1854 ();
 sg13g2_decap_8 FILLER_5_1861 ();
 sg13g2_decap_8 FILLER_5_1868 ();
 sg13g2_decap_8 FILLER_5_1875 ();
 sg13g2_decap_8 FILLER_5_1882 ();
 sg13g2_decap_8 FILLER_5_1889 ();
 sg13g2_decap_8 FILLER_5_1896 ();
 sg13g2_decap_8 FILLER_5_1903 ();
 sg13g2_decap_8 FILLER_5_1910 ();
 sg13g2_decap_8 FILLER_5_1917 ();
 sg13g2_decap_8 FILLER_5_1924 ();
 sg13g2_decap_8 FILLER_5_1931 ();
 sg13g2_decap_8 FILLER_5_1938 ();
 sg13g2_decap_8 FILLER_5_1945 ();
 sg13g2_decap_8 FILLER_5_1952 ();
 sg13g2_decap_8 FILLER_5_1959 ();
 sg13g2_decap_8 FILLER_5_1966 ();
 sg13g2_decap_8 FILLER_5_1973 ();
 sg13g2_decap_8 FILLER_5_1980 ();
 sg13g2_decap_8 FILLER_5_1987 ();
 sg13g2_decap_8 FILLER_5_1994 ();
 sg13g2_decap_8 FILLER_5_2001 ();
 sg13g2_decap_8 FILLER_5_2008 ();
 sg13g2_decap_8 FILLER_5_2015 ();
 sg13g2_decap_8 FILLER_5_2022 ();
 sg13g2_decap_8 FILLER_5_2029 ();
 sg13g2_decap_8 FILLER_5_2036 ();
 sg13g2_decap_8 FILLER_5_2043 ();
 sg13g2_decap_8 FILLER_5_2050 ();
 sg13g2_decap_8 FILLER_5_2057 ();
 sg13g2_decap_8 FILLER_5_2064 ();
 sg13g2_decap_8 FILLER_5_2071 ();
 sg13g2_decap_8 FILLER_5_2078 ();
 sg13g2_decap_8 FILLER_5_2085 ();
 sg13g2_decap_8 FILLER_5_2092 ();
 sg13g2_decap_8 FILLER_5_2099 ();
 sg13g2_decap_8 FILLER_5_2106 ();
 sg13g2_decap_8 FILLER_5_2113 ();
 sg13g2_decap_8 FILLER_5_2120 ();
 sg13g2_decap_8 FILLER_5_2127 ();
 sg13g2_decap_8 FILLER_5_2134 ();
 sg13g2_decap_8 FILLER_5_2141 ();
 sg13g2_decap_8 FILLER_5_2148 ();
 sg13g2_decap_8 FILLER_5_2155 ();
 sg13g2_decap_8 FILLER_5_2162 ();
 sg13g2_decap_8 FILLER_5_2169 ();
 sg13g2_decap_8 FILLER_5_2176 ();
 sg13g2_decap_8 FILLER_5_2183 ();
 sg13g2_decap_8 FILLER_5_2190 ();
 sg13g2_decap_8 FILLER_5_2197 ();
 sg13g2_decap_8 FILLER_5_2204 ();
 sg13g2_decap_8 FILLER_5_2211 ();
 sg13g2_decap_8 FILLER_5_2218 ();
 sg13g2_decap_8 FILLER_5_2225 ();
 sg13g2_decap_8 FILLER_5_2232 ();
 sg13g2_decap_8 FILLER_5_2239 ();
 sg13g2_decap_8 FILLER_5_2246 ();
 sg13g2_decap_8 FILLER_5_2253 ();
 sg13g2_decap_8 FILLER_5_2260 ();
 sg13g2_decap_8 FILLER_5_2267 ();
 sg13g2_decap_8 FILLER_5_2274 ();
 sg13g2_decap_8 FILLER_5_2281 ();
 sg13g2_decap_8 FILLER_5_2288 ();
 sg13g2_decap_8 FILLER_5_2295 ();
 sg13g2_decap_8 FILLER_5_2302 ();
 sg13g2_decap_8 FILLER_5_2309 ();
 sg13g2_decap_8 FILLER_5_2316 ();
 sg13g2_decap_8 FILLER_5_2323 ();
 sg13g2_decap_8 FILLER_5_2330 ();
 sg13g2_decap_8 FILLER_5_2337 ();
 sg13g2_decap_8 FILLER_5_2344 ();
 sg13g2_decap_8 FILLER_5_2351 ();
 sg13g2_decap_8 FILLER_5_2358 ();
 sg13g2_decap_8 FILLER_5_2365 ();
 sg13g2_decap_8 FILLER_5_2372 ();
 sg13g2_decap_8 FILLER_5_2379 ();
 sg13g2_decap_8 FILLER_5_2386 ();
 sg13g2_decap_8 FILLER_5_2393 ();
 sg13g2_decap_8 FILLER_5_2400 ();
 sg13g2_decap_8 FILLER_5_2407 ();
 sg13g2_decap_8 FILLER_5_2414 ();
 sg13g2_decap_8 FILLER_5_2421 ();
 sg13g2_decap_8 FILLER_5_2428 ();
 sg13g2_decap_8 FILLER_5_2435 ();
 sg13g2_decap_8 FILLER_5_2442 ();
 sg13g2_decap_8 FILLER_5_2449 ();
 sg13g2_decap_8 FILLER_5_2456 ();
 sg13g2_decap_8 FILLER_5_2463 ();
 sg13g2_decap_8 FILLER_5_2470 ();
 sg13g2_decap_8 FILLER_5_2477 ();
 sg13g2_decap_8 FILLER_5_2484 ();
 sg13g2_decap_8 FILLER_5_2491 ();
 sg13g2_decap_8 FILLER_5_2498 ();
 sg13g2_decap_8 FILLER_5_2505 ();
 sg13g2_decap_8 FILLER_5_2512 ();
 sg13g2_decap_8 FILLER_5_2519 ();
 sg13g2_decap_8 FILLER_5_2526 ();
 sg13g2_decap_8 FILLER_5_2533 ();
 sg13g2_decap_8 FILLER_5_2540 ();
 sg13g2_decap_8 FILLER_5_2547 ();
 sg13g2_decap_8 FILLER_5_2554 ();
 sg13g2_decap_8 FILLER_5_2561 ();
 sg13g2_decap_8 FILLER_5_2568 ();
 sg13g2_decap_8 FILLER_5_2575 ();
 sg13g2_decap_8 FILLER_5_2582 ();
 sg13g2_decap_8 FILLER_5_2589 ();
 sg13g2_decap_8 FILLER_5_2596 ();
 sg13g2_decap_8 FILLER_5_2603 ();
 sg13g2_decap_8 FILLER_5_2610 ();
 sg13g2_decap_8 FILLER_5_2617 ();
 sg13g2_decap_8 FILLER_5_2624 ();
 sg13g2_decap_8 FILLER_5_2631 ();
 sg13g2_decap_8 FILLER_5_2638 ();
 sg13g2_decap_8 FILLER_5_2645 ();
 sg13g2_decap_8 FILLER_5_2652 ();
 sg13g2_decap_8 FILLER_5_2659 ();
 sg13g2_decap_4 FILLER_5_2666 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_fill_1 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_253 ();
 sg13g2_decap_4 FILLER_6_264 ();
 sg13g2_decap_8 FILLER_6_271 ();
 sg13g2_decap_8 FILLER_6_278 ();
 sg13g2_decap_8 FILLER_6_285 ();
 sg13g2_decap_8 FILLER_6_292 ();
 sg13g2_decap_8 FILLER_6_299 ();
 sg13g2_decap_8 FILLER_6_306 ();
 sg13g2_decap_8 FILLER_6_313 ();
 sg13g2_decap_8 FILLER_6_320 ();
 sg13g2_decap_8 FILLER_6_327 ();
 sg13g2_decap_8 FILLER_6_334 ();
 sg13g2_decap_8 FILLER_6_341 ();
 sg13g2_decap_8 FILLER_6_348 ();
 sg13g2_decap_8 FILLER_6_355 ();
 sg13g2_decap_8 FILLER_6_362 ();
 sg13g2_decap_8 FILLER_6_369 ();
 sg13g2_decap_8 FILLER_6_376 ();
 sg13g2_decap_8 FILLER_6_383 ();
 sg13g2_decap_8 FILLER_6_390 ();
 sg13g2_decap_8 FILLER_6_397 ();
 sg13g2_decap_8 FILLER_6_404 ();
 sg13g2_decap_8 FILLER_6_411 ();
 sg13g2_decap_8 FILLER_6_418 ();
 sg13g2_decap_8 FILLER_6_425 ();
 sg13g2_decap_8 FILLER_6_432 ();
 sg13g2_decap_4 FILLER_6_439 ();
 sg13g2_fill_1 FILLER_6_443 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_4 FILLER_6_469 ();
 sg13g2_fill_1 FILLER_6_473 ();
 sg13g2_decap_8 FILLER_6_494 ();
 sg13g2_decap_8 FILLER_6_501 ();
 sg13g2_fill_1 FILLER_6_508 ();
 sg13g2_decap_8 FILLER_6_521 ();
 sg13g2_decap_8 FILLER_6_528 ();
 sg13g2_decap_8 FILLER_6_535 ();
 sg13g2_decap_8 FILLER_6_542 ();
 sg13g2_decap_8 FILLER_6_549 ();
 sg13g2_decap_8 FILLER_6_556 ();
 sg13g2_decap_8 FILLER_6_566 ();
 sg13g2_decap_8 FILLER_6_573 ();
 sg13g2_decap_8 FILLER_6_580 ();
 sg13g2_decap_4 FILLER_6_587 ();
 sg13g2_fill_1 FILLER_6_591 ();
 sg13g2_decap_8 FILLER_6_596 ();
 sg13g2_decap_8 FILLER_6_603 ();
 sg13g2_decap_4 FILLER_6_610 ();
 sg13g2_fill_1 FILLER_6_614 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_666 ();
 sg13g2_decap_8 FILLER_6_673 ();
 sg13g2_decap_8 FILLER_6_680 ();
 sg13g2_decap_8 FILLER_6_687 ();
 sg13g2_decap_8 FILLER_6_694 ();
 sg13g2_decap_8 FILLER_6_701 ();
 sg13g2_decap_8 FILLER_6_708 ();
 sg13g2_decap_8 FILLER_6_715 ();
 sg13g2_fill_2 FILLER_6_722 ();
 sg13g2_fill_1 FILLER_6_724 ();
 sg13g2_decap_8 FILLER_6_740 ();
 sg13g2_decap_8 FILLER_6_747 ();
 sg13g2_decap_8 FILLER_6_754 ();
 sg13g2_decap_8 FILLER_6_761 ();
 sg13g2_decap_8 FILLER_6_768 ();
 sg13g2_decap_8 FILLER_6_775 ();
 sg13g2_decap_8 FILLER_6_782 ();
 sg13g2_decap_4 FILLER_6_789 ();
 sg13g2_fill_2 FILLER_6_793 ();
 sg13g2_fill_2 FILLER_6_810 ();
 sg13g2_decap_8 FILLER_6_816 ();
 sg13g2_decap_8 FILLER_6_823 ();
 sg13g2_decap_8 FILLER_6_830 ();
 sg13g2_decap_8 FILLER_6_837 ();
 sg13g2_fill_2 FILLER_6_844 ();
 sg13g2_fill_1 FILLER_6_849 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_decap_8 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_6_868 ();
 sg13g2_decap_8 FILLER_6_875 ();
 sg13g2_decap_8 FILLER_6_882 ();
 sg13g2_decap_8 FILLER_6_889 ();
 sg13g2_decap_8 FILLER_6_896 ();
 sg13g2_decap_8 FILLER_6_903 ();
 sg13g2_decap_8 FILLER_6_910 ();
 sg13g2_decap_8 FILLER_6_917 ();
 sg13g2_fill_2 FILLER_6_924 ();
 sg13g2_fill_1 FILLER_6_926 ();
 sg13g2_decap_8 FILLER_6_948 ();
 sg13g2_decap_8 FILLER_6_955 ();
 sg13g2_decap_4 FILLER_6_962 ();
 sg13g2_fill_2 FILLER_6_966 ();
 sg13g2_decap_8 FILLER_6_971 ();
 sg13g2_fill_2 FILLER_6_993 ();
 sg13g2_decap_8 FILLER_6_1001 ();
 sg13g2_decap_8 FILLER_6_1008 ();
 sg13g2_decap_8 FILLER_6_1015 ();
 sg13g2_decap_8 FILLER_6_1022 ();
 sg13g2_fill_1 FILLER_6_1029 ();
 sg13g2_decap_8 FILLER_6_1033 ();
 sg13g2_decap_8 FILLER_6_1040 ();
 sg13g2_decap_8 FILLER_6_1047 ();
 sg13g2_decap_4 FILLER_6_1054 ();
 sg13g2_fill_2 FILLER_6_1058 ();
 sg13g2_decap_8 FILLER_6_1075 ();
 sg13g2_decap_8 FILLER_6_1082 ();
 sg13g2_decap_8 FILLER_6_1089 ();
 sg13g2_decap_4 FILLER_6_1096 ();
 sg13g2_decap_8 FILLER_6_1112 ();
 sg13g2_decap_8 FILLER_6_1119 ();
 sg13g2_decap_4 FILLER_6_1126 ();
 sg13g2_fill_1 FILLER_6_1130 ();
 sg13g2_decap_8 FILLER_6_1142 ();
 sg13g2_decap_8 FILLER_6_1149 ();
 sg13g2_decap_8 FILLER_6_1156 ();
 sg13g2_decap_8 FILLER_6_1163 ();
 sg13g2_decap_8 FILLER_6_1170 ();
 sg13g2_fill_2 FILLER_6_1177 ();
 sg13g2_fill_1 FILLER_6_1179 ();
 sg13g2_decap_8 FILLER_6_1189 ();
 sg13g2_decap_8 FILLER_6_1196 ();
 sg13g2_decap_8 FILLER_6_1203 ();
 sg13g2_decap_8 FILLER_6_1210 ();
 sg13g2_decap_8 FILLER_6_1217 ();
 sg13g2_decap_8 FILLER_6_1224 ();
 sg13g2_decap_8 FILLER_6_1231 ();
 sg13g2_decap_8 FILLER_6_1238 ();
 sg13g2_decap_8 FILLER_6_1261 ();
 sg13g2_decap_8 FILLER_6_1268 ();
 sg13g2_decap_8 FILLER_6_1275 ();
 sg13g2_decap_8 FILLER_6_1282 ();
 sg13g2_decap_8 FILLER_6_1289 ();
 sg13g2_decap_8 FILLER_6_1296 ();
 sg13g2_decap_8 FILLER_6_1303 ();
 sg13g2_decap_8 FILLER_6_1310 ();
 sg13g2_decap_8 FILLER_6_1317 ();
 sg13g2_decap_8 FILLER_6_1324 ();
 sg13g2_decap_8 FILLER_6_1331 ();
 sg13g2_decap_8 FILLER_6_1338 ();
 sg13g2_decap_8 FILLER_6_1345 ();
 sg13g2_decap_8 FILLER_6_1352 ();
 sg13g2_decap_8 FILLER_6_1359 ();
 sg13g2_decap_8 FILLER_6_1366 ();
 sg13g2_decap_8 FILLER_6_1373 ();
 sg13g2_decap_8 FILLER_6_1380 ();
 sg13g2_fill_2 FILLER_6_1387 ();
 sg13g2_fill_1 FILLER_6_1389 ();
 sg13g2_decap_8 FILLER_6_1394 ();
 sg13g2_decap_8 FILLER_6_1401 ();
 sg13g2_decap_8 FILLER_6_1408 ();
 sg13g2_decap_8 FILLER_6_1415 ();
 sg13g2_decap_4 FILLER_6_1422 ();
 sg13g2_fill_2 FILLER_6_1429 ();
 sg13g2_fill_2 FILLER_6_1438 ();
 sg13g2_decap_8 FILLER_6_1453 ();
 sg13g2_decap_8 FILLER_6_1460 ();
 sg13g2_decap_8 FILLER_6_1467 ();
 sg13g2_decap_8 FILLER_6_1474 ();
 sg13g2_decap_8 FILLER_6_1481 ();
 sg13g2_decap_8 FILLER_6_1488 ();
 sg13g2_decap_8 FILLER_6_1495 ();
 sg13g2_decap_8 FILLER_6_1502 ();
 sg13g2_decap_4 FILLER_6_1509 ();
 sg13g2_fill_1 FILLER_6_1513 ();
 sg13g2_decap_8 FILLER_6_1517 ();
 sg13g2_decap_8 FILLER_6_1524 ();
 sg13g2_decap_8 FILLER_6_1531 ();
 sg13g2_decap_8 FILLER_6_1538 ();
 sg13g2_decap_4 FILLER_6_1545 ();
 sg13g2_decap_8 FILLER_6_1552 ();
 sg13g2_decap_4 FILLER_6_1559 ();
 sg13g2_fill_2 FILLER_6_1563 ();
 sg13g2_decap_8 FILLER_6_1569 ();
 sg13g2_decap_8 FILLER_6_1576 ();
 sg13g2_decap_8 FILLER_6_1583 ();
 sg13g2_decap_8 FILLER_6_1590 ();
 sg13g2_decap_8 FILLER_6_1597 ();
 sg13g2_decap_8 FILLER_6_1604 ();
 sg13g2_decap_8 FILLER_6_1611 ();
 sg13g2_decap_8 FILLER_6_1618 ();
 sg13g2_decap_8 FILLER_6_1625 ();
 sg13g2_decap_8 FILLER_6_1632 ();
 sg13g2_decap_8 FILLER_6_1639 ();
 sg13g2_decap_8 FILLER_6_1646 ();
 sg13g2_fill_1 FILLER_6_1653 ();
 sg13g2_decap_8 FILLER_6_1658 ();
 sg13g2_decap_8 FILLER_6_1665 ();
 sg13g2_decap_8 FILLER_6_1672 ();
 sg13g2_decap_8 FILLER_6_1679 ();
 sg13g2_decap_8 FILLER_6_1686 ();
 sg13g2_decap_8 FILLER_6_1693 ();
 sg13g2_decap_8 FILLER_6_1700 ();
 sg13g2_decap_8 FILLER_6_1707 ();
 sg13g2_decap_8 FILLER_6_1714 ();
 sg13g2_fill_2 FILLER_6_1721 ();
 sg13g2_decap_8 FILLER_6_1736 ();
 sg13g2_decap_8 FILLER_6_1743 ();
 sg13g2_fill_2 FILLER_6_1750 ();
 sg13g2_decap_8 FILLER_6_1765 ();
 sg13g2_decap_8 FILLER_6_1772 ();
 sg13g2_decap_8 FILLER_6_1779 ();
 sg13g2_decap_8 FILLER_6_1786 ();
 sg13g2_decap_8 FILLER_6_1793 ();
 sg13g2_fill_2 FILLER_6_1800 ();
 sg13g2_fill_1 FILLER_6_1802 ();
 sg13g2_decap_8 FILLER_6_1820 ();
 sg13g2_decap_8 FILLER_6_1827 ();
 sg13g2_decap_8 FILLER_6_1834 ();
 sg13g2_decap_8 FILLER_6_1841 ();
 sg13g2_decap_8 FILLER_6_1848 ();
 sg13g2_decap_8 FILLER_6_1855 ();
 sg13g2_decap_8 FILLER_6_1862 ();
 sg13g2_decap_8 FILLER_6_1869 ();
 sg13g2_decap_8 FILLER_6_1876 ();
 sg13g2_decap_8 FILLER_6_1883 ();
 sg13g2_decap_8 FILLER_6_1890 ();
 sg13g2_decap_8 FILLER_6_1897 ();
 sg13g2_decap_8 FILLER_6_1904 ();
 sg13g2_decap_8 FILLER_6_1911 ();
 sg13g2_decap_8 FILLER_6_1918 ();
 sg13g2_decap_8 FILLER_6_1925 ();
 sg13g2_decap_8 FILLER_6_1932 ();
 sg13g2_decap_8 FILLER_6_1939 ();
 sg13g2_decap_8 FILLER_6_1946 ();
 sg13g2_decap_8 FILLER_6_1953 ();
 sg13g2_decap_8 FILLER_6_1960 ();
 sg13g2_decap_8 FILLER_6_1967 ();
 sg13g2_decap_8 FILLER_6_1974 ();
 sg13g2_decap_8 FILLER_6_1981 ();
 sg13g2_decap_8 FILLER_6_1988 ();
 sg13g2_decap_8 FILLER_6_1995 ();
 sg13g2_decap_8 FILLER_6_2002 ();
 sg13g2_decap_8 FILLER_6_2009 ();
 sg13g2_decap_8 FILLER_6_2016 ();
 sg13g2_decap_8 FILLER_6_2023 ();
 sg13g2_decap_8 FILLER_6_2030 ();
 sg13g2_decap_8 FILLER_6_2037 ();
 sg13g2_decap_8 FILLER_6_2044 ();
 sg13g2_decap_8 FILLER_6_2051 ();
 sg13g2_decap_8 FILLER_6_2058 ();
 sg13g2_decap_8 FILLER_6_2065 ();
 sg13g2_decap_8 FILLER_6_2072 ();
 sg13g2_decap_8 FILLER_6_2079 ();
 sg13g2_decap_8 FILLER_6_2086 ();
 sg13g2_decap_8 FILLER_6_2093 ();
 sg13g2_decap_8 FILLER_6_2100 ();
 sg13g2_decap_8 FILLER_6_2107 ();
 sg13g2_decap_8 FILLER_6_2114 ();
 sg13g2_decap_8 FILLER_6_2121 ();
 sg13g2_decap_8 FILLER_6_2128 ();
 sg13g2_decap_8 FILLER_6_2135 ();
 sg13g2_decap_8 FILLER_6_2142 ();
 sg13g2_decap_8 FILLER_6_2149 ();
 sg13g2_decap_8 FILLER_6_2156 ();
 sg13g2_decap_8 FILLER_6_2163 ();
 sg13g2_decap_8 FILLER_6_2170 ();
 sg13g2_decap_8 FILLER_6_2177 ();
 sg13g2_decap_8 FILLER_6_2184 ();
 sg13g2_decap_8 FILLER_6_2191 ();
 sg13g2_decap_8 FILLER_6_2198 ();
 sg13g2_decap_8 FILLER_6_2205 ();
 sg13g2_decap_8 FILLER_6_2212 ();
 sg13g2_decap_8 FILLER_6_2219 ();
 sg13g2_decap_8 FILLER_6_2226 ();
 sg13g2_decap_8 FILLER_6_2233 ();
 sg13g2_decap_8 FILLER_6_2240 ();
 sg13g2_decap_8 FILLER_6_2247 ();
 sg13g2_decap_8 FILLER_6_2254 ();
 sg13g2_decap_8 FILLER_6_2261 ();
 sg13g2_decap_8 FILLER_6_2268 ();
 sg13g2_decap_8 FILLER_6_2275 ();
 sg13g2_decap_8 FILLER_6_2282 ();
 sg13g2_decap_8 FILLER_6_2289 ();
 sg13g2_decap_8 FILLER_6_2296 ();
 sg13g2_decap_8 FILLER_6_2303 ();
 sg13g2_decap_8 FILLER_6_2310 ();
 sg13g2_decap_8 FILLER_6_2317 ();
 sg13g2_decap_8 FILLER_6_2324 ();
 sg13g2_decap_8 FILLER_6_2331 ();
 sg13g2_decap_8 FILLER_6_2338 ();
 sg13g2_decap_8 FILLER_6_2345 ();
 sg13g2_decap_8 FILLER_6_2352 ();
 sg13g2_decap_8 FILLER_6_2359 ();
 sg13g2_decap_8 FILLER_6_2366 ();
 sg13g2_decap_8 FILLER_6_2373 ();
 sg13g2_decap_8 FILLER_6_2380 ();
 sg13g2_decap_8 FILLER_6_2387 ();
 sg13g2_decap_8 FILLER_6_2394 ();
 sg13g2_decap_8 FILLER_6_2401 ();
 sg13g2_decap_8 FILLER_6_2408 ();
 sg13g2_decap_8 FILLER_6_2415 ();
 sg13g2_decap_8 FILLER_6_2422 ();
 sg13g2_decap_8 FILLER_6_2429 ();
 sg13g2_decap_8 FILLER_6_2436 ();
 sg13g2_decap_8 FILLER_6_2443 ();
 sg13g2_decap_8 FILLER_6_2450 ();
 sg13g2_decap_8 FILLER_6_2457 ();
 sg13g2_decap_8 FILLER_6_2464 ();
 sg13g2_decap_8 FILLER_6_2471 ();
 sg13g2_decap_8 FILLER_6_2478 ();
 sg13g2_decap_8 FILLER_6_2485 ();
 sg13g2_decap_8 FILLER_6_2492 ();
 sg13g2_decap_8 FILLER_6_2499 ();
 sg13g2_decap_8 FILLER_6_2506 ();
 sg13g2_decap_8 FILLER_6_2513 ();
 sg13g2_decap_8 FILLER_6_2520 ();
 sg13g2_decap_8 FILLER_6_2527 ();
 sg13g2_decap_8 FILLER_6_2534 ();
 sg13g2_decap_8 FILLER_6_2541 ();
 sg13g2_decap_8 FILLER_6_2548 ();
 sg13g2_decap_8 FILLER_6_2555 ();
 sg13g2_decap_8 FILLER_6_2562 ();
 sg13g2_decap_8 FILLER_6_2569 ();
 sg13g2_decap_8 FILLER_6_2576 ();
 sg13g2_decap_8 FILLER_6_2583 ();
 sg13g2_decap_8 FILLER_6_2590 ();
 sg13g2_decap_8 FILLER_6_2597 ();
 sg13g2_decap_8 FILLER_6_2604 ();
 sg13g2_decap_8 FILLER_6_2611 ();
 sg13g2_decap_8 FILLER_6_2618 ();
 sg13g2_decap_8 FILLER_6_2625 ();
 sg13g2_decap_8 FILLER_6_2632 ();
 sg13g2_decap_8 FILLER_6_2639 ();
 sg13g2_decap_8 FILLER_6_2646 ();
 sg13g2_decap_8 FILLER_6_2653 ();
 sg13g2_decap_8 FILLER_6_2660 ();
 sg13g2_fill_2 FILLER_6_2667 ();
 sg13g2_fill_1 FILLER_6_2669 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_4 FILLER_7_105 ();
 sg13g2_fill_1 FILLER_7_109 ();
 sg13g2_decap_8 FILLER_7_114 ();
 sg13g2_decap_8 FILLER_7_121 ();
 sg13g2_decap_8 FILLER_7_128 ();
 sg13g2_decap_8 FILLER_7_135 ();
 sg13g2_decap_8 FILLER_7_142 ();
 sg13g2_decap_8 FILLER_7_149 ();
 sg13g2_decap_8 FILLER_7_156 ();
 sg13g2_decap_8 FILLER_7_163 ();
 sg13g2_decap_8 FILLER_7_170 ();
 sg13g2_decap_8 FILLER_7_177 ();
 sg13g2_fill_2 FILLER_7_184 ();
 sg13g2_fill_1 FILLER_7_186 ();
 sg13g2_decap_8 FILLER_7_191 ();
 sg13g2_decap_8 FILLER_7_198 ();
 sg13g2_decap_8 FILLER_7_205 ();
 sg13g2_decap_8 FILLER_7_212 ();
 sg13g2_decap_8 FILLER_7_219 ();
 sg13g2_decap_8 FILLER_7_226 ();
 sg13g2_decap_8 FILLER_7_233 ();
 sg13g2_decap_8 FILLER_7_240 ();
 sg13g2_decap_8 FILLER_7_247 ();
 sg13g2_decap_8 FILLER_7_254 ();
 sg13g2_decap_8 FILLER_7_261 ();
 sg13g2_decap_8 FILLER_7_268 ();
 sg13g2_decap_8 FILLER_7_275 ();
 sg13g2_decap_8 FILLER_7_282 ();
 sg13g2_decap_8 FILLER_7_289 ();
 sg13g2_decap_8 FILLER_7_296 ();
 sg13g2_decap_8 FILLER_7_303 ();
 sg13g2_decap_8 FILLER_7_310 ();
 sg13g2_decap_8 FILLER_7_317 ();
 sg13g2_decap_8 FILLER_7_324 ();
 sg13g2_decap_8 FILLER_7_331 ();
 sg13g2_decap_8 FILLER_7_338 ();
 sg13g2_decap_8 FILLER_7_345 ();
 sg13g2_decap_8 FILLER_7_352 ();
 sg13g2_decap_8 FILLER_7_359 ();
 sg13g2_decap_8 FILLER_7_366 ();
 sg13g2_decap_8 FILLER_7_373 ();
 sg13g2_decap_8 FILLER_7_380 ();
 sg13g2_fill_2 FILLER_7_387 ();
 sg13g2_fill_1 FILLER_7_389 ();
 sg13g2_decap_8 FILLER_7_398 ();
 sg13g2_decap_8 FILLER_7_405 ();
 sg13g2_decap_8 FILLER_7_412 ();
 sg13g2_decap_8 FILLER_7_419 ();
 sg13g2_decap_8 FILLER_7_426 ();
 sg13g2_decap_8 FILLER_7_433 ();
 sg13g2_decap_8 FILLER_7_440 ();
 sg13g2_decap_8 FILLER_7_447 ();
 sg13g2_decap_8 FILLER_7_454 ();
 sg13g2_decap_8 FILLER_7_461 ();
 sg13g2_decap_8 FILLER_7_468 ();
 sg13g2_decap_8 FILLER_7_475 ();
 sg13g2_decap_8 FILLER_7_482 ();
 sg13g2_decap_8 FILLER_7_489 ();
 sg13g2_decap_8 FILLER_7_496 ();
 sg13g2_fill_2 FILLER_7_503 ();
 sg13g2_fill_1 FILLER_7_505 ();
 sg13g2_decap_8 FILLER_7_517 ();
 sg13g2_decap_4 FILLER_7_524 ();
 sg13g2_fill_1 FILLER_7_528 ();
 sg13g2_decap_8 FILLER_7_533 ();
 sg13g2_decap_8 FILLER_7_540 ();
 sg13g2_decap_8 FILLER_7_547 ();
 sg13g2_decap_4 FILLER_7_554 ();
 sg13g2_fill_2 FILLER_7_558 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_fill_2 FILLER_7_588 ();
 sg13g2_fill_1 FILLER_7_599 ();
 sg13g2_decap_8 FILLER_7_607 ();
 sg13g2_decap_4 FILLER_7_614 ();
 sg13g2_decap_8 FILLER_7_622 ();
 sg13g2_decap_8 FILLER_7_629 ();
 sg13g2_decap_8 FILLER_7_636 ();
 sg13g2_decap_8 FILLER_7_643 ();
 sg13g2_decap_4 FILLER_7_650 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_4 FILLER_7_679 ();
 sg13g2_fill_1 FILLER_7_683 ();
 sg13g2_decap_8 FILLER_7_694 ();
 sg13g2_fill_2 FILLER_7_701 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_fill_1 FILLER_7_721 ();
 sg13g2_fill_1 FILLER_7_733 ();
 sg13g2_fill_1 FILLER_7_738 ();
 sg13g2_decap_4 FILLER_7_744 ();
 sg13g2_fill_2 FILLER_7_748 ();
 sg13g2_fill_1 FILLER_7_754 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_4 FILLER_7_791 ();
 sg13g2_fill_2 FILLER_7_795 ();
 sg13g2_decap_8 FILLER_7_814 ();
 sg13g2_decap_8 FILLER_7_821 ();
 sg13g2_decap_8 FILLER_7_828 ();
 sg13g2_decap_8 FILLER_7_835 ();
 sg13g2_decap_4 FILLER_7_842 ();
 sg13g2_decap_8 FILLER_7_851 ();
 sg13g2_decap_8 FILLER_7_858 ();
 sg13g2_decap_8 FILLER_7_865 ();
 sg13g2_decap_8 FILLER_7_872 ();
 sg13g2_decap_8 FILLER_7_879 ();
 sg13g2_fill_2 FILLER_7_886 ();
 sg13g2_decap_8 FILLER_7_892 ();
 sg13g2_decap_8 FILLER_7_899 ();
 sg13g2_decap_8 FILLER_7_906 ();
 sg13g2_decap_8 FILLER_7_913 ();
 sg13g2_decap_8 FILLER_7_920 ();
 sg13g2_decap_8 FILLER_7_927 ();
 sg13g2_decap_8 FILLER_7_942 ();
 sg13g2_decap_8 FILLER_7_949 ();
 sg13g2_fill_2 FILLER_7_965 ();
 sg13g2_fill_2 FILLER_7_982 ();
 sg13g2_decap_8 FILLER_7_1002 ();
 sg13g2_decap_8 FILLER_7_1021 ();
 sg13g2_fill_2 FILLER_7_1028 ();
 sg13g2_fill_1 FILLER_7_1034 ();
 sg13g2_fill_1 FILLER_7_1050 ();
 sg13g2_decap_8 FILLER_7_1055 ();
 sg13g2_fill_1 FILLER_7_1062 ();
 sg13g2_decap_8 FILLER_7_1067 ();
 sg13g2_decap_8 FILLER_7_1074 ();
 sg13g2_decap_8 FILLER_7_1081 ();
 sg13g2_decap_8 FILLER_7_1088 ();
 sg13g2_fill_2 FILLER_7_1095 ();
 sg13g2_fill_1 FILLER_7_1097 ();
 sg13g2_decap_8 FILLER_7_1107 ();
 sg13g2_decap_8 FILLER_7_1114 ();
 sg13g2_decap_8 FILLER_7_1121 ();
 sg13g2_decap_8 FILLER_7_1128 ();
 sg13g2_decap_8 FILLER_7_1135 ();
 sg13g2_decap_8 FILLER_7_1142 ();
 sg13g2_decap_8 FILLER_7_1149 ();
 sg13g2_decap_8 FILLER_7_1156 ();
 sg13g2_decap_8 FILLER_7_1163 ();
 sg13g2_decap_8 FILLER_7_1170 ();
 sg13g2_decap_8 FILLER_7_1177 ();
 sg13g2_decap_8 FILLER_7_1184 ();
 sg13g2_decap_8 FILLER_7_1191 ();
 sg13g2_decap_8 FILLER_7_1198 ();
 sg13g2_decap_8 FILLER_7_1205 ();
 sg13g2_decap_8 FILLER_7_1212 ();
 sg13g2_decap_8 FILLER_7_1219 ();
 sg13g2_decap_8 FILLER_7_1226 ();
 sg13g2_decap_8 FILLER_7_1233 ();
 sg13g2_decap_8 FILLER_7_1240 ();
 sg13g2_decap_8 FILLER_7_1247 ();
 sg13g2_decap_8 FILLER_7_1254 ();
 sg13g2_decap_8 FILLER_7_1261 ();
 sg13g2_decap_8 FILLER_7_1271 ();
 sg13g2_decap_8 FILLER_7_1278 ();
 sg13g2_fill_2 FILLER_7_1285 ();
 sg13g2_decap_8 FILLER_7_1291 ();
 sg13g2_decap_4 FILLER_7_1298 ();
 sg13g2_fill_2 FILLER_7_1302 ();
 sg13g2_decap_8 FILLER_7_1309 ();
 sg13g2_decap_8 FILLER_7_1316 ();
 sg13g2_decap_8 FILLER_7_1323 ();
 sg13g2_decap_8 FILLER_7_1330 ();
 sg13g2_decap_8 FILLER_7_1337 ();
 sg13g2_decap_4 FILLER_7_1344 ();
 sg13g2_decap_8 FILLER_7_1357 ();
 sg13g2_decap_8 FILLER_7_1364 ();
 sg13g2_decap_8 FILLER_7_1371 ();
 sg13g2_decap_8 FILLER_7_1393 ();
 sg13g2_decap_8 FILLER_7_1400 ();
 sg13g2_decap_8 FILLER_7_1407 ();
 sg13g2_decap_8 FILLER_7_1414 ();
 sg13g2_decap_4 FILLER_7_1421 ();
 sg13g2_fill_1 FILLER_7_1425 ();
 sg13g2_fill_1 FILLER_7_1432 ();
 sg13g2_fill_1 FILLER_7_1441 ();
 sg13g2_fill_1 FILLER_7_1445 ();
 sg13g2_decap_8 FILLER_7_1453 ();
 sg13g2_decap_8 FILLER_7_1460 ();
 sg13g2_decap_8 FILLER_7_1467 ();
 sg13g2_decap_8 FILLER_7_1474 ();
 sg13g2_decap_8 FILLER_7_1481 ();
 sg13g2_decap_8 FILLER_7_1488 ();
 sg13g2_decap_8 FILLER_7_1495 ();
 sg13g2_decap_8 FILLER_7_1502 ();
 sg13g2_decap_8 FILLER_7_1509 ();
 sg13g2_decap_8 FILLER_7_1516 ();
 sg13g2_decap_8 FILLER_7_1523 ();
 sg13g2_decap_8 FILLER_7_1530 ();
 sg13g2_decap_4 FILLER_7_1537 ();
 sg13g2_fill_2 FILLER_7_1541 ();
 sg13g2_decap_8 FILLER_7_1566 ();
 sg13g2_decap_8 FILLER_7_1573 ();
 sg13g2_decap_8 FILLER_7_1580 ();
 sg13g2_decap_4 FILLER_7_1587 ();
 sg13g2_decap_8 FILLER_7_1603 ();
 sg13g2_fill_1 FILLER_7_1610 ();
 sg13g2_decap_8 FILLER_7_1615 ();
 sg13g2_decap_8 FILLER_7_1622 ();
 sg13g2_decap_8 FILLER_7_1629 ();
 sg13g2_decap_8 FILLER_7_1636 ();
 sg13g2_decap_8 FILLER_7_1643 ();
 sg13g2_decap_8 FILLER_7_1650 ();
 sg13g2_decap_8 FILLER_7_1657 ();
 sg13g2_fill_1 FILLER_7_1664 ();
 sg13g2_decap_8 FILLER_7_1668 ();
 sg13g2_decap_8 FILLER_7_1675 ();
 sg13g2_decap_8 FILLER_7_1682 ();
 sg13g2_decap_8 FILLER_7_1689 ();
 sg13g2_decap_8 FILLER_7_1696 ();
 sg13g2_decap_8 FILLER_7_1703 ();
 sg13g2_decap_8 FILLER_7_1710 ();
 sg13g2_decap_8 FILLER_7_1717 ();
 sg13g2_decap_8 FILLER_7_1724 ();
 sg13g2_decap_8 FILLER_7_1731 ();
 sg13g2_decap_8 FILLER_7_1738 ();
 sg13g2_decap_8 FILLER_7_1745 ();
 sg13g2_decap_4 FILLER_7_1752 ();
 sg13g2_fill_2 FILLER_7_1756 ();
 sg13g2_decap_8 FILLER_7_1766 ();
 sg13g2_decap_8 FILLER_7_1773 ();
 sg13g2_decap_8 FILLER_7_1780 ();
 sg13g2_decap_8 FILLER_7_1787 ();
 sg13g2_decap_8 FILLER_7_1794 ();
 sg13g2_decap_8 FILLER_7_1801 ();
 sg13g2_decap_8 FILLER_7_1808 ();
 sg13g2_decap_8 FILLER_7_1815 ();
 sg13g2_decap_8 FILLER_7_1822 ();
 sg13g2_decap_8 FILLER_7_1829 ();
 sg13g2_decap_8 FILLER_7_1836 ();
 sg13g2_decap_8 FILLER_7_1843 ();
 sg13g2_decap_8 FILLER_7_1850 ();
 sg13g2_decap_8 FILLER_7_1857 ();
 sg13g2_decap_8 FILLER_7_1864 ();
 sg13g2_decap_8 FILLER_7_1871 ();
 sg13g2_decap_8 FILLER_7_1878 ();
 sg13g2_decap_8 FILLER_7_1885 ();
 sg13g2_decap_8 FILLER_7_1892 ();
 sg13g2_decap_8 FILLER_7_1899 ();
 sg13g2_decap_8 FILLER_7_1906 ();
 sg13g2_decap_8 FILLER_7_1913 ();
 sg13g2_decap_8 FILLER_7_1920 ();
 sg13g2_decap_8 FILLER_7_1927 ();
 sg13g2_decap_8 FILLER_7_1934 ();
 sg13g2_decap_8 FILLER_7_1941 ();
 sg13g2_decap_8 FILLER_7_1948 ();
 sg13g2_decap_8 FILLER_7_1955 ();
 sg13g2_decap_8 FILLER_7_1962 ();
 sg13g2_decap_8 FILLER_7_1969 ();
 sg13g2_decap_8 FILLER_7_1976 ();
 sg13g2_decap_8 FILLER_7_1983 ();
 sg13g2_decap_8 FILLER_7_1990 ();
 sg13g2_decap_8 FILLER_7_1997 ();
 sg13g2_decap_8 FILLER_7_2004 ();
 sg13g2_decap_8 FILLER_7_2011 ();
 sg13g2_decap_8 FILLER_7_2018 ();
 sg13g2_decap_8 FILLER_7_2025 ();
 sg13g2_decap_8 FILLER_7_2032 ();
 sg13g2_decap_8 FILLER_7_2039 ();
 sg13g2_decap_8 FILLER_7_2046 ();
 sg13g2_decap_8 FILLER_7_2053 ();
 sg13g2_decap_8 FILLER_7_2060 ();
 sg13g2_decap_8 FILLER_7_2067 ();
 sg13g2_decap_8 FILLER_7_2074 ();
 sg13g2_decap_8 FILLER_7_2081 ();
 sg13g2_decap_8 FILLER_7_2088 ();
 sg13g2_decap_8 FILLER_7_2095 ();
 sg13g2_decap_8 FILLER_7_2102 ();
 sg13g2_decap_8 FILLER_7_2109 ();
 sg13g2_decap_8 FILLER_7_2116 ();
 sg13g2_decap_8 FILLER_7_2123 ();
 sg13g2_decap_8 FILLER_7_2130 ();
 sg13g2_decap_8 FILLER_7_2137 ();
 sg13g2_decap_8 FILLER_7_2144 ();
 sg13g2_decap_8 FILLER_7_2151 ();
 sg13g2_decap_8 FILLER_7_2158 ();
 sg13g2_decap_8 FILLER_7_2165 ();
 sg13g2_decap_8 FILLER_7_2172 ();
 sg13g2_decap_8 FILLER_7_2179 ();
 sg13g2_decap_8 FILLER_7_2186 ();
 sg13g2_decap_8 FILLER_7_2193 ();
 sg13g2_decap_8 FILLER_7_2200 ();
 sg13g2_decap_8 FILLER_7_2207 ();
 sg13g2_decap_8 FILLER_7_2214 ();
 sg13g2_decap_8 FILLER_7_2221 ();
 sg13g2_decap_8 FILLER_7_2228 ();
 sg13g2_decap_8 FILLER_7_2235 ();
 sg13g2_decap_8 FILLER_7_2242 ();
 sg13g2_decap_8 FILLER_7_2249 ();
 sg13g2_decap_8 FILLER_7_2256 ();
 sg13g2_decap_8 FILLER_7_2263 ();
 sg13g2_decap_8 FILLER_7_2270 ();
 sg13g2_decap_8 FILLER_7_2277 ();
 sg13g2_decap_8 FILLER_7_2284 ();
 sg13g2_decap_8 FILLER_7_2291 ();
 sg13g2_decap_8 FILLER_7_2298 ();
 sg13g2_decap_8 FILLER_7_2305 ();
 sg13g2_decap_8 FILLER_7_2312 ();
 sg13g2_decap_8 FILLER_7_2319 ();
 sg13g2_decap_8 FILLER_7_2326 ();
 sg13g2_decap_8 FILLER_7_2333 ();
 sg13g2_decap_8 FILLER_7_2340 ();
 sg13g2_decap_8 FILLER_7_2347 ();
 sg13g2_decap_8 FILLER_7_2354 ();
 sg13g2_decap_8 FILLER_7_2361 ();
 sg13g2_decap_8 FILLER_7_2368 ();
 sg13g2_decap_8 FILLER_7_2375 ();
 sg13g2_decap_8 FILLER_7_2382 ();
 sg13g2_decap_8 FILLER_7_2389 ();
 sg13g2_decap_8 FILLER_7_2396 ();
 sg13g2_decap_8 FILLER_7_2403 ();
 sg13g2_decap_8 FILLER_7_2410 ();
 sg13g2_decap_8 FILLER_7_2417 ();
 sg13g2_decap_8 FILLER_7_2424 ();
 sg13g2_decap_8 FILLER_7_2431 ();
 sg13g2_decap_8 FILLER_7_2438 ();
 sg13g2_decap_8 FILLER_7_2445 ();
 sg13g2_decap_8 FILLER_7_2452 ();
 sg13g2_decap_8 FILLER_7_2459 ();
 sg13g2_decap_8 FILLER_7_2466 ();
 sg13g2_decap_8 FILLER_7_2473 ();
 sg13g2_decap_8 FILLER_7_2480 ();
 sg13g2_decap_8 FILLER_7_2487 ();
 sg13g2_decap_8 FILLER_7_2494 ();
 sg13g2_decap_8 FILLER_7_2501 ();
 sg13g2_decap_8 FILLER_7_2508 ();
 sg13g2_decap_8 FILLER_7_2515 ();
 sg13g2_decap_8 FILLER_7_2522 ();
 sg13g2_decap_8 FILLER_7_2529 ();
 sg13g2_decap_8 FILLER_7_2536 ();
 sg13g2_decap_8 FILLER_7_2543 ();
 sg13g2_decap_8 FILLER_7_2550 ();
 sg13g2_decap_8 FILLER_7_2557 ();
 sg13g2_decap_8 FILLER_7_2564 ();
 sg13g2_decap_8 FILLER_7_2571 ();
 sg13g2_decap_8 FILLER_7_2578 ();
 sg13g2_decap_8 FILLER_7_2585 ();
 sg13g2_decap_8 FILLER_7_2592 ();
 sg13g2_decap_8 FILLER_7_2599 ();
 sg13g2_decap_8 FILLER_7_2606 ();
 sg13g2_decap_8 FILLER_7_2613 ();
 sg13g2_decap_8 FILLER_7_2620 ();
 sg13g2_decap_8 FILLER_7_2627 ();
 sg13g2_decap_8 FILLER_7_2634 ();
 sg13g2_decap_8 FILLER_7_2641 ();
 sg13g2_decap_8 FILLER_7_2648 ();
 sg13g2_decap_8 FILLER_7_2655 ();
 sg13g2_decap_8 FILLER_7_2662 ();
 sg13g2_fill_1 FILLER_7_2669 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_4 FILLER_8_98 ();
 sg13g2_fill_1 FILLER_8_102 ();
 sg13g2_decap_8 FILLER_8_129 ();
 sg13g2_decap_8 FILLER_8_136 ();
 sg13g2_decap_8 FILLER_8_143 ();
 sg13g2_decap_8 FILLER_8_150 ();
 sg13g2_decap_8 FILLER_8_157 ();
 sg13g2_decap_8 FILLER_8_164 ();
 sg13g2_decap_8 FILLER_8_171 ();
 sg13g2_fill_1 FILLER_8_178 ();
 sg13g2_fill_1 FILLER_8_213 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_fill_2 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_4 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_394 ();
 sg13g2_decap_8 FILLER_8_401 ();
 sg13g2_decap_8 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_8_415 ();
 sg13g2_decap_8 FILLER_8_422 ();
 sg13g2_decap_8 FILLER_8_429 ();
 sg13g2_decap_4 FILLER_8_436 ();
 sg13g2_fill_2 FILLER_8_440 ();
 sg13g2_decap_4 FILLER_8_447 ();
 sg13g2_fill_2 FILLER_8_451 ();
 sg13g2_decap_8 FILLER_8_477 ();
 sg13g2_decap_8 FILLER_8_484 ();
 sg13g2_decap_8 FILLER_8_491 ();
 sg13g2_decap_8 FILLER_8_503 ();
 sg13g2_fill_2 FILLER_8_510 ();
 sg13g2_decap_4 FILLER_8_519 ();
 sg13g2_fill_2 FILLER_8_523 ();
 sg13g2_decap_8 FILLER_8_529 ();
 sg13g2_decap_8 FILLER_8_536 ();
 sg13g2_decap_8 FILLER_8_543 ();
 sg13g2_fill_2 FILLER_8_550 ();
 sg13g2_decap_8 FILLER_8_561 ();
 sg13g2_decap_8 FILLER_8_568 ();
 sg13g2_decap_8 FILLER_8_575 ();
 sg13g2_decap_8 FILLER_8_582 ();
 sg13g2_decap_4 FILLER_8_589 ();
 sg13g2_fill_2 FILLER_8_593 ();
 sg13g2_fill_2 FILLER_8_603 ();
 sg13g2_fill_1 FILLER_8_605 ();
 sg13g2_decap_8 FILLER_8_611 ();
 sg13g2_decap_8 FILLER_8_621 ();
 sg13g2_decap_8 FILLER_8_628 ();
 sg13g2_decap_8 FILLER_8_635 ();
 sg13g2_decap_4 FILLER_8_649 ();
 sg13g2_fill_2 FILLER_8_653 ();
 sg13g2_decap_8 FILLER_8_659 ();
 sg13g2_decap_8 FILLER_8_666 ();
 sg13g2_decap_8 FILLER_8_673 ();
 sg13g2_decap_8 FILLER_8_680 ();
 sg13g2_fill_2 FILLER_8_687 ();
 sg13g2_fill_1 FILLER_8_689 ();
 sg13g2_decap_8 FILLER_8_694 ();
 sg13g2_decap_8 FILLER_8_701 ();
 sg13g2_decap_8 FILLER_8_708 ();
 sg13g2_decap_8 FILLER_8_715 ();
 sg13g2_fill_2 FILLER_8_722 ();
 sg13g2_fill_1 FILLER_8_724 ();
 sg13g2_decap_8 FILLER_8_734 ();
 sg13g2_decap_8 FILLER_8_741 ();
 sg13g2_decap_8 FILLER_8_748 ();
 sg13g2_fill_2 FILLER_8_755 ();
 sg13g2_fill_1 FILLER_8_757 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_4 FILLER_8_798 ();
 sg13g2_fill_2 FILLER_8_802 ();
 sg13g2_decap_4 FILLER_8_807 ();
 sg13g2_decap_8 FILLER_8_815 ();
 sg13g2_decap_8 FILLER_8_822 ();
 sg13g2_decap_8 FILLER_8_829 ();
 sg13g2_decap_8 FILLER_8_836 ();
 sg13g2_decap_8 FILLER_8_843 ();
 sg13g2_decap_4 FILLER_8_850 ();
 sg13g2_fill_1 FILLER_8_854 ();
 sg13g2_decap_8 FILLER_8_863 ();
 sg13g2_fill_1 FILLER_8_870 ();
 sg13g2_decap_8 FILLER_8_876 ();
 sg13g2_decap_8 FILLER_8_883 ();
 sg13g2_decap_8 FILLER_8_890 ();
 sg13g2_decap_8 FILLER_8_897 ();
 sg13g2_decap_8 FILLER_8_904 ();
 sg13g2_decap_8 FILLER_8_911 ();
 sg13g2_decap_8 FILLER_8_918 ();
 sg13g2_decap_8 FILLER_8_925 ();
 sg13g2_decap_8 FILLER_8_932 ();
 sg13g2_decap_8 FILLER_8_939 ();
 sg13g2_decap_8 FILLER_8_946 ();
 sg13g2_decap_8 FILLER_8_953 ();
 sg13g2_fill_2 FILLER_8_960 ();
 sg13g2_decap_8 FILLER_8_966 ();
 sg13g2_fill_2 FILLER_8_973 ();
 sg13g2_fill_1 FILLER_8_975 ();
 sg13g2_decap_8 FILLER_8_986 ();
 sg13g2_decap_8 FILLER_8_993 ();
 sg13g2_decap_4 FILLER_8_1000 ();
 sg13g2_fill_2 FILLER_8_1004 ();
 sg13g2_decap_8 FILLER_8_1014 ();
 sg13g2_decap_8 FILLER_8_1021 ();
 sg13g2_decap_4 FILLER_8_1028 ();
 sg13g2_fill_2 FILLER_8_1048 ();
 sg13g2_decap_8 FILLER_8_1054 ();
 sg13g2_decap_8 FILLER_8_1061 ();
 sg13g2_decap_8 FILLER_8_1068 ();
 sg13g2_decap_8 FILLER_8_1075 ();
 sg13g2_fill_1 FILLER_8_1082 ();
 sg13g2_decap_8 FILLER_8_1087 ();
 sg13g2_decap_8 FILLER_8_1102 ();
 sg13g2_decap_8 FILLER_8_1109 ();
 sg13g2_decap_8 FILLER_8_1116 ();
 sg13g2_decap_8 FILLER_8_1123 ();
 sg13g2_decap_8 FILLER_8_1130 ();
 sg13g2_fill_2 FILLER_8_1137 ();
 sg13g2_fill_1 FILLER_8_1139 ();
 sg13g2_decap_8 FILLER_8_1145 ();
 sg13g2_decap_8 FILLER_8_1152 ();
 sg13g2_decap_8 FILLER_8_1159 ();
 sg13g2_decap_8 FILLER_8_1166 ();
 sg13g2_decap_8 FILLER_8_1173 ();
 sg13g2_fill_2 FILLER_8_1180 ();
 sg13g2_decap_8 FILLER_8_1186 ();
 sg13g2_decap_8 FILLER_8_1193 ();
 sg13g2_decap_8 FILLER_8_1200 ();
 sg13g2_decap_8 FILLER_8_1207 ();
 sg13g2_decap_8 FILLER_8_1214 ();
 sg13g2_decap_8 FILLER_8_1221 ();
 sg13g2_decap_4 FILLER_8_1228 ();
 sg13g2_fill_1 FILLER_8_1232 ();
 sg13g2_decap_8 FILLER_8_1250 ();
 sg13g2_fill_2 FILLER_8_1257 ();
 sg13g2_decap_8 FILLER_8_1273 ();
 sg13g2_fill_1 FILLER_8_1280 ();
 sg13g2_decap_8 FILLER_8_1290 ();
 sg13g2_decap_8 FILLER_8_1297 ();
 sg13g2_decap_8 FILLER_8_1304 ();
 sg13g2_decap_8 FILLER_8_1311 ();
 sg13g2_decap_8 FILLER_8_1318 ();
 sg13g2_decap_8 FILLER_8_1325 ();
 sg13g2_decap_8 FILLER_8_1332 ();
 sg13g2_decap_8 FILLER_8_1339 ();
 sg13g2_decap_8 FILLER_8_1346 ();
 sg13g2_decap_8 FILLER_8_1353 ();
 sg13g2_decap_8 FILLER_8_1364 ();
 sg13g2_fill_2 FILLER_8_1375 ();
 sg13g2_fill_1 FILLER_8_1377 ();
 sg13g2_decap_8 FILLER_8_1386 ();
 sg13g2_decap_8 FILLER_8_1393 ();
 sg13g2_decap_8 FILLER_8_1400 ();
 sg13g2_decap_8 FILLER_8_1407 ();
 sg13g2_decap_8 FILLER_8_1414 ();
 sg13g2_decap_8 FILLER_8_1421 ();
 sg13g2_decap_4 FILLER_8_1428 ();
 sg13g2_fill_2 FILLER_8_1432 ();
 sg13g2_fill_1 FILLER_8_1438 ();
 sg13g2_fill_2 FILLER_8_1445 ();
 sg13g2_fill_2 FILLER_8_1450 ();
 sg13g2_fill_1 FILLER_8_1470 ();
 sg13g2_decap_8 FILLER_8_1479 ();
 sg13g2_decap_8 FILLER_8_1486 ();
 sg13g2_decap_8 FILLER_8_1493 ();
 sg13g2_decap_8 FILLER_8_1500 ();
 sg13g2_decap_4 FILLER_8_1507 ();
 sg13g2_decap_8 FILLER_8_1517 ();
 sg13g2_decap_8 FILLER_8_1524 ();
 sg13g2_decap_8 FILLER_8_1531 ();
 sg13g2_decap_4 FILLER_8_1538 ();
 sg13g2_fill_1 FILLER_8_1542 ();
 sg13g2_decap_8 FILLER_8_1549 ();
 sg13g2_decap_8 FILLER_8_1556 ();
 sg13g2_decap_8 FILLER_8_1563 ();
 sg13g2_fill_1 FILLER_8_1570 ();
 sg13g2_decap_8 FILLER_8_1580 ();
 sg13g2_decap_4 FILLER_8_1587 ();
 sg13g2_decap_8 FILLER_8_1595 ();
 sg13g2_fill_1 FILLER_8_1602 ();
 sg13g2_decap_8 FILLER_8_1611 ();
 sg13g2_fill_2 FILLER_8_1618 ();
 sg13g2_decap_8 FILLER_8_1624 ();
 sg13g2_decap_8 FILLER_8_1631 ();
 sg13g2_decap_8 FILLER_8_1642 ();
 sg13g2_decap_8 FILLER_8_1649 ();
 sg13g2_decap_8 FILLER_8_1656 ();
 sg13g2_fill_2 FILLER_8_1663 ();
 sg13g2_decap_8 FILLER_8_1680 ();
 sg13g2_decap_4 FILLER_8_1687 ();
 sg13g2_fill_2 FILLER_8_1691 ();
 sg13g2_decap_8 FILLER_8_1701 ();
 sg13g2_decap_8 FILLER_8_1708 ();
 sg13g2_decap_8 FILLER_8_1715 ();
 sg13g2_decap_8 FILLER_8_1722 ();
 sg13g2_decap_8 FILLER_8_1729 ();
 sg13g2_decap_8 FILLER_8_1736 ();
 sg13g2_decap_8 FILLER_8_1743 ();
 sg13g2_decap_8 FILLER_8_1750 ();
 sg13g2_decap_8 FILLER_8_1757 ();
 sg13g2_decap_8 FILLER_8_1764 ();
 sg13g2_decap_8 FILLER_8_1771 ();
 sg13g2_decap_8 FILLER_8_1778 ();
 sg13g2_decap_8 FILLER_8_1785 ();
 sg13g2_decap_8 FILLER_8_1792 ();
 sg13g2_decap_8 FILLER_8_1799 ();
 sg13g2_decap_8 FILLER_8_1806 ();
 sg13g2_decap_8 FILLER_8_1813 ();
 sg13g2_decap_8 FILLER_8_1820 ();
 sg13g2_decap_8 FILLER_8_1827 ();
 sg13g2_decap_8 FILLER_8_1834 ();
 sg13g2_decap_8 FILLER_8_1841 ();
 sg13g2_decap_8 FILLER_8_1848 ();
 sg13g2_decap_8 FILLER_8_1855 ();
 sg13g2_decap_8 FILLER_8_1862 ();
 sg13g2_decap_8 FILLER_8_1869 ();
 sg13g2_decap_8 FILLER_8_1876 ();
 sg13g2_decap_8 FILLER_8_1883 ();
 sg13g2_decap_8 FILLER_8_1890 ();
 sg13g2_decap_8 FILLER_8_1897 ();
 sg13g2_decap_8 FILLER_8_1904 ();
 sg13g2_decap_8 FILLER_8_1911 ();
 sg13g2_decap_8 FILLER_8_1918 ();
 sg13g2_decap_8 FILLER_8_1925 ();
 sg13g2_decap_8 FILLER_8_1932 ();
 sg13g2_decap_8 FILLER_8_1939 ();
 sg13g2_decap_8 FILLER_8_1946 ();
 sg13g2_decap_8 FILLER_8_1953 ();
 sg13g2_decap_8 FILLER_8_1960 ();
 sg13g2_decap_8 FILLER_8_1967 ();
 sg13g2_decap_8 FILLER_8_1974 ();
 sg13g2_decap_8 FILLER_8_1981 ();
 sg13g2_decap_8 FILLER_8_1988 ();
 sg13g2_decap_8 FILLER_8_1995 ();
 sg13g2_decap_8 FILLER_8_2002 ();
 sg13g2_decap_8 FILLER_8_2009 ();
 sg13g2_decap_8 FILLER_8_2016 ();
 sg13g2_decap_8 FILLER_8_2023 ();
 sg13g2_decap_8 FILLER_8_2030 ();
 sg13g2_decap_8 FILLER_8_2037 ();
 sg13g2_decap_8 FILLER_8_2044 ();
 sg13g2_decap_8 FILLER_8_2051 ();
 sg13g2_decap_8 FILLER_8_2058 ();
 sg13g2_decap_8 FILLER_8_2065 ();
 sg13g2_decap_8 FILLER_8_2072 ();
 sg13g2_decap_8 FILLER_8_2079 ();
 sg13g2_decap_8 FILLER_8_2086 ();
 sg13g2_decap_8 FILLER_8_2093 ();
 sg13g2_decap_8 FILLER_8_2100 ();
 sg13g2_decap_8 FILLER_8_2107 ();
 sg13g2_decap_8 FILLER_8_2114 ();
 sg13g2_decap_8 FILLER_8_2121 ();
 sg13g2_decap_8 FILLER_8_2128 ();
 sg13g2_decap_8 FILLER_8_2135 ();
 sg13g2_decap_8 FILLER_8_2142 ();
 sg13g2_decap_8 FILLER_8_2149 ();
 sg13g2_decap_8 FILLER_8_2156 ();
 sg13g2_decap_8 FILLER_8_2163 ();
 sg13g2_decap_8 FILLER_8_2170 ();
 sg13g2_decap_8 FILLER_8_2177 ();
 sg13g2_decap_8 FILLER_8_2184 ();
 sg13g2_decap_8 FILLER_8_2191 ();
 sg13g2_decap_8 FILLER_8_2198 ();
 sg13g2_decap_8 FILLER_8_2205 ();
 sg13g2_decap_8 FILLER_8_2212 ();
 sg13g2_decap_8 FILLER_8_2219 ();
 sg13g2_decap_8 FILLER_8_2226 ();
 sg13g2_decap_8 FILLER_8_2233 ();
 sg13g2_decap_8 FILLER_8_2240 ();
 sg13g2_decap_8 FILLER_8_2247 ();
 sg13g2_decap_8 FILLER_8_2254 ();
 sg13g2_decap_8 FILLER_8_2261 ();
 sg13g2_decap_8 FILLER_8_2268 ();
 sg13g2_decap_8 FILLER_8_2275 ();
 sg13g2_decap_8 FILLER_8_2282 ();
 sg13g2_decap_8 FILLER_8_2289 ();
 sg13g2_decap_8 FILLER_8_2296 ();
 sg13g2_decap_8 FILLER_8_2303 ();
 sg13g2_decap_8 FILLER_8_2310 ();
 sg13g2_decap_8 FILLER_8_2317 ();
 sg13g2_decap_8 FILLER_8_2324 ();
 sg13g2_decap_8 FILLER_8_2331 ();
 sg13g2_decap_8 FILLER_8_2338 ();
 sg13g2_decap_8 FILLER_8_2345 ();
 sg13g2_decap_8 FILLER_8_2352 ();
 sg13g2_decap_8 FILLER_8_2359 ();
 sg13g2_decap_8 FILLER_8_2366 ();
 sg13g2_decap_8 FILLER_8_2373 ();
 sg13g2_decap_8 FILLER_8_2380 ();
 sg13g2_decap_8 FILLER_8_2387 ();
 sg13g2_decap_8 FILLER_8_2394 ();
 sg13g2_decap_8 FILLER_8_2401 ();
 sg13g2_decap_8 FILLER_8_2408 ();
 sg13g2_decap_8 FILLER_8_2415 ();
 sg13g2_decap_8 FILLER_8_2422 ();
 sg13g2_decap_8 FILLER_8_2429 ();
 sg13g2_decap_8 FILLER_8_2436 ();
 sg13g2_decap_8 FILLER_8_2443 ();
 sg13g2_decap_8 FILLER_8_2450 ();
 sg13g2_decap_8 FILLER_8_2457 ();
 sg13g2_decap_8 FILLER_8_2464 ();
 sg13g2_decap_8 FILLER_8_2471 ();
 sg13g2_decap_8 FILLER_8_2478 ();
 sg13g2_decap_8 FILLER_8_2485 ();
 sg13g2_decap_8 FILLER_8_2492 ();
 sg13g2_decap_8 FILLER_8_2499 ();
 sg13g2_decap_8 FILLER_8_2506 ();
 sg13g2_decap_8 FILLER_8_2513 ();
 sg13g2_decap_8 FILLER_8_2520 ();
 sg13g2_decap_8 FILLER_8_2527 ();
 sg13g2_decap_8 FILLER_8_2534 ();
 sg13g2_decap_8 FILLER_8_2541 ();
 sg13g2_decap_8 FILLER_8_2548 ();
 sg13g2_decap_8 FILLER_8_2555 ();
 sg13g2_decap_8 FILLER_8_2562 ();
 sg13g2_decap_8 FILLER_8_2569 ();
 sg13g2_decap_8 FILLER_8_2576 ();
 sg13g2_decap_8 FILLER_8_2583 ();
 sg13g2_decap_8 FILLER_8_2590 ();
 sg13g2_decap_8 FILLER_8_2597 ();
 sg13g2_decap_8 FILLER_8_2604 ();
 sg13g2_decap_8 FILLER_8_2611 ();
 sg13g2_decap_8 FILLER_8_2618 ();
 sg13g2_decap_8 FILLER_8_2625 ();
 sg13g2_decap_8 FILLER_8_2632 ();
 sg13g2_decap_8 FILLER_8_2639 ();
 sg13g2_decap_8 FILLER_8_2646 ();
 sg13g2_decap_8 FILLER_8_2653 ();
 sg13g2_decap_8 FILLER_8_2660 ();
 sg13g2_fill_2 FILLER_8_2667 ();
 sg13g2_fill_1 FILLER_8_2669 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_fill_2 FILLER_9_357 ();
 sg13g2_fill_1 FILLER_9_359 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_418 ();
 sg13g2_decap_8 FILLER_9_425 ();
 sg13g2_decap_8 FILLER_9_432 ();
 sg13g2_decap_8 FILLER_9_439 ();
 sg13g2_fill_2 FILLER_9_446 ();
 sg13g2_decap_8 FILLER_9_451 ();
 sg13g2_decap_8 FILLER_9_458 ();
 sg13g2_decap_8 FILLER_9_465 ();
 sg13g2_decap_8 FILLER_9_472 ();
 sg13g2_decap_8 FILLER_9_479 ();
 sg13g2_decap_8 FILLER_9_486 ();
 sg13g2_decap_8 FILLER_9_493 ();
 sg13g2_decap_8 FILLER_9_512 ();
 sg13g2_decap_8 FILLER_9_519 ();
 sg13g2_decap_8 FILLER_9_526 ();
 sg13g2_decap_8 FILLER_9_533 ();
 sg13g2_decap_8 FILLER_9_540 ();
 sg13g2_decap_8 FILLER_9_547 ();
 sg13g2_decap_8 FILLER_9_554 ();
 sg13g2_decap_8 FILLER_9_561 ();
 sg13g2_decap_8 FILLER_9_568 ();
 sg13g2_decap_8 FILLER_9_603 ();
 sg13g2_decap_8 FILLER_9_615 ();
 sg13g2_decap_8 FILLER_9_622 ();
 sg13g2_decap_8 FILLER_9_629 ();
 sg13g2_decap_8 FILLER_9_636 ();
 sg13g2_decap_8 FILLER_9_643 ();
 sg13g2_decap_8 FILLER_9_650 ();
 sg13g2_decap_8 FILLER_9_657 ();
 sg13g2_decap_8 FILLER_9_664 ();
 sg13g2_decap_4 FILLER_9_671 ();
 sg13g2_fill_2 FILLER_9_675 ();
 sg13g2_decap_8 FILLER_9_696 ();
 sg13g2_decap_8 FILLER_9_703 ();
 sg13g2_decap_8 FILLER_9_710 ();
 sg13g2_decap_8 FILLER_9_717 ();
 sg13g2_decap_4 FILLER_9_724 ();
 sg13g2_decap_8 FILLER_9_740 ();
 sg13g2_decap_8 FILLER_9_747 ();
 sg13g2_decap_8 FILLER_9_754 ();
 sg13g2_fill_1 FILLER_9_761 ();
 sg13g2_decap_8 FILLER_9_766 ();
 sg13g2_decap_8 FILLER_9_773 ();
 sg13g2_decap_8 FILLER_9_780 ();
 sg13g2_decap_8 FILLER_9_787 ();
 sg13g2_decap_8 FILLER_9_794 ();
 sg13g2_decap_8 FILLER_9_801 ();
 sg13g2_decap_8 FILLER_9_808 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_833 ();
 sg13g2_decap_8 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_859 ();
 sg13g2_decap_8 FILLER_9_866 ();
 sg13g2_decap_8 FILLER_9_873 ();
 sg13g2_decap_8 FILLER_9_880 ();
 sg13g2_fill_1 FILLER_9_887 ();
 sg13g2_decap_8 FILLER_9_893 ();
 sg13g2_decap_8 FILLER_9_900 ();
 sg13g2_decap_8 FILLER_9_907 ();
 sg13g2_decap_8 FILLER_9_914 ();
 sg13g2_decap_8 FILLER_9_921 ();
 sg13g2_decap_4 FILLER_9_928 ();
 sg13g2_decap_8 FILLER_9_935 ();
 sg13g2_decap_8 FILLER_9_942 ();
 sg13g2_decap_8 FILLER_9_949 ();
 sg13g2_decap_4 FILLER_9_956 ();
 sg13g2_fill_2 FILLER_9_960 ();
 sg13g2_decap_8 FILLER_9_972 ();
 sg13g2_decap_8 FILLER_9_985 ();
 sg13g2_decap_8 FILLER_9_992 ();
 sg13g2_fill_1 FILLER_9_1011 ();
 sg13g2_decap_8 FILLER_9_1018 ();
 sg13g2_decap_8 FILLER_9_1025 ();
 sg13g2_decap_8 FILLER_9_1032 ();
 sg13g2_decap_4 FILLER_9_1039 ();
 sg13g2_fill_1 FILLER_9_1043 ();
 sg13g2_fill_2 FILLER_9_1048 ();
 sg13g2_fill_1 FILLER_9_1050 ();
 sg13g2_decap_8 FILLER_9_1055 ();
 sg13g2_decap_8 FILLER_9_1062 ();
 sg13g2_decap_8 FILLER_9_1069 ();
 sg13g2_decap_8 FILLER_9_1076 ();
 sg13g2_fill_1 FILLER_9_1083 ();
 sg13g2_decap_8 FILLER_9_1089 ();
 sg13g2_fill_2 FILLER_9_1096 ();
 sg13g2_fill_2 FILLER_9_1101 ();
 sg13g2_decap_8 FILLER_9_1107 ();
 sg13g2_decap_8 FILLER_9_1114 ();
 sg13g2_decap_4 FILLER_9_1121 ();
 sg13g2_decap_4 FILLER_9_1129 ();
 sg13g2_fill_2 FILLER_9_1133 ();
 sg13g2_fill_1 FILLER_9_1150 ();
 sg13g2_decap_8 FILLER_9_1159 ();
 sg13g2_decap_8 FILLER_9_1166 ();
 sg13g2_decap_8 FILLER_9_1173 ();
 sg13g2_decap_8 FILLER_9_1180 ();
 sg13g2_decap_8 FILLER_9_1187 ();
 sg13g2_decap_8 FILLER_9_1194 ();
 sg13g2_decap_8 FILLER_9_1201 ();
 sg13g2_decap_8 FILLER_9_1208 ();
 sg13g2_decap_8 FILLER_9_1215 ();
 sg13g2_decap_8 FILLER_9_1222 ();
 sg13g2_decap_8 FILLER_9_1229 ();
 sg13g2_fill_2 FILLER_9_1236 ();
 sg13g2_fill_1 FILLER_9_1238 ();
 sg13g2_decap_8 FILLER_9_1248 ();
 sg13g2_decap_8 FILLER_9_1270 ();
 sg13g2_decap_8 FILLER_9_1277 ();
 sg13g2_decap_8 FILLER_9_1284 ();
 sg13g2_fill_2 FILLER_9_1291 ();
 sg13g2_decap_8 FILLER_9_1298 ();
 sg13g2_decap_8 FILLER_9_1305 ();
 sg13g2_decap_8 FILLER_9_1312 ();
 sg13g2_decap_8 FILLER_9_1319 ();
 sg13g2_decap_8 FILLER_9_1326 ();
 sg13g2_decap_8 FILLER_9_1333 ();
 sg13g2_decap_8 FILLER_9_1340 ();
 sg13g2_decap_8 FILLER_9_1347 ();
 sg13g2_decap_8 FILLER_9_1354 ();
 sg13g2_decap_8 FILLER_9_1361 ();
 sg13g2_decap_4 FILLER_9_1368 ();
 sg13g2_decap_4 FILLER_9_1377 ();
 sg13g2_fill_1 FILLER_9_1381 ();
 sg13g2_decap_8 FILLER_9_1391 ();
 sg13g2_decap_8 FILLER_9_1398 ();
 sg13g2_decap_8 FILLER_9_1405 ();
 sg13g2_decap_8 FILLER_9_1412 ();
 sg13g2_decap_8 FILLER_9_1419 ();
 sg13g2_decap_4 FILLER_9_1426 ();
 sg13g2_fill_2 FILLER_9_1430 ();
 sg13g2_fill_2 FILLER_9_1450 ();
 sg13g2_decap_8 FILLER_9_1460 ();
 sg13g2_decap_8 FILLER_9_1467 ();
 sg13g2_fill_1 FILLER_9_1474 ();
 sg13g2_fill_1 FILLER_9_1478 ();
 sg13g2_decap_4 FILLER_9_1483 ();
 sg13g2_decap_8 FILLER_9_1495 ();
 sg13g2_decap_8 FILLER_9_1502 ();
 sg13g2_decap_8 FILLER_9_1509 ();
 sg13g2_decap_8 FILLER_9_1516 ();
 sg13g2_decap_8 FILLER_9_1523 ();
 sg13g2_decap_8 FILLER_9_1530 ();
 sg13g2_decap_8 FILLER_9_1555 ();
 sg13g2_fill_2 FILLER_9_1562 ();
 sg13g2_fill_1 FILLER_9_1564 ();
 sg13g2_decap_8 FILLER_9_1582 ();
 sg13g2_decap_8 FILLER_9_1589 ();
 sg13g2_decap_4 FILLER_9_1596 ();
 sg13g2_decap_8 FILLER_9_1604 ();
 sg13g2_decap_8 FILLER_9_1611 ();
 sg13g2_decap_8 FILLER_9_1618 ();
 sg13g2_decap_8 FILLER_9_1625 ();
 sg13g2_decap_4 FILLER_9_1632 ();
 sg13g2_decap_8 FILLER_9_1647 ();
 sg13g2_fill_1 FILLER_9_1654 ();
 sg13g2_decap_8 FILLER_9_1677 ();
 sg13g2_decap_8 FILLER_9_1684 ();
 sg13g2_decap_8 FILLER_9_1691 ();
 sg13g2_decap_8 FILLER_9_1698 ();
 sg13g2_decap_8 FILLER_9_1705 ();
 sg13g2_decap_8 FILLER_9_1712 ();
 sg13g2_decap_8 FILLER_9_1719 ();
 sg13g2_decap_8 FILLER_9_1726 ();
 sg13g2_decap_8 FILLER_9_1733 ();
 sg13g2_decap_8 FILLER_9_1740 ();
 sg13g2_decap_4 FILLER_9_1747 ();
 sg13g2_decap_8 FILLER_9_1754 ();
 sg13g2_decap_8 FILLER_9_1761 ();
 sg13g2_decap_8 FILLER_9_1768 ();
 sg13g2_decap_8 FILLER_9_1775 ();
 sg13g2_decap_8 FILLER_9_1782 ();
 sg13g2_decap_8 FILLER_9_1789 ();
 sg13g2_decap_8 FILLER_9_1796 ();
 sg13g2_decap_8 FILLER_9_1803 ();
 sg13g2_decap_8 FILLER_9_1810 ();
 sg13g2_decap_8 FILLER_9_1817 ();
 sg13g2_decap_8 FILLER_9_1824 ();
 sg13g2_decap_8 FILLER_9_1831 ();
 sg13g2_decap_8 FILLER_9_1838 ();
 sg13g2_decap_8 FILLER_9_1845 ();
 sg13g2_decap_8 FILLER_9_1852 ();
 sg13g2_decap_8 FILLER_9_1859 ();
 sg13g2_decap_8 FILLER_9_1866 ();
 sg13g2_decap_8 FILLER_9_1873 ();
 sg13g2_decap_8 FILLER_9_1880 ();
 sg13g2_decap_8 FILLER_9_1887 ();
 sg13g2_decap_8 FILLER_9_1894 ();
 sg13g2_decap_8 FILLER_9_1901 ();
 sg13g2_decap_8 FILLER_9_1908 ();
 sg13g2_decap_8 FILLER_9_1915 ();
 sg13g2_decap_8 FILLER_9_1922 ();
 sg13g2_decap_8 FILLER_9_1929 ();
 sg13g2_decap_8 FILLER_9_1936 ();
 sg13g2_decap_8 FILLER_9_1943 ();
 sg13g2_decap_8 FILLER_9_1950 ();
 sg13g2_decap_8 FILLER_9_1957 ();
 sg13g2_decap_8 FILLER_9_1964 ();
 sg13g2_decap_8 FILLER_9_1971 ();
 sg13g2_decap_8 FILLER_9_1978 ();
 sg13g2_decap_8 FILLER_9_1985 ();
 sg13g2_decap_8 FILLER_9_1992 ();
 sg13g2_decap_8 FILLER_9_1999 ();
 sg13g2_decap_8 FILLER_9_2006 ();
 sg13g2_decap_8 FILLER_9_2013 ();
 sg13g2_decap_8 FILLER_9_2020 ();
 sg13g2_decap_8 FILLER_9_2027 ();
 sg13g2_decap_8 FILLER_9_2034 ();
 sg13g2_decap_8 FILLER_9_2041 ();
 sg13g2_decap_8 FILLER_9_2048 ();
 sg13g2_decap_8 FILLER_9_2055 ();
 sg13g2_decap_8 FILLER_9_2062 ();
 sg13g2_decap_8 FILLER_9_2069 ();
 sg13g2_decap_8 FILLER_9_2076 ();
 sg13g2_decap_8 FILLER_9_2083 ();
 sg13g2_decap_8 FILLER_9_2090 ();
 sg13g2_decap_8 FILLER_9_2097 ();
 sg13g2_decap_8 FILLER_9_2104 ();
 sg13g2_decap_8 FILLER_9_2111 ();
 sg13g2_decap_8 FILLER_9_2118 ();
 sg13g2_decap_8 FILLER_9_2125 ();
 sg13g2_decap_8 FILLER_9_2132 ();
 sg13g2_decap_8 FILLER_9_2139 ();
 sg13g2_decap_8 FILLER_9_2146 ();
 sg13g2_decap_8 FILLER_9_2153 ();
 sg13g2_decap_8 FILLER_9_2160 ();
 sg13g2_decap_8 FILLER_9_2167 ();
 sg13g2_decap_8 FILLER_9_2174 ();
 sg13g2_decap_8 FILLER_9_2181 ();
 sg13g2_decap_8 FILLER_9_2188 ();
 sg13g2_decap_8 FILLER_9_2195 ();
 sg13g2_decap_8 FILLER_9_2202 ();
 sg13g2_decap_8 FILLER_9_2209 ();
 sg13g2_decap_8 FILLER_9_2216 ();
 sg13g2_decap_8 FILLER_9_2223 ();
 sg13g2_decap_8 FILLER_9_2230 ();
 sg13g2_decap_8 FILLER_9_2237 ();
 sg13g2_decap_8 FILLER_9_2244 ();
 sg13g2_decap_8 FILLER_9_2251 ();
 sg13g2_decap_8 FILLER_9_2258 ();
 sg13g2_decap_8 FILLER_9_2265 ();
 sg13g2_decap_8 FILLER_9_2272 ();
 sg13g2_decap_8 FILLER_9_2279 ();
 sg13g2_decap_8 FILLER_9_2286 ();
 sg13g2_decap_8 FILLER_9_2293 ();
 sg13g2_decap_8 FILLER_9_2300 ();
 sg13g2_decap_8 FILLER_9_2307 ();
 sg13g2_decap_8 FILLER_9_2314 ();
 sg13g2_decap_8 FILLER_9_2321 ();
 sg13g2_decap_8 FILLER_9_2328 ();
 sg13g2_decap_8 FILLER_9_2335 ();
 sg13g2_decap_8 FILLER_9_2342 ();
 sg13g2_decap_8 FILLER_9_2349 ();
 sg13g2_decap_8 FILLER_9_2356 ();
 sg13g2_decap_8 FILLER_9_2363 ();
 sg13g2_decap_8 FILLER_9_2370 ();
 sg13g2_decap_8 FILLER_9_2377 ();
 sg13g2_decap_8 FILLER_9_2384 ();
 sg13g2_decap_8 FILLER_9_2391 ();
 sg13g2_decap_8 FILLER_9_2398 ();
 sg13g2_decap_8 FILLER_9_2405 ();
 sg13g2_decap_8 FILLER_9_2412 ();
 sg13g2_decap_8 FILLER_9_2419 ();
 sg13g2_decap_8 FILLER_9_2426 ();
 sg13g2_decap_8 FILLER_9_2433 ();
 sg13g2_decap_8 FILLER_9_2440 ();
 sg13g2_decap_8 FILLER_9_2447 ();
 sg13g2_decap_8 FILLER_9_2454 ();
 sg13g2_decap_8 FILLER_9_2461 ();
 sg13g2_decap_8 FILLER_9_2468 ();
 sg13g2_decap_8 FILLER_9_2475 ();
 sg13g2_decap_8 FILLER_9_2482 ();
 sg13g2_decap_8 FILLER_9_2489 ();
 sg13g2_decap_8 FILLER_9_2496 ();
 sg13g2_decap_8 FILLER_9_2503 ();
 sg13g2_decap_8 FILLER_9_2510 ();
 sg13g2_decap_8 FILLER_9_2517 ();
 sg13g2_decap_8 FILLER_9_2524 ();
 sg13g2_decap_8 FILLER_9_2531 ();
 sg13g2_decap_8 FILLER_9_2538 ();
 sg13g2_decap_8 FILLER_9_2545 ();
 sg13g2_decap_8 FILLER_9_2552 ();
 sg13g2_decap_8 FILLER_9_2559 ();
 sg13g2_decap_8 FILLER_9_2566 ();
 sg13g2_decap_8 FILLER_9_2573 ();
 sg13g2_decap_8 FILLER_9_2580 ();
 sg13g2_decap_8 FILLER_9_2587 ();
 sg13g2_decap_8 FILLER_9_2594 ();
 sg13g2_decap_8 FILLER_9_2601 ();
 sg13g2_decap_8 FILLER_9_2608 ();
 sg13g2_decap_8 FILLER_9_2615 ();
 sg13g2_decap_8 FILLER_9_2622 ();
 sg13g2_decap_8 FILLER_9_2629 ();
 sg13g2_decap_8 FILLER_9_2636 ();
 sg13g2_decap_8 FILLER_9_2643 ();
 sg13g2_decap_8 FILLER_9_2650 ();
 sg13g2_decap_8 FILLER_9_2657 ();
 sg13g2_decap_4 FILLER_9_2664 ();
 sg13g2_fill_2 FILLER_9_2668 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_4 FILLER_10_238 ();
 sg13g2_fill_2 FILLER_10_242 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_455 ();
 sg13g2_decap_8 FILLER_10_462 ();
 sg13g2_decap_8 FILLER_10_469 ();
 sg13g2_decap_8 FILLER_10_476 ();
 sg13g2_fill_1 FILLER_10_483 ();
 sg13g2_decap_4 FILLER_10_488 ();
 sg13g2_fill_2 FILLER_10_492 ();
 sg13g2_decap_8 FILLER_10_513 ();
 sg13g2_decap_8 FILLER_10_520 ();
 sg13g2_decap_8 FILLER_10_527 ();
 sg13g2_decap_8 FILLER_10_534 ();
 sg13g2_decap_8 FILLER_10_541 ();
 sg13g2_decap_8 FILLER_10_548 ();
 sg13g2_decap_8 FILLER_10_555 ();
 sg13g2_decap_8 FILLER_10_562 ();
 sg13g2_decap_8 FILLER_10_569 ();
 sg13g2_decap_8 FILLER_10_576 ();
 sg13g2_decap_8 FILLER_10_583 ();
 sg13g2_decap_4 FILLER_10_590 ();
 sg13g2_fill_1 FILLER_10_594 ();
 sg13g2_decap_8 FILLER_10_607 ();
 sg13g2_decap_4 FILLER_10_614 ();
 sg13g2_decap_8 FILLER_10_621 ();
 sg13g2_decap_8 FILLER_10_628 ();
 sg13g2_decap_8 FILLER_10_635 ();
 sg13g2_decap_8 FILLER_10_642 ();
 sg13g2_decap_8 FILLER_10_649 ();
 sg13g2_decap_8 FILLER_10_656 ();
 sg13g2_decap_8 FILLER_10_663 ();
 sg13g2_decap_8 FILLER_10_670 ();
 sg13g2_decap_8 FILLER_10_677 ();
 sg13g2_fill_2 FILLER_10_684 ();
 sg13g2_decap_8 FILLER_10_690 ();
 sg13g2_decap_8 FILLER_10_697 ();
 sg13g2_decap_8 FILLER_10_704 ();
 sg13g2_decap_8 FILLER_10_711 ();
 sg13g2_decap_8 FILLER_10_718 ();
 sg13g2_decap_8 FILLER_10_725 ();
 sg13g2_decap_8 FILLER_10_732 ();
 sg13g2_decap_8 FILLER_10_739 ();
 sg13g2_decap_8 FILLER_10_746 ();
 sg13g2_decap_4 FILLER_10_753 ();
 sg13g2_fill_2 FILLER_10_757 ();
 sg13g2_fill_1 FILLER_10_769 ();
 sg13g2_decap_8 FILLER_10_779 ();
 sg13g2_decap_8 FILLER_10_786 ();
 sg13g2_decap_8 FILLER_10_793 ();
 sg13g2_decap_8 FILLER_10_800 ();
 sg13g2_decap_8 FILLER_10_807 ();
 sg13g2_decap_8 FILLER_10_814 ();
 sg13g2_decap_8 FILLER_10_821 ();
 sg13g2_decap_8 FILLER_10_828 ();
 sg13g2_decap_8 FILLER_10_835 ();
 sg13g2_decap_4 FILLER_10_842 ();
 sg13g2_decap_4 FILLER_10_851 ();
 sg13g2_fill_1 FILLER_10_855 ();
 sg13g2_decap_8 FILLER_10_871 ();
 sg13g2_decap_8 FILLER_10_878 ();
 sg13g2_decap_8 FILLER_10_885 ();
 sg13g2_fill_1 FILLER_10_892 ();
 sg13g2_decap_8 FILLER_10_898 ();
 sg13g2_decap_8 FILLER_10_905 ();
 sg13g2_decap_8 FILLER_10_912 ();
 sg13g2_decap_8 FILLER_10_919 ();
 sg13g2_fill_2 FILLER_10_926 ();
 sg13g2_fill_1 FILLER_10_928 ();
 sg13g2_decap_8 FILLER_10_937 ();
 sg13g2_decap_8 FILLER_10_944 ();
 sg13g2_decap_4 FILLER_10_951 ();
 sg13g2_fill_2 FILLER_10_955 ();
 sg13g2_decap_8 FILLER_10_964 ();
 sg13g2_decap_8 FILLER_10_971 ();
 sg13g2_decap_4 FILLER_10_978 ();
 sg13g2_fill_1 FILLER_10_982 ();
 sg13g2_decap_8 FILLER_10_988 ();
 sg13g2_decap_8 FILLER_10_995 ();
 sg13g2_decap_4 FILLER_10_1002 ();
 sg13g2_fill_2 FILLER_10_1006 ();
 sg13g2_decap_8 FILLER_10_1012 ();
 sg13g2_decap_8 FILLER_10_1019 ();
 sg13g2_decap_8 FILLER_10_1026 ();
 sg13g2_decap_8 FILLER_10_1033 ();
 sg13g2_decap_8 FILLER_10_1040 ();
 sg13g2_decap_8 FILLER_10_1047 ();
 sg13g2_decap_8 FILLER_10_1054 ();
 sg13g2_decap_8 FILLER_10_1061 ();
 sg13g2_decap_8 FILLER_10_1068 ();
 sg13g2_decap_8 FILLER_10_1075 ();
 sg13g2_decap_8 FILLER_10_1082 ();
 sg13g2_decap_8 FILLER_10_1089 ();
 sg13g2_decap_8 FILLER_10_1096 ();
 sg13g2_decap_8 FILLER_10_1103 ();
 sg13g2_decap_8 FILLER_10_1110 ();
 sg13g2_decap_8 FILLER_10_1117 ();
 sg13g2_decap_8 FILLER_10_1124 ();
 sg13g2_decap_8 FILLER_10_1131 ();
 sg13g2_decap_4 FILLER_10_1138 ();
 sg13g2_fill_2 FILLER_10_1142 ();
 sg13g2_fill_1 FILLER_10_1147 ();
 sg13g2_decap_8 FILLER_10_1155 ();
 sg13g2_decap_8 FILLER_10_1162 ();
 sg13g2_decap_8 FILLER_10_1169 ();
 sg13g2_decap_4 FILLER_10_1176 ();
 sg13g2_decap_8 FILLER_10_1188 ();
 sg13g2_fill_2 FILLER_10_1195 ();
 sg13g2_fill_1 FILLER_10_1197 ();
 sg13g2_fill_1 FILLER_10_1218 ();
 sg13g2_decap_8 FILLER_10_1231 ();
 sg13g2_decap_8 FILLER_10_1238 ();
 sg13g2_decap_8 FILLER_10_1245 ();
 sg13g2_fill_1 FILLER_10_1252 ();
 sg13g2_fill_2 FILLER_10_1256 ();
 sg13g2_decap_8 FILLER_10_1262 ();
 sg13g2_decap_8 FILLER_10_1269 ();
 sg13g2_decap_8 FILLER_10_1276 ();
 sg13g2_fill_1 FILLER_10_1283 ();
 sg13g2_decap_8 FILLER_10_1287 ();
 sg13g2_fill_1 FILLER_10_1294 ();
 sg13g2_decap_8 FILLER_10_1310 ();
 sg13g2_decap_8 FILLER_10_1317 ();
 sg13g2_decap_8 FILLER_10_1324 ();
 sg13g2_decap_4 FILLER_10_1331 ();
 sg13g2_decap_8 FILLER_10_1339 ();
 sg13g2_decap_8 FILLER_10_1346 ();
 sg13g2_decap_8 FILLER_10_1353 ();
 sg13g2_decap_8 FILLER_10_1360 ();
 sg13g2_decap_8 FILLER_10_1367 ();
 sg13g2_decap_8 FILLER_10_1374 ();
 sg13g2_decap_8 FILLER_10_1381 ();
 sg13g2_decap_8 FILLER_10_1388 ();
 sg13g2_decap_8 FILLER_10_1395 ();
 sg13g2_decap_8 FILLER_10_1402 ();
 sg13g2_decap_8 FILLER_10_1409 ();
 sg13g2_decap_8 FILLER_10_1416 ();
 sg13g2_decap_8 FILLER_10_1423 ();
 sg13g2_decap_8 FILLER_10_1430 ();
 sg13g2_decap_8 FILLER_10_1437 ();
 sg13g2_decap_8 FILLER_10_1444 ();
 sg13g2_decap_8 FILLER_10_1451 ();
 sg13g2_decap_8 FILLER_10_1458 ();
 sg13g2_decap_8 FILLER_10_1465 ();
 sg13g2_decap_8 FILLER_10_1472 ();
 sg13g2_decap_8 FILLER_10_1479 ();
 sg13g2_decap_8 FILLER_10_1486 ();
 sg13g2_decap_8 FILLER_10_1493 ();
 sg13g2_decap_8 FILLER_10_1500 ();
 sg13g2_decap_8 FILLER_10_1507 ();
 sg13g2_decap_8 FILLER_10_1514 ();
 sg13g2_decap_8 FILLER_10_1521 ();
 sg13g2_decap_8 FILLER_10_1528 ();
 sg13g2_decap_8 FILLER_10_1535 ();
 sg13g2_fill_1 FILLER_10_1542 ();
 sg13g2_decap_8 FILLER_10_1551 ();
 sg13g2_decap_8 FILLER_10_1558 ();
 sg13g2_decap_4 FILLER_10_1565 ();
 sg13g2_fill_2 FILLER_10_1569 ();
 sg13g2_decap_8 FILLER_10_1575 ();
 sg13g2_decap_8 FILLER_10_1582 ();
 sg13g2_decap_8 FILLER_10_1589 ();
 sg13g2_decap_8 FILLER_10_1596 ();
 sg13g2_decap_8 FILLER_10_1603 ();
 sg13g2_decap_8 FILLER_10_1610 ();
 sg13g2_decap_8 FILLER_10_1617 ();
 sg13g2_fill_2 FILLER_10_1624 ();
 sg13g2_fill_1 FILLER_10_1626 ();
 sg13g2_decap_8 FILLER_10_1633 ();
 sg13g2_fill_1 FILLER_10_1640 ();
 sg13g2_decap_4 FILLER_10_1660 ();
 sg13g2_fill_1 FILLER_10_1664 ();
 sg13g2_fill_1 FILLER_10_1668 ();
 sg13g2_decap_8 FILLER_10_1693 ();
 sg13g2_decap_8 FILLER_10_1700 ();
 sg13g2_decap_8 FILLER_10_1707 ();
 sg13g2_decap_8 FILLER_10_1714 ();
 sg13g2_decap_8 FILLER_10_1721 ();
 sg13g2_decap_8 FILLER_10_1728 ();
 sg13g2_decap_8 FILLER_10_1735 ();
 sg13g2_decap_8 FILLER_10_1742 ();
 sg13g2_fill_2 FILLER_10_1749 ();
 sg13g2_decap_8 FILLER_10_1768 ();
 sg13g2_decap_8 FILLER_10_1775 ();
 sg13g2_fill_2 FILLER_10_1782 ();
 sg13g2_decap_8 FILLER_10_1805 ();
 sg13g2_decap_8 FILLER_10_1812 ();
 sg13g2_decap_8 FILLER_10_1819 ();
 sg13g2_decap_8 FILLER_10_1826 ();
 sg13g2_decap_8 FILLER_10_1833 ();
 sg13g2_decap_8 FILLER_10_1840 ();
 sg13g2_decap_8 FILLER_10_1847 ();
 sg13g2_decap_8 FILLER_10_1854 ();
 sg13g2_decap_8 FILLER_10_1861 ();
 sg13g2_decap_8 FILLER_10_1868 ();
 sg13g2_decap_8 FILLER_10_1875 ();
 sg13g2_decap_8 FILLER_10_1882 ();
 sg13g2_decap_8 FILLER_10_1889 ();
 sg13g2_decap_8 FILLER_10_1896 ();
 sg13g2_decap_8 FILLER_10_1903 ();
 sg13g2_decap_8 FILLER_10_1910 ();
 sg13g2_decap_8 FILLER_10_1917 ();
 sg13g2_decap_8 FILLER_10_1924 ();
 sg13g2_decap_8 FILLER_10_1931 ();
 sg13g2_decap_8 FILLER_10_1938 ();
 sg13g2_decap_8 FILLER_10_1945 ();
 sg13g2_decap_8 FILLER_10_1952 ();
 sg13g2_decap_8 FILLER_10_1959 ();
 sg13g2_decap_8 FILLER_10_1966 ();
 sg13g2_decap_8 FILLER_10_1973 ();
 sg13g2_decap_8 FILLER_10_1980 ();
 sg13g2_decap_8 FILLER_10_1987 ();
 sg13g2_decap_8 FILLER_10_1994 ();
 sg13g2_decap_8 FILLER_10_2001 ();
 sg13g2_decap_8 FILLER_10_2008 ();
 sg13g2_decap_8 FILLER_10_2015 ();
 sg13g2_decap_8 FILLER_10_2022 ();
 sg13g2_decap_8 FILLER_10_2029 ();
 sg13g2_decap_8 FILLER_10_2036 ();
 sg13g2_decap_8 FILLER_10_2043 ();
 sg13g2_decap_8 FILLER_10_2050 ();
 sg13g2_decap_8 FILLER_10_2057 ();
 sg13g2_decap_8 FILLER_10_2064 ();
 sg13g2_decap_8 FILLER_10_2071 ();
 sg13g2_decap_8 FILLER_10_2078 ();
 sg13g2_decap_8 FILLER_10_2085 ();
 sg13g2_decap_8 FILLER_10_2092 ();
 sg13g2_decap_8 FILLER_10_2099 ();
 sg13g2_decap_8 FILLER_10_2106 ();
 sg13g2_decap_8 FILLER_10_2113 ();
 sg13g2_decap_8 FILLER_10_2120 ();
 sg13g2_decap_8 FILLER_10_2127 ();
 sg13g2_decap_8 FILLER_10_2134 ();
 sg13g2_decap_8 FILLER_10_2141 ();
 sg13g2_decap_8 FILLER_10_2148 ();
 sg13g2_decap_8 FILLER_10_2155 ();
 sg13g2_decap_8 FILLER_10_2162 ();
 sg13g2_decap_8 FILLER_10_2169 ();
 sg13g2_decap_8 FILLER_10_2176 ();
 sg13g2_decap_8 FILLER_10_2183 ();
 sg13g2_decap_8 FILLER_10_2190 ();
 sg13g2_decap_8 FILLER_10_2197 ();
 sg13g2_decap_8 FILLER_10_2204 ();
 sg13g2_decap_8 FILLER_10_2211 ();
 sg13g2_decap_8 FILLER_10_2218 ();
 sg13g2_decap_8 FILLER_10_2225 ();
 sg13g2_decap_8 FILLER_10_2232 ();
 sg13g2_decap_8 FILLER_10_2239 ();
 sg13g2_decap_8 FILLER_10_2246 ();
 sg13g2_decap_8 FILLER_10_2253 ();
 sg13g2_decap_8 FILLER_10_2260 ();
 sg13g2_decap_8 FILLER_10_2267 ();
 sg13g2_decap_8 FILLER_10_2274 ();
 sg13g2_decap_8 FILLER_10_2281 ();
 sg13g2_decap_8 FILLER_10_2288 ();
 sg13g2_decap_8 FILLER_10_2295 ();
 sg13g2_decap_8 FILLER_10_2302 ();
 sg13g2_decap_8 FILLER_10_2309 ();
 sg13g2_decap_8 FILLER_10_2316 ();
 sg13g2_decap_8 FILLER_10_2323 ();
 sg13g2_decap_8 FILLER_10_2330 ();
 sg13g2_decap_8 FILLER_10_2337 ();
 sg13g2_decap_8 FILLER_10_2344 ();
 sg13g2_decap_8 FILLER_10_2351 ();
 sg13g2_decap_8 FILLER_10_2358 ();
 sg13g2_decap_8 FILLER_10_2365 ();
 sg13g2_decap_8 FILLER_10_2372 ();
 sg13g2_decap_8 FILLER_10_2379 ();
 sg13g2_decap_8 FILLER_10_2386 ();
 sg13g2_decap_8 FILLER_10_2393 ();
 sg13g2_decap_8 FILLER_10_2400 ();
 sg13g2_decap_8 FILLER_10_2407 ();
 sg13g2_decap_8 FILLER_10_2414 ();
 sg13g2_decap_8 FILLER_10_2421 ();
 sg13g2_decap_8 FILLER_10_2428 ();
 sg13g2_decap_8 FILLER_10_2435 ();
 sg13g2_decap_8 FILLER_10_2442 ();
 sg13g2_decap_8 FILLER_10_2449 ();
 sg13g2_decap_8 FILLER_10_2456 ();
 sg13g2_decap_8 FILLER_10_2463 ();
 sg13g2_decap_8 FILLER_10_2470 ();
 sg13g2_decap_8 FILLER_10_2477 ();
 sg13g2_decap_8 FILLER_10_2484 ();
 sg13g2_decap_8 FILLER_10_2491 ();
 sg13g2_decap_8 FILLER_10_2498 ();
 sg13g2_decap_8 FILLER_10_2505 ();
 sg13g2_decap_8 FILLER_10_2512 ();
 sg13g2_decap_8 FILLER_10_2519 ();
 sg13g2_decap_8 FILLER_10_2526 ();
 sg13g2_decap_8 FILLER_10_2533 ();
 sg13g2_decap_8 FILLER_10_2540 ();
 sg13g2_decap_8 FILLER_10_2547 ();
 sg13g2_decap_8 FILLER_10_2554 ();
 sg13g2_decap_8 FILLER_10_2561 ();
 sg13g2_decap_8 FILLER_10_2568 ();
 sg13g2_decap_8 FILLER_10_2575 ();
 sg13g2_decap_8 FILLER_10_2582 ();
 sg13g2_decap_8 FILLER_10_2589 ();
 sg13g2_decap_8 FILLER_10_2596 ();
 sg13g2_decap_8 FILLER_10_2603 ();
 sg13g2_decap_8 FILLER_10_2610 ();
 sg13g2_decap_8 FILLER_10_2617 ();
 sg13g2_decap_8 FILLER_10_2624 ();
 sg13g2_decap_8 FILLER_10_2631 ();
 sg13g2_decap_8 FILLER_10_2638 ();
 sg13g2_decap_8 FILLER_10_2645 ();
 sg13g2_decap_8 FILLER_10_2652 ();
 sg13g2_decap_8 FILLER_10_2659 ();
 sg13g2_decap_4 FILLER_10_2666 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_fill_2 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_76 ();
 sg13g2_decap_8 FILLER_11_83 ();
 sg13g2_decap_8 FILLER_11_90 ();
 sg13g2_decap_8 FILLER_11_97 ();
 sg13g2_decap_8 FILLER_11_104 ();
 sg13g2_decap_8 FILLER_11_111 ();
 sg13g2_decap_8 FILLER_11_118 ();
 sg13g2_decap_8 FILLER_11_125 ();
 sg13g2_decap_8 FILLER_11_132 ();
 sg13g2_decap_8 FILLER_11_139 ();
 sg13g2_decap_8 FILLER_11_146 ();
 sg13g2_decap_8 FILLER_11_153 ();
 sg13g2_decap_8 FILLER_11_160 ();
 sg13g2_decap_8 FILLER_11_167 ();
 sg13g2_decap_8 FILLER_11_174 ();
 sg13g2_decap_8 FILLER_11_181 ();
 sg13g2_decap_8 FILLER_11_188 ();
 sg13g2_decap_8 FILLER_11_195 ();
 sg13g2_decap_8 FILLER_11_202 ();
 sg13g2_decap_8 FILLER_11_209 ();
 sg13g2_decap_8 FILLER_11_216 ();
 sg13g2_decap_8 FILLER_11_223 ();
 sg13g2_decap_8 FILLER_11_230 ();
 sg13g2_decap_8 FILLER_11_237 ();
 sg13g2_decap_8 FILLER_11_244 ();
 sg13g2_decap_8 FILLER_11_251 ();
 sg13g2_decap_8 FILLER_11_258 ();
 sg13g2_decap_4 FILLER_11_265 ();
 sg13g2_fill_2 FILLER_11_269 ();
 sg13g2_decap_8 FILLER_11_275 ();
 sg13g2_decap_8 FILLER_11_282 ();
 sg13g2_decap_8 FILLER_11_289 ();
 sg13g2_decap_8 FILLER_11_296 ();
 sg13g2_decap_8 FILLER_11_303 ();
 sg13g2_decap_8 FILLER_11_310 ();
 sg13g2_decap_8 FILLER_11_317 ();
 sg13g2_decap_4 FILLER_11_324 ();
 sg13g2_decap_8 FILLER_11_353 ();
 sg13g2_decap_8 FILLER_11_360 ();
 sg13g2_decap_8 FILLER_11_367 ();
 sg13g2_decap_8 FILLER_11_374 ();
 sg13g2_decap_8 FILLER_11_381 ();
 sg13g2_decap_8 FILLER_11_388 ();
 sg13g2_decap_8 FILLER_11_395 ();
 sg13g2_decap_8 FILLER_11_402 ();
 sg13g2_decap_8 FILLER_11_409 ();
 sg13g2_fill_2 FILLER_11_416 ();
 sg13g2_fill_1 FILLER_11_418 ();
 sg13g2_decap_8 FILLER_11_423 ();
 sg13g2_decap_8 FILLER_11_430 ();
 sg13g2_decap_8 FILLER_11_437 ();
 sg13g2_decap_8 FILLER_11_444 ();
 sg13g2_fill_2 FILLER_11_451 ();
 sg13g2_fill_1 FILLER_11_453 ();
 sg13g2_decap_8 FILLER_11_457 ();
 sg13g2_decap_8 FILLER_11_464 ();
 sg13g2_fill_2 FILLER_11_471 ();
 sg13g2_decap_8 FILLER_11_477 ();
 sg13g2_decap_8 FILLER_11_484 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_decap_8 FILLER_11_518 ();
 sg13g2_decap_8 FILLER_11_525 ();
 sg13g2_decap_8 FILLER_11_532 ();
 sg13g2_decap_4 FILLER_11_539 ();
 sg13g2_fill_1 FILLER_11_543 ();
 sg13g2_decap_8 FILLER_11_548 ();
 sg13g2_decap_8 FILLER_11_555 ();
 sg13g2_decap_4 FILLER_11_562 ();
 sg13g2_fill_2 FILLER_11_566 ();
 sg13g2_decap_8 FILLER_11_583 ();
 sg13g2_decap_8 FILLER_11_590 ();
 sg13g2_decap_8 FILLER_11_597 ();
 sg13g2_decap_8 FILLER_11_604 ();
 sg13g2_decap_8 FILLER_11_611 ();
 sg13g2_decap_8 FILLER_11_622 ();
 sg13g2_decap_8 FILLER_11_629 ();
 sg13g2_decap_8 FILLER_11_636 ();
 sg13g2_decap_8 FILLER_11_648 ();
 sg13g2_decap_8 FILLER_11_655 ();
 sg13g2_fill_1 FILLER_11_662 ();
 sg13g2_decap_8 FILLER_11_667 ();
 sg13g2_decap_8 FILLER_11_674 ();
 sg13g2_decap_8 FILLER_11_681 ();
 sg13g2_decap_8 FILLER_11_688 ();
 sg13g2_decap_8 FILLER_11_695 ();
 sg13g2_decap_8 FILLER_11_702 ();
 sg13g2_decap_8 FILLER_11_709 ();
 sg13g2_decap_8 FILLER_11_716 ();
 sg13g2_decap_8 FILLER_11_723 ();
 sg13g2_decap_8 FILLER_11_730 ();
 sg13g2_decap_8 FILLER_11_737 ();
 sg13g2_decap_8 FILLER_11_744 ();
 sg13g2_decap_4 FILLER_11_751 ();
 sg13g2_fill_1 FILLER_11_755 ();
 sg13g2_fill_1 FILLER_11_766 ();
 sg13g2_decap_4 FILLER_11_779 ();
 sg13g2_decap_8 FILLER_11_798 ();
 sg13g2_decap_8 FILLER_11_805 ();
 sg13g2_decap_8 FILLER_11_812 ();
 sg13g2_decap_8 FILLER_11_819 ();
 sg13g2_decap_8 FILLER_11_830 ();
 sg13g2_decap_8 FILLER_11_837 ();
 sg13g2_decap_8 FILLER_11_844 ();
 sg13g2_fill_2 FILLER_11_851 ();
 sg13g2_fill_1 FILLER_11_853 ();
 sg13g2_decap_8 FILLER_11_863 ();
 sg13g2_decap_8 FILLER_11_870 ();
 sg13g2_decap_8 FILLER_11_877 ();
 sg13g2_decap_8 FILLER_11_884 ();
 sg13g2_decap_8 FILLER_11_891 ();
 sg13g2_decap_8 FILLER_11_898 ();
 sg13g2_decap_8 FILLER_11_905 ();
 sg13g2_decap_8 FILLER_11_912 ();
 sg13g2_decap_8 FILLER_11_919 ();
 sg13g2_decap_4 FILLER_11_926 ();
 sg13g2_fill_2 FILLER_11_930 ();
 sg13g2_decap_8 FILLER_11_935 ();
 sg13g2_decap_8 FILLER_11_942 ();
 sg13g2_decap_8 FILLER_11_949 ();
 sg13g2_decap_4 FILLER_11_956 ();
 sg13g2_fill_2 FILLER_11_963 ();
 sg13g2_fill_1 FILLER_11_965 ();
 sg13g2_decap_8 FILLER_11_971 ();
 sg13g2_decap_8 FILLER_11_978 ();
 sg13g2_decap_8 FILLER_11_985 ();
 sg13g2_decap_8 FILLER_11_992 ();
 sg13g2_fill_2 FILLER_11_999 ();
 sg13g2_fill_2 FILLER_11_1006 ();
 sg13g2_decap_8 FILLER_11_1014 ();
 sg13g2_decap_8 FILLER_11_1021 ();
 sg13g2_decap_8 FILLER_11_1028 ();
 sg13g2_decap_8 FILLER_11_1035 ();
 sg13g2_decap_8 FILLER_11_1042 ();
 sg13g2_fill_2 FILLER_11_1049 ();
 sg13g2_fill_1 FILLER_11_1051 ();
 sg13g2_decap_8 FILLER_11_1067 ();
 sg13g2_decap_8 FILLER_11_1074 ();
 sg13g2_decap_8 FILLER_11_1081 ();
 sg13g2_decap_8 FILLER_11_1088 ();
 sg13g2_decap_8 FILLER_11_1095 ();
 sg13g2_decap_8 FILLER_11_1102 ();
 sg13g2_decap_8 FILLER_11_1109 ();
 sg13g2_decap_8 FILLER_11_1116 ();
 sg13g2_decap_8 FILLER_11_1127 ();
 sg13g2_decap_8 FILLER_11_1134 ();
 sg13g2_fill_2 FILLER_11_1141 ();
 sg13g2_fill_2 FILLER_11_1149 ();
 sg13g2_decap_8 FILLER_11_1154 ();
 sg13g2_decap_8 FILLER_11_1161 ();
 sg13g2_decap_8 FILLER_11_1168 ();
 sg13g2_decap_8 FILLER_11_1175 ();
 sg13g2_decap_8 FILLER_11_1182 ();
 sg13g2_decap_8 FILLER_11_1189 ();
 sg13g2_decap_8 FILLER_11_1196 ();
 sg13g2_fill_1 FILLER_11_1203 ();
 sg13g2_fill_1 FILLER_11_1215 ();
 sg13g2_decap_8 FILLER_11_1223 ();
 sg13g2_decap_8 FILLER_11_1230 ();
 sg13g2_decap_8 FILLER_11_1237 ();
 sg13g2_decap_8 FILLER_11_1244 ();
 sg13g2_fill_2 FILLER_11_1251 ();
 sg13g2_decap_8 FILLER_11_1257 ();
 sg13g2_decap_8 FILLER_11_1264 ();
 sg13g2_fill_1 FILLER_11_1271 ();
 sg13g2_decap_4 FILLER_11_1287 ();
 sg13g2_fill_2 FILLER_11_1291 ();
 sg13g2_fill_2 FILLER_11_1306 ();
 sg13g2_decap_8 FILLER_11_1323 ();
 sg13g2_decap_8 FILLER_11_1330 ();
 sg13g2_decap_8 FILLER_11_1337 ();
 sg13g2_decap_8 FILLER_11_1344 ();
 sg13g2_decap_8 FILLER_11_1351 ();
 sg13g2_decap_8 FILLER_11_1358 ();
 sg13g2_fill_2 FILLER_11_1365 ();
 sg13g2_fill_1 FILLER_11_1367 ();
 sg13g2_decap_8 FILLER_11_1371 ();
 sg13g2_decap_4 FILLER_11_1378 ();
 sg13g2_fill_1 FILLER_11_1382 ();
 sg13g2_decap_8 FILLER_11_1388 ();
 sg13g2_decap_8 FILLER_11_1395 ();
 sg13g2_decap_8 FILLER_11_1402 ();
 sg13g2_decap_8 FILLER_11_1409 ();
 sg13g2_fill_1 FILLER_11_1416 ();
 sg13g2_fill_1 FILLER_11_1420 ();
 sg13g2_decap_8 FILLER_11_1427 ();
 sg13g2_fill_2 FILLER_11_1434 ();
 sg13g2_decap_8 FILLER_11_1442 ();
 sg13g2_decap_8 FILLER_11_1449 ();
 sg13g2_decap_8 FILLER_11_1456 ();
 sg13g2_decap_8 FILLER_11_1463 ();
 sg13g2_decap_8 FILLER_11_1470 ();
 sg13g2_decap_8 FILLER_11_1477 ();
 sg13g2_decap_8 FILLER_11_1484 ();
 sg13g2_decap_8 FILLER_11_1491 ();
 sg13g2_decap_8 FILLER_11_1498 ();
 sg13g2_decap_8 FILLER_11_1505 ();
 sg13g2_decap_8 FILLER_11_1512 ();
 sg13g2_decap_8 FILLER_11_1519 ();
 sg13g2_decap_8 FILLER_11_1526 ();
 sg13g2_decap_8 FILLER_11_1533 ();
 sg13g2_decap_8 FILLER_11_1540 ();
 sg13g2_decap_8 FILLER_11_1547 ();
 sg13g2_decap_4 FILLER_11_1554 ();
 sg13g2_fill_1 FILLER_11_1570 ();
 sg13g2_decap_8 FILLER_11_1586 ();
 sg13g2_decap_8 FILLER_11_1593 ();
 sg13g2_fill_2 FILLER_11_1600 ();
 sg13g2_fill_1 FILLER_11_1602 ();
 sg13g2_decap_8 FILLER_11_1607 ();
 sg13g2_decap_8 FILLER_11_1614 ();
 sg13g2_decap_8 FILLER_11_1638 ();
 sg13g2_decap_8 FILLER_11_1645 ();
 sg13g2_decap_8 FILLER_11_1652 ();
 sg13g2_decap_8 FILLER_11_1659 ();
 sg13g2_decap_8 FILLER_11_1673 ();
 sg13g2_decap_8 FILLER_11_1680 ();
 sg13g2_decap_8 FILLER_11_1687 ();
 sg13g2_fill_2 FILLER_11_1694 ();
 sg13g2_fill_1 FILLER_11_1696 ();
 sg13g2_decap_8 FILLER_11_1701 ();
 sg13g2_decap_4 FILLER_11_1708 ();
 sg13g2_fill_2 FILLER_11_1712 ();
 sg13g2_decap_8 FILLER_11_1723 ();
 sg13g2_decap_8 FILLER_11_1730 ();
 sg13g2_decap_8 FILLER_11_1737 ();
 sg13g2_decap_8 FILLER_11_1744 ();
 sg13g2_decap_8 FILLER_11_1751 ();
 sg13g2_decap_8 FILLER_11_1758 ();
 sg13g2_decap_8 FILLER_11_1765 ();
 sg13g2_decap_4 FILLER_11_1772 ();
 sg13g2_fill_2 FILLER_11_1776 ();
 sg13g2_decap_8 FILLER_11_1795 ();
 sg13g2_fill_2 FILLER_11_1802 ();
 sg13g2_fill_1 FILLER_11_1804 ();
 sg13g2_decap_8 FILLER_11_1818 ();
 sg13g2_decap_8 FILLER_11_1825 ();
 sg13g2_decap_8 FILLER_11_1832 ();
 sg13g2_decap_8 FILLER_11_1839 ();
 sg13g2_decap_8 FILLER_11_1846 ();
 sg13g2_decap_8 FILLER_11_1853 ();
 sg13g2_decap_8 FILLER_11_1860 ();
 sg13g2_decap_8 FILLER_11_1867 ();
 sg13g2_decap_8 FILLER_11_1874 ();
 sg13g2_decap_8 FILLER_11_1881 ();
 sg13g2_decap_8 FILLER_11_1888 ();
 sg13g2_decap_8 FILLER_11_1895 ();
 sg13g2_decap_8 FILLER_11_1902 ();
 sg13g2_decap_8 FILLER_11_1909 ();
 sg13g2_decap_8 FILLER_11_1916 ();
 sg13g2_decap_8 FILLER_11_1923 ();
 sg13g2_decap_8 FILLER_11_1930 ();
 sg13g2_decap_8 FILLER_11_1937 ();
 sg13g2_decap_8 FILLER_11_1944 ();
 sg13g2_decap_8 FILLER_11_1951 ();
 sg13g2_decap_8 FILLER_11_1958 ();
 sg13g2_decap_8 FILLER_11_1965 ();
 sg13g2_decap_8 FILLER_11_1972 ();
 sg13g2_decap_8 FILLER_11_1979 ();
 sg13g2_decap_8 FILLER_11_1986 ();
 sg13g2_decap_8 FILLER_11_1993 ();
 sg13g2_decap_8 FILLER_11_2000 ();
 sg13g2_decap_8 FILLER_11_2007 ();
 sg13g2_decap_8 FILLER_11_2014 ();
 sg13g2_decap_8 FILLER_11_2021 ();
 sg13g2_decap_8 FILLER_11_2028 ();
 sg13g2_decap_8 FILLER_11_2035 ();
 sg13g2_decap_8 FILLER_11_2042 ();
 sg13g2_decap_8 FILLER_11_2049 ();
 sg13g2_decap_8 FILLER_11_2056 ();
 sg13g2_decap_8 FILLER_11_2063 ();
 sg13g2_decap_8 FILLER_11_2070 ();
 sg13g2_decap_8 FILLER_11_2077 ();
 sg13g2_decap_8 FILLER_11_2084 ();
 sg13g2_decap_8 FILLER_11_2091 ();
 sg13g2_decap_8 FILLER_11_2098 ();
 sg13g2_decap_8 FILLER_11_2105 ();
 sg13g2_decap_8 FILLER_11_2112 ();
 sg13g2_decap_8 FILLER_11_2119 ();
 sg13g2_decap_8 FILLER_11_2126 ();
 sg13g2_decap_8 FILLER_11_2133 ();
 sg13g2_decap_8 FILLER_11_2140 ();
 sg13g2_decap_8 FILLER_11_2147 ();
 sg13g2_decap_8 FILLER_11_2154 ();
 sg13g2_decap_8 FILLER_11_2161 ();
 sg13g2_decap_8 FILLER_11_2168 ();
 sg13g2_decap_8 FILLER_11_2175 ();
 sg13g2_decap_8 FILLER_11_2182 ();
 sg13g2_decap_8 FILLER_11_2189 ();
 sg13g2_decap_8 FILLER_11_2196 ();
 sg13g2_decap_8 FILLER_11_2203 ();
 sg13g2_decap_8 FILLER_11_2210 ();
 sg13g2_decap_8 FILLER_11_2217 ();
 sg13g2_decap_8 FILLER_11_2224 ();
 sg13g2_decap_8 FILLER_11_2231 ();
 sg13g2_decap_8 FILLER_11_2238 ();
 sg13g2_decap_8 FILLER_11_2245 ();
 sg13g2_decap_8 FILLER_11_2252 ();
 sg13g2_decap_8 FILLER_11_2259 ();
 sg13g2_decap_8 FILLER_11_2266 ();
 sg13g2_decap_8 FILLER_11_2273 ();
 sg13g2_decap_8 FILLER_11_2280 ();
 sg13g2_decap_8 FILLER_11_2287 ();
 sg13g2_decap_8 FILLER_11_2294 ();
 sg13g2_decap_8 FILLER_11_2301 ();
 sg13g2_decap_8 FILLER_11_2308 ();
 sg13g2_decap_8 FILLER_11_2315 ();
 sg13g2_decap_8 FILLER_11_2322 ();
 sg13g2_decap_8 FILLER_11_2329 ();
 sg13g2_decap_8 FILLER_11_2336 ();
 sg13g2_decap_8 FILLER_11_2343 ();
 sg13g2_decap_8 FILLER_11_2350 ();
 sg13g2_decap_8 FILLER_11_2357 ();
 sg13g2_decap_8 FILLER_11_2364 ();
 sg13g2_decap_8 FILLER_11_2371 ();
 sg13g2_decap_8 FILLER_11_2378 ();
 sg13g2_decap_8 FILLER_11_2385 ();
 sg13g2_decap_8 FILLER_11_2392 ();
 sg13g2_decap_8 FILLER_11_2399 ();
 sg13g2_decap_8 FILLER_11_2406 ();
 sg13g2_decap_8 FILLER_11_2413 ();
 sg13g2_decap_8 FILLER_11_2420 ();
 sg13g2_decap_8 FILLER_11_2427 ();
 sg13g2_decap_8 FILLER_11_2434 ();
 sg13g2_decap_8 FILLER_11_2441 ();
 sg13g2_decap_8 FILLER_11_2448 ();
 sg13g2_decap_8 FILLER_11_2455 ();
 sg13g2_decap_8 FILLER_11_2462 ();
 sg13g2_decap_8 FILLER_11_2469 ();
 sg13g2_decap_8 FILLER_11_2476 ();
 sg13g2_decap_8 FILLER_11_2483 ();
 sg13g2_decap_8 FILLER_11_2490 ();
 sg13g2_decap_8 FILLER_11_2497 ();
 sg13g2_decap_8 FILLER_11_2504 ();
 sg13g2_decap_8 FILLER_11_2511 ();
 sg13g2_decap_8 FILLER_11_2518 ();
 sg13g2_decap_8 FILLER_11_2525 ();
 sg13g2_decap_8 FILLER_11_2532 ();
 sg13g2_decap_8 FILLER_11_2539 ();
 sg13g2_decap_8 FILLER_11_2546 ();
 sg13g2_decap_8 FILLER_11_2553 ();
 sg13g2_decap_8 FILLER_11_2560 ();
 sg13g2_decap_8 FILLER_11_2567 ();
 sg13g2_decap_8 FILLER_11_2574 ();
 sg13g2_decap_8 FILLER_11_2581 ();
 sg13g2_decap_8 FILLER_11_2588 ();
 sg13g2_decap_8 FILLER_11_2595 ();
 sg13g2_decap_8 FILLER_11_2602 ();
 sg13g2_decap_8 FILLER_11_2609 ();
 sg13g2_decap_8 FILLER_11_2616 ();
 sg13g2_decap_8 FILLER_11_2623 ();
 sg13g2_decap_8 FILLER_11_2630 ();
 sg13g2_decap_8 FILLER_11_2637 ();
 sg13g2_decap_8 FILLER_11_2644 ();
 sg13g2_decap_8 FILLER_11_2651 ();
 sg13g2_decap_8 FILLER_11_2658 ();
 sg13g2_decap_4 FILLER_11_2665 ();
 sg13g2_fill_1 FILLER_11_2669 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_fill_2 FILLER_12_63 ();
 sg13g2_fill_1 FILLER_12_65 ();
 sg13g2_decap_8 FILLER_12_92 ();
 sg13g2_decap_8 FILLER_12_99 ();
 sg13g2_decap_8 FILLER_12_106 ();
 sg13g2_decap_8 FILLER_12_113 ();
 sg13g2_decap_8 FILLER_12_120 ();
 sg13g2_decap_8 FILLER_12_139 ();
 sg13g2_decap_8 FILLER_12_146 ();
 sg13g2_decap_8 FILLER_12_153 ();
 sg13g2_decap_8 FILLER_12_160 ();
 sg13g2_fill_2 FILLER_12_167 ();
 sg13g2_fill_1 FILLER_12_169 ();
 sg13g2_decap_8 FILLER_12_174 ();
 sg13g2_decap_8 FILLER_12_181 ();
 sg13g2_decap_8 FILLER_12_188 ();
 sg13g2_decap_8 FILLER_12_195 ();
 sg13g2_decap_8 FILLER_12_202 ();
 sg13g2_decap_8 FILLER_12_209 ();
 sg13g2_decap_8 FILLER_12_216 ();
 sg13g2_decap_8 FILLER_12_223 ();
 sg13g2_decap_8 FILLER_12_230 ();
 sg13g2_decap_8 FILLER_12_237 ();
 sg13g2_decap_8 FILLER_12_244 ();
 sg13g2_decap_8 FILLER_12_251 ();
 sg13g2_decap_4 FILLER_12_258 ();
 sg13g2_fill_2 FILLER_12_262 ();
 sg13g2_decap_8 FILLER_12_290 ();
 sg13g2_decap_8 FILLER_12_297 ();
 sg13g2_decap_8 FILLER_12_304 ();
 sg13g2_decap_8 FILLER_12_311 ();
 sg13g2_decap_8 FILLER_12_318 ();
 sg13g2_decap_8 FILLER_12_325 ();
 sg13g2_decap_8 FILLER_12_332 ();
 sg13g2_decap_8 FILLER_12_339 ();
 sg13g2_decap_8 FILLER_12_346 ();
 sg13g2_decap_8 FILLER_12_353 ();
 sg13g2_fill_2 FILLER_12_360 ();
 sg13g2_fill_1 FILLER_12_362 ();
 sg13g2_decap_8 FILLER_12_367 ();
 sg13g2_decap_8 FILLER_12_374 ();
 sg13g2_decap_8 FILLER_12_381 ();
 sg13g2_decap_8 FILLER_12_388 ();
 sg13g2_decap_8 FILLER_12_395 ();
 sg13g2_decap_8 FILLER_12_402 ();
 sg13g2_decap_8 FILLER_12_409 ();
 sg13g2_decap_8 FILLER_12_416 ();
 sg13g2_decap_4 FILLER_12_423 ();
 sg13g2_fill_1 FILLER_12_427 ();
 sg13g2_fill_2 FILLER_12_433 ();
 sg13g2_fill_1 FILLER_12_435 ();
 sg13g2_decap_8 FILLER_12_440 ();
 sg13g2_fill_1 FILLER_12_447 ();
 sg13g2_fill_2 FILLER_12_452 ();
 sg13g2_fill_2 FILLER_12_477 ();
 sg13g2_fill_1 FILLER_12_479 ();
 sg13g2_decap_8 FILLER_12_485 ();
 sg13g2_decap_8 FILLER_12_492 ();
 sg13g2_decap_4 FILLER_12_499 ();
 sg13g2_decap_8 FILLER_12_512 ();
 sg13g2_decap_8 FILLER_12_519 ();
 sg13g2_decap_8 FILLER_12_526 ();
 sg13g2_decap_8 FILLER_12_533 ();
 sg13g2_decap_4 FILLER_12_540 ();
 sg13g2_decap_8 FILLER_12_548 ();
 sg13g2_decap_8 FILLER_12_555 ();
 sg13g2_decap_8 FILLER_12_562 ();
 sg13g2_fill_2 FILLER_12_569 ();
 sg13g2_decap_4 FILLER_12_579 ();
 sg13g2_fill_1 FILLER_12_602 ();
 sg13g2_decap_8 FILLER_12_608 ();
 sg13g2_decap_8 FILLER_12_615 ();
 sg13g2_fill_2 FILLER_12_622 ();
 sg13g2_fill_1 FILLER_12_624 ();
 sg13g2_fill_2 FILLER_12_645 ();
 sg13g2_decap_8 FILLER_12_652 ();
 sg13g2_decap_4 FILLER_12_659 ();
 sg13g2_fill_1 FILLER_12_663 ();
 sg13g2_decap_8 FILLER_12_669 ();
 sg13g2_decap_8 FILLER_12_676 ();
 sg13g2_decap_4 FILLER_12_683 ();
 sg13g2_fill_1 FILLER_12_687 ();
 sg13g2_decap_8 FILLER_12_694 ();
 sg13g2_decap_8 FILLER_12_701 ();
 sg13g2_fill_2 FILLER_12_708 ();
 sg13g2_fill_1 FILLER_12_710 ();
 sg13g2_decap_8 FILLER_12_715 ();
 sg13g2_decap_8 FILLER_12_722 ();
 sg13g2_fill_2 FILLER_12_729 ();
 sg13g2_fill_1 FILLER_12_731 ();
 sg13g2_decap_8 FILLER_12_735 ();
 sg13g2_decap_8 FILLER_12_742 ();
 sg13g2_decap_4 FILLER_12_749 ();
 sg13g2_fill_1 FILLER_12_753 ();
 sg13g2_fill_1 FILLER_12_770 ();
 sg13g2_decap_8 FILLER_12_791 ();
 sg13g2_decap_8 FILLER_12_798 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_8 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_12_847 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_decap_8 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_12_868 ();
 sg13g2_decap_8 FILLER_12_875 ();
 sg13g2_decap_8 FILLER_12_882 ();
 sg13g2_fill_2 FILLER_12_889 ();
 sg13g2_fill_1 FILLER_12_891 ();
 sg13g2_fill_1 FILLER_12_907 ();
 sg13g2_decap_8 FILLER_12_917 ();
 sg13g2_decap_8 FILLER_12_924 ();
 sg13g2_decap_8 FILLER_12_931 ();
 sg13g2_decap_8 FILLER_12_938 ();
 sg13g2_decap_4 FILLER_12_945 ();
 sg13g2_fill_1 FILLER_12_949 ();
 sg13g2_decap_8 FILLER_12_958 ();
 sg13g2_decap_8 FILLER_12_965 ();
 sg13g2_decap_8 FILLER_12_972 ();
 sg13g2_decap_8 FILLER_12_979 ();
 sg13g2_decap_4 FILLER_12_986 ();
 sg13g2_fill_2 FILLER_12_990 ();
 sg13g2_fill_2 FILLER_12_1001 ();
 sg13g2_decap_8 FILLER_12_1016 ();
 sg13g2_decap_8 FILLER_12_1023 ();
 sg13g2_decap_8 FILLER_12_1030 ();
 sg13g2_decap_8 FILLER_12_1037 ();
 sg13g2_decap_4 FILLER_12_1044 ();
 sg13g2_fill_1 FILLER_12_1048 ();
 sg13g2_decap_8 FILLER_12_1063 ();
 sg13g2_decap_8 FILLER_12_1073 ();
 sg13g2_decap_8 FILLER_12_1080 ();
 sg13g2_decap_8 FILLER_12_1094 ();
 sg13g2_fill_1 FILLER_12_1101 ();
 sg13g2_decap_8 FILLER_12_1117 ();
 sg13g2_decap_8 FILLER_12_1124 ();
 sg13g2_decap_8 FILLER_12_1131 ();
 sg13g2_decap_8 FILLER_12_1138 ();
 sg13g2_decap_8 FILLER_12_1145 ();
 sg13g2_decap_8 FILLER_12_1152 ();
 sg13g2_decap_8 FILLER_12_1159 ();
 sg13g2_decap_8 FILLER_12_1166 ();
 sg13g2_decap_8 FILLER_12_1173 ();
 sg13g2_decap_8 FILLER_12_1180 ();
 sg13g2_decap_8 FILLER_12_1187 ();
 sg13g2_decap_8 FILLER_12_1194 ();
 sg13g2_decap_4 FILLER_12_1201 ();
 sg13g2_fill_2 FILLER_12_1205 ();
 sg13g2_decap_8 FILLER_12_1210 ();
 sg13g2_decap_8 FILLER_12_1217 ();
 sg13g2_decap_8 FILLER_12_1224 ();
 sg13g2_fill_1 FILLER_12_1231 ();
 sg13g2_fill_2 FILLER_12_1241 ();
 sg13g2_decap_8 FILLER_12_1255 ();
 sg13g2_decap_8 FILLER_12_1262 ();
 sg13g2_decap_4 FILLER_12_1269 ();
 sg13g2_fill_2 FILLER_12_1273 ();
 sg13g2_decap_8 FILLER_12_1279 ();
 sg13g2_decap_8 FILLER_12_1286 ();
 sg13g2_decap_8 FILLER_12_1293 ();
 sg13g2_decap_4 FILLER_12_1305 ();
 sg13g2_fill_2 FILLER_12_1309 ();
 sg13g2_decap_8 FILLER_12_1315 ();
 sg13g2_fill_2 FILLER_12_1322 ();
 sg13g2_fill_2 FILLER_12_1327 ();
 sg13g2_fill_1 FILLER_12_1329 ();
 sg13g2_decap_8 FILLER_12_1345 ();
 sg13g2_decap_8 FILLER_12_1352 ();
 sg13g2_decap_8 FILLER_12_1359 ();
 sg13g2_fill_2 FILLER_12_1366 ();
 sg13g2_fill_2 FILLER_12_1371 ();
 sg13g2_fill_2 FILLER_12_1380 ();
 sg13g2_decap_8 FILLER_12_1392 ();
 sg13g2_decap_8 FILLER_12_1399 ();
 sg13g2_decap_4 FILLER_12_1406 ();
 sg13g2_fill_1 FILLER_12_1420 ();
 sg13g2_decap_8 FILLER_12_1436 ();
 sg13g2_decap_8 FILLER_12_1443 ();
 sg13g2_decap_8 FILLER_12_1450 ();
 sg13g2_decap_8 FILLER_12_1457 ();
 sg13g2_decap_8 FILLER_12_1464 ();
 sg13g2_decap_8 FILLER_12_1471 ();
 sg13g2_decap_8 FILLER_12_1478 ();
 sg13g2_decap_8 FILLER_12_1485 ();
 sg13g2_decap_8 FILLER_12_1492 ();
 sg13g2_decap_8 FILLER_12_1499 ();
 sg13g2_decap_8 FILLER_12_1506 ();
 sg13g2_fill_1 FILLER_12_1513 ();
 sg13g2_decap_8 FILLER_12_1518 ();
 sg13g2_decap_8 FILLER_12_1525 ();
 sg13g2_decap_8 FILLER_12_1532 ();
 sg13g2_decap_8 FILLER_12_1539 ();
 sg13g2_decap_8 FILLER_12_1546 ();
 sg13g2_fill_2 FILLER_12_1553 ();
 sg13g2_decap_8 FILLER_12_1562 ();
 sg13g2_fill_2 FILLER_12_1569 ();
 sg13g2_decap_8 FILLER_12_1577 ();
 sg13g2_decap_8 FILLER_12_1584 ();
 sg13g2_decap_8 FILLER_12_1591 ();
 sg13g2_fill_2 FILLER_12_1598 ();
 sg13g2_fill_1 FILLER_12_1600 ();
 sg13g2_decap_8 FILLER_12_1605 ();
 sg13g2_decap_8 FILLER_12_1612 ();
 sg13g2_decap_8 FILLER_12_1619 ();
 sg13g2_fill_1 FILLER_12_1626 ();
 sg13g2_fill_2 FILLER_12_1633 ();
 sg13g2_decap_8 FILLER_12_1647 ();
 sg13g2_decap_8 FILLER_12_1654 ();
 sg13g2_decap_8 FILLER_12_1661 ();
 sg13g2_fill_1 FILLER_12_1668 ();
 sg13g2_decap_8 FILLER_12_1678 ();
 sg13g2_decap_8 FILLER_12_1685 ();
 sg13g2_decap_8 FILLER_12_1692 ();
 sg13g2_decap_8 FILLER_12_1699 ();
 sg13g2_decap_8 FILLER_12_1706 ();
 sg13g2_decap_8 FILLER_12_1713 ();
 sg13g2_decap_8 FILLER_12_1720 ();
 sg13g2_decap_8 FILLER_12_1727 ();
 sg13g2_decap_8 FILLER_12_1734 ();
 sg13g2_decap_8 FILLER_12_1741 ();
 sg13g2_decap_8 FILLER_12_1748 ();
 sg13g2_decap_8 FILLER_12_1755 ();
 sg13g2_decap_8 FILLER_12_1762 ();
 sg13g2_decap_8 FILLER_12_1769 ();
 sg13g2_decap_8 FILLER_12_1776 ();
 sg13g2_decap_8 FILLER_12_1783 ();
 sg13g2_decap_8 FILLER_12_1790 ();
 sg13g2_decap_8 FILLER_12_1797 ();
 sg13g2_decap_8 FILLER_12_1804 ();
 sg13g2_decap_8 FILLER_12_1811 ();
 sg13g2_decap_8 FILLER_12_1818 ();
 sg13g2_decap_8 FILLER_12_1825 ();
 sg13g2_decap_8 FILLER_12_1832 ();
 sg13g2_decap_8 FILLER_12_1839 ();
 sg13g2_decap_8 FILLER_12_1846 ();
 sg13g2_decap_8 FILLER_12_1853 ();
 sg13g2_decap_8 FILLER_12_1860 ();
 sg13g2_decap_8 FILLER_12_1867 ();
 sg13g2_decap_8 FILLER_12_1874 ();
 sg13g2_decap_8 FILLER_12_1881 ();
 sg13g2_decap_8 FILLER_12_1888 ();
 sg13g2_decap_8 FILLER_12_1895 ();
 sg13g2_decap_8 FILLER_12_1902 ();
 sg13g2_decap_8 FILLER_12_1909 ();
 sg13g2_decap_8 FILLER_12_1916 ();
 sg13g2_decap_8 FILLER_12_1923 ();
 sg13g2_decap_8 FILLER_12_1930 ();
 sg13g2_decap_8 FILLER_12_1937 ();
 sg13g2_decap_8 FILLER_12_1944 ();
 sg13g2_decap_8 FILLER_12_1951 ();
 sg13g2_decap_8 FILLER_12_1958 ();
 sg13g2_decap_8 FILLER_12_1965 ();
 sg13g2_decap_8 FILLER_12_1972 ();
 sg13g2_decap_8 FILLER_12_1979 ();
 sg13g2_decap_8 FILLER_12_1986 ();
 sg13g2_decap_8 FILLER_12_1993 ();
 sg13g2_decap_8 FILLER_12_2000 ();
 sg13g2_decap_8 FILLER_12_2007 ();
 sg13g2_decap_8 FILLER_12_2014 ();
 sg13g2_decap_8 FILLER_12_2021 ();
 sg13g2_decap_8 FILLER_12_2028 ();
 sg13g2_decap_8 FILLER_12_2035 ();
 sg13g2_decap_8 FILLER_12_2042 ();
 sg13g2_decap_8 FILLER_12_2049 ();
 sg13g2_decap_8 FILLER_12_2056 ();
 sg13g2_decap_8 FILLER_12_2063 ();
 sg13g2_decap_8 FILLER_12_2070 ();
 sg13g2_decap_8 FILLER_12_2077 ();
 sg13g2_decap_8 FILLER_12_2084 ();
 sg13g2_decap_8 FILLER_12_2091 ();
 sg13g2_decap_8 FILLER_12_2098 ();
 sg13g2_decap_8 FILLER_12_2105 ();
 sg13g2_decap_8 FILLER_12_2112 ();
 sg13g2_decap_8 FILLER_12_2119 ();
 sg13g2_decap_8 FILLER_12_2126 ();
 sg13g2_decap_8 FILLER_12_2133 ();
 sg13g2_decap_8 FILLER_12_2140 ();
 sg13g2_decap_8 FILLER_12_2147 ();
 sg13g2_decap_8 FILLER_12_2154 ();
 sg13g2_decap_8 FILLER_12_2161 ();
 sg13g2_decap_8 FILLER_12_2168 ();
 sg13g2_decap_8 FILLER_12_2175 ();
 sg13g2_decap_8 FILLER_12_2182 ();
 sg13g2_decap_8 FILLER_12_2189 ();
 sg13g2_decap_8 FILLER_12_2196 ();
 sg13g2_decap_8 FILLER_12_2203 ();
 sg13g2_decap_8 FILLER_12_2210 ();
 sg13g2_decap_8 FILLER_12_2217 ();
 sg13g2_decap_8 FILLER_12_2224 ();
 sg13g2_decap_8 FILLER_12_2231 ();
 sg13g2_decap_8 FILLER_12_2238 ();
 sg13g2_decap_8 FILLER_12_2245 ();
 sg13g2_decap_8 FILLER_12_2252 ();
 sg13g2_decap_8 FILLER_12_2259 ();
 sg13g2_decap_8 FILLER_12_2266 ();
 sg13g2_decap_8 FILLER_12_2273 ();
 sg13g2_decap_8 FILLER_12_2280 ();
 sg13g2_decap_8 FILLER_12_2287 ();
 sg13g2_decap_8 FILLER_12_2294 ();
 sg13g2_decap_8 FILLER_12_2301 ();
 sg13g2_decap_8 FILLER_12_2308 ();
 sg13g2_decap_8 FILLER_12_2315 ();
 sg13g2_decap_8 FILLER_12_2322 ();
 sg13g2_decap_8 FILLER_12_2329 ();
 sg13g2_decap_8 FILLER_12_2336 ();
 sg13g2_decap_8 FILLER_12_2343 ();
 sg13g2_decap_8 FILLER_12_2350 ();
 sg13g2_decap_8 FILLER_12_2357 ();
 sg13g2_decap_8 FILLER_12_2364 ();
 sg13g2_decap_8 FILLER_12_2371 ();
 sg13g2_decap_8 FILLER_12_2378 ();
 sg13g2_decap_8 FILLER_12_2385 ();
 sg13g2_decap_8 FILLER_12_2392 ();
 sg13g2_decap_8 FILLER_12_2399 ();
 sg13g2_decap_8 FILLER_12_2406 ();
 sg13g2_decap_8 FILLER_12_2413 ();
 sg13g2_decap_8 FILLER_12_2420 ();
 sg13g2_decap_8 FILLER_12_2427 ();
 sg13g2_decap_8 FILLER_12_2434 ();
 sg13g2_decap_8 FILLER_12_2441 ();
 sg13g2_decap_8 FILLER_12_2448 ();
 sg13g2_decap_8 FILLER_12_2455 ();
 sg13g2_decap_8 FILLER_12_2462 ();
 sg13g2_decap_8 FILLER_12_2469 ();
 sg13g2_decap_8 FILLER_12_2476 ();
 sg13g2_decap_8 FILLER_12_2483 ();
 sg13g2_decap_8 FILLER_12_2490 ();
 sg13g2_decap_8 FILLER_12_2497 ();
 sg13g2_decap_8 FILLER_12_2504 ();
 sg13g2_decap_8 FILLER_12_2511 ();
 sg13g2_decap_8 FILLER_12_2518 ();
 sg13g2_decap_8 FILLER_12_2525 ();
 sg13g2_decap_8 FILLER_12_2532 ();
 sg13g2_decap_8 FILLER_12_2539 ();
 sg13g2_decap_8 FILLER_12_2546 ();
 sg13g2_decap_8 FILLER_12_2553 ();
 sg13g2_decap_8 FILLER_12_2560 ();
 sg13g2_decap_8 FILLER_12_2567 ();
 sg13g2_decap_8 FILLER_12_2574 ();
 sg13g2_decap_8 FILLER_12_2581 ();
 sg13g2_decap_8 FILLER_12_2588 ();
 sg13g2_decap_8 FILLER_12_2595 ();
 sg13g2_decap_8 FILLER_12_2602 ();
 sg13g2_decap_8 FILLER_12_2609 ();
 sg13g2_decap_8 FILLER_12_2616 ();
 sg13g2_decap_8 FILLER_12_2623 ();
 sg13g2_decap_8 FILLER_12_2630 ();
 sg13g2_decap_8 FILLER_12_2637 ();
 sg13g2_decap_8 FILLER_12_2644 ();
 sg13g2_decap_8 FILLER_12_2651 ();
 sg13g2_decap_8 FILLER_12_2658 ();
 sg13g2_decap_4 FILLER_12_2665 ();
 sg13g2_fill_1 FILLER_12_2669 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_4 FILLER_13_119 ();
 sg13g2_fill_1 FILLER_13_123 ();
 sg13g2_decap_8 FILLER_13_132 ();
 sg13g2_decap_8 FILLER_13_139 ();
 sg13g2_decap_8 FILLER_13_146 ();
 sg13g2_decap_8 FILLER_13_153 ();
 sg13g2_fill_2 FILLER_13_160 ();
 sg13g2_fill_1 FILLER_13_162 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_4 FILLER_13_350 ();
 sg13g2_fill_2 FILLER_13_354 ();
 sg13g2_decap_8 FILLER_13_382 ();
 sg13g2_decap_8 FILLER_13_389 ();
 sg13g2_decap_8 FILLER_13_396 ();
 sg13g2_decap_8 FILLER_13_403 ();
 sg13g2_decap_8 FILLER_13_410 ();
 sg13g2_decap_8 FILLER_13_417 ();
 sg13g2_decap_8 FILLER_13_424 ();
 sg13g2_decap_8 FILLER_13_431 ();
 sg13g2_decap_8 FILLER_13_438 ();
 sg13g2_decap_8 FILLER_13_445 ();
 sg13g2_decap_8 FILLER_13_452 ();
 sg13g2_decap_8 FILLER_13_459 ();
 sg13g2_decap_8 FILLER_13_466 ();
 sg13g2_fill_1 FILLER_13_473 ();
 sg13g2_decap_8 FILLER_13_486 ();
 sg13g2_decap_8 FILLER_13_493 ();
 sg13g2_decap_8 FILLER_13_500 ();
 sg13g2_decap_4 FILLER_13_507 ();
 sg13g2_decap_8 FILLER_13_516 ();
 sg13g2_decap_8 FILLER_13_523 ();
 sg13g2_decap_8 FILLER_13_530 ();
 sg13g2_decap_8 FILLER_13_537 ();
 sg13g2_decap_8 FILLER_13_544 ();
 sg13g2_decap_8 FILLER_13_551 ();
 sg13g2_decap_8 FILLER_13_558 ();
 sg13g2_decap_8 FILLER_13_565 ();
 sg13g2_decap_8 FILLER_13_572 ();
 sg13g2_decap_8 FILLER_13_579 ();
 sg13g2_decap_8 FILLER_13_586 ();
 sg13g2_fill_1 FILLER_13_598 ();
 sg13g2_decap_8 FILLER_13_605 ();
 sg13g2_decap_4 FILLER_13_612 ();
 sg13g2_fill_2 FILLER_13_616 ();
 sg13g2_fill_2 FILLER_13_622 ();
 sg13g2_decap_8 FILLER_13_629 ();
 sg13g2_decap_4 FILLER_13_636 ();
 sg13g2_fill_2 FILLER_13_640 ();
 sg13g2_decap_8 FILLER_13_654 ();
 sg13g2_decap_8 FILLER_13_661 ();
 sg13g2_decap_8 FILLER_13_668 ();
 sg13g2_decap_8 FILLER_13_675 ();
 sg13g2_decap_8 FILLER_13_682 ();
 sg13g2_decap_8 FILLER_13_689 ();
 sg13g2_decap_8 FILLER_13_696 ();
 sg13g2_decap_8 FILLER_13_703 ();
 sg13g2_decap_8 FILLER_13_710 ();
 sg13g2_fill_1 FILLER_13_717 ();
 sg13g2_decap_4 FILLER_13_721 ();
 sg13g2_fill_2 FILLER_13_725 ();
 sg13g2_decap_8 FILLER_13_737 ();
 sg13g2_decap_8 FILLER_13_744 ();
 sg13g2_fill_2 FILLER_13_751 ();
 sg13g2_fill_1 FILLER_13_753 ();
 sg13g2_decap_8 FILLER_13_758 ();
 sg13g2_decap_8 FILLER_13_765 ();
 sg13g2_fill_2 FILLER_13_772 ();
 sg13g2_decap_4 FILLER_13_780 ();
 sg13g2_fill_1 FILLER_13_784 ();
 sg13g2_decap_8 FILLER_13_789 ();
 sg13g2_decap_8 FILLER_13_796 ();
 sg13g2_decap_8 FILLER_13_803 ();
 sg13g2_fill_1 FILLER_13_810 ();
 sg13g2_decap_8 FILLER_13_834 ();
 sg13g2_decap_8 FILLER_13_841 ();
 sg13g2_decap_4 FILLER_13_848 ();
 sg13g2_fill_2 FILLER_13_852 ();
 sg13g2_decap_8 FILLER_13_859 ();
 sg13g2_decap_8 FILLER_13_866 ();
 sg13g2_decap_4 FILLER_13_873 ();
 sg13g2_fill_2 FILLER_13_877 ();
 sg13g2_fill_2 FILLER_13_906 ();
 sg13g2_decap_8 FILLER_13_927 ();
 sg13g2_decap_8 FILLER_13_934 ();
 sg13g2_decap_8 FILLER_13_941 ();
 sg13g2_fill_2 FILLER_13_948 ();
 sg13g2_fill_1 FILLER_13_950 ();
 sg13g2_decap_8 FILLER_13_956 ();
 sg13g2_decap_8 FILLER_13_963 ();
 sg13g2_decap_8 FILLER_13_970 ();
 sg13g2_decap_4 FILLER_13_977 ();
 sg13g2_fill_1 FILLER_13_981 ();
 sg13g2_decap_4 FILLER_13_986 ();
 sg13g2_fill_2 FILLER_13_990 ();
 sg13g2_decap_8 FILLER_13_1003 ();
 sg13g2_decap_8 FILLER_13_1010 ();
 sg13g2_decap_8 FILLER_13_1017 ();
 sg13g2_decap_8 FILLER_13_1024 ();
 sg13g2_decap_8 FILLER_13_1031 ();
 sg13g2_decap_8 FILLER_13_1038 ();
 sg13g2_decap_8 FILLER_13_1045 ();
 sg13g2_decap_8 FILLER_13_1052 ();
 sg13g2_decap_8 FILLER_13_1059 ();
 sg13g2_decap_4 FILLER_13_1066 ();
 sg13g2_fill_1 FILLER_13_1074 ();
 sg13g2_fill_1 FILLER_13_1080 ();
 sg13g2_decap_4 FILLER_13_1084 ();
 sg13g2_decap_8 FILLER_13_1092 ();
 sg13g2_decap_4 FILLER_13_1099 ();
 sg13g2_fill_2 FILLER_13_1103 ();
 sg13g2_decap_8 FILLER_13_1109 ();
 sg13g2_decap_8 FILLER_13_1116 ();
 sg13g2_fill_1 FILLER_13_1123 ();
 sg13g2_decap_8 FILLER_13_1127 ();
 sg13g2_decap_8 FILLER_13_1134 ();
 sg13g2_fill_2 FILLER_13_1141 ();
 sg13g2_decap_8 FILLER_13_1147 ();
 sg13g2_fill_1 FILLER_13_1154 ();
 sg13g2_decap_4 FILLER_13_1175 ();
 sg13g2_decap_8 FILLER_13_1186 ();
 sg13g2_decap_8 FILLER_13_1193 ();
 sg13g2_fill_1 FILLER_13_1200 ();
 sg13g2_fill_2 FILLER_13_1228 ();
 sg13g2_fill_1 FILLER_13_1237 ();
 sg13g2_fill_1 FILLER_13_1242 ();
 sg13g2_fill_1 FILLER_13_1252 ();
 sg13g2_decap_8 FILLER_13_1258 ();
 sg13g2_decap_8 FILLER_13_1265 ();
 sg13g2_decap_8 FILLER_13_1272 ();
 sg13g2_decap_8 FILLER_13_1279 ();
 sg13g2_decap_8 FILLER_13_1286 ();
 sg13g2_decap_8 FILLER_13_1293 ();
 sg13g2_decap_8 FILLER_13_1303 ();
 sg13g2_fill_1 FILLER_13_1310 ();
 sg13g2_decap_4 FILLER_13_1319 ();
 sg13g2_fill_1 FILLER_13_1323 ();
 sg13g2_decap_4 FILLER_13_1328 ();
 sg13g2_fill_1 FILLER_13_1332 ();
 sg13g2_decap_8 FILLER_13_1338 ();
 sg13g2_decap_8 FILLER_13_1345 ();
 sg13g2_decap_8 FILLER_13_1352 ();
 sg13g2_decap_4 FILLER_13_1359 ();
 sg13g2_fill_2 FILLER_13_1363 ();
 sg13g2_decap_8 FILLER_13_1376 ();
 sg13g2_decap_8 FILLER_13_1387 ();
 sg13g2_decap_8 FILLER_13_1394 ();
 sg13g2_decap_8 FILLER_13_1401 ();
 sg13g2_decap_8 FILLER_13_1408 ();
 sg13g2_fill_2 FILLER_13_1415 ();
 sg13g2_decap_8 FILLER_13_1422 ();
 sg13g2_decap_4 FILLER_13_1429 ();
 sg13g2_fill_2 FILLER_13_1433 ();
 sg13g2_decap_8 FILLER_13_1455 ();
 sg13g2_decap_4 FILLER_13_1462 ();
 sg13g2_decap_8 FILLER_13_1471 ();
 sg13g2_decap_8 FILLER_13_1478 ();
 sg13g2_decap_8 FILLER_13_1485 ();
 sg13g2_decap_8 FILLER_13_1492 ();
 sg13g2_decap_8 FILLER_13_1499 ();
 sg13g2_decap_8 FILLER_13_1506 ();
 sg13g2_decap_8 FILLER_13_1513 ();
 sg13g2_decap_8 FILLER_13_1520 ();
 sg13g2_fill_2 FILLER_13_1542 ();
 sg13g2_decap_8 FILLER_13_1547 ();
 sg13g2_decap_4 FILLER_13_1554 ();
 sg13g2_fill_1 FILLER_13_1558 ();
 sg13g2_decap_8 FILLER_13_1562 ();
 sg13g2_decap_8 FILLER_13_1569 ();
 sg13g2_decap_8 FILLER_13_1576 ();
 sg13g2_decap_8 FILLER_13_1583 ();
 sg13g2_decap_8 FILLER_13_1590 ();
 sg13g2_decap_8 FILLER_13_1597 ();
 sg13g2_decap_8 FILLER_13_1604 ();
 sg13g2_decap_8 FILLER_13_1611 ();
 sg13g2_decap_8 FILLER_13_1618 ();
 sg13g2_fill_2 FILLER_13_1625 ();
 sg13g2_decap_4 FILLER_13_1630 ();
 sg13g2_fill_1 FILLER_13_1634 ();
 sg13g2_decap_8 FILLER_13_1639 ();
 sg13g2_decap_8 FILLER_13_1646 ();
 sg13g2_decap_8 FILLER_13_1653 ();
 sg13g2_decap_8 FILLER_13_1660 ();
 sg13g2_decap_4 FILLER_13_1667 ();
 sg13g2_decap_8 FILLER_13_1675 ();
 sg13g2_decap_8 FILLER_13_1682 ();
 sg13g2_decap_8 FILLER_13_1689 ();
 sg13g2_decap_4 FILLER_13_1696 ();
 sg13g2_fill_2 FILLER_13_1700 ();
 sg13g2_decap_8 FILLER_13_1706 ();
 sg13g2_decap_8 FILLER_13_1713 ();
 sg13g2_decap_8 FILLER_13_1720 ();
 sg13g2_decap_8 FILLER_13_1727 ();
 sg13g2_decap_8 FILLER_13_1734 ();
 sg13g2_decap_8 FILLER_13_1741 ();
 sg13g2_decap_8 FILLER_13_1748 ();
 sg13g2_decap_8 FILLER_13_1755 ();
 sg13g2_decap_8 FILLER_13_1762 ();
 sg13g2_decap_8 FILLER_13_1769 ();
 sg13g2_decap_8 FILLER_13_1776 ();
 sg13g2_decap_8 FILLER_13_1783 ();
 sg13g2_decap_8 FILLER_13_1790 ();
 sg13g2_decap_8 FILLER_13_1797 ();
 sg13g2_fill_1 FILLER_13_1804 ();
 sg13g2_decap_8 FILLER_13_1809 ();
 sg13g2_decap_8 FILLER_13_1816 ();
 sg13g2_decap_8 FILLER_13_1823 ();
 sg13g2_decap_8 FILLER_13_1830 ();
 sg13g2_decap_8 FILLER_13_1865 ();
 sg13g2_decap_8 FILLER_13_1872 ();
 sg13g2_decap_8 FILLER_13_1879 ();
 sg13g2_decap_8 FILLER_13_1886 ();
 sg13g2_decap_8 FILLER_13_1893 ();
 sg13g2_decap_8 FILLER_13_1900 ();
 sg13g2_decap_8 FILLER_13_1907 ();
 sg13g2_decap_8 FILLER_13_1914 ();
 sg13g2_decap_8 FILLER_13_1921 ();
 sg13g2_decap_8 FILLER_13_1928 ();
 sg13g2_decap_8 FILLER_13_1935 ();
 sg13g2_decap_8 FILLER_13_1942 ();
 sg13g2_decap_8 FILLER_13_1949 ();
 sg13g2_decap_8 FILLER_13_1956 ();
 sg13g2_decap_8 FILLER_13_1963 ();
 sg13g2_decap_8 FILLER_13_1970 ();
 sg13g2_decap_8 FILLER_13_1977 ();
 sg13g2_decap_8 FILLER_13_1984 ();
 sg13g2_decap_8 FILLER_13_1991 ();
 sg13g2_decap_8 FILLER_13_1998 ();
 sg13g2_decap_8 FILLER_13_2005 ();
 sg13g2_decap_8 FILLER_13_2012 ();
 sg13g2_decap_8 FILLER_13_2019 ();
 sg13g2_decap_8 FILLER_13_2026 ();
 sg13g2_decap_8 FILLER_13_2033 ();
 sg13g2_decap_8 FILLER_13_2040 ();
 sg13g2_decap_8 FILLER_13_2047 ();
 sg13g2_decap_8 FILLER_13_2054 ();
 sg13g2_decap_8 FILLER_13_2061 ();
 sg13g2_decap_8 FILLER_13_2068 ();
 sg13g2_decap_8 FILLER_13_2075 ();
 sg13g2_decap_8 FILLER_13_2082 ();
 sg13g2_decap_8 FILLER_13_2089 ();
 sg13g2_decap_8 FILLER_13_2096 ();
 sg13g2_decap_8 FILLER_13_2103 ();
 sg13g2_decap_8 FILLER_13_2110 ();
 sg13g2_decap_8 FILLER_13_2117 ();
 sg13g2_decap_8 FILLER_13_2124 ();
 sg13g2_decap_8 FILLER_13_2131 ();
 sg13g2_decap_8 FILLER_13_2138 ();
 sg13g2_decap_8 FILLER_13_2145 ();
 sg13g2_decap_8 FILLER_13_2152 ();
 sg13g2_decap_8 FILLER_13_2159 ();
 sg13g2_decap_8 FILLER_13_2166 ();
 sg13g2_decap_8 FILLER_13_2173 ();
 sg13g2_decap_8 FILLER_13_2180 ();
 sg13g2_decap_8 FILLER_13_2187 ();
 sg13g2_decap_8 FILLER_13_2194 ();
 sg13g2_decap_8 FILLER_13_2201 ();
 sg13g2_decap_8 FILLER_13_2208 ();
 sg13g2_decap_8 FILLER_13_2215 ();
 sg13g2_decap_8 FILLER_13_2222 ();
 sg13g2_decap_8 FILLER_13_2229 ();
 sg13g2_decap_8 FILLER_13_2236 ();
 sg13g2_decap_8 FILLER_13_2243 ();
 sg13g2_decap_8 FILLER_13_2250 ();
 sg13g2_decap_8 FILLER_13_2257 ();
 sg13g2_decap_8 FILLER_13_2264 ();
 sg13g2_decap_8 FILLER_13_2271 ();
 sg13g2_decap_8 FILLER_13_2278 ();
 sg13g2_decap_8 FILLER_13_2285 ();
 sg13g2_decap_8 FILLER_13_2292 ();
 sg13g2_decap_8 FILLER_13_2299 ();
 sg13g2_decap_8 FILLER_13_2306 ();
 sg13g2_decap_8 FILLER_13_2313 ();
 sg13g2_decap_8 FILLER_13_2320 ();
 sg13g2_decap_8 FILLER_13_2327 ();
 sg13g2_decap_8 FILLER_13_2334 ();
 sg13g2_decap_8 FILLER_13_2341 ();
 sg13g2_decap_8 FILLER_13_2348 ();
 sg13g2_decap_8 FILLER_13_2355 ();
 sg13g2_decap_8 FILLER_13_2362 ();
 sg13g2_decap_8 FILLER_13_2369 ();
 sg13g2_decap_8 FILLER_13_2376 ();
 sg13g2_decap_8 FILLER_13_2383 ();
 sg13g2_decap_8 FILLER_13_2390 ();
 sg13g2_decap_8 FILLER_13_2397 ();
 sg13g2_decap_8 FILLER_13_2404 ();
 sg13g2_decap_8 FILLER_13_2411 ();
 sg13g2_decap_8 FILLER_13_2418 ();
 sg13g2_decap_8 FILLER_13_2425 ();
 sg13g2_decap_8 FILLER_13_2432 ();
 sg13g2_decap_8 FILLER_13_2439 ();
 sg13g2_decap_8 FILLER_13_2446 ();
 sg13g2_decap_8 FILLER_13_2453 ();
 sg13g2_decap_8 FILLER_13_2460 ();
 sg13g2_decap_8 FILLER_13_2467 ();
 sg13g2_decap_8 FILLER_13_2474 ();
 sg13g2_decap_8 FILLER_13_2481 ();
 sg13g2_decap_8 FILLER_13_2488 ();
 sg13g2_decap_8 FILLER_13_2495 ();
 sg13g2_decap_8 FILLER_13_2502 ();
 sg13g2_decap_8 FILLER_13_2509 ();
 sg13g2_decap_8 FILLER_13_2516 ();
 sg13g2_decap_8 FILLER_13_2523 ();
 sg13g2_decap_8 FILLER_13_2530 ();
 sg13g2_decap_8 FILLER_13_2537 ();
 sg13g2_decap_8 FILLER_13_2544 ();
 sg13g2_decap_8 FILLER_13_2551 ();
 sg13g2_decap_8 FILLER_13_2558 ();
 sg13g2_decap_8 FILLER_13_2565 ();
 sg13g2_decap_8 FILLER_13_2572 ();
 sg13g2_decap_8 FILLER_13_2579 ();
 sg13g2_decap_8 FILLER_13_2586 ();
 sg13g2_decap_8 FILLER_13_2593 ();
 sg13g2_decap_8 FILLER_13_2600 ();
 sg13g2_decap_8 FILLER_13_2607 ();
 sg13g2_decap_8 FILLER_13_2614 ();
 sg13g2_decap_8 FILLER_13_2621 ();
 sg13g2_decap_8 FILLER_13_2628 ();
 sg13g2_decap_8 FILLER_13_2635 ();
 sg13g2_decap_8 FILLER_13_2642 ();
 sg13g2_decap_8 FILLER_13_2649 ();
 sg13g2_decap_8 FILLER_13_2656 ();
 sg13g2_decap_8 FILLER_13_2663 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_fill_2 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_decap_8 FILLER_14_427 ();
 sg13g2_decap_8 FILLER_14_434 ();
 sg13g2_decap_8 FILLER_14_441 ();
 sg13g2_decap_8 FILLER_14_448 ();
 sg13g2_decap_8 FILLER_14_455 ();
 sg13g2_decap_8 FILLER_14_462 ();
 sg13g2_fill_2 FILLER_14_469 ();
 sg13g2_fill_1 FILLER_14_471 ();
 sg13g2_fill_2 FILLER_14_478 ();
 sg13g2_decap_8 FILLER_14_484 ();
 sg13g2_decap_8 FILLER_14_491 ();
 sg13g2_decap_8 FILLER_14_498 ();
 sg13g2_decap_8 FILLER_14_505 ();
 sg13g2_decap_8 FILLER_14_512 ();
 sg13g2_decap_8 FILLER_14_519 ();
 sg13g2_decap_8 FILLER_14_526 ();
 sg13g2_decap_4 FILLER_14_553 ();
 sg13g2_decap_8 FILLER_14_561 ();
 sg13g2_decap_8 FILLER_14_568 ();
 sg13g2_decap_8 FILLER_14_575 ();
 sg13g2_decap_8 FILLER_14_582 ();
 sg13g2_decap_8 FILLER_14_589 ();
 sg13g2_decap_8 FILLER_14_596 ();
 sg13g2_decap_4 FILLER_14_603 ();
 sg13g2_fill_1 FILLER_14_607 ();
 sg13g2_decap_8 FILLER_14_612 ();
 sg13g2_decap_8 FILLER_14_619 ();
 sg13g2_decap_8 FILLER_14_626 ();
 sg13g2_decap_8 FILLER_14_633 ();
 sg13g2_decap_8 FILLER_14_640 ();
 sg13g2_decap_8 FILLER_14_647 ();
 sg13g2_decap_8 FILLER_14_654 ();
 sg13g2_fill_2 FILLER_14_661 ();
 sg13g2_decap_8 FILLER_14_675 ();
 sg13g2_decap_8 FILLER_14_682 ();
 sg13g2_decap_8 FILLER_14_689 ();
 sg13g2_decap_8 FILLER_14_696 ();
 sg13g2_decap_8 FILLER_14_703 ();
 sg13g2_decap_8 FILLER_14_710 ();
 sg13g2_decap_8 FILLER_14_717 ();
 sg13g2_decap_8 FILLER_14_724 ();
 sg13g2_fill_1 FILLER_14_731 ();
 sg13g2_decap_8 FILLER_14_735 ();
 sg13g2_decap_8 FILLER_14_742 ();
 sg13g2_decap_8 FILLER_14_749 ();
 sg13g2_decap_8 FILLER_14_756 ();
 sg13g2_decap_8 FILLER_14_763 ();
 sg13g2_decap_8 FILLER_14_770 ();
 sg13g2_decap_4 FILLER_14_777 ();
 sg13g2_fill_1 FILLER_14_781 ();
 sg13g2_decap_8 FILLER_14_786 ();
 sg13g2_decap_8 FILLER_14_793 ();
 sg13g2_decap_8 FILLER_14_800 ();
 sg13g2_decap_8 FILLER_14_807 ();
 sg13g2_decap_8 FILLER_14_814 ();
 sg13g2_fill_2 FILLER_14_821 ();
 sg13g2_decap_8 FILLER_14_827 ();
 sg13g2_decap_4 FILLER_14_834 ();
 sg13g2_decap_8 FILLER_14_850 ();
 sg13g2_fill_2 FILLER_14_857 ();
 sg13g2_fill_1 FILLER_14_859 ();
 sg13g2_decap_8 FILLER_14_865 ();
 sg13g2_decap_8 FILLER_14_872 ();
 sg13g2_decap_4 FILLER_14_879 ();
 sg13g2_decap_8 FILLER_14_900 ();
 sg13g2_fill_1 FILLER_14_907 ();
 sg13g2_decap_8 FILLER_14_918 ();
 sg13g2_decap_8 FILLER_14_925 ();
 sg13g2_decap_8 FILLER_14_932 ();
 sg13g2_decap_8 FILLER_14_939 ();
 sg13g2_decap_8 FILLER_14_946 ();
 sg13g2_decap_8 FILLER_14_953 ();
 sg13g2_decap_8 FILLER_14_960 ();
 sg13g2_decap_8 FILLER_14_967 ();
 sg13g2_decap_8 FILLER_14_974 ();
 sg13g2_decap_4 FILLER_14_981 ();
 sg13g2_fill_2 FILLER_14_985 ();
 sg13g2_decap_8 FILLER_14_996 ();
 sg13g2_decap_8 FILLER_14_1003 ();
 sg13g2_decap_8 FILLER_14_1010 ();
 sg13g2_decap_8 FILLER_14_1017 ();
 sg13g2_decap_8 FILLER_14_1024 ();
 sg13g2_decap_8 FILLER_14_1031 ();
 sg13g2_decap_8 FILLER_14_1038 ();
 sg13g2_decap_8 FILLER_14_1045 ();
 sg13g2_decap_8 FILLER_14_1052 ();
 sg13g2_decap_8 FILLER_14_1059 ();
 sg13g2_decap_8 FILLER_14_1066 ();
 sg13g2_decap_8 FILLER_14_1073 ();
 sg13g2_decap_4 FILLER_14_1080 ();
 sg13g2_fill_2 FILLER_14_1084 ();
 sg13g2_decap_8 FILLER_14_1091 ();
 sg13g2_decap_8 FILLER_14_1098 ();
 sg13g2_decap_8 FILLER_14_1108 ();
 sg13g2_decap_4 FILLER_14_1115 ();
 sg13g2_fill_1 FILLER_14_1119 ();
 sg13g2_decap_8 FILLER_14_1129 ();
 sg13g2_decap_8 FILLER_14_1136 ();
 sg13g2_decap_8 FILLER_14_1143 ();
 sg13g2_decap_8 FILLER_14_1150 ();
 sg13g2_decap_8 FILLER_14_1157 ();
 sg13g2_decap_8 FILLER_14_1169 ();
 sg13g2_decap_8 FILLER_14_1176 ();
 sg13g2_decap_8 FILLER_14_1183 ();
 sg13g2_decap_8 FILLER_14_1190 ();
 sg13g2_decap_8 FILLER_14_1197 ();
 sg13g2_decap_8 FILLER_14_1204 ();
 sg13g2_decap_4 FILLER_14_1211 ();
 sg13g2_fill_1 FILLER_14_1215 ();
 sg13g2_decap_4 FILLER_14_1220 ();
 sg13g2_fill_1 FILLER_14_1224 ();
 sg13g2_decap_8 FILLER_14_1234 ();
 sg13g2_decap_4 FILLER_14_1241 ();
 sg13g2_fill_1 FILLER_14_1245 ();
 sg13g2_decap_8 FILLER_14_1251 ();
 sg13g2_decap_4 FILLER_14_1258 ();
 sg13g2_fill_1 FILLER_14_1262 ();
 sg13g2_fill_2 FILLER_14_1268 ();
 sg13g2_decap_8 FILLER_14_1274 ();
 sg13g2_decap_8 FILLER_14_1281 ();
 sg13g2_decap_8 FILLER_14_1288 ();
 sg13g2_decap_8 FILLER_14_1295 ();
 sg13g2_decap_8 FILLER_14_1302 ();
 sg13g2_fill_2 FILLER_14_1309 ();
 sg13g2_decap_8 FILLER_14_1316 ();
 sg13g2_decap_8 FILLER_14_1323 ();
 sg13g2_fill_2 FILLER_14_1330 ();
 sg13g2_fill_1 FILLER_14_1332 ();
 sg13g2_decap_8 FILLER_14_1342 ();
 sg13g2_decap_8 FILLER_14_1349 ();
 sg13g2_decap_8 FILLER_14_1356 ();
 sg13g2_decap_4 FILLER_14_1363 ();
 sg13g2_fill_1 FILLER_14_1367 ();
 sg13g2_decap_8 FILLER_14_1377 ();
 sg13g2_decap_8 FILLER_14_1384 ();
 sg13g2_decap_8 FILLER_14_1391 ();
 sg13g2_decap_8 FILLER_14_1398 ();
 sg13g2_decap_8 FILLER_14_1405 ();
 sg13g2_fill_1 FILLER_14_1412 ();
 sg13g2_fill_1 FILLER_14_1416 ();
 sg13g2_fill_1 FILLER_14_1428 ();
 sg13g2_fill_1 FILLER_14_1434 ();
 sg13g2_decap_8 FILLER_14_1440 ();
 sg13g2_decap_8 FILLER_14_1447 ();
 sg13g2_decap_4 FILLER_14_1454 ();
 sg13g2_decap_8 FILLER_14_1461 ();
 sg13g2_decap_8 FILLER_14_1472 ();
 sg13g2_decap_8 FILLER_14_1479 ();
 sg13g2_decap_8 FILLER_14_1486 ();
 sg13g2_decap_8 FILLER_14_1493 ();
 sg13g2_decap_8 FILLER_14_1500 ();
 sg13g2_decap_8 FILLER_14_1507 ();
 sg13g2_decap_4 FILLER_14_1514 ();
 sg13g2_fill_1 FILLER_14_1518 ();
 sg13g2_fill_1 FILLER_14_1526 ();
 sg13g2_decap_8 FILLER_14_1531 ();
 sg13g2_decap_8 FILLER_14_1538 ();
 sg13g2_decap_4 FILLER_14_1545 ();
 sg13g2_fill_2 FILLER_14_1549 ();
 sg13g2_fill_2 FILLER_14_1563 ();
 sg13g2_fill_1 FILLER_14_1565 ();
 sg13g2_decap_8 FILLER_14_1570 ();
 sg13g2_decap_8 FILLER_14_1577 ();
 sg13g2_decap_8 FILLER_14_1584 ();
 sg13g2_decap_8 FILLER_14_1591 ();
 sg13g2_decap_8 FILLER_14_1598 ();
 sg13g2_decap_8 FILLER_14_1605 ();
 sg13g2_decap_4 FILLER_14_1616 ();
 sg13g2_decap_8 FILLER_14_1624 ();
 sg13g2_decap_8 FILLER_14_1631 ();
 sg13g2_decap_8 FILLER_14_1638 ();
 sg13g2_decap_8 FILLER_14_1645 ();
 sg13g2_fill_2 FILLER_14_1652 ();
 sg13g2_decap_8 FILLER_14_1666 ();
 sg13g2_decap_4 FILLER_14_1673 ();
 sg13g2_fill_2 FILLER_14_1677 ();
 sg13g2_decap_8 FILLER_14_1694 ();
 sg13g2_decap_8 FILLER_14_1701 ();
 sg13g2_decap_8 FILLER_14_1708 ();
 sg13g2_decap_4 FILLER_14_1715 ();
 sg13g2_fill_2 FILLER_14_1719 ();
 sg13g2_decap_8 FILLER_14_1742 ();
 sg13g2_decap_8 FILLER_14_1749 ();
 sg13g2_decap_8 FILLER_14_1756 ();
 sg13g2_decap_8 FILLER_14_1763 ();
 sg13g2_decap_8 FILLER_14_1770 ();
 sg13g2_decap_8 FILLER_14_1777 ();
 sg13g2_decap_4 FILLER_14_1784 ();
 sg13g2_decap_8 FILLER_14_1793 ();
 sg13g2_decap_8 FILLER_14_1800 ();
 sg13g2_decap_8 FILLER_14_1807 ();
 sg13g2_decap_4 FILLER_14_1814 ();
 sg13g2_fill_1 FILLER_14_1818 ();
 sg13g2_decap_8 FILLER_14_1823 ();
 sg13g2_fill_2 FILLER_14_1830 ();
 sg13g2_decap_8 FILLER_14_1837 ();
 sg13g2_decap_4 FILLER_14_1844 ();
 sg13g2_fill_2 FILLER_14_1848 ();
 sg13g2_decap_8 FILLER_14_1854 ();
 sg13g2_decap_8 FILLER_14_1861 ();
 sg13g2_decap_8 FILLER_14_1868 ();
 sg13g2_decap_8 FILLER_14_1875 ();
 sg13g2_decap_8 FILLER_14_1882 ();
 sg13g2_decap_8 FILLER_14_1889 ();
 sg13g2_decap_8 FILLER_14_1896 ();
 sg13g2_decap_8 FILLER_14_1903 ();
 sg13g2_decap_8 FILLER_14_1910 ();
 sg13g2_decap_8 FILLER_14_1917 ();
 sg13g2_decap_8 FILLER_14_1924 ();
 sg13g2_decap_8 FILLER_14_1931 ();
 sg13g2_decap_8 FILLER_14_1938 ();
 sg13g2_decap_8 FILLER_14_1945 ();
 sg13g2_decap_8 FILLER_14_1952 ();
 sg13g2_decap_8 FILLER_14_1959 ();
 sg13g2_decap_8 FILLER_14_1966 ();
 sg13g2_decap_8 FILLER_14_1973 ();
 sg13g2_decap_8 FILLER_14_1980 ();
 sg13g2_decap_8 FILLER_14_1987 ();
 sg13g2_decap_8 FILLER_14_1994 ();
 sg13g2_decap_8 FILLER_14_2001 ();
 sg13g2_decap_8 FILLER_14_2008 ();
 sg13g2_decap_8 FILLER_14_2015 ();
 sg13g2_decap_8 FILLER_14_2022 ();
 sg13g2_decap_8 FILLER_14_2029 ();
 sg13g2_decap_8 FILLER_14_2036 ();
 sg13g2_decap_8 FILLER_14_2043 ();
 sg13g2_decap_8 FILLER_14_2050 ();
 sg13g2_decap_8 FILLER_14_2057 ();
 sg13g2_decap_8 FILLER_14_2064 ();
 sg13g2_decap_8 FILLER_14_2071 ();
 sg13g2_decap_8 FILLER_14_2078 ();
 sg13g2_decap_8 FILLER_14_2085 ();
 sg13g2_decap_8 FILLER_14_2092 ();
 sg13g2_decap_8 FILLER_14_2099 ();
 sg13g2_decap_8 FILLER_14_2106 ();
 sg13g2_decap_8 FILLER_14_2113 ();
 sg13g2_decap_8 FILLER_14_2120 ();
 sg13g2_decap_8 FILLER_14_2127 ();
 sg13g2_decap_8 FILLER_14_2134 ();
 sg13g2_decap_8 FILLER_14_2141 ();
 sg13g2_decap_8 FILLER_14_2148 ();
 sg13g2_decap_8 FILLER_14_2155 ();
 sg13g2_decap_8 FILLER_14_2162 ();
 sg13g2_decap_8 FILLER_14_2169 ();
 sg13g2_decap_8 FILLER_14_2176 ();
 sg13g2_decap_8 FILLER_14_2183 ();
 sg13g2_decap_8 FILLER_14_2190 ();
 sg13g2_decap_8 FILLER_14_2197 ();
 sg13g2_decap_8 FILLER_14_2204 ();
 sg13g2_decap_8 FILLER_14_2211 ();
 sg13g2_decap_8 FILLER_14_2218 ();
 sg13g2_decap_8 FILLER_14_2225 ();
 sg13g2_decap_8 FILLER_14_2232 ();
 sg13g2_decap_8 FILLER_14_2239 ();
 sg13g2_decap_8 FILLER_14_2246 ();
 sg13g2_decap_8 FILLER_14_2253 ();
 sg13g2_decap_8 FILLER_14_2260 ();
 sg13g2_decap_8 FILLER_14_2267 ();
 sg13g2_decap_8 FILLER_14_2274 ();
 sg13g2_decap_8 FILLER_14_2281 ();
 sg13g2_decap_8 FILLER_14_2288 ();
 sg13g2_decap_8 FILLER_14_2295 ();
 sg13g2_decap_8 FILLER_14_2302 ();
 sg13g2_decap_8 FILLER_14_2309 ();
 sg13g2_decap_8 FILLER_14_2316 ();
 sg13g2_decap_8 FILLER_14_2323 ();
 sg13g2_decap_8 FILLER_14_2330 ();
 sg13g2_decap_8 FILLER_14_2337 ();
 sg13g2_decap_8 FILLER_14_2344 ();
 sg13g2_decap_8 FILLER_14_2351 ();
 sg13g2_decap_8 FILLER_14_2358 ();
 sg13g2_decap_8 FILLER_14_2365 ();
 sg13g2_decap_8 FILLER_14_2372 ();
 sg13g2_decap_8 FILLER_14_2379 ();
 sg13g2_decap_8 FILLER_14_2386 ();
 sg13g2_decap_8 FILLER_14_2393 ();
 sg13g2_decap_8 FILLER_14_2400 ();
 sg13g2_decap_8 FILLER_14_2407 ();
 sg13g2_decap_8 FILLER_14_2414 ();
 sg13g2_decap_8 FILLER_14_2421 ();
 sg13g2_decap_8 FILLER_14_2428 ();
 sg13g2_decap_8 FILLER_14_2435 ();
 sg13g2_decap_8 FILLER_14_2442 ();
 sg13g2_decap_8 FILLER_14_2449 ();
 sg13g2_decap_8 FILLER_14_2456 ();
 sg13g2_decap_8 FILLER_14_2463 ();
 sg13g2_decap_8 FILLER_14_2470 ();
 sg13g2_decap_8 FILLER_14_2477 ();
 sg13g2_decap_8 FILLER_14_2484 ();
 sg13g2_decap_8 FILLER_14_2491 ();
 sg13g2_decap_8 FILLER_14_2498 ();
 sg13g2_decap_8 FILLER_14_2505 ();
 sg13g2_decap_8 FILLER_14_2512 ();
 sg13g2_decap_8 FILLER_14_2519 ();
 sg13g2_decap_8 FILLER_14_2526 ();
 sg13g2_decap_8 FILLER_14_2533 ();
 sg13g2_decap_8 FILLER_14_2540 ();
 sg13g2_decap_8 FILLER_14_2547 ();
 sg13g2_decap_8 FILLER_14_2554 ();
 sg13g2_decap_8 FILLER_14_2561 ();
 sg13g2_decap_8 FILLER_14_2568 ();
 sg13g2_decap_8 FILLER_14_2575 ();
 sg13g2_decap_8 FILLER_14_2582 ();
 sg13g2_decap_8 FILLER_14_2589 ();
 sg13g2_decap_8 FILLER_14_2596 ();
 sg13g2_decap_8 FILLER_14_2603 ();
 sg13g2_decap_8 FILLER_14_2610 ();
 sg13g2_decap_8 FILLER_14_2617 ();
 sg13g2_decap_8 FILLER_14_2624 ();
 sg13g2_decap_8 FILLER_14_2631 ();
 sg13g2_decap_8 FILLER_14_2638 ();
 sg13g2_decap_8 FILLER_14_2645 ();
 sg13g2_decap_8 FILLER_14_2652 ();
 sg13g2_decap_8 FILLER_14_2659 ();
 sg13g2_decap_4 FILLER_14_2666 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_fill_1 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_68 ();
 sg13g2_decap_8 FILLER_15_75 ();
 sg13g2_decap_8 FILLER_15_82 ();
 sg13g2_decap_8 FILLER_15_89 ();
 sg13g2_decap_8 FILLER_15_96 ();
 sg13g2_decap_8 FILLER_15_103 ();
 sg13g2_decap_8 FILLER_15_110 ();
 sg13g2_decap_8 FILLER_15_121 ();
 sg13g2_decap_8 FILLER_15_128 ();
 sg13g2_decap_8 FILLER_15_135 ();
 sg13g2_decap_8 FILLER_15_142 ();
 sg13g2_decap_8 FILLER_15_149 ();
 sg13g2_decap_8 FILLER_15_156 ();
 sg13g2_decap_8 FILLER_15_163 ();
 sg13g2_decap_8 FILLER_15_170 ();
 sg13g2_decap_8 FILLER_15_177 ();
 sg13g2_decap_8 FILLER_15_184 ();
 sg13g2_decap_8 FILLER_15_191 ();
 sg13g2_decap_8 FILLER_15_198 ();
 sg13g2_decap_8 FILLER_15_205 ();
 sg13g2_decap_8 FILLER_15_212 ();
 sg13g2_decap_8 FILLER_15_219 ();
 sg13g2_fill_1 FILLER_15_226 ();
 sg13g2_decap_4 FILLER_15_232 ();
 sg13g2_fill_1 FILLER_15_239 ();
 sg13g2_decap_8 FILLER_15_244 ();
 sg13g2_decap_8 FILLER_15_251 ();
 sg13g2_decap_8 FILLER_15_258 ();
 sg13g2_decap_8 FILLER_15_265 ();
 sg13g2_decap_8 FILLER_15_272 ();
 sg13g2_fill_2 FILLER_15_279 ();
 sg13g2_decap_8 FILLER_15_286 ();
 sg13g2_decap_8 FILLER_15_293 ();
 sg13g2_decap_8 FILLER_15_300 ();
 sg13g2_decap_8 FILLER_15_307 ();
 sg13g2_decap_8 FILLER_15_314 ();
 sg13g2_decap_8 FILLER_15_321 ();
 sg13g2_decap_8 FILLER_15_328 ();
 sg13g2_decap_8 FILLER_15_335 ();
 sg13g2_decap_8 FILLER_15_342 ();
 sg13g2_decap_8 FILLER_15_349 ();
 sg13g2_decap_8 FILLER_15_356 ();
 sg13g2_decap_8 FILLER_15_363 ();
 sg13g2_decap_8 FILLER_15_370 ();
 sg13g2_decap_8 FILLER_15_377 ();
 sg13g2_decap_8 FILLER_15_384 ();
 sg13g2_decap_8 FILLER_15_391 ();
 sg13g2_decap_8 FILLER_15_398 ();
 sg13g2_decap_8 FILLER_15_405 ();
 sg13g2_decap_8 FILLER_15_412 ();
 sg13g2_decap_8 FILLER_15_419 ();
 sg13g2_fill_2 FILLER_15_426 ();
 sg13g2_fill_1 FILLER_15_428 ();
 sg13g2_decap_8 FILLER_15_433 ();
 sg13g2_fill_2 FILLER_15_440 ();
 sg13g2_fill_1 FILLER_15_442 ();
 sg13g2_decap_8 FILLER_15_447 ();
 sg13g2_decap_4 FILLER_15_454 ();
 sg13g2_fill_2 FILLER_15_458 ();
 sg13g2_decap_8 FILLER_15_479 ();
 sg13g2_decap_8 FILLER_15_486 ();
 sg13g2_decap_8 FILLER_15_493 ();
 sg13g2_decap_8 FILLER_15_500 ();
 sg13g2_decap_8 FILLER_15_507 ();
 sg13g2_decap_8 FILLER_15_514 ();
 sg13g2_decap_8 FILLER_15_521 ();
 sg13g2_decap_8 FILLER_15_528 ();
 sg13g2_decap_8 FILLER_15_535 ();
 sg13g2_decap_4 FILLER_15_542 ();
 sg13g2_fill_2 FILLER_15_546 ();
 sg13g2_decap_8 FILLER_15_567 ();
 sg13g2_decap_8 FILLER_15_574 ();
 sg13g2_decap_4 FILLER_15_581 ();
 sg13g2_fill_1 FILLER_15_585 ();
 sg13g2_fill_1 FILLER_15_598 ();
 sg13g2_decap_4 FILLER_15_604 ();
 sg13g2_fill_1 FILLER_15_608 ();
 sg13g2_decap_8 FILLER_15_615 ();
 sg13g2_decap_8 FILLER_15_622 ();
 sg13g2_decap_8 FILLER_15_629 ();
 sg13g2_decap_8 FILLER_15_636 ();
 sg13g2_decap_8 FILLER_15_643 ();
 sg13g2_fill_1 FILLER_15_650 ();
 sg13g2_decap_8 FILLER_15_670 ();
 sg13g2_decap_8 FILLER_15_677 ();
 sg13g2_decap_8 FILLER_15_684 ();
 sg13g2_decap_8 FILLER_15_691 ();
 sg13g2_decap_8 FILLER_15_698 ();
 sg13g2_decap_8 FILLER_15_705 ();
 sg13g2_decap_8 FILLER_15_712 ();
 sg13g2_decap_8 FILLER_15_719 ();
 sg13g2_decap_8 FILLER_15_726 ();
 sg13g2_fill_1 FILLER_15_733 ();
 sg13g2_decap_8 FILLER_15_751 ();
 sg13g2_decap_8 FILLER_15_758 ();
 sg13g2_decap_8 FILLER_15_765 ();
 sg13g2_decap_8 FILLER_15_772 ();
 sg13g2_decap_8 FILLER_15_779 ();
 sg13g2_decap_8 FILLER_15_786 ();
 sg13g2_decap_8 FILLER_15_793 ();
 sg13g2_decap_8 FILLER_15_800 ();
 sg13g2_decap_8 FILLER_15_807 ();
 sg13g2_decap_8 FILLER_15_814 ();
 sg13g2_decap_4 FILLER_15_821 ();
 sg13g2_fill_1 FILLER_15_825 ();
 sg13g2_decap_8 FILLER_15_849 ();
 sg13g2_decap_8 FILLER_15_856 ();
 sg13g2_decap_8 FILLER_15_863 ();
 sg13g2_decap_8 FILLER_15_870 ();
 sg13g2_decap_8 FILLER_15_877 ();
 sg13g2_fill_1 FILLER_15_884 ();
 sg13g2_fill_2 FILLER_15_890 ();
 sg13g2_decap_8 FILLER_15_904 ();
 sg13g2_decap_8 FILLER_15_923 ();
 sg13g2_decap_8 FILLER_15_930 ();
 sg13g2_decap_8 FILLER_15_937 ();
 sg13g2_decap_8 FILLER_15_944 ();
 sg13g2_decap_4 FILLER_15_951 ();
 sg13g2_decap_8 FILLER_15_964 ();
 sg13g2_decap_8 FILLER_15_971 ();
 sg13g2_decap_8 FILLER_15_978 ();
 sg13g2_decap_8 FILLER_15_985 ();
 sg13g2_decap_8 FILLER_15_992 ();
 sg13g2_decap_8 FILLER_15_999 ();
 sg13g2_decap_8 FILLER_15_1006 ();
 sg13g2_decap_8 FILLER_15_1013 ();
 sg13g2_decap_8 FILLER_15_1020 ();
 sg13g2_decap_8 FILLER_15_1027 ();
 sg13g2_decap_8 FILLER_15_1034 ();
 sg13g2_decap_8 FILLER_15_1041 ();
 sg13g2_decap_8 FILLER_15_1048 ();
 sg13g2_decap_8 FILLER_15_1055 ();
 sg13g2_decap_8 FILLER_15_1062 ();
 sg13g2_decap_8 FILLER_15_1069 ();
 sg13g2_decap_8 FILLER_15_1076 ();
 sg13g2_fill_1 FILLER_15_1083 ();
 sg13g2_decap_8 FILLER_15_1093 ();
 sg13g2_decap_8 FILLER_15_1100 ();
 sg13g2_decap_8 FILLER_15_1107 ();
 sg13g2_decap_8 FILLER_15_1114 ();
 sg13g2_decap_8 FILLER_15_1121 ();
 sg13g2_fill_2 FILLER_15_1128 ();
 sg13g2_fill_1 FILLER_15_1130 ();
 sg13g2_fill_1 FILLER_15_1146 ();
 sg13g2_decap_8 FILLER_15_1152 ();
 sg13g2_decap_8 FILLER_15_1159 ();
 sg13g2_decap_8 FILLER_15_1166 ();
 sg13g2_decap_8 FILLER_15_1173 ();
 sg13g2_fill_1 FILLER_15_1180 ();
 sg13g2_fill_2 FILLER_15_1187 ();
 sg13g2_decap_8 FILLER_15_1193 ();
 sg13g2_decap_8 FILLER_15_1200 ();
 sg13g2_decap_8 FILLER_15_1207 ();
 sg13g2_fill_2 FILLER_15_1214 ();
 sg13g2_decap_8 FILLER_15_1219 ();
 sg13g2_decap_8 FILLER_15_1226 ();
 sg13g2_decap_8 FILLER_15_1233 ();
 sg13g2_decap_8 FILLER_15_1240 ();
 sg13g2_decap_8 FILLER_15_1247 ();
 sg13g2_decap_8 FILLER_15_1254 ();
 sg13g2_decap_8 FILLER_15_1261 ();
 sg13g2_decap_8 FILLER_15_1268 ();
 sg13g2_decap_8 FILLER_15_1275 ();
 sg13g2_decap_8 FILLER_15_1282 ();
 sg13g2_decap_8 FILLER_15_1289 ();
 sg13g2_decap_8 FILLER_15_1296 ();
 sg13g2_decap_8 FILLER_15_1303 ();
 sg13g2_decap_8 FILLER_15_1310 ();
 sg13g2_decap_8 FILLER_15_1317 ();
 sg13g2_decap_8 FILLER_15_1324 ();
 sg13g2_decap_8 FILLER_15_1331 ();
 sg13g2_decap_8 FILLER_15_1338 ();
 sg13g2_decap_8 FILLER_15_1358 ();
 sg13g2_decap_8 FILLER_15_1365 ();
 sg13g2_decap_8 FILLER_15_1372 ();
 sg13g2_fill_2 FILLER_15_1379 ();
 sg13g2_fill_1 FILLER_15_1381 ();
 sg13g2_decap_8 FILLER_15_1394 ();
 sg13g2_decap_8 FILLER_15_1401 ();
 sg13g2_decap_8 FILLER_15_1408 ();
 sg13g2_fill_1 FILLER_15_1415 ();
 sg13g2_decap_8 FILLER_15_1419 ();
 sg13g2_decap_8 FILLER_15_1426 ();
 sg13g2_decap_8 FILLER_15_1433 ();
 sg13g2_decap_8 FILLER_15_1440 ();
 sg13g2_decap_8 FILLER_15_1447 ();
 sg13g2_decap_8 FILLER_15_1454 ();
 sg13g2_decap_8 FILLER_15_1461 ();
 sg13g2_decap_8 FILLER_15_1468 ();
 sg13g2_decap_8 FILLER_15_1475 ();
 sg13g2_decap_8 FILLER_15_1482 ();
 sg13g2_decap_8 FILLER_15_1489 ();
 sg13g2_decap_8 FILLER_15_1496 ();
 sg13g2_decap_8 FILLER_15_1503 ();
 sg13g2_decap_4 FILLER_15_1510 ();
 sg13g2_fill_2 FILLER_15_1514 ();
 sg13g2_decap_8 FILLER_15_1526 ();
 sg13g2_decap_8 FILLER_15_1533 ();
 sg13g2_decap_8 FILLER_15_1540 ();
 sg13g2_decap_8 FILLER_15_1547 ();
 sg13g2_decap_8 FILLER_15_1554 ();
 sg13g2_decap_8 FILLER_15_1561 ();
 sg13g2_decap_8 FILLER_15_1568 ();
 sg13g2_decap_8 FILLER_15_1575 ();
 sg13g2_decap_8 FILLER_15_1582 ();
 sg13g2_decap_4 FILLER_15_1589 ();
 sg13g2_decap_8 FILLER_15_1602 ();
 sg13g2_decap_8 FILLER_15_1609 ();
 sg13g2_decap_4 FILLER_15_1616 ();
 sg13g2_fill_1 FILLER_15_1620 ();
 sg13g2_decap_8 FILLER_15_1625 ();
 sg13g2_decap_8 FILLER_15_1632 ();
 sg13g2_decap_4 FILLER_15_1639 ();
 sg13g2_decap_8 FILLER_15_1661 ();
 sg13g2_decap_8 FILLER_15_1668 ();
 sg13g2_decap_4 FILLER_15_1675 ();
 sg13g2_decap_8 FILLER_15_1689 ();
 sg13g2_decap_8 FILLER_15_1696 ();
 sg13g2_decap_8 FILLER_15_1703 ();
 sg13g2_decap_4 FILLER_15_1710 ();
 sg13g2_decap_4 FILLER_15_1746 ();
 sg13g2_decap_8 FILLER_15_1759 ();
 sg13g2_decap_8 FILLER_15_1766 ();
 sg13g2_decap_8 FILLER_15_1773 ();
 sg13g2_decap_8 FILLER_15_1780 ();
 sg13g2_decap_8 FILLER_15_1787 ();
 sg13g2_fill_2 FILLER_15_1794 ();
 sg13g2_fill_2 FILLER_15_1809 ();
 sg13g2_decap_8 FILLER_15_1816 ();
 sg13g2_decap_8 FILLER_15_1823 ();
 sg13g2_decap_8 FILLER_15_1830 ();
 sg13g2_decap_8 FILLER_15_1837 ();
 sg13g2_decap_8 FILLER_15_1844 ();
 sg13g2_decap_8 FILLER_15_1851 ();
 sg13g2_decap_8 FILLER_15_1858 ();
 sg13g2_decap_8 FILLER_15_1865 ();
 sg13g2_decap_8 FILLER_15_1872 ();
 sg13g2_decap_8 FILLER_15_1879 ();
 sg13g2_decap_8 FILLER_15_1886 ();
 sg13g2_decap_8 FILLER_15_1893 ();
 sg13g2_decap_8 FILLER_15_1900 ();
 sg13g2_decap_8 FILLER_15_1907 ();
 sg13g2_decap_8 FILLER_15_1914 ();
 sg13g2_decap_8 FILLER_15_1921 ();
 sg13g2_decap_8 FILLER_15_1928 ();
 sg13g2_decap_8 FILLER_15_1935 ();
 sg13g2_decap_8 FILLER_15_1942 ();
 sg13g2_decap_8 FILLER_15_1949 ();
 sg13g2_decap_8 FILLER_15_1956 ();
 sg13g2_decap_8 FILLER_15_1963 ();
 sg13g2_decap_8 FILLER_15_1970 ();
 sg13g2_decap_8 FILLER_15_1977 ();
 sg13g2_decap_8 FILLER_15_1984 ();
 sg13g2_decap_8 FILLER_15_1991 ();
 sg13g2_decap_8 FILLER_15_1998 ();
 sg13g2_decap_8 FILLER_15_2005 ();
 sg13g2_decap_8 FILLER_15_2012 ();
 sg13g2_decap_8 FILLER_15_2019 ();
 sg13g2_decap_8 FILLER_15_2026 ();
 sg13g2_decap_8 FILLER_15_2033 ();
 sg13g2_decap_8 FILLER_15_2040 ();
 sg13g2_decap_8 FILLER_15_2047 ();
 sg13g2_decap_8 FILLER_15_2054 ();
 sg13g2_decap_8 FILLER_15_2061 ();
 sg13g2_decap_8 FILLER_15_2068 ();
 sg13g2_decap_8 FILLER_15_2075 ();
 sg13g2_decap_8 FILLER_15_2082 ();
 sg13g2_decap_8 FILLER_15_2089 ();
 sg13g2_decap_8 FILLER_15_2096 ();
 sg13g2_decap_8 FILLER_15_2103 ();
 sg13g2_decap_8 FILLER_15_2110 ();
 sg13g2_decap_8 FILLER_15_2117 ();
 sg13g2_decap_8 FILLER_15_2124 ();
 sg13g2_decap_8 FILLER_15_2131 ();
 sg13g2_decap_8 FILLER_15_2138 ();
 sg13g2_decap_8 FILLER_15_2145 ();
 sg13g2_decap_8 FILLER_15_2152 ();
 sg13g2_decap_8 FILLER_15_2159 ();
 sg13g2_decap_8 FILLER_15_2166 ();
 sg13g2_decap_8 FILLER_15_2173 ();
 sg13g2_decap_8 FILLER_15_2180 ();
 sg13g2_decap_8 FILLER_15_2187 ();
 sg13g2_decap_8 FILLER_15_2194 ();
 sg13g2_decap_8 FILLER_15_2201 ();
 sg13g2_decap_8 FILLER_15_2208 ();
 sg13g2_decap_8 FILLER_15_2215 ();
 sg13g2_decap_8 FILLER_15_2222 ();
 sg13g2_decap_8 FILLER_15_2229 ();
 sg13g2_decap_8 FILLER_15_2236 ();
 sg13g2_decap_8 FILLER_15_2243 ();
 sg13g2_decap_8 FILLER_15_2250 ();
 sg13g2_decap_8 FILLER_15_2257 ();
 sg13g2_decap_8 FILLER_15_2264 ();
 sg13g2_decap_8 FILLER_15_2271 ();
 sg13g2_decap_8 FILLER_15_2278 ();
 sg13g2_decap_8 FILLER_15_2285 ();
 sg13g2_decap_8 FILLER_15_2292 ();
 sg13g2_decap_8 FILLER_15_2299 ();
 sg13g2_decap_8 FILLER_15_2306 ();
 sg13g2_decap_8 FILLER_15_2313 ();
 sg13g2_decap_8 FILLER_15_2320 ();
 sg13g2_decap_8 FILLER_15_2327 ();
 sg13g2_decap_8 FILLER_15_2334 ();
 sg13g2_decap_8 FILLER_15_2341 ();
 sg13g2_decap_8 FILLER_15_2348 ();
 sg13g2_decap_8 FILLER_15_2355 ();
 sg13g2_decap_8 FILLER_15_2362 ();
 sg13g2_decap_8 FILLER_15_2369 ();
 sg13g2_decap_8 FILLER_15_2376 ();
 sg13g2_decap_8 FILLER_15_2383 ();
 sg13g2_decap_8 FILLER_15_2390 ();
 sg13g2_decap_8 FILLER_15_2397 ();
 sg13g2_decap_8 FILLER_15_2404 ();
 sg13g2_decap_8 FILLER_15_2411 ();
 sg13g2_decap_8 FILLER_15_2418 ();
 sg13g2_decap_8 FILLER_15_2425 ();
 sg13g2_decap_8 FILLER_15_2432 ();
 sg13g2_decap_8 FILLER_15_2439 ();
 sg13g2_decap_8 FILLER_15_2446 ();
 sg13g2_decap_8 FILLER_15_2453 ();
 sg13g2_decap_8 FILLER_15_2460 ();
 sg13g2_decap_8 FILLER_15_2467 ();
 sg13g2_decap_8 FILLER_15_2474 ();
 sg13g2_decap_8 FILLER_15_2481 ();
 sg13g2_decap_8 FILLER_15_2488 ();
 sg13g2_decap_8 FILLER_15_2495 ();
 sg13g2_decap_8 FILLER_15_2502 ();
 sg13g2_decap_8 FILLER_15_2509 ();
 sg13g2_decap_8 FILLER_15_2516 ();
 sg13g2_decap_8 FILLER_15_2523 ();
 sg13g2_decap_8 FILLER_15_2530 ();
 sg13g2_decap_8 FILLER_15_2537 ();
 sg13g2_decap_8 FILLER_15_2544 ();
 sg13g2_decap_8 FILLER_15_2551 ();
 sg13g2_decap_8 FILLER_15_2558 ();
 sg13g2_decap_8 FILLER_15_2565 ();
 sg13g2_decap_8 FILLER_15_2572 ();
 sg13g2_decap_8 FILLER_15_2579 ();
 sg13g2_decap_8 FILLER_15_2586 ();
 sg13g2_decap_8 FILLER_15_2593 ();
 sg13g2_decap_8 FILLER_15_2600 ();
 sg13g2_decap_8 FILLER_15_2607 ();
 sg13g2_decap_8 FILLER_15_2614 ();
 sg13g2_decap_8 FILLER_15_2621 ();
 sg13g2_decap_8 FILLER_15_2628 ();
 sg13g2_decap_8 FILLER_15_2635 ();
 sg13g2_decap_8 FILLER_15_2642 ();
 sg13g2_decap_8 FILLER_15_2649 ();
 sg13g2_decap_8 FILLER_15_2656 ();
 sg13g2_decap_8 FILLER_15_2663 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_fill_1 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_decap_8 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_420 ();
 sg13g2_fill_2 FILLER_16_427 ();
 sg13g2_decap_8 FILLER_16_437 ();
 sg13g2_decap_8 FILLER_16_444 ();
 sg13g2_decap_8 FILLER_16_451 ();
 sg13g2_decap_8 FILLER_16_458 ();
 sg13g2_decap_8 FILLER_16_465 ();
 sg13g2_decap_8 FILLER_16_472 ();
 sg13g2_decap_8 FILLER_16_479 ();
 sg13g2_decap_8 FILLER_16_486 ();
 sg13g2_decap_8 FILLER_16_493 ();
 sg13g2_decap_8 FILLER_16_500 ();
 sg13g2_decap_8 FILLER_16_507 ();
 sg13g2_decap_8 FILLER_16_514 ();
 sg13g2_decap_8 FILLER_16_521 ();
 sg13g2_decap_8 FILLER_16_528 ();
 sg13g2_decap_8 FILLER_16_535 ();
 sg13g2_decap_8 FILLER_16_542 ();
 sg13g2_decap_8 FILLER_16_549 ();
 sg13g2_decap_8 FILLER_16_556 ();
 sg13g2_decap_8 FILLER_16_563 ();
 sg13g2_decap_8 FILLER_16_574 ();
 sg13g2_decap_8 FILLER_16_581 ();
 sg13g2_fill_1 FILLER_16_588 ();
 sg13g2_decap_8 FILLER_16_593 ();
 sg13g2_decap_8 FILLER_16_600 ();
 sg13g2_decap_8 FILLER_16_607 ();
 sg13g2_decap_4 FILLER_16_614 ();
 sg13g2_fill_1 FILLER_16_618 ();
 sg13g2_decap_8 FILLER_16_624 ();
 sg13g2_decap_8 FILLER_16_631 ();
 sg13g2_decap_8 FILLER_16_638 ();
 sg13g2_decap_8 FILLER_16_660 ();
 sg13g2_decap_4 FILLER_16_667 ();
 sg13g2_decap_8 FILLER_16_676 ();
 sg13g2_decap_8 FILLER_16_683 ();
 sg13g2_decap_8 FILLER_16_690 ();
 sg13g2_decap_8 FILLER_16_697 ();
 sg13g2_decap_4 FILLER_16_704 ();
 sg13g2_decap_8 FILLER_16_723 ();
 sg13g2_fill_1 FILLER_16_730 ();
 sg13g2_fill_1 FILLER_16_736 ();
 sg13g2_decap_8 FILLER_16_752 ();
 sg13g2_fill_1 FILLER_16_759 ();
 sg13g2_decap_8 FILLER_16_764 ();
 sg13g2_decap_8 FILLER_16_771 ();
 sg13g2_decap_8 FILLER_16_778 ();
 sg13g2_decap_8 FILLER_16_785 ();
 sg13g2_fill_1 FILLER_16_792 ();
 sg13g2_decap_4 FILLER_16_796 ();
 sg13g2_fill_2 FILLER_16_800 ();
 sg13g2_decap_8 FILLER_16_806 ();
 sg13g2_decap_8 FILLER_16_813 ();
 sg13g2_decap_8 FILLER_16_820 ();
 sg13g2_decap_8 FILLER_16_827 ();
 sg13g2_decap_8 FILLER_16_834 ();
 sg13g2_decap_8 FILLER_16_841 ();
 sg13g2_decap_8 FILLER_16_848 ();
 sg13g2_decap_8 FILLER_16_855 ();
 sg13g2_decap_8 FILLER_16_877 ();
 sg13g2_decap_4 FILLER_16_884 ();
 sg13g2_decap_8 FILLER_16_892 ();
 sg13g2_decap_8 FILLER_16_899 ();
 sg13g2_decap_8 FILLER_16_906 ();
 sg13g2_decap_8 FILLER_16_913 ();
 sg13g2_fill_1 FILLER_16_920 ();
 sg13g2_decap_8 FILLER_16_942 ();
 sg13g2_fill_2 FILLER_16_949 ();
 sg13g2_fill_1 FILLER_16_951 ();
 sg13g2_decap_8 FILLER_16_959 ();
 sg13g2_decap_8 FILLER_16_966 ();
 sg13g2_decap_8 FILLER_16_973 ();
 sg13g2_decap_8 FILLER_16_980 ();
 sg13g2_fill_1 FILLER_16_987 ();
 sg13g2_decap_8 FILLER_16_1003 ();
 sg13g2_fill_1 FILLER_16_1010 ();
 sg13g2_decap_8 FILLER_16_1015 ();
 sg13g2_decap_8 FILLER_16_1022 ();
 sg13g2_fill_2 FILLER_16_1029 ();
 sg13g2_decap_8 FILLER_16_1034 ();
 sg13g2_fill_2 FILLER_16_1041 ();
 sg13g2_fill_1 FILLER_16_1043 ();
 sg13g2_decap_8 FILLER_16_1064 ();
 sg13g2_fill_1 FILLER_16_1071 ();
 sg13g2_decap_8 FILLER_16_1076 ();
 sg13g2_fill_1 FILLER_16_1083 ();
 sg13g2_decap_8 FILLER_16_1087 ();
 sg13g2_decap_8 FILLER_16_1094 ();
 sg13g2_decap_8 FILLER_16_1101 ();
 sg13g2_decap_8 FILLER_16_1108 ();
 sg13g2_decap_8 FILLER_16_1115 ();
 sg13g2_decap_8 FILLER_16_1122 ();
 sg13g2_decap_4 FILLER_16_1129 ();
 sg13g2_fill_1 FILLER_16_1133 ();
 sg13g2_decap_8 FILLER_16_1138 ();
 sg13g2_decap_8 FILLER_16_1145 ();
 sg13g2_decap_8 FILLER_16_1152 ();
 sg13g2_decap_8 FILLER_16_1159 ();
 sg13g2_decap_8 FILLER_16_1166 ();
 sg13g2_decap_8 FILLER_16_1173 ();
 sg13g2_fill_1 FILLER_16_1180 ();
 sg13g2_decap_8 FILLER_16_1190 ();
 sg13g2_decap_8 FILLER_16_1197 ();
 sg13g2_decap_8 FILLER_16_1204 ();
 sg13g2_decap_8 FILLER_16_1211 ();
 sg13g2_decap_8 FILLER_16_1218 ();
 sg13g2_decap_8 FILLER_16_1225 ();
 sg13g2_decap_8 FILLER_16_1232 ();
 sg13g2_decap_8 FILLER_16_1239 ();
 sg13g2_decap_8 FILLER_16_1246 ();
 sg13g2_decap_8 FILLER_16_1253 ();
 sg13g2_decap_8 FILLER_16_1260 ();
 sg13g2_fill_2 FILLER_16_1267 ();
 sg13g2_fill_1 FILLER_16_1269 ();
 sg13g2_decap_8 FILLER_16_1275 ();
 sg13g2_decap_8 FILLER_16_1282 ();
 sg13g2_decap_8 FILLER_16_1289 ();
 sg13g2_decap_8 FILLER_16_1296 ();
 sg13g2_decap_8 FILLER_16_1303 ();
 sg13g2_decap_8 FILLER_16_1310 ();
 sg13g2_fill_1 FILLER_16_1329 ();
 sg13g2_fill_1 FILLER_16_1341 ();
 sg13g2_decap_8 FILLER_16_1364 ();
 sg13g2_decap_8 FILLER_16_1375 ();
 sg13g2_fill_1 FILLER_16_1386 ();
 sg13g2_decap_8 FILLER_16_1391 ();
 sg13g2_decap_8 FILLER_16_1398 ();
 sg13g2_decap_8 FILLER_16_1405 ();
 sg13g2_decap_8 FILLER_16_1412 ();
 sg13g2_decap_4 FILLER_16_1419 ();
 sg13g2_decap_8 FILLER_16_1427 ();
 sg13g2_decap_4 FILLER_16_1434 ();
 sg13g2_fill_2 FILLER_16_1438 ();
 sg13g2_decap_8 FILLER_16_1444 ();
 sg13g2_decap_8 FILLER_16_1451 ();
 sg13g2_decap_8 FILLER_16_1458 ();
 sg13g2_decap_8 FILLER_16_1465 ();
 sg13g2_decap_8 FILLER_16_1472 ();
 sg13g2_decap_8 FILLER_16_1479 ();
 sg13g2_decap_8 FILLER_16_1486 ();
 sg13g2_decap_8 FILLER_16_1493 ();
 sg13g2_decap_8 FILLER_16_1500 ();
 sg13g2_fill_2 FILLER_16_1507 ();
 sg13g2_fill_1 FILLER_16_1509 ();
 sg13g2_fill_2 FILLER_16_1516 ();
 sg13g2_fill_1 FILLER_16_1518 ();
 sg13g2_decap_8 FILLER_16_1522 ();
 sg13g2_decap_8 FILLER_16_1529 ();
 sg13g2_decap_4 FILLER_16_1536 ();
 sg13g2_fill_1 FILLER_16_1540 ();
 sg13g2_decap_8 FILLER_16_1545 ();
 sg13g2_fill_1 FILLER_16_1552 ();
 sg13g2_decap_8 FILLER_16_1561 ();
 sg13g2_decap_8 FILLER_16_1568 ();
 sg13g2_decap_8 FILLER_16_1575 ();
 sg13g2_decap_8 FILLER_16_1582 ();
 sg13g2_fill_2 FILLER_16_1589 ();
 sg13g2_decap_8 FILLER_16_1595 ();
 sg13g2_decap_8 FILLER_16_1602 ();
 sg13g2_decap_8 FILLER_16_1609 ();
 sg13g2_decap_8 FILLER_16_1616 ();
 sg13g2_fill_2 FILLER_16_1623 ();
 sg13g2_decap_8 FILLER_16_1640 ();
 sg13g2_decap_8 FILLER_16_1647 ();
 sg13g2_decap_8 FILLER_16_1657 ();
 sg13g2_decap_8 FILLER_16_1664 ();
 sg13g2_decap_8 FILLER_16_1671 ();
 sg13g2_decap_8 FILLER_16_1678 ();
 sg13g2_fill_1 FILLER_16_1685 ();
 sg13g2_decap_8 FILLER_16_1689 ();
 sg13g2_decap_8 FILLER_16_1696 ();
 sg13g2_decap_8 FILLER_16_1703 ();
 sg13g2_decap_4 FILLER_16_1710 ();
 sg13g2_fill_2 FILLER_16_1714 ();
 sg13g2_decap_8 FILLER_16_1721 ();
 sg13g2_decap_8 FILLER_16_1728 ();
 sg13g2_decap_8 FILLER_16_1735 ();
 sg13g2_decap_8 FILLER_16_1742 ();
 sg13g2_decap_8 FILLER_16_1749 ();
 sg13g2_decap_8 FILLER_16_1756 ();
 sg13g2_decap_8 FILLER_16_1763 ();
 sg13g2_decap_8 FILLER_16_1770 ();
 sg13g2_decap_8 FILLER_16_1777 ();
 sg13g2_decap_8 FILLER_16_1784 ();
 sg13g2_decap_8 FILLER_16_1791 ();
 sg13g2_decap_8 FILLER_16_1798 ();
 sg13g2_decap_8 FILLER_16_1805 ();
 sg13g2_decap_8 FILLER_16_1812 ();
 sg13g2_decap_8 FILLER_16_1819 ();
 sg13g2_decap_8 FILLER_16_1826 ();
 sg13g2_fill_2 FILLER_16_1833 ();
 sg13g2_decap_8 FILLER_16_1840 ();
 sg13g2_decap_8 FILLER_16_1847 ();
 sg13g2_decap_8 FILLER_16_1854 ();
 sg13g2_decap_8 FILLER_16_1861 ();
 sg13g2_decap_8 FILLER_16_1868 ();
 sg13g2_decap_8 FILLER_16_1875 ();
 sg13g2_decap_8 FILLER_16_1882 ();
 sg13g2_decap_8 FILLER_16_1889 ();
 sg13g2_decap_8 FILLER_16_1896 ();
 sg13g2_decap_8 FILLER_16_1903 ();
 sg13g2_decap_8 FILLER_16_1910 ();
 sg13g2_decap_8 FILLER_16_1917 ();
 sg13g2_decap_8 FILLER_16_1924 ();
 sg13g2_decap_8 FILLER_16_1931 ();
 sg13g2_decap_8 FILLER_16_1938 ();
 sg13g2_decap_8 FILLER_16_1945 ();
 sg13g2_decap_8 FILLER_16_1952 ();
 sg13g2_decap_8 FILLER_16_1959 ();
 sg13g2_decap_8 FILLER_16_1966 ();
 sg13g2_decap_8 FILLER_16_1973 ();
 sg13g2_decap_8 FILLER_16_1980 ();
 sg13g2_decap_8 FILLER_16_1987 ();
 sg13g2_decap_8 FILLER_16_1994 ();
 sg13g2_decap_8 FILLER_16_2001 ();
 sg13g2_decap_8 FILLER_16_2008 ();
 sg13g2_decap_8 FILLER_16_2015 ();
 sg13g2_decap_8 FILLER_16_2022 ();
 sg13g2_decap_8 FILLER_16_2029 ();
 sg13g2_decap_8 FILLER_16_2036 ();
 sg13g2_decap_8 FILLER_16_2043 ();
 sg13g2_decap_8 FILLER_16_2050 ();
 sg13g2_decap_8 FILLER_16_2057 ();
 sg13g2_decap_8 FILLER_16_2064 ();
 sg13g2_decap_8 FILLER_16_2071 ();
 sg13g2_decap_8 FILLER_16_2078 ();
 sg13g2_decap_8 FILLER_16_2085 ();
 sg13g2_decap_8 FILLER_16_2092 ();
 sg13g2_decap_8 FILLER_16_2099 ();
 sg13g2_decap_8 FILLER_16_2106 ();
 sg13g2_decap_8 FILLER_16_2113 ();
 sg13g2_decap_8 FILLER_16_2120 ();
 sg13g2_decap_8 FILLER_16_2127 ();
 sg13g2_decap_8 FILLER_16_2134 ();
 sg13g2_decap_8 FILLER_16_2141 ();
 sg13g2_decap_8 FILLER_16_2148 ();
 sg13g2_decap_8 FILLER_16_2155 ();
 sg13g2_decap_8 FILLER_16_2162 ();
 sg13g2_decap_8 FILLER_16_2169 ();
 sg13g2_decap_8 FILLER_16_2176 ();
 sg13g2_decap_8 FILLER_16_2183 ();
 sg13g2_decap_8 FILLER_16_2190 ();
 sg13g2_decap_8 FILLER_16_2197 ();
 sg13g2_decap_8 FILLER_16_2204 ();
 sg13g2_decap_8 FILLER_16_2211 ();
 sg13g2_decap_8 FILLER_16_2218 ();
 sg13g2_decap_8 FILLER_16_2225 ();
 sg13g2_decap_8 FILLER_16_2232 ();
 sg13g2_decap_8 FILLER_16_2239 ();
 sg13g2_decap_8 FILLER_16_2246 ();
 sg13g2_decap_8 FILLER_16_2253 ();
 sg13g2_decap_8 FILLER_16_2260 ();
 sg13g2_decap_8 FILLER_16_2267 ();
 sg13g2_decap_8 FILLER_16_2274 ();
 sg13g2_decap_8 FILLER_16_2281 ();
 sg13g2_decap_8 FILLER_16_2288 ();
 sg13g2_decap_8 FILLER_16_2295 ();
 sg13g2_decap_8 FILLER_16_2302 ();
 sg13g2_decap_8 FILLER_16_2309 ();
 sg13g2_decap_8 FILLER_16_2316 ();
 sg13g2_decap_8 FILLER_16_2323 ();
 sg13g2_decap_8 FILLER_16_2330 ();
 sg13g2_decap_8 FILLER_16_2337 ();
 sg13g2_decap_8 FILLER_16_2344 ();
 sg13g2_decap_8 FILLER_16_2351 ();
 sg13g2_decap_8 FILLER_16_2358 ();
 sg13g2_decap_8 FILLER_16_2365 ();
 sg13g2_decap_8 FILLER_16_2372 ();
 sg13g2_decap_8 FILLER_16_2379 ();
 sg13g2_decap_8 FILLER_16_2386 ();
 sg13g2_decap_8 FILLER_16_2393 ();
 sg13g2_decap_8 FILLER_16_2400 ();
 sg13g2_decap_8 FILLER_16_2407 ();
 sg13g2_decap_8 FILLER_16_2414 ();
 sg13g2_decap_8 FILLER_16_2421 ();
 sg13g2_decap_8 FILLER_16_2428 ();
 sg13g2_decap_8 FILLER_16_2435 ();
 sg13g2_decap_8 FILLER_16_2442 ();
 sg13g2_decap_8 FILLER_16_2449 ();
 sg13g2_decap_8 FILLER_16_2456 ();
 sg13g2_decap_8 FILLER_16_2463 ();
 sg13g2_decap_8 FILLER_16_2470 ();
 sg13g2_decap_8 FILLER_16_2477 ();
 sg13g2_decap_8 FILLER_16_2484 ();
 sg13g2_decap_8 FILLER_16_2491 ();
 sg13g2_decap_8 FILLER_16_2498 ();
 sg13g2_decap_8 FILLER_16_2505 ();
 sg13g2_decap_8 FILLER_16_2512 ();
 sg13g2_decap_8 FILLER_16_2519 ();
 sg13g2_decap_8 FILLER_16_2526 ();
 sg13g2_decap_8 FILLER_16_2533 ();
 sg13g2_decap_8 FILLER_16_2540 ();
 sg13g2_decap_8 FILLER_16_2547 ();
 sg13g2_decap_8 FILLER_16_2554 ();
 sg13g2_decap_8 FILLER_16_2561 ();
 sg13g2_decap_8 FILLER_16_2568 ();
 sg13g2_decap_8 FILLER_16_2575 ();
 sg13g2_decap_8 FILLER_16_2582 ();
 sg13g2_decap_8 FILLER_16_2589 ();
 sg13g2_decap_8 FILLER_16_2596 ();
 sg13g2_decap_8 FILLER_16_2603 ();
 sg13g2_decap_8 FILLER_16_2610 ();
 sg13g2_decap_8 FILLER_16_2617 ();
 sg13g2_decap_8 FILLER_16_2624 ();
 sg13g2_decap_8 FILLER_16_2631 ();
 sg13g2_decap_8 FILLER_16_2638 ();
 sg13g2_decap_8 FILLER_16_2645 ();
 sg13g2_decap_8 FILLER_16_2652 ();
 sg13g2_decap_8 FILLER_16_2659 ();
 sg13g2_decap_4 FILLER_16_2666 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_4 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_50 ();
 sg13g2_decap_8 FILLER_17_57 ();
 sg13g2_decap_8 FILLER_17_64 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_fill_1 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_100 ();
 sg13g2_decap_8 FILLER_17_107 ();
 sg13g2_decap_8 FILLER_17_114 ();
 sg13g2_fill_1 FILLER_17_121 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_4 FILLER_17_252 ();
 sg13g2_fill_2 FILLER_17_256 ();
 sg13g2_decap_8 FILLER_17_279 ();
 sg13g2_decap_8 FILLER_17_286 ();
 sg13g2_decap_8 FILLER_17_293 ();
 sg13g2_decap_8 FILLER_17_300 ();
 sg13g2_decap_8 FILLER_17_307 ();
 sg13g2_decap_8 FILLER_17_314 ();
 sg13g2_decap_8 FILLER_17_321 ();
 sg13g2_decap_8 FILLER_17_328 ();
 sg13g2_decap_8 FILLER_17_335 ();
 sg13g2_decap_8 FILLER_17_342 ();
 sg13g2_decap_8 FILLER_17_349 ();
 sg13g2_decap_8 FILLER_17_356 ();
 sg13g2_decap_8 FILLER_17_363 ();
 sg13g2_decap_8 FILLER_17_370 ();
 sg13g2_decap_8 FILLER_17_377 ();
 sg13g2_decap_8 FILLER_17_384 ();
 sg13g2_decap_8 FILLER_17_391 ();
 sg13g2_decap_8 FILLER_17_398 ();
 sg13g2_decap_8 FILLER_17_405 ();
 sg13g2_decap_8 FILLER_17_412 ();
 sg13g2_decap_8 FILLER_17_419 ();
 sg13g2_decap_8 FILLER_17_426 ();
 sg13g2_decap_8 FILLER_17_433 ();
 sg13g2_decap_8 FILLER_17_440 ();
 sg13g2_decap_8 FILLER_17_447 ();
 sg13g2_decap_8 FILLER_17_454 ();
 sg13g2_decap_8 FILLER_17_461 ();
 sg13g2_decap_8 FILLER_17_468 ();
 sg13g2_decap_8 FILLER_17_475 ();
 sg13g2_decap_8 FILLER_17_482 ();
 sg13g2_fill_1 FILLER_17_489 ();
 sg13g2_decap_8 FILLER_17_494 ();
 sg13g2_decap_4 FILLER_17_501 ();
 sg13g2_decap_8 FILLER_17_513 ();
 sg13g2_decap_8 FILLER_17_520 ();
 sg13g2_decap_8 FILLER_17_527 ();
 sg13g2_decap_8 FILLER_17_534 ();
 sg13g2_decap_8 FILLER_17_541 ();
 sg13g2_fill_2 FILLER_17_548 ();
 sg13g2_fill_1 FILLER_17_550 ();
 sg13g2_decap_8 FILLER_17_554 ();
 sg13g2_decap_8 FILLER_17_561 ();
 sg13g2_decap_8 FILLER_17_568 ();
 sg13g2_decap_8 FILLER_17_602 ();
 sg13g2_decap_8 FILLER_17_609 ();
 sg13g2_decap_8 FILLER_17_616 ();
 sg13g2_decap_8 FILLER_17_623 ();
 sg13g2_decap_8 FILLER_17_630 ();
 sg13g2_decap_8 FILLER_17_637 ();
 sg13g2_decap_4 FILLER_17_644 ();
 sg13g2_decap_8 FILLER_17_654 ();
 sg13g2_decap_8 FILLER_17_661 ();
 sg13g2_decap_8 FILLER_17_668 ();
 sg13g2_decap_8 FILLER_17_675 ();
 sg13g2_decap_8 FILLER_17_682 ();
 sg13g2_decap_8 FILLER_17_689 ();
 sg13g2_decap_4 FILLER_17_696 ();
 sg13g2_fill_1 FILLER_17_700 ();
 sg13g2_decap_4 FILLER_17_706 ();
 sg13g2_fill_1 FILLER_17_710 ();
 sg13g2_decap_8 FILLER_17_716 ();
 sg13g2_decap_4 FILLER_17_723 ();
 sg13g2_fill_1 FILLER_17_727 ();
 sg13g2_decap_4 FILLER_17_751 ();
 sg13g2_fill_2 FILLER_17_755 ();
 sg13g2_fill_1 FILLER_17_792 ();
 sg13g2_fill_1 FILLER_17_799 ();
 sg13g2_decap_8 FILLER_17_808 ();
 sg13g2_decap_8 FILLER_17_815 ();
 sg13g2_decap_8 FILLER_17_822 ();
 sg13g2_decap_8 FILLER_17_829 ();
 sg13g2_decap_8 FILLER_17_836 ();
 sg13g2_decap_8 FILLER_17_843 ();
 sg13g2_fill_1 FILLER_17_850 ();
 sg13g2_fill_2 FILLER_17_859 ();
 sg13g2_fill_1 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_17_874 ();
 sg13g2_fill_1 FILLER_17_881 ();
 sg13g2_decap_8 FILLER_17_887 ();
 sg13g2_decap_8 FILLER_17_894 ();
 sg13g2_decap_8 FILLER_17_901 ();
 sg13g2_decap_8 FILLER_17_908 ();
 sg13g2_decap_4 FILLER_17_915 ();
 sg13g2_decap_8 FILLER_17_938 ();
 sg13g2_decap_8 FILLER_17_945 ();
 sg13g2_decap_8 FILLER_17_952 ();
 sg13g2_decap_8 FILLER_17_959 ();
 sg13g2_decap_8 FILLER_17_966 ();
 sg13g2_decap_4 FILLER_17_973 ();
 sg13g2_fill_1 FILLER_17_977 ();
 sg13g2_decap_8 FILLER_17_983 ();
 sg13g2_fill_1 FILLER_17_990 ();
 sg13g2_decap_8 FILLER_17_996 ();
 sg13g2_decap_8 FILLER_17_1003 ();
 sg13g2_decap_8 FILLER_17_1010 ();
 sg13g2_decap_8 FILLER_17_1017 ();
 sg13g2_decap_8 FILLER_17_1024 ();
 sg13g2_decap_8 FILLER_17_1031 ();
 sg13g2_decap_8 FILLER_17_1038 ();
 sg13g2_decap_8 FILLER_17_1045 ();
 sg13g2_fill_1 FILLER_17_1052 ();
 sg13g2_decap_8 FILLER_17_1057 ();
 sg13g2_decap_4 FILLER_17_1064 ();
 sg13g2_decap_8 FILLER_17_1071 ();
 sg13g2_decap_8 FILLER_17_1078 ();
 sg13g2_decap_8 FILLER_17_1085 ();
 sg13g2_decap_8 FILLER_17_1092 ();
 sg13g2_decap_8 FILLER_17_1099 ();
 sg13g2_decap_8 FILLER_17_1106 ();
 sg13g2_decap_8 FILLER_17_1113 ();
 sg13g2_decap_8 FILLER_17_1120 ();
 sg13g2_decap_8 FILLER_17_1127 ();
 sg13g2_decap_8 FILLER_17_1134 ();
 sg13g2_fill_2 FILLER_17_1141 ();
 sg13g2_fill_1 FILLER_17_1143 ();
 sg13g2_decap_8 FILLER_17_1159 ();
 sg13g2_decap_8 FILLER_17_1166 ();
 sg13g2_decap_8 FILLER_17_1173 ();
 sg13g2_decap_8 FILLER_17_1180 ();
 sg13g2_decap_8 FILLER_17_1187 ();
 sg13g2_decap_8 FILLER_17_1194 ();
 sg13g2_decap_8 FILLER_17_1201 ();
 sg13g2_decap_8 FILLER_17_1208 ();
 sg13g2_decap_8 FILLER_17_1215 ();
 sg13g2_decap_8 FILLER_17_1222 ();
 sg13g2_decap_8 FILLER_17_1229 ();
 sg13g2_decap_8 FILLER_17_1236 ();
 sg13g2_decap_8 FILLER_17_1243 ();
 sg13g2_decap_8 FILLER_17_1250 ();
 sg13g2_decap_8 FILLER_17_1257 ();
 sg13g2_decap_8 FILLER_17_1264 ();
 sg13g2_decap_8 FILLER_17_1271 ();
 sg13g2_decap_8 FILLER_17_1278 ();
 sg13g2_decap_8 FILLER_17_1285 ();
 sg13g2_decap_8 FILLER_17_1292 ();
 sg13g2_decap_8 FILLER_17_1299 ();
 sg13g2_decap_4 FILLER_17_1306 ();
 sg13g2_fill_2 FILLER_17_1310 ();
 sg13g2_fill_2 FILLER_17_1343 ();
 sg13g2_decap_8 FILLER_17_1354 ();
 sg13g2_decap_8 FILLER_17_1361 ();
 sg13g2_decap_8 FILLER_17_1368 ();
 sg13g2_decap_8 FILLER_17_1375 ();
 sg13g2_decap_8 FILLER_17_1382 ();
 sg13g2_decap_8 FILLER_17_1389 ();
 sg13g2_decap_8 FILLER_17_1396 ();
 sg13g2_decap_8 FILLER_17_1403 ();
 sg13g2_decap_8 FILLER_17_1410 ();
 sg13g2_decap_8 FILLER_17_1417 ();
 sg13g2_decap_8 FILLER_17_1424 ();
 sg13g2_fill_2 FILLER_17_1431 ();
 sg13g2_fill_1 FILLER_17_1433 ();
 sg13g2_decap_8 FILLER_17_1438 ();
 sg13g2_decap_4 FILLER_17_1445 ();
 sg13g2_fill_2 FILLER_17_1449 ();
 sg13g2_decap_4 FILLER_17_1455 ();
 sg13g2_decap_8 FILLER_17_1474 ();
 sg13g2_decap_8 FILLER_17_1481 ();
 sg13g2_decap_8 FILLER_17_1488 ();
 sg13g2_decap_8 FILLER_17_1495 ();
 sg13g2_decap_8 FILLER_17_1502 ();
 sg13g2_fill_1 FILLER_17_1509 ();
 sg13g2_decap_4 FILLER_17_1519 ();
 sg13g2_fill_2 FILLER_17_1523 ();
 sg13g2_decap_8 FILLER_17_1530 ();
 sg13g2_decap_8 FILLER_17_1537 ();
 sg13g2_decap_8 FILLER_17_1544 ();
 sg13g2_decap_8 FILLER_17_1551 ();
 sg13g2_decap_8 FILLER_17_1558 ();
 sg13g2_decap_8 FILLER_17_1565 ();
 sg13g2_decap_8 FILLER_17_1572 ();
 sg13g2_decap_8 FILLER_17_1579 ();
 sg13g2_decap_8 FILLER_17_1586 ();
 sg13g2_decap_8 FILLER_17_1593 ();
 sg13g2_decap_4 FILLER_17_1600 ();
 sg13g2_fill_1 FILLER_17_1604 ();
 sg13g2_decap_8 FILLER_17_1609 ();
 sg13g2_decap_8 FILLER_17_1616 ();
 sg13g2_fill_2 FILLER_17_1623 ();
 sg13g2_decap_8 FILLER_17_1629 ();
 sg13g2_decap_8 FILLER_17_1636 ();
 sg13g2_decap_8 FILLER_17_1643 ();
 sg13g2_decap_8 FILLER_17_1650 ();
 sg13g2_decap_8 FILLER_17_1657 ();
 sg13g2_decap_8 FILLER_17_1664 ();
 sg13g2_decap_8 FILLER_17_1671 ();
 sg13g2_decap_4 FILLER_17_1678 ();
 sg13g2_fill_1 FILLER_17_1682 ();
 sg13g2_decap_8 FILLER_17_1689 ();
 sg13g2_decap_8 FILLER_17_1696 ();
 sg13g2_decap_8 FILLER_17_1703 ();
 sg13g2_decap_4 FILLER_17_1710 ();
 sg13g2_fill_1 FILLER_17_1714 ();
 sg13g2_decap_8 FILLER_17_1719 ();
 sg13g2_decap_8 FILLER_17_1726 ();
 sg13g2_decap_8 FILLER_17_1733 ();
 sg13g2_decap_8 FILLER_17_1740 ();
 sg13g2_decap_8 FILLER_17_1747 ();
 sg13g2_decap_8 FILLER_17_1754 ();
 sg13g2_decap_8 FILLER_17_1761 ();
 sg13g2_decap_8 FILLER_17_1768 ();
 sg13g2_decap_8 FILLER_17_1775 ();
 sg13g2_decap_8 FILLER_17_1782 ();
 sg13g2_decap_8 FILLER_17_1789 ();
 sg13g2_decap_8 FILLER_17_1796 ();
 sg13g2_decap_8 FILLER_17_1803 ();
 sg13g2_decap_8 FILLER_17_1810 ();
 sg13g2_decap_8 FILLER_17_1817 ();
 sg13g2_decap_8 FILLER_17_1824 ();
 sg13g2_decap_8 FILLER_17_1831 ();
 sg13g2_decap_8 FILLER_17_1838 ();
 sg13g2_decap_8 FILLER_17_1845 ();
 sg13g2_decap_8 FILLER_17_1852 ();
 sg13g2_decap_8 FILLER_17_1859 ();
 sg13g2_decap_8 FILLER_17_1866 ();
 sg13g2_decap_8 FILLER_17_1873 ();
 sg13g2_decap_8 FILLER_17_1880 ();
 sg13g2_decap_8 FILLER_17_1887 ();
 sg13g2_decap_8 FILLER_17_1894 ();
 sg13g2_decap_8 FILLER_17_1901 ();
 sg13g2_decap_8 FILLER_17_1908 ();
 sg13g2_decap_8 FILLER_17_1915 ();
 sg13g2_decap_8 FILLER_17_1922 ();
 sg13g2_decap_8 FILLER_17_1929 ();
 sg13g2_decap_8 FILLER_17_1936 ();
 sg13g2_decap_8 FILLER_17_1943 ();
 sg13g2_decap_8 FILLER_17_1950 ();
 sg13g2_decap_8 FILLER_17_1957 ();
 sg13g2_decap_8 FILLER_17_1964 ();
 sg13g2_decap_8 FILLER_17_1971 ();
 sg13g2_decap_8 FILLER_17_1978 ();
 sg13g2_decap_8 FILLER_17_1985 ();
 sg13g2_decap_8 FILLER_17_1992 ();
 sg13g2_decap_8 FILLER_17_1999 ();
 sg13g2_decap_8 FILLER_17_2006 ();
 sg13g2_decap_8 FILLER_17_2013 ();
 sg13g2_decap_8 FILLER_17_2020 ();
 sg13g2_decap_8 FILLER_17_2027 ();
 sg13g2_decap_8 FILLER_17_2034 ();
 sg13g2_decap_8 FILLER_17_2041 ();
 sg13g2_decap_8 FILLER_17_2048 ();
 sg13g2_decap_8 FILLER_17_2055 ();
 sg13g2_decap_8 FILLER_17_2062 ();
 sg13g2_decap_8 FILLER_17_2069 ();
 sg13g2_decap_8 FILLER_17_2076 ();
 sg13g2_decap_8 FILLER_17_2083 ();
 sg13g2_decap_8 FILLER_17_2090 ();
 sg13g2_decap_8 FILLER_17_2097 ();
 sg13g2_decap_8 FILLER_17_2104 ();
 sg13g2_decap_8 FILLER_17_2111 ();
 sg13g2_decap_8 FILLER_17_2118 ();
 sg13g2_decap_8 FILLER_17_2125 ();
 sg13g2_decap_8 FILLER_17_2132 ();
 sg13g2_decap_8 FILLER_17_2139 ();
 sg13g2_decap_8 FILLER_17_2146 ();
 sg13g2_decap_8 FILLER_17_2153 ();
 sg13g2_decap_8 FILLER_17_2160 ();
 sg13g2_decap_8 FILLER_17_2167 ();
 sg13g2_decap_8 FILLER_17_2174 ();
 sg13g2_decap_8 FILLER_17_2181 ();
 sg13g2_decap_8 FILLER_17_2188 ();
 sg13g2_decap_8 FILLER_17_2195 ();
 sg13g2_decap_8 FILLER_17_2202 ();
 sg13g2_decap_8 FILLER_17_2209 ();
 sg13g2_decap_8 FILLER_17_2216 ();
 sg13g2_decap_8 FILLER_17_2223 ();
 sg13g2_decap_8 FILLER_17_2230 ();
 sg13g2_decap_8 FILLER_17_2237 ();
 sg13g2_decap_8 FILLER_17_2244 ();
 sg13g2_decap_8 FILLER_17_2251 ();
 sg13g2_decap_8 FILLER_17_2258 ();
 sg13g2_decap_8 FILLER_17_2265 ();
 sg13g2_decap_8 FILLER_17_2272 ();
 sg13g2_decap_8 FILLER_17_2279 ();
 sg13g2_decap_8 FILLER_17_2286 ();
 sg13g2_decap_8 FILLER_17_2293 ();
 sg13g2_decap_8 FILLER_17_2300 ();
 sg13g2_decap_8 FILLER_17_2307 ();
 sg13g2_decap_8 FILLER_17_2314 ();
 sg13g2_decap_8 FILLER_17_2321 ();
 sg13g2_decap_8 FILLER_17_2328 ();
 sg13g2_decap_8 FILLER_17_2335 ();
 sg13g2_decap_8 FILLER_17_2342 ();
 sg13g2_decap_8 FILLER_17_2349 ();
 sg13g2_decap_8 FILLER_17_2356 ();
 sg13g2_decap_8 FILLER_17_2363 ();
 sg13g2_decap_8 FILLER_17_2370 ();
 sg13g2_decap_8 FILLER_17_2377 ();
 sg13g2_decap_8 FILLER_17_2384 ();
 sg13g2_decap_8 FILLER_17_2391 ();
 sg13g2_decap_8 FILLER_17_2398 ();
 sg13g2_decap_8 FILLER_17_2405 ();
 sg13g2_decap_8 FILLER_17_2412 ();
 sg13g2_decap_8 FILLER_17_2419 ();
 sg13g2_decap_8 FILLER_17_2426 ();
 sg13g2_decap_8 FILLER_17_2433 ();
 sg13g2_decap_8 FILLER_17_2440 ();
 sg13g2_decap_8 FILLER_17_2447 ();
 sg13g2_decap_8 FILLER_17_2454 ();
 sg13g2_decap_8 FILLER_17_2461 ();
 sg13g2_decap_8 FILLER_17_2468 ();
 sg13g2_decap_8 FILLER_17_2475 ();
 sg13g2_decap_8 FILLER_17_2482 ();
 sg13g2_decap_8 FILLER_17_2489 ();
 sg13g2_decap_8 FILLER_17_2496 ();
 sg13g2_decap_8 FILLER_17_2503 ();
 sg13g2_decap_8 FILLER_17_2510 ();
 sg13g2_decap_8 FILLER_17_2517 ();
 sg13g2_decap_8 FILLER_17_2524 ();
 sg13g2_decap_8 FILLER_17_2531 ();
 sg13g2_decap_8 FILLER_17_2538 ();
 sg13g2_decap_8 FILLER_17_2545 ();
 sg13g2_decap_8 FILLER_17_2552 ();
 sg13g2_decap_8 FILLER_17_2559 ();
 sg13g2_decap_8 FILLER_17_2566 ();
 sg13g2_decap_8 FILLER_17_2573 ();
 sg13g2_decap_8 FILLER_17_2580 ();
 sg13g2_decap_8 FILLER_17_2587 ();
 sg13g2_decap_8 FILLER_17_2594 ();
 sg13g2_decap_8 FILLER_17_2601 ();
 sg13g2_decap_8 FILLER_17_2608 ();
 sg13g2_decap_8 FILLER_17_2615 ();
 sg13g2_decap_8 FILLER_17_2622 ();
 sg13g2_decap_8 FILLER_17_2629 ();
 sg13g2_decap_8 FILLER_17_2636 ();
 sg13g2_decap_8 FILLER_17_2643 ();
 sg13g2_decap_8 FILLER_17_2650 ();
 sg13g2_decap_8 FILLER_17_2657 ();
 sg13g2_decap_4 FILLER_17_2664 ();
 sg13g2_fill_2 FILLER_17_2668 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_4 FILLER_18_42 ();
 sg13g2_fill_2 FILLER_18_46 ();
 sg13g2_decap_8 FILLER_18_78 ();
 sg13g2_decap_8 FILLER_18_85 ();
 sg13g2_decap_8 FILLER_18_92 ();
 sg13g2_decap_8 FILLER_18_99 ();
 sg13g2_decap_8 FILLER_18_106 ();
 sg13g2_decap_8 FILLER_18_113 ();
 sg13g2_decap_8 FILLER_18_120 ();
 sg13g2_decap_8 FILLER_18_135 ();
 sg13g2_decap_8 FILLER_18_142 ();
 sg13g2_decap_8 FILLER_18_149 ();
 sg13g2_decap_8 FILLER_18_156 ();
 sg13g2_fill_1 FILLER_18_163 ();
 sg13g2_decap_8 FILLER_18_169 ();
 sg13g2_decap_8 FILLER_18_176 ();
 sg13g2_decap_8 FILLER_18_183 ();
 sg13g2_decap_8 FILLER_18_190 ();
 sg13g2_decap_8 FILLER_18_197 ();
 sg13g2_decap_8 FILLER_18_204 ();
 sg13g2_decap_8 FILLER_18_211 ();
 sg13g2_decap_8 FILLER_18_218 ();
 sg13g2_decap_8 FILLER_18_225 ();
 sg13g2_decap_8 FILLER_18_232 ();
 sg13g2_decap_8 FILLER_18_239 ();
 sg13g2_decap_8 FILLER_18_246 ();
 sg13g2_decap_8 FILLER_18_253 ();
 sg13g2_fill_2 FILLER_18_260 ();
 sg13g2_fill_1 FILLER_18_262 ();
 sg13g2_fill_1 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_270 ();
 sg13g2_decap_8 FILLER_18_277 ();
 sg13g2_decap_8 FILLER_18_284 ();
 sg13g2_decap_8 FILLER_18_291 ();
 sg13g2_decap_8 FILLER_18_298 ();
 sg13g2_decap_8 FILLER_18_305 ();
 sg13g2_decap_8 FILLER_18_312 ();
 sg13g2_decap_8 FILLER_18_319 ();
 sg13g2_decap_8 FILLER_18_326 ();
 sg13g2_decap_8 FILLER_18_333 ();
 sg13g2_decap_4 FILLER_18_340 ();
 sg13g2_fill_2 FILLER_18_344 ();
 sg13g2_fill_2 FILLER_18_350 ();
 sg13g2_fill_1 FILLER_18_352 ();
 sg13g2_decap_8 FILLER_18_379 ();
 sg13g2_decap_8 FILLER_18_386 ();
 sg13g2_decap_8 FILLER_18_393 ();
 sg13g2_decap_8 FILLER_18_400 ();
 sg13g2_decap_8 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_18_414 ();
 sg13g2_decap_8 FILLER_18_421 ();
 sg13g2_decap_8 FILLER_18_428 ();
 sg13g2_decap_8 FILLER_18_444 ();
 sg13g2_decap_8 FILLER_18_451 ();
 sg13g2_decap_8 FILLER_18_458 ();
 sg13g2_decap_8 FILLER_18_465 ();
 sg13g2_fill_1 FILLER_18_472 ();
 sg13g2_decap_8 FILLER_18_477 ();
 sg13g2_decap_8 FILLER_18_484 ();
 sg13g2_decap_8 FILLER_18_491 ();
 sg13g2_fill_2 FILLER_18_498 ();
 sg13g2_fill_1 FILLER_18_500 ();
 sg13g2_decap_8 FILLER_18_506 ();
 sg13g2_decap_8 FILLER_18_513 ();
 sg13g2_decap_8 FILLER_18_520 ();
 sg13g2_decap_4 FILLER_18_527 ();
 sg13g2_fill_2 FILLER_18_535 ();
 sg13g2_fill_1 FILLER_18_537 ();
 sg13g2_fill_2 FILLER_18_566 ();
 sg13g2_fill_1 FILLER_18_568 ();
 sg13g2_decap_8 FILLER_18_585 ();
 sg13g2_decap_8 FILLER_18_600 ();
 sg13g2_decap_8 FILLER_18_607 ();
 sg13g2_decap_8 FILLER_18_614 ();
 sg13g2_decap_8 FILLER_18_621 ();
 sg13g2_decap_8 FILLER_18_628 ();
 sg13g2_decap_8 FILLER_18_635 ();
 sg13g2_fill_2 FILLER_18_642 ();
 sg13g2_fill_2 FILLER_18_648 ();
 sg13g2_fill_1 FILLER_18_650 ();
 sg13g2_decap_8 FILLER_18_654 ();
 sg13g2_fill_1 FILLER_18_661 ();
 sg13g2_decap_8 FILLER_18_681 ();
 sg13g2_decap_8 FILLER_18_698 ();
 sg13g2_decap_8 FILLER_18_705 ();
 sg13g2_decap_8 FILLER_18_712 ();
 sg13g2_decap_4 FILLER_18_719 ();
 sg13g2_fill_1 FILLER_18_733 ();
 sg13g2_decap_8 FILLER_18_741 ();
 sg13g2_decap_8 FILLER_18_748 ();
 sg13g2_decap_8 FILLER_18_755 ();
 sg13g2_fill_2 FILLER_18_762 ();
 sg13g2_fill_1 FILLER_18_764 ();
 sg13g2_fill_1 FILLER_18_785 ();
 sg13g2_decap_8 FILLER_18_808 ();
 sg13g2_decap_8 FILLER_18_815 ();
 sg13g2_decap_4 FILLER_18_822 ();
 sg13g2_fill_1 FILLER_18_826 ();
 sg13g2_decap_8 FILLER_18_831 ();
 sg13g2_decap_8 FILLER_18_838 ();
 sg13g2_decap_4 FILLER_18_845 ();
 sg13g2_decap_8 FILLER_18_878 ();
 sg13g2_decap_8 FILLER_18_885 ();
 sg13g2_decap_8 FILLER_18_892 ();
 sg13g2_decap_8 FILLER_18_899 ();
 sg13g2_decap_4 FILLER_18_906 ();
 sg13g2_decap_8 FILLER_18_916 ();
 sg13g2_decap_8 FILLER_18_923 ();
 sg13g2_decap_8 FILLER_18_939 ();
 sg13g2_decap_8 FILLER_18_946 ();
 sg13g2_decap_8 FILLER_18_953 ();
 sg13g2_decap_8 FILLER_18_960 ();
 sg13g2_decap_8 FILLER_18_967 ();
 sg13g2_decap_8 FILLER_18_974 ();
 sg13g2_decap_8 FILLER_18_981 ();
 sg13g2_decap_8 FILLER_18_988 ();
 sg13g2_decap_8 FILLER_18_999 ();
 sg13g2_decap_8 FILLER_18_1006 ();
 sg13g2_decap_8 FILLER_18_1013 ();
 sg13g2_decap_8 FILLER_18_1020 ();
 sg13g2_decap_8 FILLER_18_1027 ();
 sg13g2_decap_8 FILLER_18_1034 ();
 sg13g2_decap_8 FILLER_18_1041 ();
 sg13g2_decap_4 FILLER_18_1048 ();
 sg13g2_fill_1 FILLER_18_1052 ();
 sg13g2_decap_8 FILLER_18_1059 ();
 sg13g2_fill_2 FILLER_18_1066 ();
 sg13g2_fill_1 FILLER_18_1073 ();
 sg13g2_decap_8 FILLER_18_1080 ();
 sg13g2_decap_4 FILLER_18_1087 ();
 sg13g2_fill_2 FILLER_18_1091 ();
 sg13g2_fill_2 FILLER_18_1098 ();
 sg13g2_decap_8 FILLER_18_1105 ();
 sg13g2_decap_8 FILLER_18_1119 ();
 sg13g2_decap_8 FILLER_18_1126 ();
 sg13g2_decap_8 FILLER_18_1133 ();
 sg13g2_decap_8 FILLER_18_1140 ();
 sg13g2_decap_4 FILLER_18_1151 ();
 sg13g2_fill_1 FILLER_18_1155 ();
 sg13g2_decap_8 FILLER_18_1160 ();
 sg13g2_decap_8 FILLER_18_1167 ();
 sg13g2_decap_4 FILLER_18_1174 ();
 sg13g2_fill_2 FILLER_18_1178 ();
 sg13g2_decap_8 FILLER_18_1195 ();
 sg13g2_decap_8 FILLER_18_1202 ();
 sg13g2_decap_8 FILLER_18_1209 ();
 sg13g2_decap_8 FILLER_18_1216 ();
 sg13g2_decap_4 FILLER_18_1223 ();
 sg13g2_fill_1 FILLER_18_1227 ();
 sg13g2_decap_4 FILLER_18_1232 ();
 sg13g2_decap_8 FILLER_18_1240 ();
 sg13g2_decap_8 FILLER_18_1247 ();
 sg13g2_decap_8 FILLER_18_1254 ();
 sg13g2_decap_8 FILLER_18_1261 ();
 sg13g2_decap_8 FILLER_18_1268 ();
 sg13g2_decap_8 FILLER_18_1275 ();
 sg13g2_decap_8 FILLER_18_1282 ();
 sg13g2_decap_8 FILLER_18_1289 ();
 sg13g2_decap_8 FILLER_18_1296 ();
 sg13g2_decap_8 FILLER_18_1303 ();
 sg13g2_fill_2 FILLER_18_1310 ();
 sg13g2_fill_1 FILLER_18_1312 ();
 sg13g2_decap_8 FILLER_18_1327 ();
 sg13g2_decap_8 FILLER_18_1334 ();
 sg13g2_fill_1 FILLER_18_1341 ();
 sg13g2_decap_8 FILLER_18_1353 ();
 sg13g2_decap_4 FILLER_18_1360 ();
 sg13g2_decap_8 FILLER_18_1369 ();
 sg13g2_decap_8 FILLER_18_1376 ();
 sg13g2_decap_8 FILLER_18_1383 ();
 sg13g2_decap_8 FILLER_18_1390 ();
 sg13g2_decap_8 FILLER_18_1397 ();
 sg13g2_fill_2 FILLER_18_1404 ();
 sg13g2_fill_1 FILLER_18_1406 ();
 sg13g2_fill_2 FILLER_18_1412 ();
 sg13g2_fill_1 FILLER_18_1414 ();
 sg13g2_decap_8 FILLER_18_1420 ();
 sg13g2_decap_8 FILLER_18_1427 ();
 sg13g2_decap_8 FILLER_18_1434 ();
 sg13g2_decap_8 FILLER_18_1441 ();
 sg13g2_decap_8 FILLER_18_1448 ();
 sg13g2_decap_4 FILLER_18_1455 ();
 sg13g2_decap_4 FILLER_18_1464 ();
 sg13g2_fill_1 FILLER_18_1468 ();
 sg13g2_decap_8 FILLER_18_1475 ();
 sg13g2_decap_8 FILLER_18_1482 ();
 sg13g2_decap_8 FILLER_18_1489 ();
 sg13g2_decap_8 FILLER_18_1496 ();
 sg13g2_decap_8 FILLER_18_1503 ();
 sg13g2_decap_8 FILLER_18_1510 ();
 sg13g2_decap_8 FILLER_18_1517 ();
 sg13g2_decap_8 FILLER_18_1524 ();
 sg13g2_decap_8 FILLER_18_1531 ();
 sg13g2_decap_8 FILLER_18_1538 ();
 sg13g2_decap_8 FILLER_18_1545 ();
 sg13g2_decap_8 FILLER_18_1552 ();
 sg13g2_decap_8 FILLER_18_1559 ();
 sg13g2_decap_8 FILLER_18_1566 ();
 sg13g2_decap_8 FILLER_18_1573 ();
 sg13g2_decap_8 FILLER_18_1592 ();
 sg13g2_decap_4 FILLER_18_1599 ();
 sg13g2_fill_2 FILLER_18_1603 ();
 sg13g2_decap_4 FILLER_18_1620 ();
 sg13g2_fill_1 FILLER_18_1624 ();
 sg13g2_decap_8 FILLER_18_1631 ();
 sg13g2_decap_8 FILLER_18_1638 ();
 sg13g2_decap_8 FILLER_18_1645 ();
 sg13g2_decap_8 FILLER_18_1652 ();
 sg13g2_decap_4 FILLER_18_1659 ();
 sg13g2_fill_1 FILLER_18_1663 ();
 sg13g2_fill_2 FILLER_18_1679 ();
 sg13g2_fill_1 FILLER_18_1681 ();
 sg13g2_fill_1 FILLER_18_1685 ();
 sg13g2_fill_2 FILLER_18_1694 ();
 sg13g2_decap_8 FILLER_18_1711 ();
 sg13g2_decap_8 FILLER_18_1718 ();
 sg13g2_decap_8 FILLER_18_1725 ();
 sg13g2_decap_8 FILLER_18_1732 ();
 sg13g2_decap_8 FILLER_18_1739 ();
 sg13g2_decap_8 FILLER_18_1746 ();
 sg13g2_decap_8 FILLER_18_1753 ();
 sg13g2_decap_8 FILLER_18_1760 ();
 sg13g2_decap_8 FILLER_18_1767 ();
 sg13g2_decap_8 FILLER_18_1774 ();
 sg13g2_decap_8 FILLER_18_1781 ();
 sg13g2_decap_8 FILLER_18_1788 ();
 sg13g2_decap_8 FILLER_18_1795 ();
 sg13g2_decap_8 FILLER_18_1802 ();
 sg13g2_decap_8 FILLER_18_1809 ();
 sg13g2_decap_8 FILLER_18_1816 ();
 sg13g2_decap_8 FILLER_18_1823 ();
 sg13g2_decap_8 FILLER_18_1830 ();
 sg13g2_decap_8 FILLER_18_1837 ();
 sg13g2_decap_8 FILLER_18_1844 ();
 sg13g2_decap_8 FILLER_18_1851 ();
 sg13g2_decap_8 FILLER_18_1858 ();
 sg13g2_decap_8 FILLER_18_1865 ();
 sg13g2_decap_8 FILLER_18_1872 ();
 sg13g2_decap_8 FILLER_18_1879 ();
 sg13g2_decap_8 FILLER_18_1886 ();
 sg13g2_decap_8 FILLER_18_1893 ();
 sg13g2_decap_8 FILLER_18_1900 ();
 sg13g2_decap_8 FILLER_18_1907 ();
 sg13g2_decap_8 FILLER_18_1914 ();
 sg13g2_decap_8 FILLER_18_1921 ();
 sg13g2_decap_8 FILLER_18_1928 ();
 sg13g2_decap_8 FILLER_18_1935 ();
 sg13g2_decap_8 FILLER_18_1942 ();
 sg13g2_decap_8 FILLER_18_1949 ();
 sg13g2_decap_8 FILLER_18_1956 ();
 sg13g2_decap_8 FILLER_18_1963 ();
 sg13g2_decap_8 FILLER_18_1970 ();
 sg13g2_decap_8 FILLER_18_1977 ();
 sg13g2_decap_8 FILLER_18_1984 ();
 sg13g2_decap_8 FILLER_18_1991 ();
 sg13g2_decap_8 FILLER_18_1998 ();
 sg13g2_decap_8 FILLER_18_2005 ();
 sg13g2_decap_8 FILLER_18_2012 ();
 sg13g2_decap_8 FILLER_18_2019 ();
 sg13g2_decap_8 FILLER_18_2026 ();
 sg13g2_decap_8 FILLER_18_2033 ();
 sg13g2_decap_8 FILLER_18_2040 ();
 sg13g2_decap_8 FILLER_18_2047 ();
 sg13g2_decap_8 FILLER_18_2054 ();
 sg13g2_decap_8 FILLER_18_2061 ();
 sg13g2_decap_8 FILLER_18_2068 ();
 sg13g2_decap_8 FILLER_18_2075 ();
 sg13g2_decap_8 FILLER_18_2082 ();
 sg13g2_decap_8 FILLER_18_2089 ();
 sg13g2_decap_8 FILLER_18_2096 ();
 sg13g2_decap_8 FILLER_18_2103 ();
 sg13g2_decap_8 FILLER_18_2110 ();
 sg13g2_decap_8 FILLER_18_2117 ();
 sg13g2_decap_8 FILLER_18_2124 ();
 sg13g2_decap_8 FILLER_18_2131 ();
 sg13g2_decap_8 FILLER_18_2138 ();
 sg13g2_decap_8 FILLER_18_2145 ();
 sg13g2_decap_8 FILLER_18_2152 ();
 sg13g2_decap_8 FILLER_18_2159 ();
 sg13g2_decap_8 FILLER_18_2166 ();
 sg13g2_decap_8 FILLER_18_2173 ();
 sg13g2_decap_8 FILLER_18_2180 ();
 sg13g2_decap_8 FILLER_18_2187 ();
 sg13g2_decap_8 FILLER_18_2194 ();
 sg13g2_decap_8 FILLER_18_2201 ();
 sg13g2_decap_8 FILLER_18_2208 ();
 sg13g2_decap_8 FILLER_18_2215 ();
 sg13g2_decap_8 FILLER_18_2222 ();
 sg13g2_decap_8 FILLER_18_2229 ();
 sg13g2_decap_8 FILLER_18_2236 ();
 sg13g2_decap_8 FILLER_18_2243 ();
 sg13g2_decap_8 FILLER_18_2250 ();
 sg13g2_decap_8 FILLER_18_2257 ();
 sg13g2_decap_8 FILLER_18_2264 ();
 sg13g2_decap_8 FILLER_18_2271 ();
 sg13g2_decap_8 FILLER_18_2278 ();
 sg13g2_decap_8 FILLER_18_2285 ();
 sg13g2_decap_8 FILLER_18_2292 ();
 sg13g2_decap_8 FILLER_18_2299 ();
 sg13g2_decap_8 FILLER_18_2306 ();
 sg13g2_decap_8 FILLER_18_2313 ();
 sg13g2_decap_8 FILLER_18_2320 ();
 sg13g2_decap_8 FILLER_18_2327 ();
 sg13g2_decap_8 FILLER_18_2334 ();
 sg13g2_decap_8 FILLER_18_2341 ();
 sg13g2_decap_8 FILLER_18_2348 ();
 sg13g2_decap_8 FILLER_18_2355 ();
 sg13g2_decap_8 FILLER_18_2362 ();
 sg13g2_decap_8 FILLER_18_2369 ();
 sg13g2_decap_8 FILLER_18_2376 ();
 sg13g2_decap_8 FILLER_18_2383 ();
 sg13g2_decap_8 FILLER_18_2390 ();
 sg13g2_decap_8 FILLER_18_2397 ();
 sg13g2_decap_8 FILLER_18_2404 ();
 sg13g2_decap_8 FILLER_18_2411 ();
 sg13g2_decap_8 FILLER_18_2418 ();
 sg13g2_decap_8 FILLER_18_2425 ();
 sg13g2_decap_8 FILLER_18_2432 ();
 sg13g2_decap_8 FILLER_18_2439 ();
 sg13g2_decap_8 FILLER_18_2446 ();
 sg13g2_decap_8 FILLER_18_2453 ();
 sg13g2_decap_8 FILLER_18_2460 ();
 sg13g2_decap_8 FILLER_18_2467 ();
 sg13g2_decap_8 FILLER_18_2474 ();
 sg13g2_decap_8 FILLER_18_2481 ();
 sg13g2_decap_8 FILLER_18_2488 ();
 sg13g2_decap_8 FILLER_18_2495 ();
 sg13g2_decap_8 FILLER_18_2502 ();
 sg13g2_decap_8 FILLER_18_2509 ();
 sg13g2_decap_8 FILLER_18_2516 ();
 sg13g2_decap_8 FILLER_18_2523 ();
 sg13g2_decap_8 FILLER_18_2530 ();
 sg13g2_decap_8 FILLER_18_2537 ();
 sg13g2_decap_8 FILLER_18_2544 ();
 sg13g2_decap_8 FILLER_18_2551 ();
 sg13g2_decap_8 FILLER_18_2558 ();
 sg13g2_decap_8 FILLER_18_2565 ();
 sg13g2_decap_8 FILLER_18_2572 ();
 sg13g2_decap_8 FILLER_18_2579 ();
 sg13g2_decap_8 FILLER_18_2586 ();
 sg13g2_decap_8 FILLER_18_2593 ();
 sg13g2_decap_8 FILLER_18_2600 ();
 sg13g2_decap_8 FILLER_18_2607 ();
 sg13g2_decap_8 FILLER_18_2614 ();
 sg13g2_decap_8 FILLER_18_2621 ();
 sg13g2_decap_8 FILLER_18_2628 ();
 sg13g2_decap_8 FILLER_18_2635 ();
 sg13g2_decap_8 FILLER_18_2642 ();
 sg13g2_decap_8 FILLER_18_2649 ();
 sg13g2_decap_8 FILLER_18_2656 ();
 sg13g2_decap_8 FILLER_18_2663 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_fill_2 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_85 ();
 sg13g2_decap_8 FILLER_19_96 ();
 sg13g2_decap_8 FILLER_19_103 ();
 sg13g2_decap_8 FILLER_19_110 ();
 sg13g2_decap_8 FILLER_19_117 ();
 sg13g2_decap_8 FILLER_19_124 ();
 sg13g2_decap_8 FILLER_19_131 ();
 sg13g2_fill_1 FILLER_19_138 ();
 sg13g2_decap_8 FILLER_19_144 ();
 sg13g2_fill_1 FILLER_19_151 ();
 sg13g2_decap_8 FILLER_19_157 ();
 sg13g2_decap_4 FILLER_19_164 ();
 sg13g2_fill_2 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_174 ();
 sg13g2_decap_8 FILLER_19_181 ();
 sg13g2_fill_1 FILLER_19_188 ();
 sg13g2_decap_8 FILLER_19_193 ();
 sg13g2_decap_8 FILLER_19_200 ();
 sg13g2_decap_8 FILLER_19_207 ();
 sg13g2_decap_8 FILLER_19_214 ();
 sg13g2_decap_8 FILLER_19_221 ();
 sg13g2_decap_8 FILLER_19_228 ();
 sg13g2_decap_8 FILLER_19_235 ();
 sg13g2_decap_8 FILLER_19_242 ();
 sg13g2_fill_1 FILLER_19_249 ();
 sg13g2_fill_1 FILLER_19_255 ();
 sg13g2_fill_2 FILLER_19_261 ();
 sg13g2_decap_8 FILLER_19_275 ();
 sg13g2_decap_8 FILLER_19_282 ();
 sg13g2_decap_8 FILLER_19_289 ();
 sg13g2_decap_8 FILLER_19_296 ();
 sg13g2_decap_8 FILLER_19_303 ();
 sg13g2_decap_8 FILLER_19_310 ();
 sg13g2_decap_8 FILLER_19_317 ();
 sg13g2_decap_8 FILLER_19_324 ();
 sg13g2_decap_8 FILLER_19_331 ();
 sg13g2_decap_8 FILLER_19_338 ();
 sg13g2_decap_8 FILLER_19_345 ();
 sg13g2_fill_2 FILLER_19_352 ();
 sg13g2_fill_1 FILLER_19_354 ();
 sg13g2_decap_4 FILLER_19_359 ();
 sg13g2_fill_1 FILLER_19_363 ();
 sg13g2_decap_8 FILLER_19_370 ();
 sg13g2_fill_2 FILLER_19_377 ();
 sg13g2_fill_1 FILLER_19_379 ();
 sg13g2_decap_8 FILLER_19_388 ();
 sg13g2_decap_8 FILLER_19_395 ();
 sg13g2_decap_8 FILLER_19_402 ();
 sg13g2_decap_8 FILLER_19_409 ();
 sg13g2_decap_8 FILLER_19_416 ();
 sg13g2_decap_8 FILLER_19_423 ();
 sg13g2_decap_8 FILLER_19_430 ();
 sg13g2_decap_8 FILLER_19_437 ();
 sg13g2_decap_8 FILLER_19_444 ();
 sg13g2_decap_8 FILLER_19_451 ();
 sg13g2_decap_8 FILLER_19_458 ();
 sg13g2_fill_1 FILLER_19_465 ();
 sg13g2_decap_8 FILLER_19_482 ();
 sg13g2_decap_8 FILLER_19_489 ();
 sg13g2_decap_8 FILLER_19_496 ();
 sg13g2_decap_8 FILLER_19_503 ();
 sg13g2_decap_8 FILLER_19_510 ();
 sg13g2_decap_8 FILLER_19_517 ();
 sg13g2_decap_8 FILLER_19_524 ();
 sg13g2_decap_8 FILLER_19_531 ();
 sg13g2_decap_8 FILLER_19_538 ();
 sg13g2_fill_1 FILLER_19_545 ();
 sg13g2_decap_8 FILLER_19_550 ();
 sg13g2_decap_8 FILLER_19_557 ();
 sg13g2_decap_8 FILLER_19_564 ();
 sg13g2_decap_4 FILLER_19_571 ();
 sg13g2_fill_1 FILLER_19_575 ();
 sg13g2_decap_8 FILLER_19_583 ();
 sg13g2_fill_2 FILLER_19_590 ();
 sg13g2_fill_2 FILLER_19_596 ();
 sg13g2_decap_8 FILLER_19_602 ();
 sg13g2_decap_8 FILLER_19_609 ();
 sg13g2_decap_8 FILLER_19_616 ();
 sg13g2_decap_8 FILLER_19_623 ();
 sg13g2_decap_8 FILLER_19_630 ();
 sg13g2_decap_8 FILLER_19_637 ();
 sg13g2_decap_8 FILLER_19_644 ();
 sg13g2_decap_8 FILLER_19_654 ();
 sg13g2_decap_8 FILLER_19_661 ();
 sg13g2_fill_1 FILLER_19_668 ();
 sg13g2_decap_8 FILLER_19_675 ();
 sg13g2_decap_8 FILLER_19_682 ();
 sg13g2_decap_8 FILLER_19_689 ();
 sg13g2_decap_8 FILLER_19_696 ();
 sg13g2_decap_8 FILLER_19_703 ();
 sg13g2_decap_8 FILLER_19_710 ();
 sg13g2_decap_8 FILLER_19_717 ();
 sg13g2_decap_8 FILLER_19_724 ();
 sg13g2_decap_8 FILLER_19_749 ();
 sg13g2_decap_8 FILLER_19_756 ();
 sg13g2_decap_8 FILLER_19_763 ();
 sg13g2_decap_8 FILLER_19_770 ();
 sg13g2_decap_4 FILLER_19_777 ();
 sg13g2_decap_8 FILLER_19_788 ();
 sg13g2_fill_1 FILLER_19_795 ();
 sg13g2_decap_8 FILLER_19_801 ();
 sg13g2_decap_8 FILLER_19_808 ();
 sg13g2_decap_8 FILLER_19_815 ();
 sg13g2_decap_8 FILLER_19_822 ();
 sg13g2_decap_8 FILLER_19_829 ();
 sg13g2_decap_8 FILLER_19_836 ();
 sg13g2_decap_8 FILLER_19_843 ();
 sg13g2_decap_8 FILLER_19_850 ();
 sg13g2_decap_8 FILLER_19_857 ();
 sg13g2_decap_8 FILLER_19_864 ();
 sg13g2_decap_8 FILLER_19_871 ();
 sg13g2_decap_8 FILLER_19_878 ();
 sg13g2_decap_8 FILLER_19_885 ();
 sg13g2_decap_8 FILLER_19_892 ();
 sg13g2_decap_4 FILLER_19_899 ();
 sg13g2_fill_1 FILLER_19_903 ();
 sg13g2_fill_1 FILLER_19_914 ();
 sg13g2_decap_4 FILLER_19_920 ();
 sg13g2_fill_1 FILLER_19_924 ();
 sg13g2_decap_8 FILLER_19_929 ();
 sg13g2_decap_8 FILLER_19_936 ();
 sg13g2_decap_4 FILLER_19_943 ();
 sg13g2_fill_1 FILLER_19_947 ();
 sg13g2_decap_8 FILLER_19_957 ();
 sg13g2_fill_2 FILLER_19_964 ();
 sg13g2_fill_1 FILLER_19_966 ();
 sg13g2_decap_8 FILLER_19_971 ();
 sg13g2_decap_8 FILLER_19_978 ();
 sg13g2_decap_4 FILLER_19_985 ();
 sg13g2_fill_1 FILLER_19_989 ();
 sg13g2_decap_4 FILLER_19_1005 ();
 sg13g2_fill_2 FILLER_19_1009 ();
 sg13g2_decap_8 FILLER_19_1014 ();
 sg13g2_decap_8 FILLER_19_1021 ();
 sg13g2_decap_8 FILLER_19_1028 ();
 sg13g2_decap_8 FILLER_19_1035 ();
 sg13g2_decap_8 FILLER_19_1042 ();
 sg13g2_decap_8 FILLER_19_1049 ();
 sg13g2_decap_8 FILLER_19_1056 ();
 sg13g2_decap_8 FILLER_19_1063 ();
 sg13g2_decap_8 FILLER_19_1070 ();
 sg13g2_decap_8 FILLER_19_1077 ();
 sg13g2_decap_8 FILLER_19_1084 ();
 sg13g2_decap_4 FILLER_19_1091 ();
 sg13g2_fill_1 FILLER_19_1095 ();
 sg13g2_fill_1 FILLER_19_1101 ();
 sg13g2_decap_8 FILLER_19_1107 ();
 sg13g2_decap_8 FILLER_19_1114 ();
 sg13g2_decap_8 FILLER_19_1121 ();
 sg13g2_decap_8 FILLER_19_1128 ();
 sg13g2_decap_8 FILLER_19_1135 ();
 sg13g2_fill_2 FILLER_19_1142 ();
 sg13g2_fill_1 FILLER_19_1144 ();
 sg13g2_decap_8 FILLER_19_1149 ();
 sg13g2_decap_8 FILLER_19_1156 ();
 sg13g2_decap_8 FILLER_19_1163 ();
 sg13g2_decap_8 FILLER_19_1170 ();
 sg13g2_fill_2 FILLER_19_1177 ();
 sg13g2_fill_1 FILLER_19_1179 ();
 sg13g2_decap_8 FILLER_19_1190 ();
 sg13g2_decap_8 FILLER_19_1197 ();
 sg13g2_decap_8 FILLER_19_1204 ();
 sg13g2_decap_8 FILLER_19_1211 ();
 sg13g2_decap_8 FILLER_19_1218 ();
 sg13g2_decap_8 FILLER_19_1225 ();
 sg13g2_decap_8 FILLER_19_1232 ();
 sg13g2_decap_8 FILLER_19_1239 ();
 sg13g2_decap_4 FILLER_19_1246 ();
 sg13g2_fill_2 FILLER_19_1250 ();
 sg13g2_fill_1 FILLER_19_1256 ();
 sg13g2_decap_4 FILLER_19_1262 ();
 sg13g2_fill_1 FILLER_19_1266 ();
 sg13g2_fill_1 FILLER_19_1271 ();
 sg13g2_decap_8 FILLER_19_1276 ();
 sg13g2_decap_8 FILLER_19_1283 ();
 sg13g2_decap_8 FILLER_19_1290 ();
 sg13g2_decap_8 FILLER_19_1297 ();
 sg13g2_decap_8 FILLER_19_1304 ();
 sg13g2_decap_8 FILLER_19_1311 ();
 sg13g2_fill_2 FILLER_19_1318 ();
 sg13g2_decap_8 FILLER_19_1326 ();
 sg13g2_decap_8 FILLER_19_1333 ();
 sg13g2_decap_8 FILLER_19_1340 ();
 sg13g2_decap_8 FILLER_19_1347 ();
 sg13g2_decap_8 FILLER_19_1354 ();
 sg13g2_decap_8 FILLER_19_1361 ();
 sg13g2_decap_8 FILLER_19_1368 ();
 sg13g2_decap_8 FILLER_19_1375 ();
 sg13g2_fill_1 FILLER_19_1385 ();
 sg13g2_decap_8 FILLER_19_1395 ();
 sg13g2_decap_8 FILLER_19_1402 ();
 sg13g2_decap_8 FILLER_19_1409 ();
 sg13g2_decap_8 FILLER_19_1416 ();
 sg13g2_decap_8 FILLER_19_1423 ();
 sg13g2_decap_8 FILLER_19_1430 ();
 sg13g2_decap_8 FILLER_19_1437 ();
 sg13g2_decap_4 FILLER_19_1444 ();
 sg13g2_fill_1 FILLER_19_1448 ();
 sg13g2_decap_8 FILLER_19_1453 ();
 sg13g2_decap_4 FILLER_19_1460 ();
 sg13g2_fill_2 FILLER_19_1464 ();
 sg13g2_decap_8 FILLER_19_1482 ();
 sg13g2_decap_8 FILLER_19_1489 ();
 sg13g2_decap_8 FILLER_19_1496 ();
 sg13g2_decap_8 FILLER_19_1503 ();
 sg13g2_decap_8 FILLER_19_1510 ();
 sg13g2_fill_1 FILLER_19_1517 ();
 sg13g2_decap_8 FILLER_19_1522 ();
 sg13g2_decap_8 FILLER_19_1529 ();
 sg13g2_fill_2 FILLER_19_1536 ();
 sg13g2_fill_1 FILLER_19_1538 ();
 sg13g2_fill_2 FILLER_19_1542 ();
 sg13g2_decap_8 FILLER_19_1557 ();
 sg13g2_decap_8 FILLER_19_1564 ();
 sg13g2_decap_8 FILLER_19_1571 ();
 sg13g2_fill_2 FILLER_19_1578 ();
 sg13g2_decap_8 FILLER_19_1585 ();
 sg13g2_decap_4 FILLER_19_1592 ();
 sg13g2_fill_2 FILLER_19_1596 ();
 sg13g2_fill_1 FILLER_19_1604 ();
 sg13g2_decap_8 FILLER_19_1615 ();
 sg13g2_decap_8 FILLER_19_1622 ();
 sg13g2_decap_8 FILLER_19_1629 ();
 sg13g2_decap_8 FILLER_19_1636 ();
 sg13g2_decap_8 FILLER_19_1643 ();
 sg13g2_decap_8 FILLER_19_1650 ();
 sg13g2_decap_8 FILLER_19_1657 ();
 sg13g2_fill_2 FILLER_19_1664 ();
 sg13g2_fill_1 FILLER_19_1666 ();
 sg13g2_decap_8 FILLER_19_1671 ();
 sg13g2_decap_4 FILLER_19_1678 ();
 sg13g2_decap_8 FILLER_19_1687 ();
 sg13g2_fill_2 FILLER_19_1694 ();
 sg13g2_decap_8 FILLER_19_1700 ();
 sg13g2_decap_8 FILLER_19_1707 ();
 sg13g2_decap_8 FILLER_19_1714 ();
 sg13g2_decap_4 FILLER_19_1721 ();
 sg13g2_decap_8 FILLER_19_1733 ();
 sg13g2_decap_8 FILLER_19_1740 ();
 sg13g2_decap_8 FILLER_19_1747 ();
 sg13g2_decap_8 FILLER_19_1754 ();
 sg13g2_decap_8 FILLER_19_1761 ();
 sg13g2_decap_8 FILLER_19_1768 ();
 sg13g2_decap_4 FILLER_19_1775 ();
 sg13g2_decap_8 FILLER_19_1784 ();
 sg13g2_decap_8 FILLER_19_1791 ();
 sg13g2_decap_8 FILLER_19_1798 ();
 sg13g2_decap_8 FILLER_19_1805 ();
 sg13g2_decap_8 FILLER_19_1812 ();
 sg13g2_decap_8 FILLER_19_1819 ();
 sg13g2_decap_8 FILLER_19_1839 ();
 sg13g2_decap_8 FILLER_19_1846 ();
 sg13g2_decap_8 FILLER_19_1853 ();
 sg13g2_decap_8 FILLER_19_1860 ();
 sg13g2_decap_8 FILLER_19_1880 ();
 sg13g2_decap_8 FILLER_19_1887 ();
 sg13g2_decap_8 FILLER_19_1894 ();
 sg13g2_decap_8 FILLER_19_1901 ();
 sg13g2_decap_8 FILLER_19_1908 ();
 sg13g2_decap_8 FILLER_19_1915 ();
 sg13g2_decap_8 FILLER_19_1922 ();
 sg13g2_decap_8 FILLER_19_1929 ();
 sg13g2_decap_8 FILLER_19_1936 ();
 sg13g2_decap_8 FILLER_19_1943 ();
 sg13g2_decap_8 FILLER_19_1950 ();
 sg13g2_decap_8 FILLER_19_1957 ();
 sg13g2_decap_8 FILLER_19_1964 ();
 sg13g2_decap_8 FILLER_19_1971 ();
 sg13g2_decap_8 FILLER_19_1978 ();
 sg13g2_decap_8 FILLER_19_1985 ();
 sg13g2_decap_8 FILLER_19_1992 ();
 sg13g2_decap_8 FILLER_19_1999 ();
 sg13g2_decap_8 FILLER_19_2006 ();
 sg13g2_decap_8 FILLER_19_2013 ();
 sg13g2_decap_8 FILLER_19_2020 ();
 sg13g2_decap_8 FILLER_19_2027 ();
 sg13g2_decap_8 FILLER_19_2034 ();
 sg13g2_decap_8 FILLER_19_2041 ();
 sg13g2_decap_8 FILLER_19_2048 ();
 sg13g2_decap_8 FILLER_19_2055 ();
 sg13g2_decap_8 FILLER_19_2062 ();
 sg13g2_decap_8 FILLER_19_2069 ();
 sg13g2_decap_8 FILLER_19_2076 ();
 sg13g2_decap_8 FILLER_19_2083 ();
 sg13g2_decap_8 FILLER_19_2090 ();
 sg13g2_decap_8 FILLER_19_2097 ();
 sg13g2_decap_8 FILLER_19_2104 ();
 sg13g2_decap_8 FILLER_19_2111 ();
 sg13g2_decap_8 FILLER_19_2118 ();
 sg13g2_decap_8 FILLER_19_2125 ();
 sg13g2_decap_8 FILLER_19_2132 ();
 sg13g2_decap_8 FILLER_19_2139 ();
 sg13g2_decap_8 FILLER_19_2146 ();
 sg13g2_decap_8 FILLER_19_2153 ();
 sg13g2_decap_8 FILLER_19_2160 ();
 sg13g2_decap_8 FILLER_19_2167 ();
 sg13g2_decap_8 FILLER_19_2174 ();
 sg13g2_decap_8 FILLER_19_2181 ();
 sg13g2_decap_8 FILLER_19_2188 ();
 sg13g2_decap_8 FILLER_19_2195 ();
 sg13g2_decap_8 FILLER_19_2202 ();
 sg13g2_decap_8 FILLER_19_2209 ();
 sg13g2_decap_8 FILLER_19_2216 ();
 sg13g2_decap_8 FILLER_19_2223 ();
 sg13g2_decap_8 FILLER_19_2230 ();
 sg13g2_decap_8 FILLER_19_2237 ();
 sg13g2_decap_8 FILLER_19_2244 ();
 sg13g2_decap_8 FILLER_19_2251 ();
 sg13g2_decap_8 FILLER_19_2258 ();
 sg13g2_decap_8 FILLER_19_2265 ();
 sg13g2_decap_8 FILLER_19_2272 ();
 sg13g2_decap_8 FILLER_19_2279 ();
 sg13g2_decap_8 FILLER_19_2286 ();
 sg13g2_decap_8 FILLER_19_2293 ();
 sg13g2_decap_8 FILLER_19_2300 ();
 sg13g2_decap_8 FILLER_19_2307 ();
 sg13g2_decap_8 FILLER_19_2314 ();
 sg13g2_decap_8 FILLER_19_2321 ();
 sg13g2_decap_8 FILLER_19_2328 ();
 sg13g2_decap_8 FILLER_19_2335 ();
 sg13g2_decap_8 FILLER_19_2342 ();
 sg13g2_decap_8 FILLER_19_2349 ();
 sg13g2_decap_8 FILLER_19_2356 ();
 sg13g2_decap_8 FILLER_19_2363 ();
 sg13g2_decap_8 FILLER_19_2370 ();
 sg13g2_decap_8 FILLER_19_2377 ();
 sg13g2_decap_8 FILLER_19_2384 ();
 sg13g2_decap_8 FILLER_19_2391 ();
 sg13g2_decap_8 FILLER_19_2398 ();
 sg13g2_decap_8 FILLER_19_2405 ();
 sg13g2_decap_8 FILLER_19_2412 ();
 sg13g2_decap_8 FILLER_19_2419 ();
 sg13g2_decap_8 FILLER_19_2426 ();
 sg13g2_decap_8 FILLER_19_2433 ();
 sg13g2_decap_8 FILLER_19_2440 ();
 sg13g2_decap_8 FILLER_19_2447 ();
 sg13g2_decap_8 FILLER_19_2454 ();
 sg13g2_decap_8 FILLER_19_2461 ();
 sg13g2_decap_8 FILLER_19_2468 ();
 sg13g2_decap_8 FILLER_19_2475 ();
 sg13g2_decap_8 FILLER_19_2482 ();
 sg13g2_decap_8 FILLER_19_2489 ();
 sg13g2_decap_8 FILLER_19_2496 ();
 sg13g2_decap_8 FILLER_19_2503 ();
 sg13g2_decap_8 FILLER_19_2510 ();
 sg13g2_decap_8 FILLER_19_2517 ();
 sg13g2_decap_8 FILLER_19_2524 ();
 sg13g2_decap_8 FILLER_19_2531 ();
 sg13g2_decap_8 FILLER_19_2538 ();
 sg13g2_decap_8 FILLER_19_2545 ();
 sg13g2_decap_8 FILLER_19_2552 ();
 sg13g2_decap_8 FILLER_19_2559 ();
 sg13g2_decap_8 FILLER_19_2566 ();
 sg13g2_decap_8 FILLER_19_2573 ();
 sg13g2_decap_8 FILLER_19_2580 ();
 sg13g2_decap_8 FILLER_19_2587 ();
 sg13g2_decap_8 FILLER_19_2594 ();
 sg13g2_decap_8 FILLER_19_2601 ();
 sg13g2_decap_8 FILLER_19_2608 ();
 sg13g2_decap_8 FILLER_19_2615 ();
 sg13g2_decap_8 FILLER_19_2622 ();
 sg13g2_decap_8 FILLER_19_2629 ();
 sg13g2_decap_8 FILLER_19_2636 ();
 sg13g2_decap_8 FILLER_19_2643 ();
 sg13g2_decap_8 FILLER_19_2650 ();
 sg13g2_decap_8 FILLER_19_2657 ();
 sg13g2_decap_4 FILLER_19_2664 ();
 sg13g2_fill_2 FILLER_19_2668 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_4 FILLER_20_84 ();
 sg13g2_fill_2 FILLER_20_88 ();
 sg13g2_decap_8 FILLER_20_100 ();
 sg13g2_decap_8 FILLER_20_107 ();
 sg13g2_decap_8 FILLER_20_114 ();
 sg13g2_decap_8 FILLER_20_121 ();
 sg13g2_decap_4 FILLER_20_128 ();
 sg13g2_fill_1 FILLER_20_136 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_4 FILLER_20_175 ();
 sg13g2_fill_2 FILLER_20_179 ();
 sg13g2_decap_8 FILLER_20_207 ();
 sg13g2_decap_8 FILLER_20_214 ();
 sg13g2_decap_8 FILLER_20_221 ();
 sg13g2_decap_8 FILLER_20_228 ();
 sg13g2_fill_2 FILLER_20_235 ();
 sg13g2_fill_1 FILLER_20_247 ();
 sg13g2_decap_8 FILLER_20_279 ();
 sg13g2_decap_4 FILLER_20_286 ();
 sg13g2_fill_2 FILLER_20_290 ();
 sg13g2_decap_8 FILLER_20_303 ();
 sg13g2_decap_8 FILLER_20_310 ();
 sg13g2_decap_8 FILLER_20_317 ();
 sg13g2_decap_8 FILLER_20_324 ();
 sg13g2_decap_8 FILLER_20_331 ();
 sg13g2_decap_8 FILLER_20_338 ();
 sg13g2_decap_8 FILLER_20_345 ();
 sg13g2_decap_8 FILLER_20_352 ();
 sg13g2_decap_8 FILLER_20_359 ();
 sg13g2_decap_8 FILLER_20_366 ();
 sg13g2_decap_8 FILLER_20_373 ();
 sg13g2_decap_8 FILLER_20_380 ();
 sg13g2_decap_8 FILLER_20_387 ();
 sg13g2_decap_8 FILLER_20_394 ();
 sg13g2_decap_8 FILLER_20_401 ();
 sg13g2_decap_8 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_20_415 ();
 sg13g2_decap_8 FILLER_20_422 ();
 sg13g2_decap_8 FILLER_20_429 ();
 sg13g2_decap_8 FILLER_20_436 ();
 sg13g2_decap_8 FILLER_20_443 ();
 sg13g2_decap_8 FILLER_20_450 ();
 sg13g2_fill_2 FILLER_20_470 ();
 sg13g2_decap_8 FILLER_20_482 ();
 sg13g2_decap_8 FILLER_20_489 ();
 sg13g2_decap_8 FILLER_20_496 ();
 sg13g2_fill_2 FILLER_20_503 ();
 sg13g2_decap_8 FILLER_20_509 ();
 sg13g2_fill_2 FILLER_20_516 ();
 sg13g2_fill_1 FILLER_20_518 ();
 sg13g2_decap_8 FILLER_20_524 ();
 sg13g2_decap_8 FILLER_20_531 ();
 sg13g2_decap_8 FILLER_20_538 ();
 sg13g2_decap_8 FILLER_20_545 ();
 sg13g2_decap_8 FILLER_20_552 ();
 sg13g2_decap_8 FILLER_20_559 ();
 sg13g2_decap_8 FILLER_20_566 ();
 sg13g2_decap_4 FILLER_20_573 ();
 sg13g2_fill_2 FILLER_20_577 ();
 sg13g2_decap_8 FILLER_20_582 ();
 sg13g2_fill_2 FILLER_20_589 ();
 sg13g2_fill_1 FILLER_20_591 ();
 sg13g2_decap_8 FILLER_20_601 ();
 sg13g2_decap_8 FILLER_20_608 ();
 sg13g2_decap_8 FILLER_20_615 ();
 sg13g2_decap_8 FILLER_20_622 ();
 sg13g2_decap_8 FILLER_20_629 ();
 sg13g2_decap_8 FILLER_20_636 ();
 sg13g2_decap_8 FILLER_20_643 ();
 sg13g2_decap_8 FILLER_20_650 ();
 sg13g2_decap_8 FILLER_20_657 ();
 sg13g2_decap_8 FILLER_20_664 ();
 sg13g2_decap_8 FILLER_20_671 ();
 sg13g2_decap_8 FILLER_20_678 ();
 sg13g2_decap_8 FILLER_20_685 ();
 sg13g2_decap_8 FILLER_20_692 ();
 sg13g2_decap_8 FILLER_20_699 ();
 sg13g2_decap_8 FILLER_20_706 ();
 sg13g2_decap_8 FILLER_20_713 ();
 sg13g2_decap_8 FILLER_20_720 ();
 sg13g2_decap_8 FILLER_20_727 ();
 sg13g2_fill_2 FILLER_20_734 ();
 sg13g2_fill_1 FILLER_20_736 ();
 sg13g2_decap_4 FILLER_20_740 ();
 sg13g2_fill_1 FILLER_20_744 ();
 sg13g2_fill_2 FILLER_20_748 ();
 sg13g2_fill_1 FILLER_20_750 ();
 sg13g2_decap_8 FILLER_20_757 ();
 sg13g2_decap_8 FILLER_20_764 ();
 sg13g2_decap_8 FILLER_20_771 ();
 sg13g2_decap_8 FILLER_20_778 ();
 sg13g2_decap_8 FILLER_20_785 ();
 sg13g2_fill_1 FILLER_20_792 ();
 sg13g2_decap_8 FILLER_20_808 ();
 sg13g2_fill_2 FILLER_20_815 ();
 sg13g2_decap_8 FILLER_20_820 ();
 sg13g2_decap_8 FILLER_20_827 ();
 sg13g2_decap_8 FILLER_20_834 ();
 sg13g2_decap_8 FILLER_20_841 ();
 sg13g2_decap_8 FILLER_20_848 ();
 sg13g2_fill_1 FILLER_20_873 ();
 sg13g2_decap_8 FILLER_20_886 ();
 sg13g2_decap_8 FILLER_20_893 ();
 sg13g2_decap_8 FILLER_20_900 ();
 sg13g2_fill_2 FILLER_20_907 ();
 sg13g2_decap_8 FILLER_20_913 ();
 sg13g2_decap_8 FILLER_20_920 ();
 sg13g2_decap_8 FILLER_20_927 ();
 sg13g2_decap_8 FILLER_20_934 ();
 sg13g2_decap_8 FILLER_20_941 ();
 sg13g2_decap_8 FILLER_20_948 ();
 sg13g2_decap_8 FILLER_20_955 ();
 sg13g2_decap_8 FILLER_20_962 ();
 sg13g2_decap_8 FILLER_20_969 ();
 sg13g2_decap_8 FILLER_20_976 ();
 sg13g2_fill_1 FILLER_20_983 ();
 sg13g2_decap_8 FILLER_20_1001 ();
 sg13g2_decap_8 FILLER_20_1018 ();
 sg13g2_decap_4 FILLER_20_1025 ();
 sg13g2_fill_2 FILLER_20_1029 ();
 sg13g2_decap_8 FILLER_20_1055 ();
 sg13g2_decap_8 FILLER_20_1062 ();
 sg13g2_decap_4 FILLER_20_1069 ();
 sg13g2_fill_2 FILLER_20_1073 ();
 sg13g2_decap_8 FILLER_20_1078 ();
 sg13g2_decap_8 FILLER_20_1085 ();
 sg13g2_decap_8 FILLER_20_1092 ();
 sg13g2_decap_8 FILLER_20_1099 ();
 sg13g2_decap_8 FILLER_20_1106 ();
 sg13g2_decap_8 FILLER_20_1113 ();
 sg13g2_decap_8 FILLER_20_1120 ();
 sg13g2_decap_8 FILLER_20_1127 ();
 sg13g2_decap_8 FILLER_20_1134 ();
 sg13g2_decap_8 FILLER_20_1141 ();
 sg13g2_decap_8 FILLER_20_1148 ();
 sg13g2_fill_2 FILLER_20_1155 ();
 sg13g2_fill_1 FILLER_20_1157 ();
 sg13g2_decap_8 FILLER_20_1161 ();
 sg13g2_decap_8 FILLER_20_1168 ();
 sg13g2_decap_8 FILLER_20_1175 ();
 sg13g2_fill_1 FILLER_20_1182 ();
 sg13g2_decap_8 FILLER_20_1189 ();
 sg13g2_decap_8 FILLER_20_1196 ();
 sg13g2_decap_8 FILLER_20_1203 ();
 sg13g2_decap_8 FILLER_20_1210 ();
 sg13g2_decap_8 FILLER_20_1217 ();
 sg13g2_decap_8 FILLER_20_1224 ();
 sg13g2_decap_8 FILLER_20_1231 ();
 sg13g2_decap_4 FILLER_20_1238 ();
 sg13g2_decap_8 FILLER_20_1246 ();
 sg13g2_decap_8 FILLER_20_1253 ();
 sg13g2_decap_8 FILLER_20_1260 ();
 sg13g2_decap_8 FILLER_20_1267 ();
 sg13g2_decap_8 FILLER_20_1274 ();
 sg13g2_decap_8 FILLER_20_1281 ();
 sg13g2_decap_8 FILLER_20_1288 ();
 sg13g2_decap_8 FILLER_20_1295 ();
 sg13g2_decap_8 FILLER_20_1302 ();
 sg13g2_decap_8 FILLER_20_1309 ();
 sg13g2_fill_2 FILLER_20_1316 ();
 sg13g2_fill_1 FILLER_20_1318 ();
 sg13g2_decap_8 FILLER_20_1334 ();
 sg13g2_decap_8 FILLER_20_1341 ();
 sg13g2_decap_4 FILLER_20_1348 ();
 sg13g2_decap_8 FILLER_20_1355 ();
 sg13g2_decap_8 FILLER_20_1362 ();
 sg13g2_decap_4 FILLER_20_1369 ();
 sg13g2_fill_1 FILLER_20_1382 ();
 sg13g2_decap_8 FILLER_20_1395 ();
 sg13g2_decap_8 FILLER_20_1402 ();
 sg13g2_decap_8 FILLER_20_1409 ();
 sg13g2_decap_8 FILLER_20_1416 ();
 sg13g2_decap_8 FILLER_20_1423 ();
 sg13g2_decap_8 FILLER_20_1430 ();
 sg13g2_decap_8 FILLER_20_1437 ();
 sg13g2_decap_8 FILLER_20_1444 ();
 sg13g2_decap_4 FILLER_20_1451 ();
 sg13g2_decap_8 FILLER_20_1460 ();
 sg13g2_fill_2 FILLER_20_1467 ();
 sg13g2_decap_8 FILLER_20_1473 ();
 sg13g2_decap_8 FILLER_20_1480 ();
 sg13g2_decap_8 FILLER_20_1487 ();
 sg13g2_decap_8 FILLER_20_1494 ();
 sg13g2_decap_8 FILLER_20_1501 ();
 sg13g2_decap_8 FILLER_20_1508 ();
 sg13g2_decap_8 FILLER_20_1515 ();
 sg13g2_decap_4 FILLER_20_1522 ();
 sg13g2_fill_1 FILLER_20_1526 ();
 sg13g2_decap_8 FILLER_20_1531 ();
 sg13g2_fill_1 FILLER_20_1538 ();
 sg13g2_decap_8 FILLER_20_1555 ();
 sg13g2_fill_1 FILLER_20_1562 ();
 sg13g2_decap_8 FILLER_20_1567 ();
 sg13g2_decap_8 FILLER_20_1574 ();
 sg13g2_decap_8 FILLER_20_1581 ();
 sg13g2_decap_8 FILLER_20_1588 ();
 sg13g2_fill_2 FILLER_20_1595 ();
 sg13g2_fill_1 FILLER_20_1597 ();
 sg13g2_decap_8 FILLER_20_1608 ();
 sg13g2_decap_8 FILLER_20_1615 ();
 sg13g2_decap_4 FILLER_20_1622 ();
 sg13g2_decap_8 FILLER_20_1644 ();
 sg13g2_decap_8 FILLER_20_1651 ();
 sg13g2_decap_8 FILLER_20_1658 ();
 sg13g2_decap_4 FILLER_20_1665 ();
 sg13g2_fill_1 FILLER_20_1678 ();
 sg13g2_decap_8 FILLER_20_1683 ();
 sg13g2_decap_8 FILLER_20_1690 ();
 sg13g2_decap_8 FILLER_20_1697 ();
 sg13g2_decap_8 FILLER_20_1704 ();
 sg13g2_fill_1 FILLER_20_1711 ();
 sg13g2_decap_8 FILLER_20_1721 ();
 sg13g2_decap_8 FILLER_20_1728 ();
 sg13g2_decap_8 FILLER_20_1735 ();
 sg13g2_decap_8 FILLER_20_1742 ();
 sg13g2_decap_8 FILLER_20_1749 ();
 sg13g2_decap_8 FILLER_20_1756 ();
 sg13g2_decap_8 FILLER_20_1763 ();
 sg13g2_decap_8 FILLER_20_1770 ();
 sg13g2_decap_8 FILLER_20_1785 ();
 sg13g2_decap_8 FILLER_20_1792 ();
 sg13g2_decap_4 FILLER_20_1799 ();
 sg13g2_fill_2 FILLER_20_1803 ();
 sg13g2_decap_8 FILLER_20_1817 ();
 sg13g2_decap_8 FILLER_20_1824 ();
 sg13g2_decap_8 FILLER_20_1831 ();
 sg13g2_decap_8 FILLER_20_1838 ();
 sg13g2_decap_8 FILLER_20_1845 ();
 sg13g2_decap_8 FILLER_20_1852 ();
 sg13g2_decap_8 FILLER_20_1859 ();
 sg13g2_decap_8 FILLER_20_1866 ();
 sg13g2_decap_8 FILLER_20_1873 ();
 sg13g2_decap_8 FILLER_20_1880 ();
 sg13g2_decap_8 FILLER_20_1887 ();
 sg13g2_decap_8 FILLER_20_1894 ();
 sg13g2_decap_8 FILLER_20_1901 ();
 sg13g2_decap_8 FILLER_20_1908 ();
 sg13g2_decap_8 FILLER_20_1915 ();
 sg13g2_decap_8 FILLER_20_1922 ();
 sg13g2_decap_8 FILLER_20_1929 ();
 sg13g2_decap_8 FILLER_20_1936 ();
 sg13g2_decap_8 FILLER_20_1943 ();
 sg13g2_decap_8 FILLER_20_1950 ();
 sg13g2_decap_8 FILLER_20_1957 ();
 sg13g2_decap_8 FILLER_20_1964 ();
 sg13g2_decap_8 FILLER_20_1971 ();
 sg13g2_decap_8 FILLER_20_1978 ();
 sg13g2_decap_8 FILLER_20_1985 ();
 sg13g2_decap_8 FILLER_20_1992 ();
 sg13g2_decap_8 FILLER_20_1999 ();
 sg13g2_decap_8 FILLER_20_2006 ();
 sg13g2_decap_8 FILLER_20_2013 ();
 sg13g2_decap_8 FILLER_20_2020 ();
 sg13g2_decap_8 FILLER_20_2027 ();
 sg13g2_decap_8 FILLER_20_2034 ();
 sg13g2_decap_8 FILLER_20_2041 ();
 sg13g2_decap_8 FILLER_20_2048 ();
 sg13g2_decap_8 FILLER_20_2055 ();
 sg13g2_decap_8 FILLER_20_2062 ();
 sg13g2_decap_8 FILLER_20_2069 ();
 sg13g2_decap_8 FILLER_20_2076 ();
 sg13g2_decap_8 FILLER_20_2083 ();
 sg13g2_decap_8 FILLER_20_2090 ();
 sg13g2_decap_8 FILLER_20_2097 ();
 sg13g2_decap_8 FILLER_20_2104 ();
 sg13g2_decap_8 FILLER_20_2111 ();
 sg13g2_decap_8 FILLER_20_2118 ();
 sg13g2_decap_8 FILLER_20_2125 ();
 sg13g2_decap_8 FILLER_20_2132 ();
 sg13g2_decap_8 FILLER_20_2139 ();
 sg13g2_decap_8 FILLER_20_2146 ();
 sg13g2_decap_8 FILLER_20_2153 ();
 sg13g2_decap_8 FILLER_20_2160 ();
 sg13g2_decap_8 FILLER_20_2167 ();
 sg13g2_decap_8 FILLER_20_2174 ();
 sg13g2_decap_8 FILLER_20_2181 ();
 sg13g2_decap_8 FILLER_20_2188 ();
 sg13g2_decap_8 FILLER_20_2195 ();
 sg13g2_decap_8 FILLER_20_2202 ();
 sg13g2_decap_8 FILLER_20_2209 ();
 sg13g2_decap_8 FILLER_20_2216 ();
 sg13g2_decap_8 FILLER_20_2223 ();
 sg13g2_decap_8 FILLER_20_2230 ();
 sg13g2_decap_8 FILLER_20_2237 ();
 sg13g2_decap_8 FILLER_20_2244 ();
 sg13g2_decap_8 FILLER_20_2251 ();
 sg13g2_decap_8 FILLER_20_2258 ();
 sg13g2_decap_8 FILLER_20_2265 ();
 sg13g2_decap_8 FILLER_20_2272 ();
 sg13g2_decap_8 FILLER_20_2279 ();
 sg13g2_decap_8 FILLER_20_2286 ();
 sg13g2_decap_8 FILLER_20_2293 ();
 sg13g2_decap_8 FILLER_20_2300 ();
 sg13g2_decap_8 FILLER_20_2307 ();
 sg13g2_decap_8 FILLER_20_2314 ();
 sg13g2_decap_8 FILLER_20_2321 ();
 sg13g2_decap_8 FILLER_20_2328 ();
 sg13g2_decap_8 FILLER_20_2335 ();
 sg13g2_decap_8 FILLER_20_2342 ();
 sg13g2_decap_8 FILLER_20_2349 ();
 sg13g2_decap_8 FILLER_20_2356 ();
 sg13g2_decap_8 FILLER_20_2363 ();
 sg13g2_decap_8 FILLER_20_2370 ();
 sg13g2_decap_8 FILLER_20_2377 ();
 sg13g2_decap_8 FILLER_20_2384 ();
 sg13g2_decap_8 FILLER_20_2391 ();
 sg13g2_decap_8 FILLER_20_2398 ();
 sg13g2_decap_8 FILLER_20_2405 ();
 sg13g2_decap_8 FILLER_20_2412 ();
 sg13g2_decap_8 FILLER_20_2419 ();
 sg13g2_decap_8 FILLER_20_2426 ();
 sg13g2_decap_8 FILLER_20_2433 ();
 sg13g2_decap_8 FILLER_20_2440 ();
 sg13g2_decap_8 FILLER_20_2447 ();
 sg13g2_decap_8 FILLER_20_2454 ();
 sg13g2_decap_8 FILLER_20_2461 ();
 sg13g2_decap_8 FILLER_20_2468 ();
 sg13g2_decap_8 FILLER_20_2475 ();
 sg13g2_decap_8 FILLER_20_2482 ();
 sg13g2_decap_8 FILLER_20_2489 ();
 sg13g2_decap_8 FILLER_20_2496 ();
 sg13g2_decap_8 FILLER_20_2503 ();
 sg13g2_decap_8 FILLER_20_2510 ();
 sg13g2_decap_8 FILLER_20_2517 ();
 sg13g2_decap_8 FILLER_20_2524 ();
 sg13g2_decap_8 FILLER_20_2531 ();
 sg13g2_decap_8 FILLER_20_2538 ();
 sg13g2_decap_8 FILLER_20_2545 ();
 sg13g2_decap_8 FILLER_20_2552 ();
 sg13g2_decap_8 FILLER_20_2559 ();
 sg13g2_decap_8 FILLER_20_2566 ();
 sg13g2_decap_8 FILLER_20_2573 ();
 sg13g2_decap_8 FILLER_20_2580 ();
 sg13g2_decap_8 FILLER_20_2587 ();
 sg13g2_decap_8 FILLER_20_2594 ();
 sg13g2_decap_8 FILLER_20_2601 ();
 sg13g2_decap_8 FILLER_20_2608 ();
 sg13g2_decap_8 FILLER_20_2615 ();
 sg13g2_decap_8 FILLER_20_2622 ();
 sg13g2_decap_8 FILLER_20_2629 ();
 sg13g2_decap_8 FILLER_20_2636 ();
 sg13g2_decap_8 FILLER_20_2643 ();
 sg13g2_decap_8 FILLER_20_2650 ();
 sg13g2_decap_8 FILLER_20_2657 ();
 sg13g2_decap_4 FILLER_20_2664 ();
 sg13g2_fill_2 FILLER_20_2668 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_fill_1 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_92 ();
 sg13g2_decap_8 FILLER_21_99 ();
 sg13g2_decap_4 FILLER_21_106 ();
 sg13g2_decap_8 FILLER_21_115 ();
 sg13g2_decap_8 FILLER_21_122 ();
 sg13g2_decap_8 FILLER_21_129 ();
 sg13g2_decap_8 FILLER_21_136 ();
 sg13g2_decap_8 FILLER_21_143 ();
 sg13g2_decap_8 FILLER_21_150 ();
 sg13g2_decap_8 FILLER_21_157 ();
 sg13g2_decap_8 FILLER_21_164 ();
 sg13g2_decap_8 FILLER_21_171 ();
 sg13g2_decap_4 FILLER_21_178 ();
 sg13g2_fill_2 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_188 ();
 sg13g2_decap_8 FILLER_21_195 ();
 sg13g2_decap_8 FILLER_21_202 ();
 sg13g2_decap_8 FILLER_21_209 ();
 sg13g2_decap_8 FILLER_21_216 ();
 sg13g2_decap_8 FILLER_21_223 ();
 sg13g2_decap_8 FILLER_21_230 ();
 sg13g2_decap_8 FILLER_21_237 ();
 sg13g2_decap_8 FILLER_21_244 ();
 sg13g2_decap_8 FILLER_21_251 ();
 sg13g2_decap_8 FILLER_21_258 ();
 sg13g2_decap_8 FILLER_21_265 ();
 sg13g2_decap_8 FILLER_21_272 ();
 sg13g2_decap_8 FILLER_21_279 ();
 sg13g2_decap_8 FILLER_21_286 ();
 sg13g2_decap_8 FILLER_21_293 ();
 sg13g2_decap_8 FILLER_21_300 ();
 sg13g2_decap_8 FILLER_21_307 ();
 sg13g2_decap_8 FILLER_21_314 ();
 sg13g2_decap_8 FILLER_21_321 ();
 sg13g2_decap_8 FILLER_21_328 ();
 sg13g2_decap_8 FILLER_21_335 ();
 sg13g2_decap_4 FILLER_21_342 ();
 sg13g2_fill_2 FILLER_21_346 ();
 sg13g2_fill_1 FILLER_21_360 ();
 sg13g2_decap_8 FILLER_21_368 ();
 sg13g2_decap_8 FILLER_21_375 ();
 sg13g2_decap_8 FILLER_21_382 ();
 sg13g2_decap_8 FILLER_21_389 ();
 sg13g2_decap_8 FILLER_21_396 ();
 sg13g2_decap_8 FILLER_21_403 ();
 sg13g2_decap_8 FILLER_21_410 ();
 sg13g2_decap_8 FILLER_21_417 ();
 sg13g2_decap_8 FILLER_21_424 ();
 sg13g2_decap_4 FILLER_21_431 ();
 sg13g2_fill_2 FILLER_21_435 ();
 sg13g2_decap_4 FILLER_21_443 ();
 sg13g2_fill_1 FILLER_21_447 ();
 sg13g2_decap_8 FILLER_21_471 ();
 sg13g2_decap_8 FILLER_21_478 ();
 sg13g2_decap_8 FILLER_21_485 ();
 sg13g2_decap_8 FILLER_21_492 ();
 sg13g2_fill_1 FILLER_21_499 ();
 sg13g2_decap_8 FILLER_21_504 ();
 sg13g2_decap_8 FILLER_21_515 ();
 sg13g2_decap_8 FILLER_21_522 ();
 sg13g2_decap_8 FILLER_21_529 ();
 sg13g2_decap_8 FILLER_21_536 ();
 sg13g2_decap_8 FILLER_21_543 ();
 sg13g2_decap_8 FILLER_21_550 ();
 sg13g2_decap_8 FILLER_21_557 ();
 sg13g2_decap_8 FILLER_21_564 ();
 sg13g2_decap_8 FILLER_21_571 ();
 sg13g2_decap_8 FILLER_21_578 ();
 sg13g2_fill_2 FILLER_21_585 ();
 sg13g2_decap_8 FILLER_21_602 ();
 sg13g2_fill_2 FILLER_21_609 ();
 sg13g2_fill_1 FILLER_21_611 ();
 sg13g2_decap_8 FILLER_21_624 ();
 sg13g2_decap_8 FILLER_21_631 ();
 sg13g2_decap_8 FILLER_21_638 ();
 sg13g2_decap_8 FILLER_21_645 ();
 sg13g2_decap_8 FILLER_21_652 ();
 sg13g2_decap_8 FILLER_21_674 ();
 sg13g2_decap_8 FILLER_21_681 ();
 sg13g2_fill_2 FILLER_21_688 ();
 sg13g2_decap_8 FILLER_21_694 ();
 sg13g2_decap_8 FILLER_21_701 ();
 sg13g2_decap_8 FILLER_21_708 ();
 sg13g2_decap_4 FILLER_21_715 ();
 sg13g2_fill_2 FILLER_21_728 ();
 sg13g2_fill_1 FILLER_21_739 ();
 sg13g2_fill_2 FILLER_21_743 ();
 sg13g2_fill_1 FILLER_21_750 ();
 sg13g2_decap_8 FILLER_21_761 ();
 sg13g2_decap_8 FILLER_21_768 ();
 sg13g2_decap_8 FILLER_21_775 ();
 sg13g2_decap_8 FILLER_21_782 ();
 sg13g2_decap_8 FILLER_21_789 ();
 sg13g2_decap_8 FILLER_21_796 ();
 sg13g2_decap_8 FILLER_21_803 ();
 sg13g2_decap_8 FILLER_21_810 ();
 sg13g2_decap_8 FILLER_21_821 ();
 sg13g2_decap_8 FILLER_21_828 ();
 sg13g2_decap_4 FILLER_21_835 ();
 sg13g2_fill_1 FILLER_21_839 ();
 sg13g2_decap_8 FILLER_21_845 ();
 sg13g2_decap_8 FILLER_21_852 ();
 sg13g2_decap_8 FILLER_21_859 ();
 sg13g2_decap_4 FILLER_21_866 ();
 sg13g2_decap_8 FILLER_21_879 ();
 sg13g2_decap_8 FILLER_21_886 ();
 sg13g2_decap_8 FILLER_21_893 ();
 sg13g2_decap_8 FILLER_21_900 ();
 sg13g2_fill_2 FILLER_21_907 ();
 sg13g2_fill_1 FILLER_21_909 ();
 sg13g2_fill_2 FILLER_21_916 ();
 sg13g2_decap_8 FILLER_21_927 ();
 sg13g2_decap_8 FILLER_21_934 ();
 sg13g2_decap_8 FILLER_21_941 ();
 sg13g2_decap_8 FILLER_21_948 ();
 sg13g2_decap_8 FILLER_21_955 ();
 sg13g2_decap_8 FILLER_21_962 ();
 sg13g2_decap_8 FILLER_21_969 ();
 sg13g2_decap_8 FILLER_21_976 ();
 sg13g2_decap_8 FILLER_21_983 ();
 sg13g2_fill_2 FILLER_21_990 ();
 sg13g2_fill_1 FILLER_21_992 ();
 sg13g2_fill_1 FILLER_21_996 ();
 sg13g2_decap_8 FILLER_21_1001 ();
 sg13g2_decap_8 FILLER_21_1008 ();
 sg13g2_decap_8 FILLER_21_1015 ();
 sg13g2_decap_8 FILLER_21_1022 ();
 sg13g2_decap_4 FILLER_21_1029 ();
 sg13g2_fill_1 FILLER_21_1039 ();
 sg13g2_decap_8 FILLER_21_1051 ();
 sg13g2_decap_8 FILLER_21_1058 ();
 sg13g2_decap_8 FILLER_21_1065 ();
 sg13g2_decap_8 FILLER_21_1072 ();
 sg13g2_decap_8 FILLER_21_1079 ();
 sg13g2_decap_8 FILLER_21_1086 ();
 sg13g2_decap_8 FILLER_21_1093 ();
 sg13g2_decap_8 FILLER_21_1100 ();
 sg13g2_decap_8 FILLER_21_1107 ();
 sg13g2_decap_8 FILLER_21_1114 ();
 sg13g2_decap_8 FILLER_21_1121 ();
 sg13g2_decap_4 FILLER_21_1128 ();
 sg13g2_fill_2 FILLER_21_1132 ();
 sg13g2_decap_8 FILLER_21_1138 ();
 sg13g2_decap_8 FILLER_21_1145 ();
 sg13g2_decap_4 FILLER_21_1152 ();
 sg13g2_fill_2 FILLER_21_1156 ();
 sg13g2_decap_8 FILLER_21_1163 ();
 sg13g2_decap_8 FILLER_21_1170 ();
 sg13g2_decap_8 FILLER_21_1177 ();
 sg13g2_decap_4 FILLER_21_1184 ();
 sg13g2_fill_1 FILLER_21_1188 ();
 sg13g2_decap_8 FILLER_21_1193 ();
 sg13g2_decap_4 FILLER_21_1200 ();
 sg13g2_decap_8 FILLER_21_1218 ();
 sg13g2_decap_8 FILLER_21_1225 ();
 sg13g2_decap_8 FILLER_21_1232 ();
 sg13g2_decap_4 FILLER_21_1239 ();
 sg13g2_fill_1 FILLER_21_1243 ();
 sg13g2_decap_8 FILLER_21_1250 ();
 sg13g2_decap_4 FILLER_21_1257 ();
 sg13g2_decap_8 FILLER_21_1265 ();
 sg13g2_decap_8 FILLER_21_1272 ();
 sg13g2_decap_8 FILLER_21_1279 ();
 sg13g2_decap_8 FILLER_21_1286 ();
 sg13g2_decap_8 FILLER_21_1293 ();
 sg13g2_decap_8 FILLER_21_1300 ();
 sg13g2_decap_4 FILLER_21_1307 ();
 sg13g2_fill_2 FILLER_21_1311 ();
 sg13g2_decap_8 FILLER_21_1329 ();
 sg13g2_decap_8 FILLER_21_1336 ();
 sg13g2_decap_4 FILLER_21_1343 ();
 sg13g2_fill_2 FILLER_21_1347 ();
 sg13g2_decap_8 FILLER_21_1361 ();
 sg13g2_decap_4 FILLER_21_1368 ();
 sg13g2_fill_1 FILLER_21_1372 ();
 sg13g2_decap_8 FILLER_21_1377 ();
 sg13g2_decap_8 FILLER_21_1384 ();
 sg13g2_decap_8 FILLER_21_1391 ();
 sg13g2_decap_8 FILLER_21_1398 ();
 sg13g2_decap_8 FILLER_21_1405 ();
 sg13g2_decap_8 FILLER_21_1412 ();
 sg13g2_decap_8 FILLER_21_1419 ();
 sg13g2_decap_8 FILLER_21_1426 ();
 sg13g2_decap_8 FILLER_21_1433 ();
 sg13g2_decap_8 FILLER_21_1444 ();
 sg13g2_decap_8 FILLER_21_1451 ();
 sg13g2_decap_8 FILLER_21_1458 ();
 sg13g2_decap_8 FILLER_21_1465 ();
 sg13g2_decap_8 FILLER_21_1476 ();
 sg13g2_decap_8 FILLER_21_1483 ();
 sg13g2_decap_8 FILLER_21_1490 ();
 sg13g2_decap_8 FILLER_21_1497 ();
 sg13g2_decap_4 FILLER_21_1504 ();
 sg13g2_fill_1 FILLER_21_1508 ();
 sg13g2_decap_8 FILLER_21_1521 ();
 sg13g2_decap_8 FILLER_21_1528 ();
 sg13g2_decap_8 FILLER_21_1535 ();
 sg13g2_decap_8 FILLER_21_1542 ();
 sg13g2_decap_8 FILLER_21_1549 ();
 sg13g2_decap_8 FILLER_21_1556 ();
 sg13g2_decap_4 FILLER_21_1563 ();
 sg13g2_fill_2 FILLER_21_1567 ();
 sg13g2_decap_4 FILLER_21_1573 ();
 sg13g2_fill_2 FILLER_21_1577 ();
 sg13g2_decap_8 FILLER_21_1583 ();
 sg13g2_decap_8 FILLER_21_1590 ();
 sg13g2_fill_1 FILLER_21_1597 ();
 sg13g2_decap_8 FILLER_21_1604 ();
 sg13g2_decap_4 FILLER_21_1611 ();
 sg13g2_fill_2 FILLER_21_1615 ();
 sg13g2_decap_8 FILLER_21_1641 ();
 sg13g2_decap_4 FILLER_21_1648 ();
 sg13g2_decap_8 FILLER_21_1658 ();
 sg13g2_decap_8 FILLER_21_1665 ();
 sg13g2_fill_2 FILLER_21_1672 ();
 sg13g2_decap_8 FILLER_21_1689 ();
 sg13g2_fill_2 FILLER_21_1696 ();
 sg13g2_fill_1 FILLER_21_1698 ();
 sg13g2_fill_2 FILLER_21_1702 ();
 sg13g2_decap_8 FILLER_21_1719 ();
 sg13g2_decap_4 FILLER_21_1726 ();
 sg13g2_fill_1 FILLER_21_1730 ();
 sg13g2_decap_8 FILLER_21_1735 ();
 sg13g2_decap_4 FILLER_21_1742 ();
 sg13g2_fill_1 FILLER_21_1746 ();
 sg13g2_decap_8 FILLER_21_1753 ();
 sg13g2_decap_8 FILLER_21_1760 ();
 sg13g2_decap_8 FILLER_21_1767 ();
 sg13g2_decap_8 FILLER_21_1774 ();
 sg13g2_decap_8 FILLER_21_1781 ();
 sg13g2_decap_8 FILLER_21_1788 ();
 sg13g2_decap_8 FILLER_21_1795 ();
 sg13g2_decap_8 FILLER_21_1802 ();
 sg13g2_decap_8 FILLER_21_1809 ();
 sg13g2_decap_8 FILLER_21_1816 ();
 sg13g2_decap_8 FILLER_21_1823 ();
 sg13g2_decap_8 FILLER_21_1830 ();
 sg13g2_decap_8 FILLER_21_1837 ();
 sg13g2_decap_8 FILLER_21_1844 ();
 sg13g2_decap_8 FILLER_21_1851 ();
 sg13g2_decap_8 FILLER_21_1858 ();
 sg13g2_decap_8 FILLER_21_1865 ();
 sg13g2_decap_8 FILLER_21_1872 ();
 sg13g2_decap_8 FILLER_21_1879 ();
 sg13g2_decap_8 FILLER_21_1886 ();
 sg13g2_decap_8 FILLER_21_1893 ();
 sg13g2_decap_8 FILLER_21_1900 ();
 sg13g2_decap_8 FILLER_21_1907 ();
 sg13g2_decap_8 FILLER_21_1914 ();
 sg13g2_decap_8 FILLER_21_1921 ();
 sg13g2_decap_8 FILLER_21_1928 ();
 sg13g2_decap_8 FILLER_21_1935 ();
 sg13g2_decap_8 FILLER_21_1942 ();
 sg13g2_decap_8 FILLER_21_1949 ();
 sg13g2_decap_8 FILLER_21_1956 ();
 sg13g2_decap_8 FILLER_21_1963 ();
 sg13g2_decap_8 FILLER_21_1970 ();
 sg13g2_decap_8 FILLER_21_1977 ();
 sg13g2_decap_8 FILLER_21_1984 ();
 sg13g2_decap_8 FILLER_21_1991 ();
 sg13g2_decap_8 FILLER_21_1998 ();
 sg13g2_decap_8 FILLER_21_2005 ();
 sg13g2_decap_8 FILLER_21_2012 ();
 sg13g2_decap_8 FILLER_21_2019 ();
 sg13g2_decap_8 FILLER_21_2026 ();
 sg13g2_decap_8 FILLER_21_2033 ();
 sg13g2_decap_8 FILLER_21_2040 ();
 sg13g2_decap_8 FILLER_21_2047 ();
 sg13g2_decap_8 FILLER_21_2054 ();
 sg13g2_decap_8 FILLER_21_2061 ();
 sg13g2_decap_8 FILLER_21_2068 ();
 sg13g2_decap_8 FILLER_21_2075 ();
 sg13g2_decap_8 FILLER_21_2082 ();
 sg13g2_decap_8 FILLER_21_2089 ();
 sg13g2_decap_8 FILLER_21_2096 ();
 sg13g2_decap_8 FILLER_21_2103 ();
 sg13g2_decap_8 FILLER_21_2110 ();
 sg13g2_decap_8 FILLER_21_2117 ();
 sg13g2_decap_8 FILLER_21_2124 ();
 sg13g2_decap_8 FILLER_21_2131 ();
 sg13g2_decap_8 FILLER_21_2138 ();
 sg13g2_decap_8 FILLER_21_2145 ();
 sg13g2_decap_8 FILLER_21_2152 ();
 sg13g2_decap_8 FILLER_21_2159 ();
 sg13g2_decap_8 FILLER_21_2166 ();
 sg13g2_decap_8 FILLER_21_2173 ();
 sg13g2_decap_8 FILLER_21_2180 ();
 sg13g2_decap_8 FILLER_21_2187 ();
 sg13g2_decap_8 FILLER_21_2194 ();
 sg13g2_decap_8 FILLER_21_2201 ();
 sg13g2_decap_8 FILLER_21_2208 ();
 sg13g2_decap_8 FILLER_21_2215 ();
 sg13g2_decap_8 FILLER_21_2222 ();
 sg13g2_decap_8 FILLER_21_2229 ();
 sg13g2_decap_8 FILLER_21_2236 ();
 sg13g2_decap_8 FILLER_21_2243 ();
 sg13g2_decap_8 FILLER_21_2250 ();
 sg13g2_decap_8 FILLER_21_2257 ();
 sg13g2_decap_8 FILLER_21_2264 ();
 sg13g2_decap_8 FILLER_21_2271 ();
 sg13g2_decap_8 FILLER_21_2278 ();
 sg13g2_decap_8 FILLER_21_2285 ();
 sg13g2_decap_8 FILLER_21_2292 ();
 sg13g2_decap_8 FILLER_21_2299 ();
 sg13g2_decap_8 FILLER_21_2306 ();
 sg13g2_decap_8 FILLER_21_2313 ();
 sg13g2_decap_8 FILLER_21_2320 ();
 sg13g2_decap_8 FILLER_21_2327 ();
 sg13g2_decap_8 FILLER_21_2334 ();
 sg13g2_decap_8 FILLER_21_2341 ();
 sg13g2_decap_8 FILLER_21_2348 ();
 sg13g2_decap_8 FILLER_21_2355 ();
 sg13g2_decap_8 FILLER_21_2362 ();
 sg13g2_decap_8 FILLER_21_2369 ();
 sg13g2_decap_8 FILLER_21_2376 ();
 sg13g2_decap_8 FILLER_21_2383 ();
 sg13g2_decap_8 FILLER_21_2390 ();
 sg13g2_decap_8 FILLER_21_2397 ();
 sg13g2_decap_8 FILLER_21_2404 ();
 sg13g2_decap_8 FILLER_21_2411 ();
 sg13g2_decap_8 FILLER_21_2418 ();
 sg13g2_decap_8 FILLER_21_2425 ();
 sg13g2_decap_8 FILLER_21_2432 ();
 sg13g2_decap_8 FILLER_21_2439 ();
 sg13g2_decap_8 FILLER_21_2446 ();
 sg13g2_decap_8 FILLER_21_2453 ();
 sg13g2_decap_8 FILLER_21_2460 ();
 sg13g2_decap_8 FILLER_21_2467 ();
 sg13g2_decap_8 FILLER_21_2474 ();
 sg13g2_decap_8 FILLER_21_2481 ();
 sg13g2_decap_8 FILLER_21_2488 ();
 sg13g2_decap_8 FILLER_21_2495 ();
 sg13g2_decap_8 FILLER_21_2502 ();
 sg13g2_decap_8 FILLER_21_2509 ();
 sg13g2_decap_8 FILLER_21_2516 ();
 sg13g2_decap_8 FILLER_21_2523 ();
 sg13g2_decap_8 FILLER_21_2530 ();
 sg13g2_decap_8 FILLER_21_2537 ();
 sg13g2_decap_8 FILLER_21_2544 ();
 sg13g2_decap_8 FILLER_21_2551 ();
 sg13g2_decap_8 FILLER_21_2558 ();
 sg13g2_decap_8 FILLER_21_2565 ();
 sg13g2_decap_8 FILLER_21_2572 ();
 sg13g2_decap_8 FILLER_21_2579 ();
 sg13g2_decap_8 FILLER_21_2586 ();
 sg13g2_decap_8 FILLER_21_2593 ();
 sg13g2_decap_8 FILLER_21_2600 ();
 sg13g2_decap_8 FILLER_21_2607 ();
 sg13g2_decap_8 FILLER_21_2614 ();
 sg13g2_decap_8 FILLER_21_2621 ();
 sg13g2_decap_8 FILLER_21_2628 ();
 sg13g2_decap_8 FILLER_21_2635 ();
 sg13g2_decap_8 FILLER_21_2642 ();
 sg13g2_decap_8 FILLER_21_2649 ();
 sg13g2_decap_8 FILLER_21_2656 ();
 sg13g2_decap_8 FILLER_21_2663 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_4 FILLER_22_49 ();
 sg13g2_fill_2 FILLER_22_53 ();
 sg13g2_decap_8 FILLER_22_59 ();
 sg13g2_fill_1 FILLER_22_66 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_fill_2 FILLER_22_336 ();
 sg13g2_fill_1 FILLER_22_338 ();
 sg13g2_fill_1 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_349 ();
 sg13g2_fill_1 FILLER_22_356 ();
 sg13g2_fill_2 FILLER_22_361 ();
 sg13g2_fill_1 FILLER_22_363 ();
 sg13g2_decap_8 FILLER_22_370 ();
 sg13g2_decap_8 FILLER_22_377 ();
 sg13g2_decap_8 FILLER_22_384 ();
 sg13g2_decap_8 FILLER_22_391 ();
 sg13g2_decap_8 FILLER_22_398 ();
 sg13g2_decap_8 FILLER_22_405 ();
 sg13g2_decap_8 FILLER_22_420 ();
 sg13g2_decap_4 FILLER_22_427 ();
 sg13g2_decap_4 FILLER_22_444 ();
 sg13g2_fill_1 FILLER_22_448 ();
 sg13g2_decap_8 FILLER_22_454 ();
 sg13g2_decap_8 FILLER_22_461 ();
 sg13g2_decap_8 FILLER_22_471 ();
 sg13g2_decap_8 FILLER_22_478 ();
 sg13g2_decap_8 FILLER_22_485 ();
 sg13g2_decap_8 FILLER_22_492 ();
 sg13g2_decap_8 FILLER_22_499 ();
 sg13g2_decap_8 FILLER_22_506 ();
 sg13g2_decap_8 FILLER_22_513 ();
 sg13g2_decap_8 FILLER_22_520 ();
 sg13g2_decap_4 FILLER_22_527 ();
 sg13g2_fill_1 FILLER_22_531 ();
 sg13g2_decap_8 FILLER_22_548 ();
 sg13g2_decap_8 FILLER_22_555 ();
 sg13g2_decap_4 FILLER_22_562 ();
 sg13g2_fill_1 FILLER_22_566 ();
 sg13g2_decap_4 FILLER_22_570 ();
 sg13g2_fill_2 FILLER_22_574 ();
 sg13g2_decap_8 FILLER_22_580 ();
 sg13g2_fill_2 FILLER_22_587 ();
 sg13g2_fill_1 FILLER_22_589 ();
 sg13g2_decap_4 FILLER_22_595 ();
 sg13g2_fill_1 FILLER_22_599 ();
 sg13g2_decap_8 FILLER_22_620 ();
 sg13g2_decap_8 FILLER_22_627 ();
 sg13g2_decap_8 FILLER_22_634 ();
 sg13g2_decap_8 FILLER_22_641 ();
 sg13g2_decap_8 FILLER_22_648 ();
 sg13g2_decap_4 FILLER_22_655 ();
 sg13g2_decap_8 FILLER_22_669 ();
 sg13g2_fill_2 FILLER_22_676 ();
 sg13g2_fill_1 FILLER_22_690 ();
 sg13g2_decap_8 FILLER_22_699 ();
 sg13g2_decap_8 FILLER_22_706 ();
 sg13g2_decap_8 FILLER_22_713 ();
 sg13g2_decap_4 FILLER_22_720 ();
 sg13g2_fill_1 FILLER_22_724 ();
 sg13g2_fill_1 FILLER_22_729 ();
 sg13g2_fill_2 FILLER_22_734 ();
 sg13g2_fill_1 FILLER_22_736 ();
 sg13g2_fill_2 FILLER_22_746 ();
 sg13g2_decap_8 FILLER_22_755 ();
 sg13g2_decap_8 FILLER_22_762 ();
 sg13g2_decap_8 FILLER_22_769 ();
 sg13g2_decap_4 FILLER_22_776 ();
 sg13g2_fill_1 FILLER_22_780 ();
 sg13g2_decap_8 FILLER_22_784 ();
 sg13g2_decap_8 FILLER_22_791 ();
 sg13g2_decap_8 FILLER_22_798 ();
 sg13g2_decap_8 FILLER_22_805 ();
 sg13g2_fill_1 FILLER_22_812 ();
 sg13g2_decap_8 FILLER_22_821 ();
 sg13g2_decap_8 FILLER_22_828 ();
 sg13g2_fill_2 FILLER_22_835 ();
 sg13g2_decap_8 FILLER_22_841 ();
 sg13g2_decap_8 FILLER_22_860 ();
 sg13g2_decap_8 FILLER_22_867 ();
 sg13g2_decap_8 FILLER_22_874 ();
 sg13g2_decap_8 FILLER_22_881 ();
 sg13g2_decap_8 FILLER_22_888 ();
 sg13g2_decap_8 FILLER_22_895 ();
 sg13g2_fill_2 FILLER_22_902 ();
 sg13g2_fill_1 FILLER_22_904 ();
 sg13g2_fill_2 FILLER_22_916 ();
 sg13g2_decap_8 FILLER_22_930 ();
 sg13g2_decap_8 FILLER_22_937 ();
 sg13g2_decap_8 FILLER_22_944 ();
 sg13g2_decap_8 FILLER_22_951 ();
 sg13g2_decap_8 FILLER_22_958 ();
 sg13g2_fill_2 FILLER_22_965 ();
 sg13g2_decap_4 FILLER_22_972 ();
 sg13g2_decap_8 FILLER_22_983 ();
 sg13g2_decap_8 FILLER_22_990 ();
 sg13g2_decap_8 FILLER_22_997 ();
 sg13g2_decap_8 FILLER_22_1004 ();
 sg13g2_decap_8 FILLER_22_1016 ();
 sg13g2_decap_8 FILLER_22_1023 ();
 sg13g2_decap_8 FILLER_22_1030 ();
 sg13g2_decap_8 FILLER_22_1037 ();
 sg13g2_decap_8 FILLER_22_1048 ();
 sg13g2_decap_8 FILLER_22_1055 ();
 sg13g2_decap_8 FILLER_22_1062 ();
 sg13g2_decap_4 FILLER_22_1069 ();
 sg13g2_decap_8 FILLER_22_1077 ();
 sg13g2_decap_8 FILLER_22_1084 ();
 sg13g2_fill_2 FILLER_22_1091 ();
 sg13g2_fill_2 FILLER_22_1096 ();
 sg13g2_decap_8 FILLER_22_1105 ();
 sg13g2_decap_4 FILLER_22_1112 ();
 sg13g2_fill_1 FILLER_22_1116 ();
 sg13g2_decap_8 FILLER_22_1120 ();
 sg13g2_decap_8 FILLER_22_1127 ();
 sg13g2_decap_8 FILLER_22_1139 ();
 sg13g2_decap_8 FILLER_22_1149 ();
 sg13g2_decap_8 FILLER_22_1156 ();
 sg13g2_decap_8 FILLER_22_1163 ();
 sg13g2_decap_8 FILLER_22_1170 ();
 sg13g2_decap_4 FILLER_22_1177 ();
 sg13g2_fill_1 FILLER_22_1181 ();
 sg13g2_decap_8 FILLER_22_1186 ();
 sg13g2_decap_8 FILLER_22_1193 ();
 sg13g2_decap_8 FILLER_22_1200 ();
 sg13g2_decap_8 FILLER_22_1212 ();
 sg13g2_decap_8 FILLER_22_1219 ();
 sg13g2_decap_8 FILLER_22_1226 ();
 sg13g2_decap_8 FILLER_22_1233 ();
 sg13g2_decap_8 FILLER_22_1240 ();
 sg13g2_decap_8 FILLER_22_1247 ();
 sg13g2_decap_8 FILLER_22_1254 ();
 sg13g2_decap_8 FILLER_22_1261 ();
 sg13g2_fill_2 FILLER_22_1268 ();
 sg13g2_decap_8 FILLER_22_1274 ();
 sg13g2_decap_8 FILLER_22_1281 ();
 sg13g2_decap_8 FILLER_22_1288 ();
 sg13g2_decap_8 FILLER_22_1295 ();
 sg13g2_decap_8 FILLER_22_1302 ();
 sg13g2_decap_8 FILLER_22_1309 ();
 sg13g2_decap_4 FILLER_22_1316 ();
 sg13g2_fill_2 FILLER_22_1320 ();
 sg13g2_decap_8 FILLER_22_1325 ();
 sg13g2_decap_8 FILLER_22_1332 ();
 sg13g2_decap_8 FILLER_22_1339 ();
 sg13g2_decap_4 FILLER_22_1346 ();
 sg13g2_fill_2 FILLER_22_1350 ();
 sg13g2_fill_1 FILLER_22_1356 ();
 sg13g2_fill_1 FILLER_22_1375 ();
 sg13g2_decap_8 FILLER_22_1387 ();
 sg13g2_decap_4 FILLER_22_1394 ();
 sg13g2_decap_8 FILLER_22_1407 ();
 sg13g2_fill_2 FILLER_22_1414 ();
 sg13g2_fill_1 FILLER_22_1416 ();
 sg13g2_decap_8 FILLER_22_1432 ();
 sg13g2_fill_1 FILLER_22_1439 ();
 sg13g2_decap_8 FILLER_22_1455 ();
 sg13g2_fill_2 FILLER_22_1462 ();
 sg13g2_fill_2 FILLER_22_1470 ();
 sg13g2_fill_1 FILLER_22_1472 ();
 sg13g2_decap_8 FILLER_22_1479 ();
 sg13g2_decap_8 FILLER_22_1486 ();
 sg13g2_decap_8 FILLER_22_1493 ();
 sg13g2_decap_4 FILLER_22_1500 ();
 sg13g2_fill_2 FILLER_22_1504 ();
 sg13g2_decap_8 FILLER_22_1526 ();
 sg13g2_decap_8 FILLER_22_1533 ();
 sg13g2_decap_8 FILLER_22_1540 ();
 sg13g2_decap_8 FILLER_22_1547 ();
 sg13g2_decap_8 FILLER_22_1554 ();
 sg13g2_decap_8 FILLER_22_1561 ();
 sg13g2_decap_8 FILLER_22_1568 ();
 sg13g2_decap_8 FILLER_22_1575 ();
 sg13g2_decap_8 FILLER_22_1582 ();
 sg13g2_decap_8 FILLER_22_1589 ();
 sg13g2_decap_8 FILLER_22_1596 ();
 sg13g2_decap_8 FILLER_22_1603 ();
 sg13g2_decap_8 FILLER_22_1610 ();
 sg13g2_decap_8 FILLER_22_1617 ();
 sg13g2_decap_8 FILLER_22_1624 ();
 sg13g2_decap_8 FILLER_22_1631 ();
 sg13g2_decap_8 FILLER_22_1638 ();
 sg13g2_decap_8 FILLER_22_1645 ();
 sg13g2_decap_8 FILLER_22_1652 ();
 sg13g2_decap_8 FILLER_22_1659 ();
 sg13g2_decap_8 FILLER_22_1666 ();
 sg13g2_fill_1 FILLER_22_1673 ();
 sg13g2_decap_8 FILLER_22_1678 ();
 sg13g2_decap_8 FILLER_22_1685 ();
 sg13g2_decap_4 FILLER_22_1692 ();
 sg13g2_fill_2 FILLER_22_1696 ();
 sg13g2_fill_2 FILLER_22_1702 ();
 sg13g2_decap_8 FILLER_22_1710 ();
 sg13g2_decap_8 FILLER_22_1717 ();
 sg13g2_decap_8 FILLER_22_1724 ();
 sg13g2_fill_2 FILLER_22_1731 ();
 sg13g2_fill_1 FILLER_22_1733 ();
 sg13g2_decap_8 FILLER_22_1740 ();
 sg13g2_decap_8 FILLER_22_1747 ();
 sg13g2_decap_8 FILLER_22_1754 ();
 sg13g2_decap_8 FILLER_22_1761 ();
 sg13g2_fill_2 FILLER_22_1768 ();
 sg13g2_fill_1 FILLER_22_1770 ();
 sg13g2_decap_8 FILLER_22_1786 ();
 sg13g2_decap_8 FILLER_22_1793 ();
 sg13g2_decap_8 FILLER_22_1800 ();
 sg13g2_decap_8 FILLER_22_1807 ();
 sg13g2_decap_8 FILLER_22_1814 ();
 sg13g2_decap_8 FILLER_22_1821 ();
 sg13g2_decap_8 FILLER_22_1828 ();
 sg13g2_decap_8 FILLER_22_1835 ();
 sg13g2_decap_8 FILLER_22_1842 ();
 sg13g2_decap_8 FILLER_22_1849 ();
 sg13g2_decap_8 FILLER_22_1856 ();
 sg13g2_decap_8 FILLER_22_1863 ();
 sg13g2_decap_8 FILLER_22_1870 ();
 sg13g2_decap_8 FILLER_22_1877 ();
 sg13g2_decap_8 FILLER_22_1884 ();
 sg13g2_decap_8 FILLER_22_1891 ();
 sg13g2_decap_8 FILLER_22_1898 ();
 sg13g2_decap_8 FILLER_22_1905 ();
 sg13g2_decap_8 FILLER_22_1912 ();
 sg13g2_decap_8 FILLER_22_1919 ();
 sg13g2_decap_8 FILLER_22_1926 ();
 sg13g2_decap_8 FILLER_22_1933 ();
 sg13g2_decap_8 FILLER_22_1940 ();
 sg13g2_decap_8 FILLER_22_1947 ();
 sg13g2_decap_8 FILLER_22_1954 ();
 sg13g2_decap_8 FILLER_22_1961 ();
 sg13g2_decap_8 FILLER_22_1968 ();
 sg13g2_decap_8 FILLER_22_1975 ();
 sg13g2_decap_8 FILLER_22_1982 ();
 sg13g2_decap_8 FILLER_22_1989 ();
 sg13g2_decap_8 FILLER_22_1996 ();
 sg13g2_decap_8 FILLER_22_2003 ();
 sg13g2_decap_8 FILLER_22_2010 ();
 sg13g2_decap_8 FILLER_22_2017 ();
 sg13g2_decap_8 FILLER_22_2024 ();
 sg13g2_decap_8 FILLER_22_2031 ();
 sg13g2_decap_8 FILLER_22_2038 ();
 sg13g2_decap_8 FILLER_22_2045 ();
 sg13g2_decap_8 FILLER_22_2052 ();
 sg13g2_decap_8 FILLER_22_2059 ();
 sg13g2_decap_8 FILLER_22_2066 ();
 sg13g2_decap_8 FILLER_22_2073 ();
 sg13g2_decap_8 FILLER_22_2080 ();
 sg13g2_decap_8 FILLER_22_2087 ();
 sg13g2_decap_8 FILLER_22_2094 ();
 sg13g2_decap_8 FILLER_22_2101 ();
 sg13g2_decap_8 FILLER_22_2108 ();
 sg13g2_decap_8 FILLER_22_2115 ();
 sg13g2_decap_8 FILLER_22_2122 ();
 sg13g2_decap_8 FILLER_22_2129 ();
 sg13g2_decap_8 FILLER_22_2136 ();
 sg13g2_decap_8 FILLER_22_2143 ();
 sg13g2_decap_8 FILLER_22_2150 ();
 sg13g2_decap_8 FILLER_22_2157 ();
 sg13g2_decap_8 FILLER_22_2164 ();
 sg13g2_decap_8 FILLER_22_2171 ();
 sg13g2_decap_8 FILLER_22_2178 ();
 sg13g2_decap_8 FILLER_22_2185 ();
 sg13g2_decap_8 FILLER_22_2192 ();
 sg13g2_decap_8 FILLER_22_2199 ();
 sg13g2_decap_8 FILLER_22_2206 ();
 sg13g2_decap_8 FILLER_22_2213 ();
 sg13g2_decap_8 FILLER_22_2220 ();
 sg13g2_decap_8 FILLER_22_2227 ();
 sg13g2_decap_8 FILLER_22_2234 ();
 sg13g2_decap_8 FILLER_22_2241 ();
 sg13g2_decap_8 FILLER_22_2248 ();
 sg13g2_decap_8 FILLER_22_2255 ();
 sg13g2_decap_8 FILLER_22_2262 ();
 sg13g2_decap_8 FILLER_22_2269 ();
 sg13g2_decap_8 FILLER_22_2276 ();
 sg13g2_decap_8 FILLER_22_2283 ();
 sg13g2_decap_8 FILLER_22_2290 ();
 sg13g2_decap_8 FILLER_22_2297 ();
 sg13g2_decap_8 FILLER_22_2304 ();
 sg13g2_decap_8 FILLER_22_2311 ();
 sg13g2_decap_8 FILLER_22_2318 ();
 sg13g2_decap_8 FILLER_22_2325 ();
 sg13g2_decap_8 FILLER_22_2332 ();
 sg13g2_decap_8 FILLER_22_2339 ();
 sg13g2_decap_8 FILLER_22_2346 ();
 sg13g2_decap_8 FILLER_22_2353 ();
 sg13g2_decap_8 FILLER_22_2360 ();
 sg13g2_decap_8 FILLER_22_2367 ();
 sg13g2_decap_8 FILLER_22_2374 ();
 sg13g2_decap_8 FILLER_22_2381 ();
 sg13g2_decap_8 FILLER_22_2388 ();
 sg13g2_decap_8 FILLER_22_2395 ();
 sg13g2_decap_8 FILLER_22_2402 ();
 sg13g2_decap_8 FILLER_22_2409 ();
 sg13g2_decap_8 FILLER_22_2416 ();
 sg13g2_decap_8 FILLER_22_2423 ();
 sg13g2_decap_8 FILLER_22_2430 ();
 sg13g2_decap_8 FILLER_22_2437 ();
 sg13g2_decap_8 FILLER_22_2444 ();
 sg13g2_decap_8 FILLER_22_2451 ();
 sg13g2_decap_8 FILLER_22_2458 ();
 sg13g2_decap_8 FILLER_22_2465 ();
 sg13g2_decap_8 FILLER_22_2472 ();
 sg13g2_decap_8 FILLER_22_2479 ();
 sg13g2_decap_8 FILLER_22_2486 ();
 sg13g2_decap_8 FILLER_22_2493 ();
 sg13g2_decap_8 FILLER_22_2500 ();
 sg13g2_decap_8 FILLER_22_2507 ();
 sg13g2_decap_8 FILLER_22_2514 ();
 sg13g2_decap_8 FILLER_22_2521 ();
 sg13g2_decap_8 FILLER_22_2528 ();
 sg13g2_decap_8 FILLER_22_2535 ();
 sg13g2_decap_8 FILLER_22_2542 ();
 sg13g2_decap_8 FILLER_22_2549 ();
 sg13g2_decap_8 FILLER_22_2556 ();
 sg13g2_decap_8 FILLER_22_2563 ();
 sg13g2_decap_8 FILLER_22_2570 ();
 sg13g2_decap_8 FILLER_22_2577 ();
 sg13g2_decap_8 FILLER_22_2584 ();
 sg13g2_decap_8 FILLER_22_2591 ();
 sg13g2_decap_8 FILLER_22_2598 ();
 sg13g2_decap_8 FILLER_22_2605 ();
 sg13g2_decap_8 FILLER_22_2612 ();
 sg13g2_decap_8 FILLER_22_2619 ();
 sg13g2_decap_8 FILLER_22_2626 ();
 sg13g2_decap_8 FILLER_22_2633 ();
 sg13g2_decap_8 FILLER_22_2640 ();
 sg13g2_decap_8 FILLER_22_2647 ();
 sg13g2_decap_8 FILLER_22_2654 ();
 sg13g2_decap_8 FILLER_22_2661 ();
 sg13g2_fill_2 FILLER_22_2668 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_4 FILLER_23_259 ();
 sg13g2_fill_1 FILLER_23_263 ();
 sg13g2_decap_8 FILLER_23_278 ();
 sg13g2_decap_8 FILLER_23_285 ();
 sg13g2_decap_8 FILLER_23_292 ();
 sg13g2_decap_8 FILLER_23_299 ();
 sg13g2_decap_8 FILLER_23_306 ();
 sg13g2_decap_8 FILLER_23_313 ();
 sg13g2_decap_8 FILLER_23_320 ();
 sg13g2_decap_8 FILLER_23_327 ();
 sg13g2_decap_8 FILLER_23_334 ();
 sg13g2_decap_8 FILLER_23_341 ();
 sg13g2_decap_8 FILLER_23_348 ();
 sg13g2_fill_2 FILLER_23_355 ();
 sg13g2_fill_1 FILLER_23_360 ();
 sg13g2_fill_2 FILLER_23_376 ();
 sg13g2_fill_1 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_394 ();
 sg13g2_decap_8 FILLER_23_401 ();
 sg13g2_decap_8 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_23_415 ();
 sg13g2_decap_8 FILLER_23_422 ();
 sg13g2_decap_8 FILLER_23_429 ();
 sg13g2_fill_1 FILLER_23_436 ();
 sg13g2_decap_8 FILLER_23_440 ();
 sg13g2_decap_4 FILLER_23_447 ();
 sg13g2_fill_2 FILLER_23_451 ();
 sg13g2_decap_8 FILLER_23_477 ();
 sg13g2_decap_8 FILLER_23_484 ();
 sg13g2_decap_8 FILLER_23_491 ();
 sg13g2_decap_8 FILLER_23_498 ();
 sg13g2_decap_8 FILLER_23_505 ();
 sg13g2_decap_8 FILLER_23_512 ();
 sg13g2_decap_8 FILLER_23_519 ();
 sg13g2_decap_8 FILLER_23_526 ();
 sg13g2_decap_8 FILLER_23_533 ();
 sg13g2_fill_2 FILLER_23_540 ();
 sg13g2_decap_8 FILLER_23_557 ();
 sg13g2_fill_2 FILLER_23_564 ();
 sg13g2_fill_1 FILLER_23_566 ();
 sg13g2_decap_8 FILLER_23_579 ();
 sg13g2_decap_4 FILLER_23_586 ();
 sg13g2_decap_4 FILLER_23_593 ();
 sg13g2_decap_8 FILLER_23_600 ();
 sg13g2_decap_4 FILLER_23_612 ();
 sg13g2_fill_2 FILLER_23_616 ();
 sg13g2_decap_4 FILLER_23_627 ();
 sg13g2_fill_2 FILLER_23_631 ();
 sg13g2_decap_8 FILLER_23_637 ();
 sg13g2_fill_2 FILLER_23_644 ();
 sg13g2_fill_1 FILLER_23_646 ();
 sg13g2_fill_1 FILLER_23_651 ();
 sg13g2_fill_1 FILLER_23_657 ();
 sg13g2_decap_8 FILLER_23_662 ();
 sg13g2_decap_8 FILLER_23_669 ();
 sg13g2_decap_8 FILLER_23_676 ();
 sg13g2_fill_1 FILLER_23_683 ();
 sg13g2_decap_8 FILLER_23_695 ();
 sg13g2_decap_8 FILLER_23_702 ();
 sg13g2_decap_8 FILLER_23_709 ();
 sg13g2_decap_8 FILLER_23_716 ();
 sg13g2_fill_2 FILLER_23_723 ();
 sg13g2_decap_8 FILLER_23_728 ();
 sg13g2_decap_4 FILLER_23_735 ();
 sg13g2_fill_1 FILLER_23_739 ();
 sg13g2_decap_8 FILLER_23_743 ();
 sg13g2_decap_8 FILLER_23_750 ();
 sg13g2_decap_8 FILLER_23_757 ();
 sg13g2_decap_8 FILLER_23_764 ();
 sg13g2_decap_8 FILLER_23_771 ();
 sg13g2_decap_8 FILLER_23_778 ();
 sg13g2_decap_8 FILLER_23_785 ();
 sg13g2_decap_8 FILLER_23_792 ();
 sg13g2_decap_8 FILLER_23_799 ();
 sg13g2_fill_2 FILLER_23_806 ();
 sg13g2_fill_1 FILLER_23_808 ();
 sg13g2_fill_2 FILLER_23_817 ();
 sg13g2_fill_1 FILLER_23_819 ();
 sg13g2_decap_8 FILLER_23_824 ();
 sg13g2_decap_4 FILLER_23_831 ();
 sg13g2_fill_1 FILLER_23_835 ();
 sg13g2_decap_8 FILLER_23_856 ();
 sg13g2_decap_8 FILLER_23_863 ();
 sg13g2_decap_8 FILLER_23_870 ();
 sg13g2_decap_8 FILLER_23_877 ();
 sg13g2_decap_8 FILLER_23_884 ();
 sg13g2_fill_1 FILLER_23_891 ();
 sg13g2_fill_2 FILLER_23_923 ();
 sg13g2_decap_8 FILLER_23_928 ();
 sg13g2_decap_8 FILLER_23_941 ();
 sg13g2_decap_8 FILLER_23_948 ();
 sg13g2_decap_8 FILLER_23_955 ();
 sg13g2_decap_8 FILLER_23_962 ();
 sg13g2_decap_8 FILLER_23_969 ();
 sg13g2_decap_4 FILLER_23_976 ();
 sg13g2_decap_8 FILLER_23_985 ();
 sg13g2_decap_4 FILLER_23_992 ();
 sg13g2_decap_8 FILLER_23_1000 ();
 sg13g2_decap_8 FILLER_23_1007 ();
 sg13g2_decap_8 FILLER_23_1014 ();
 sg13g2_decap_8 FILLER_23_1021 ();
 sg13g2_decap_8 FILLER_23_1028 ();
 sg13g2_decap_8 FILLER_23_1035 ();
 sg13g2_fill_2 FILLER_23_1042 ();
 sg13g2_decap_8 FILLER_23_1050 ();
 sg13g2_decap_8 FILLER_23_1057 ();
 sg13g2_decap_8 FILLER_23_1064 ();
 sg13g2_decap_8 FILLER_23_1071 ();
 sg13g2_decap_8 FILLER_23_1078 ();
 sg13g2_decap_4 FILLER_23_1085 ();
 sg13g2_fill_1 FILLER_23_1089 ();
 sg13g2_decap_8 FILLER_23_1100 ();
 sg13g2_decap_8 FILLER_23_1107 ();
 sg13g2_decap_4 FILLER_23_1122 ();
 sg13g2_fill_2 FILLER_23_1126 ();
 sg13g2_decap_4 FILLER_23_1137 ();
 sg13g2_fill_2 FILLER_23_1141 ();
 sg13g2_decap_8 FILLER_23_1158 ();
 sg13g2_decap_8 FILLER_23_1165 ();
 sg13g2_decap_8 FILLER_23_1172 ();
 sg13g2_decap_8 FILLER_23_1179 ();
 sg13g2_decap_4 FILLER_23_1186 ();
 sg13g2_fill_2 FILLER_23_1193 ();
 sg13g2_fill_1 FILLER_23_1195 ();
 sg13g2_decap_8 FILLER_23_1200 ();
 sg13g2_decap_8 FILLER_23_1207 ();
 sg13g2_decap_8 FILLER_23_1214 ();
 sg13g2_decap_4 FILLER_23_1221 ();
 sg13g2_decap_8 FILLER_23_1255 ();
 sg13g2_decap_8 FILLER_23_1262 ();
 sg13g2_decap_8 FILLER_23_1269 ();
 sg13g2_decap_8 FILLER_23_1276 ();
 sg13g2_decap_8 FILLER_23_1283 ();
 sg13g2_decap_8 FILLER_23_1290 ();
 sg13g2_decap_8 FILLER_23_1297 ();
 sg13g2_decap_8 FILLER_23_1304 ();
 sg13g2_decap_8 FILLER_23_1311 ();
 sg13g2_decap_8 FILLER_23_1318 ();
 sg13g2_decap_4 FILLER_23_1325 ();
 sg13g2_decap_8 FILLER_23_1334 ();
 sg13g2_decap_8 FILLER_23_1341 ();
 sg13g2_fill_2 FILLER_23_1352 ();
 sg13g2_decap_4 FILLER_23_1362 ();
 sg13g2_fill_1 FILLER_23_1366 ();
 sg13g2_decap_8 FILLER_23_1388 ();
 sg13g2_fill_2 FILLER_23_1395 ();
 sg13g2_fill_1 FILLER_23_1397 ();
 sg13g2_fill_2 FILLER_23_1403 ();
 sg13g2_fill_1 FILLER_23_1405 ();
 sg13g2_fill_1 FILLER_23_1412 ();
 sg13g2_decap_4 FILLER_23_1423 ();
 sg13g2_fill_1 FILLER_23_1427 ();
 sg13g2_decap_4 FILLER_23_1434 ();
 sg13g2_fill_2 FILLER_23_1438 ();
 sg13g2_decap_8 FILLER_23_1445 ();
 sg13g2_decap_8 FILLER_23_1452 ();
 sg13g2_fill_2 FILLER_23_1459 ();
 sg13g2_fill_1 FILLER_23_1472 ();
 sg13g2_decap_8 FILLER_23_1484 ();
 sg13g2_decap_8 FILLER_23_1491 ();
 sg13g2_decap_4 FILLER_23_1498 ();
 sg13g2_fill_1 FILLER_23_1502 ();
 sg13g2_decap_8 FILLER_23_1516 ();
 sg13g2_decap_4 FILLER_23_1523 ();
 sg13g2_decap_8 FILLER_23_1531 ();
 sg13g2_decap_8 FILLER_23_1538 ();
 sg13g2_fill_2 FILLER_23_1545 ();
 sg13g2_fill_1 FILLER_23_1547 ();
 sg13g2_decap_8 FILLER_23_1554 ();
 sg13g2_decap_8 FILLER_23_1561 ();
 sg13g2_decap_8 FILLER_23_1568 ();
 sg13g2_decap_8 FILLER_23_1575 ();
 sg13g2_decap_8 FILLER_23_1582 ();
 sg13g2_decap_8 FILLER_23_1589 ();
 sg13g2_decap_8 FILLER_23_1596 ();
 sg13g2_decap_8 FILLER_23_1603 ();
 sg13g2_decap_8 FILLER_23_1610 ();
 sg13g2_decap_8 FILLER_23_1617 ();
 sg13g2_fill_1 FILLER_23_1624 ();
 sg13g2_decap_8 FILLER_23_1634 ();
 sg13g2_decap_8 FILLER_23_1641 ();
 sg13g2_decap_8 FILLER_23_1648 ();
 sg13g2_decap_8 FILLER_23_1655 ();
 sg13g2_decap_8 FILLER_23_1662 ();
 sg13g2_decap_8 FILLER_23_1669 ();
 sg13g2_decap_8 FILLER_23_1676 ();
 sg13g2_decap_8 FILLER_23_1683 ();
 sg13g2_decap_4 FILLER_23_1690 ();
 sg13g2_fill_1 FILLER_23_1694 ();
 sg13g2_decap_8 FILLER_23_1700 ();
 sg13g2_decap_8 FILLER_23_1707 ();
 sg13g2_decap_8 FILLER_23_1714 ();
 sg13g2_decap_8 FILLER_23_1721 ();
 sg13g2_decap_8 FILLER_23_1728 ();
 sg13g2_fill_2 FILLER_23_1735 ();
 sg13g2_decap_8 FILLER_23_1752 ();
 sg13g2_decap_8 FILLER_23_1759 ();
 sg13g2_decap_4 FILLER_23_1766 ();
 sg13g2_fill_1 FILLER_23_1770 ();
 sg13g2_decap_8 FILLER_23_1779 ();
 sg13g2_decap_8 FILLER_23_1786 ();
 sg13g2_decap_8 FILLER_23_1793 ();
 sg13g2_decap_8 FILLER_23_1800 ();
 sg13g2_decap_8 FILLER_23_1807 ();
 sg13g2_fill_1 FILLER_23_1814 ();
 sg13g2_fill_1 FILLER_23_1823 ();
 sg13g2_decap_8 FILLER_23_1828 ();
 sg13g2_decap_8 FILLER_23_1835 ();
 sg13g2_fill_2 FILLER_23_1842 ();
 sg13g2_fill_1 FILLER_23_1844 ();
 sg13g2_fill_1 FILLER_23_1850 ();
 sg13g2_decap_4 FILLER_23_1855 ();
 sg13g2_decap_8 FILLER_23_1863 ();
 sg13g2_decap_8 FILLER_23_1870 ();
 sg13g2_decap_8 FILLER_23_1877 ();
 sg13g2_decap_8 FILLER_23_1884 ();
 sg13g2_decap_8 FILLER_23_1891 ();
 sg13g2_fill_2 FILLER_23_1898 ();
 sg13g2_decap_8 FILLER_23_1913 ();
 sg13g2_decap_8 FILLER_23_1920 ();
 sg13g2_decap_8 FILLER_23_1927 ();
 sg13g2_decap_8 FILLER_23_1934 ();
 sg13g2_decap_8 FILLER_23_1941 ();
 sg13g2_decap_8 FILLER_23_1948 ();
 sg13g2_decap_8 FILLER_23_1955 ();
 sg13g2_decap_8 FILLER_23_1962 ();
 sg13g2_decap_8 FILLER_23_1969 ();
 sg13g2_decap_8 FILLER_23_1976 ();
 sg13g2_decap_8 FILLER_23_1983 ();
 sg13g2_decap_8 FILLER_23_1990 ();
 sg13g2_decap_8 FILLER_23_1997 ();
 sg13g2_decap_8 FILLER_23_2004 ();
 sg13g2_decap_8 FILLER_23_2011 ();
 sg13g2_decap_8 FILLER_23_2018 ();
 sg13g2_decap_8 FILLER_23_2025 ();
 sg13g2_decap_8 FILLER_23_2032 ();
 sg13g2_decap_8 FILLER_23_2039 ();
 sg13g2_decap_8 FILLER_23_2046 ();
 sg13g2_decap_8 FILLER_23_2053 ();
 sg13g2_decap_8 FILLER_23_2060 ();
 sg13g2_decap_8 FILLER_23_2067 ();
 sg13g2_decap_8 FILLER_23_2074 ();
 sg13g2_decap_8 FILLER_23_2081 ();
 sg13g2_decap_8 FILLER_23_2088 ();
 sg13g2_decap_8 FILLER_23_2095 ();
 sg13g2_decap_8 FILLER_23_2102 ();
 sg13g2_decap_8 FILLER_23_2109 ();
 sg13g2_decap_8 FILLER_23_2116 ();
 sg13g2_decap_8 FILLER_23_2123 ();
 sg13g2_decap_8 FILLER_23_2130 ();
 sg13g2_decap_8 FILLER_23_2137 ();
 sg13g2_decap_8 FILLER_23_2144 ();
 sg13g2_decap_8 FILLER_23_2151 ();
 sg13g2_decap_8 FILLER_23_2158 ();
 sg13g2_decap_8 FILLER_23_2165 ();
 sg13g2_decap_8 FILLER_23_2172 ();
 sg13g2_decap_8 FILLER_23_2179 ();
 sg13g2_decap_8 FILLER_23_2186 ();
 sg13g2_decap_8 FILLER_23_2193 ();
 sg13g2_decap_8 FILLER_23_2200 ();
 sg13g2_decap_8 FILLER_23_2207 ();
 sg13g2_decap_8 FILLER_23_2214 ();
 sg13g2_decap_8 FILLER_23_2221 ();
 sg13g2_decap_8 FILLER_23_2228 ();
 sg13g2_decap_8 FILLER_23_2235 ();
 sg13g2_decap_8 FILLER_23_2242 ();
 sg13g2_decap_8 FILLER_23_2249 ();
 sg13g2_decap_8 FILLER_23_2256 ();
 sg13g2_decap_8 FILLER_23_2263 ();
 sg13g2_decap_8 FILLER_23_2270 ();
 sg13g2_decap_8 FILLER_23_2277 ();
 sg13g2_decap_8 FILLER_23_2284 ();
 sg13g2_decap_8 FILLER_23_2291 ();
 sg13g2_decap_8 FILLER_23_2298 ();
 sg13g2_decap_8 FILLER_23_2305 ();
 sg13g2_decap_8 FILLER_23_2312 ();
 sg13g2_decap_8 FILLER_23_2319 ();
 sg13g2_decap_8 FILLER_23_2326 ();
 sg13g2_decap_8 FILLER_23_2333 ();
 sg13g2_decap_8 FILLER_23_2340 ();
 sg13g2_decap_8 FILLER_23_2347 ();
 sg13g2_decap_8 FILLER_23_2354 ();
 sg13g2_decap_8 FILLER_23_2361 ();
 sg13g2_decap_8 FILLER_23_2368 ();
 sg13g2_decap_8 FILLER_23_2375 ();
 sg13g2_decap_8 FILLER_23_2382 ();
 sg13g2_decap_8 FILLER_23_2389 ();
 sg13g2_decap_8 FILLER_23_2396 ();
 sg13g2_decap_8 FILLER_23_2403 ();
 sg13g2_decap_8 FILLER_23_2410 ();
 sg13g2_decap_8 FILLER_23_2417 ();
 sg13g2_decap_8 FILLER_23_2424 ();
 sg13g2_decap_8 FILLER_23_2431 ();
 sg13g2_decap_8 FILLER_23_2438 ();
 sg13g2_decap_8 FILLER_23_2445 ();
 sg13g2_decap_8 FILLER_23_2452 ();
 sg13g2_decap_8 FILLER_23_2459 ();
 sg13g2_decap_8 FILLER_23_2466 ();
 sg13g2_decap_8 FILLER_23_2473 ();
 sg13g2_decap_8 FILLER_23_2480 ();
 sg13g2_decap_8 FILLER_23_2487 ();
 sg13g2_decap_8 FILLER_23_2494 ();
 sg13g2_decap_8 FILLER_23_2501 ();
 sg13g2_decap_8 FILLER_23_2508 ();
 sg13g2_decap_8 FILLER_23_2515 ();
 sg13g2_decap_8 FILLER_23_2522 ();
 sg13g2_decap_8 FILLER_23_2529 ();
 sg13g2_decap_8 FILLER_23_2536 ();
 sg13g2_decap_8 FILLER_23_2543 ();
 sg13g2_decap_8 FILLER_23_2550 ();
 sg13g2_decap_8 FILLER_23_2557 ();
 sg13g2_decap_8 FILLER_23_2564 ();
 sg13g2_decap_8 FILLER_23_2571 ();
 sg13g2_decap_8 FILLER_23_2578 ();
 sg13g2_decap_8 FILLER_23_2585 ();
 sg13g2_decap_8 FILLER_23_2592 ();
 sg13g2_decap_8 FILLER_23_2599 ();
 sg13g2_decap_8 FILLER_23_2606 ();
 sg13g2_decap_8 FILLER_23_2613 ();
 sg13g2_decap_8 FILLER_23_2620 ();
 sg13g2_decap_8 FILLER_23_2627 ();
 sg13g2_decap_8 FILLER_23_2634 ();
 sg13g2_decap_8 FILLER_23_2641 ();
 sg13g2_decap_8 FILLER_23_2648 ();
 sg13g2_decap_8 FILLER_23_2655 ();
 sg13g2_decap_8 FILLER_23_2662 ();
 sg13g2_fill_1 FILLER_23_2669 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_193 ();
 sg13g2_decap_8 FILLER_24_200 ();
 sg13g2_decap_8 FILLER_24_207 ();
 sg13g2_decap_8 FILLER_24_214 ();
 sg13g2_decap_8 FILLER_24_221 ();
 sg13g2_decap_8 FILLER_24_228 ();
 sg13g2_decap_8 FILLER_24_235 ();
 sg13g2_decap_4 FILLER_24_247 ();
 sg13g2_fill_1 FILLER_24_251 ();
 sg13g2_decap_8 FILLER_24_256 ();
 sg13g2_decap_4 FILLER_24_263 ();
 sg13g2_fill_1 FILLER_24_267 ();
 sg13g2_decap_8 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_decap_8 FILLER_24_370 ();
 sg13g2_decap_4 FILLER_24_377 ();
 sg13g2_fill_1 FILLER_24_381 ();
 sg13g2_decap_8 FILLER_24_390 ();
 sg13g2_decap_8 FILLER_24_397 ();
 sg13g2_decap_8 FILLER_24_404 ();
 sg13g2_decap_4 FILLER_24_411 ();
 sg13g2_fill_2 FILLER_24_415 ();
 sg13g2_decap_8 FILLER_24_421 ();
 sg13g2_decap_8 FILLER_24_428 ();
 sg13g2_decap_8 FILLER_24_435 ();
 sg13g2_decap_8 FILLER_24_442 ();
 sg13g2_decap_8 FILLER_24_449 ();
 sg13g2_fill_2 FILLER_24_456 ();
 sg13g2_decap_8 FILLER_24_482 ();
 sg13g2_decap_8 FILLER_24_489 ();
 sg13g2_decap_8 FILLER_24_496 ();
 sg13g2_decap_8 FILLER_24_503 ();
 sg13g2_decap_8 FILLER_24_510 ();
 sg13g2_decap_8 FILLER_24_517 ();
 sg13g2_decap_8 FILLER_24_524 ();
 sg13g2_decap_8 FILLER_24_531 ();
 sg13g2_decap_8 FILLER_24_538 ();
 sg13g2_decap_8 FILLER_24_549 ();
 sg13g2_decap_8 FILLER_24_556 ();
 sg13g2_decap_8 FILLER_24_563 ();
 sg13g2_decap_8 FILLER_24_570 ();
 sg13g2_decap_8 FILLER_24_577 ();
 sg13g2_decap_8 FILLER_24_584 ();
 sg13g2_decap_8 FILLER_24_591 ();
 sg13g2_decap_4 FILLER_24_598 ();
 sg13g2_fill_2 FILLER_24_602 ();
 sg13g2_decap_8 FILLER_24_619 ();
 sg13g2_decap_8 FILLER_24_626 ();
 sg13g2_decap_8 FILLER_24_633 ();
 sg13g2_decap_8 FILLER_24_640 ();
 sg13g2_decap_8 FILLER_24_647 ();
 sg13g2_decap_8 FILLER_24_654 ();
 sg13g2_decap_8 FILLER_24_661 ();
 sg13g2_decap_8 FILLER_24_668 ();
 sg13g2_fill_2 FILLER_24_675 ();
 sg13g2_fill_1 FILLER_24_677 ();
 sg13g2_decap_8 FILLER_24_697 ();
 sg13g2_decap_8 FILLER_24_704 ();
 sg13g2_fill_1 FILLER_24_711 ();
 sg13g2_decap_8 FILLER_24_716 ();
 sg13g2_fill_2 FILLER_24_723 ();
 sg13g2_decap_8 FILLER_24_744 ();
 sg13g2_decap_8 FILLER_24_751 ();
 sg13g2_decap_8 FILLER_24_758 ();
 sg13g2_decap_8 FILLER_24_765 ();
 sg13g2_decap_8 FILLER_24_772 ();
 sg13g2_decap_8 FILLER_24_779 ();
 sg13g2_decap_8 FILLER_24_786 ();
 sg13g2_decap_8 FILLER_24_793 ();
 sg13g2_decap_8 FILLER_24_800 ();
 sg13g2_decap_8 FILLER_24_807 ();
 sg13g2_decap_8 FILLER_24_814 ();
 sg13g2_decap_8 FILLER_24_821 ();
 sg13g2_decap_8 FILLER_24_828 ();
 sg13g2_decap_8 FILLER_24_835 ();
 sg13g2_decap_8 FILLER_24_842 ();
 sg13g2_decap_8 FILLER_24_849 ();
 sg13g2_decap_8 FILLER_24_856 ();
 sg13g2_decap_8 FILLER_24_863 ();
 sg13g2_decap_8 FILLER_24_870 ();
 sg13g2_decap_8 FILLER_24_877 ();
 sg13g2_decap_8 FILLER_24_884 ();
 sg13g2_decap_4 FILLER_24_891 ();
 sg13g2_decap_8 FILLER_24_925 ();
 sg13g2_decap_8 FILLER_24_932 ();
 sg13g2_decap_8 FILLER_24_939 ();
 sg13g2_decap_8 FILLER_24_946 ();
 sg13g2_decap_8 FILLER_24_953 ();
 sg13g2_decap_8 FILLER_24_960 ();
 sg13g2_decap_8 FILLER_24_967 ();
 sg13g2_decap_8 FILLER_24_974 ();
 sg13g2_decap_8 FILLER_24_981 ();
 sg13g2_decap_8 FILLER_24_988 ();
 sg13g2_decap_8 FILLER_24_1004 ();
 sg13g2_decap_8 FILLER_24_1011 ();
 sg13g2_decap_8 FILLER_24_1018 ();
 sg13g2_decap_8 FILLER_24_1025 ();
 sg13g2_decap_4 FILLER_24_1032 ();
 sg13g2_fill_2 FILLER_24_1036 ();
 sg13g2_decap_8 FILLER_24_1043 ();
 sg13g2_decap_8 FILLER_24_1050 ();
 sg13g2_decap_4 FILLER_24_1057 ();
 sg13g2_fill_1 FILLER_24_1061 ();
 sg13g2_decap_8 FILLER_24_1067 ();
 sg13g2_decap_8 FILLER_24_1074 ();
 sg13g2_decap_8 FILLER_24_1081 ();
 sg13g2_decap_4 FILLER_24_1088 ();
 sg13g2_fill_1 FILLER_24_1092 ();
 sg13g2_decap_8 FILLER_24_1101 ();
 sg13g2_decap_8 FILLER_24_1108 ();
 sg13g2_decap_8 FILLER_24_1115 ();
 sg13g2_decap_8 FILLER_24_1122 ();
 sg13g2_decap_8 FILLER_24_1129 ();
 sg13g2_fill_2 FILLER_24_1136 ();
 sg13g2_fill_1 FILLER_24_1138 ();
 sg13g2_decap_8 FILLER_24_1152 ();
 sg13g2_decap_8 FILLER_24_1159 ();
 sg13g2_decap_8 FILLER_24_1166 ();
 sg13g2_decap_8 FILLER_24_1173 ();
 sg13g2_decap_8 FILLER_24_1180 ();
 sg13g2_fill_2 FILLER_24_1187 ();
 sg13g2_fill_1 FILLER_24_1189 ();
 sg13g2_decap_8 FILLER_24_1194 ();
 sg13g2_decap_8 FILLER_24_1201 ();
 sg13g2_decap_8 FILLER_24_1208 ();
 sg13g2_decap_8 FILLER_24_1215 ();
 sg13g2_decap_8 FILLER_24_1222 ();
 sg13g2_decap_4 FILLER_24_1229 ();
 sg13g2_fill_1 FILLER_24_1233 ();
 sg13g2_fill_1 FILLER_24_1242 ();
 sg13g2_decap_8 FILLER_24_1247 ();
 sg13g2_decap_8 FILLER_24_1254 ();
 sg13g2_decap_8 FILLER_24_1261 ();
 sg13g2_decap_8 FILLER_24_1268 ();
 sg13g2_fill_2 FILLER_24_1275 ();
 sg13g2_decap_8 FILLER_24_1281 ();
 sg13g2_decap_4 FILLER_24_1288 ();
 sg13g2_decap_8 FILLER_24_1297 ();
 sg13g2_decap_8 FILLER_24_1304 ();
 sg13g2_decap_8 FILLER_24_1311 ();
 sg13g2_decap_4 FILLER_24_1318 ();
 sg13g2_fill_2 FILLER_24_1322 ();
 sg13g2_decap_8 FILLER_24_1330 ();
 sg13g2_decap_8 FILLER_24_1337 ();
 sg13g2_decap_8 FILLER_24_1344 ();
 sg13g2_decap_8 FILLER_24_1351 ();
 sg13g2_fill_1 FILLER_24_1358 ();
 sg13g2_fill_1 FILLER_24_1375 ();
 sg13g2_decap_8 FILLER_24_1380 ();
 sg13g2_decap_8 FILLER_24_1387 ();
 sg13g2_decap_8 FILLER_24_1394 ();
 sg13g2_decap_8 FILLER_24_1401 ();
 sg13g2_decap_8 FILLER_24_1408 ();
 sg13g2_decap_8 FILLER_24_1415 ();
 sg13g2_decap_8 FILLER_24_1422 ();
 sg13g2_decap_8 FILLER_24_1429 ();
 sg13g2_decap_8 FILLER_24_1441 ();
 sg13g2_decap_8 FILLER_24_1448 ();
 sg13g2_decap_8 FILLER_24_1455 ();
 sg13g2_decap_8 FILLER_24_1462 ();
 sg13g2_decap_8 FILLER_24_1469 ();
 sg13g2_decap_8 FILLER_24_1476 ();
 sg13g2_decap_8 FILLER_24_1483 ();
 sg13g2_decap_8 FILLER_24_1490 ();
 sg13g2_decap_8 FILLER_24_1497 ();
 sg13g2_decap_8 FILLER_24_1504 ();
 sg13g2_decap_8 FILLER_24_1511 ();
 sg13g2_decap_8 FILLER_24_1518 ();
 sg13g2_fill_2 FILLER_24_1525 ();
 sg13g2_decap_8 FILLER_24_1531 ();
 sg13g2_decap_8 FILLER_24_1538 ();
 sg13g2_decap_8 FILLER_24_1552 ();
 sg13g2_decap_8 FILLER_24_1559 ();
 sg13g2_decap_8 FILLER_24_1566 ();
 sg13g2_decap_8 FILLER_24_1573 ();
 sg13g2_fill_1 FILLER_24_1580 ();
 sg13g2_decap_8 FILLER_24_1589 ();
 sg13g2_decap_8 FILLER_24_1596 ();
 sg13g2_decap_8 FILLER_24_1603 ();
 sg13g2_decap_8 FILLER_24_1610 ();
 sg13g2_decap_8 FILLER_24_1617 ();
 sg13g2_fill_1 FILLER_24_1624 ();
 sg13g2_decap_8 FILLER_24_1633 ();
 sg13g2_decap_8 FILLER_24_1640 ();
 sg13g2_decap_8 FILLER_24_1647 ();
 sg13g2_decap_8 FILLER_24_1654 ();
 sg13g2_decap_8 FILLER_24_1661 ();
 sg13g2_decap_8 FILLER_24_1668 ();
 sg13g2_decap_8 FILLER_24_1675 ();
 sg13g2_decap_8 FILLER_24_1682 ();
 sg13g2_decap_8 FILLER_24_1689 ();
 sg13g2_decap_8 FILLER_24_1696 ();
 sg13g2_decap_8 FILLER_24_1703 ();
 sg13g2_decap_8 FILLER_24_1710 ();
 sg13g2_decap_8 FILLER_24_1717 ();
 sg13g2_decap_8 FILLER_24_1724 ();
 sg13g2_fill_1 FILLER_24_1731 ();
 sg13g2_decap_8 FILLER_24_1741 ();
 sg13g2_decap_8 FILLER_24_1748 ();
 sg13g2_decap_8 FILLER_24_1755 ();
 sg13g2_decap_8 FILLER_24_1762 ();
 sg13g2_decap_8 FILLER_24_1769 ();
 sg13g2_decap_4 FILLER_24_1776 ();
 sg13g2_fill_2 FILLER_24_1785 ();
 sg13g2_fill_1 FILLER_24_1787 ();
 sg13g2_decap_8 FILLER_24_1792 ();
 sg13g2_decap_8 FILLER_24_1799 ();
 sg13g2_decap_8 FILLER_24_1806 ();
 sg13g2_decap_8 FILLER_24_1813 ();
 sg13g2_decap_8 FILLER_24_1820 ();
 sg13g2_decap_8 FILLER_24_1827 ();
 sg13g2_decap_8 FILLER_24_1834 ();
 sg13g2_decap_8 FILLER_24_1841 ();
 sg13g2_decap_8 FILLER_24_1848 ();
 sg13g2_fill_2 FILLER_24_1855 ();
 sg13g2_decap_8 FILLER_24_1870 ();
 sg13g2_fill_2 FILLER_24_1877 ();
 sg13g2_decap_8 FILLER_24_1884 ();
 sg13g2_decap_8 FILLER_24_1891 ();
 sg13g2_decap_8 FILLER_24_1898 ();
 sg13g2_decap_8 FILLER_24_1905 ();
 sg13g2_decap_8 FILLER_24_1912 ();
 sg13g2_decap_8 FILLER_24_1919 ();
 sg13g2_decap_8 FILLER_24_1926 ();
 sg13g2_decap_8 FILLER_24_1933 ();
 sg13g2_decap_8 FILLER_24_1940 ();
 sg13g2_decap_8 FILLER_24_1947 ();
 sg13g2_decap_8 FILLER_24_1954 ();
 sg13g2_decap_8 FILLER_24_1961 ();
 sg13g2_decap_8 FILLER_24_1968 ();
 sg13g2_decap_8 FILLER_24_1975 ();
 sg13g2_decap_8 FILLER_24_1982 ();
 sg13g2_decap_8 FILLER_24_1989 ();
 sg13g2_decap_8 FILLER_24_1996 ();
 sg13g2_decap_8 FILLER_24_2003 ();
 sg13g2_decap_8 FILLER_24_2010 ();
 sg13g2_decap_8 FILLER_24_2017 ();
 sg13g2_decap_8 FILLER_24_2024 ();
 sg13g2_decap_8 FILLER_24_2031 ();
 sg13g2_decap_8 FILLER_24_2038 ();
 sg13g2_decap_8 FILLER_24_2045 ();
 sg13g2_decap_8 FILLER_24_2052 ();
 sg13g2_decap_8 FILLER_24_2059 ();
 sg13g2_decap_8 FILLER_24_2066 ();
 sg13g2_decap_8 FILLER_24_2073 ();
 sg13g2_decap_8 FILLER_24_2080 ();
 sg13g2_decap_8 FILLER_24_2087 ();
 sg13g2_decap_8 FILLER_24_2094 ();
 sg13g2_decap_8 FILLER_24_2101 ();
 sg13g2_decap_8 FILLER_24_2108 ();
 sg13g2_decap_8 FILLER_24_2115 ();
 sg13g2_decap_8 FILLER_24_2122 ();
 sg13g2_decap_8 FILLER_24_2129 ();
 sg13g2_decap_8 FILLER_24_2136 ();
 sg13g2_decap_8 FILLER_24_2143 ();
 sg13g2_decap_8 FILLER_24_2150 ();
 sg13g2_decap_8 FILLER_24_2157 ();
 sg13g2_decap_8 FILLER_24_2164 ();
 sg13g2_decap_8 FILLER_24_2171 ();
 sg13g2_decap_8 FILLER_24_2178 ();
 sg13g2_decap_8 FILLER_24_2185 ();
 sg13g2_decap_8 FILLER_24_2192 ();
 sg13g2_decap_8 FILLER_24_2199 ();
 sg13g2_decap_8 FILLER_24_2206 ();
 sg13g2_decap_8 FILLER_24_2213 ();
 sg13g2_decap_8 FILLER_24_2220 ();
 sg13g2_decap_8 FILLER_24_2227 ();
 sg13g2_decap_8 FILLER_24_2234 ();
 sg13g2_decap_8 FILLER_24_2241 ();
 sg13g2_decap_8 FILLER_24_2248 ();
 sg13g2_decap_8 FILLER_24_2255 ();
 sg13g2_decap_8 FILLER_24_2262 ();
 sg13g2_decap_8 FILLER_24_2269 ();
 sg13g2_decap_8 FILLER_24_2276 ();
 sg13g2_decap_8 FILLER_24_2283 ();
 sg13g2_decap_8 FILLER_24_2290 ();
 sg13g2_decap_8 FILLER_24_2297 ();
 sg13g2_decap_8 FILLER_24_2304 ();
 sg13g2_decap_8 FILLER_24_2311 ();
 sg13g2_decap_8 FILLER_24_2318 ();
 sg13g2_decap_8 FILLER_24_2325 ();
 sg13g2_decap_8 FILLER_24_2332 ();
 sg13g2_decap_8 FILLER_24_2339 ();
 sg13g2_decap_8 FILLER_24_2346 ();
 sg13g2_decap_8 FILLER_24_2353 ();
 sg13g2_decap_8 FILLER_24_2360 ();
 sg13g2_decap_8 FILLER_24_2367 ();
 sg13g2_decap_8 FILLER_24_2374 ();
 sg13g2_decap_8 FILLER_24_2381 ();
 sg13g2_decap_8 FILLER_24_2388 ();
 sg13g2_decap_8 FILLER_24_2395 ();
 sg13g2_decap_8 FILLER_24_2402 ();
 sg13g2_decap_8 FILLER_24_2409 ();
 sg13g2_decap_8 FILLER_24_2416 ();
 sg13g2_decap_8 FILLER_24_2423 ();
 sg13g2_decap_8 FILLER_24_2430 ();
 sg13g2_decap_8 FILLER_24_2437 ();
 sg13g2_decap_8 FILLER_24_2444 ();
 sg13g2_decap_8 FILLER_24_2451 ();
 sg13g2_decap_8 FILLER_24_2458 ();
 sg13g2_decap_8 FILLER_24_2465 ();
 sg13g2_decap_8 FILLER_24_2472 ();
 sg13g2_decap_8 FILLER_24_2479 ();
 sg13g2_decap_8 FILLER_24_2486 ();
 sg13g2_decap_8 FILLER_24_2493 ();
 sg13g2_decap_8 FILLER_24_2500 ();
 sg13g2_decap_8 FILLER_24_2507 ();
 sg13g2_decap_8 FILLER_24_2514 ();
 sg13g2_decap_8 FILLER_24_2521 ();
 sg13g2_decap_8 FILLER_24_2528 ();
 sg13g2_decap_8 FILLER_24_2535 ();
 sg13g2_decap_8 FILLER_24_2542 ();
 sg13g2_decap_8 FILLER_24_2549 ();
 sg13g2_decap_8 FILLER_24_2556 ();
 sg13g2_decap_8 FILLER_24_2563 ();
 sg13g2_decap_8 FILLER_24_2570 ();
 sg13g2_decap_8 FILLER_24_2577 ();
 sg13g2_decap_8 FILLER_24_2584 ();
 sg13g2_decap_8 FILLER_24_2591 ();
 sg13g2_decap_8 FILLER_24_2598 ();
 sg13g2_decap_8 FILLER_24_2605 ();
 sg13g2_decap_8 FILLER_24_2612 ();
 sg13g2_decap_8 FILLER_24_2619 ();
 sg13g2_decap_8 FILLER_24_2626 ();
 sg13g2_decap_8 FILLER_24_2633 ();
 sg13g2_decap_8 FILLER_24_2640 ();
 sg13g2_decap_8 FILLER_24_2647 ();
 sg13g2_decap_8 FILLER_24_2654 ();
 sg13g2_decap_8 FILLER_24_2661 ();
 sg13g2_fill_2 FILLER_24_2668 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_208 ();
 sg13g2_decap_8 FILLER_25_215 ();
 sg13g2_decap_8 FILLER_25_222 ();
 sg13g2_decap_8 FILLER_25_229 ();
 sg13g2_decap_8 FILLER_25_236 ();
 sg13g2_decap_8 FILLER_25_243 ();
 sg13g2_fill_2 FILLER_25_250 ();
 sg13g2_fill_1 FILLER_25_252 ();
 sg13g2_fill_1 FILLER_25_257 ();
 sg13g2_fill_2 FILLER_25_263 ();
 sg13g2_decap_8 FILLER_25_270 ();
 sg13g2_decap_8 FILLER_25_277 ();
 sg13g2_decap_8 FILLER_25_284 ();
 sg13g2_decap_8 FILLER_25_291 ();
 sg13g2_decap_8 FILLER_25_298 ();
 sg13g2_fill_2 FILLER_25_305 ();
 sg13g2_fill_1 FILLER_25_307 ();
 sg13g2_decap_8 FILLER_25_312 ();
 sg13g2_decap_8 FILLER_25_319 ();
 sg13g2_decap_8 FILLER_25_326 ();
 sg13g2_decap_8 FILLER_25_333 ();
 sg13g2_decap_8 FILLER_25_340 ();
 sg13g2_decap_8 FILLER_25_347 ();
 sg13g2_decap_8 FILLER_25_354 ();
 sg13g2_decap_8 FILLER_25_361 ();
 sg13g2_decap_8 FILLER_25_368 ();
 sg13g2_decap_8 FILLER_25_375 ();
 sg13g2_decap_8 FILLER_25_382 ();
 sg13g2_decap_8 FILLER_25_389 ();
 sg13g2_decap_8 FILLER_25_396 ();
 sg13g2_decap_8 FILLER_25_403 ();
 sg13g2_decap_8 FILLER_25_410 ();
 sg13g2_decap_8 FILLER_25_417 ();
 sg13g2_decap_8 FILLER_25_424 ();
 sg13g2_decap_8 FILLER_25_431 ();
 sg13g2_decap_8 FILLER_25_438 ();
 sg13g2_decap_8 FILLER_25_445 ();
 sg13g2_fill_2 FILLER_25_452 ();
 sg13g2_decap_8 FILLER_25_459 ();
 sg13g2_decap_8 FILLER_25_466 ();
 sg13g2_decap_8 FILLER_25_473 ();
 sg13g2_decap_8 FILLER_25_480 ();
 sg13g2_decap_8 FILLER_25_487 ();
 sg13g2_decap_8 FILLER_25_494 ();
 sg13g2_decap_4 FILLER_25_501 ();
 sg13g2_decap_8 FILLER_25_509 ();
 sg13g2_decap_8 FILLER_25_516 ();
 sg13g2_decap_8 FILLER_25_523 ();
 sg13g2_decap_8 FILLER_25_544 ();
 sg13g2_decap_8 FILLER_25_551 ();
 sg13g2_decap_8 FILLER_25_558 ();
 sg13g2_decap_4 FILLER_25_565 ();
 sg13g2_fill_2 FILLER_25_569 ();
 sg13g2_decap_8 FILLER_25_586 ();
 sg13g2_decap_8 FILLER_25_593 ();
 sg13g2_decap_8 FILLER_25_600 ();
 sg13g2_fill_2 FILLER_25_607 ();
 sg13g2_fill_1 FILLER_25_615 ();
 sg13g2_decap_8 FILLER_25_619 ();
 sg13g2_decap_8 FILLER_25_626 ();
 sg13g2_decap_8 FILLER_25_633 ();
 sg13g2_decap_8 FILLER_25_640 ();
 sg13g2_decap_8 FILLER_25_647 ();
 sg13g2_decap_8 FILLER_25_654 ();
 sg13g2_decap_8 FILLER_25_661 ();
 sg13g2_decap_8 FILLER_25_668 ();
 sg13g2_decap_8 FILLER_25_675 ();
 sg13g2_decap_8 FILLER_25_682 ();
 sg13g2_decap_8 FILLER_25_689 ();
 sg13g2_decap_8 FILLER_25_696 ();
 sg13g2_decap_8 FILLER_25_703 ();
 sg13g2_decap_8 FILLER_25_710 ();
 sg13g2_decap_8 FILLER_25_717 ();
 sg13g2_decap_8 FILLER_25_724 ();
 sg13g2_fill_1 FILLER_25_731 ();
 sg13g2_decap_8 FILLER_25_741 ();
 sg13g2_decap_8 FILLER_25_748 ();
 sg13g2_decap_4 FILLER_25_755 ();
 sg13g2_fill_1 FILLER_25_759 ();
 sg13g2_decap_8 FILLER_25_780 ();
 sg13g2_decap_8 FILLER_25_787 ();
 sg13g2_decap_8 FILLER_25_794 ();
 sg13g2_decap_8 FILLER_25_801 ();
 sg13g2_decap_8 FILLER_25_808 ();
 sg13g2_decap_8 FILLER_25_830 ();
 sg13g2_decap_8 FILLER_25_837 ();
 sg13g2_decap_4 FILLER_25_844 ();
 sg13g2_fill_2 FILLER_25_848 ();
 sg13g2_decap_8 FILLER_25_859 ();
 sg13g2_decap_4 FILLER_25_866 ();
 sg13g2_decap_8 FILLER_25_875 ();
 sg13g2_decap_8 FILLER_25_882 ();
 sg13g2_decap_8 FILLER_25_889 ();
 sg13g2_decap_8 FILLER_25_896 ();
 sg13g2_decap_8 FILLER_25_903 ();
 sg13g2_decap_8 FILLER_25_910 ();
 sg13g2_decap_8 FILLER_25_917 ();
 sg13g2_decap_8 FILLER_25_924 ();
 sg13g2_decap_8 FILLER_25_931 ();
 sg13g2_decap_8 FILLER_25_938 ();
 sg13g2_decap_8 FILLER_25_945 ();
 sg13g2_decap_8 FILLER_25_952 ();
 sg13g2_decap_8 FILLER_25_959 ();
 sg13g2_decap_8 FILLER_25_966 ();
 sg13g2_decap_8 FILLER_25_973 ();
 sg13g2_decap_8 FILLER_25_980 ();
 sg13g2_decap_4 FILLER_25_987 ();
 sg13g2_fill_1 FILLER_25_991 ();
 sg13g2_decap_8 FILLER_25_1001 ();
 sg13g2_decap_8 FILLER_25_1008 ();
 sg13g2_decap_8 FILLER_25_1015 ();
 sg13g2_decap_8 FILLER_25_1022 ();
 sg13g2_decap_4 FILLER_25_1029 ();
 sg13g2_fill_1 FILLER_25_1033 ();
 sg13g2_decap_8 FILLER_25_1037 ();
 sg13g2_decap_8 FILLER_25_1044 ();
 sg13g2_decap_8 FILLER_25_1051 ();
 sg13g2_decap_8 FILLER_25_1058 ();
 sg13g2_fill_1 FILLER_25_1065 ();
 sg13g2_decap_8 FILLER_25_1071 ();
 sg13g2_decap_8 FILLER_25_1078 ();
 sg13g2_decap_8 FILLER_25_1085 ();
 sg13g2_decap_8 FILLER_25_1092 ();
 sg13g2_decap_8 FILLER_25_1099 ();
 sg13g2_decap_8 FILLER_25_1106 ();
 sg13g2_decap_8 FILLER_25_1113 ();
 sg13g2_decap_8 FILLER_25_1120 ();
 sg13g2_decap_8 FILLER_25_1127 ();
 sg13g2_decap_8 FILLER_25_1134 ();
 sg13g2_decap_4 FILLER_25_1141 ();
 sg13g2_fill_1 FILLER_25_1145 ();
 sg13g2_decap_8 FILLER_25_1158 ();
 sg13g2_decap_8 FILLER_25_1165 ();
 sg13g2_decap_8 FILLER_25_1172 ();
 sg13g2_decap_8 FILLER_25_1179 ();
 sg13g2_decap_4 FILLER_25_1186 ();
 sg13g2_decap_8 FILLER_25_1198 ();
 sg13g2_decap_8 FILLER_25_1205 ();
 sg13g2_decap_8 FILLER_25_1212 ();
 sg13g2_decap_4 FILLER_25_1219 ();
 sg13g2_fill_2 FILLER_25_1223 ();
 sg13g2_decap_8 FILLER_25_1233 ();
 sg13g2_decap_8 FILLER_25_1240 ();
 sg13g2_decap_8 FILLER_25_1247 ();
 sg13g2_decap_8 FILLER_25_1254 ();
 sg13g2_decap_8 FILLER_25_1261 ();
 sg13g2_decap_4 FILLER_25_1268 ();
 sg13g2_fill_1 FILLER_25_1272 ();
 sg13g2_decap_4 FILLER_25_1281 ();
 sg13g2_decap_8 FILLER_25_1295 ();
 sg13g2_decap_8 FILLER_25_1302 ();
 sg13g2_decap_8 FILLER_25_1309 ();
 sg13g2_decap_8 FILLER_25_1316 ();
 sg13g2_decap_8 FILLER_25_1323 ();
 sg13g2_decap_8 FILLER_25_1330 ();
 sg13g2_fill_2 FILLER_25_1337 ();
 sg13g2_fill_1 FILLER_25_1339 ();
 sg13g2_decap_8 FILLER_25_1344 ();
 sg13g2_decap_8 FILLER_25_1351 ();
 sg13g2_decap_8 FILLER_25_1358 ();
 sg13g2_decap_8 FILLER_25_1365 ();
 sg13g2_decap_8 FILLER_25_1372 ();
 sg13g2_decap_8 FILLER_25_1379 ();
 sg13g2_decap_8 FILLER_25_1386 ();
 sg13g2_decap_8 FILLER_25_1393 ();
 sg13g2_decap_8 FILLER_25_1400 ();
 sg13g2_decap_8 FILLER_25_1407 ();
 sg13g2_decap_8 FILLER_25_1414 ();
 sg13g2_decap_8 FILLER_25_1421 ();
 sg13g2_decap_8 FILLER_25_1428 ();
 sg13g2_fill_2 FILLER_25_1435 ();
 sg13g2_fill_1 FILLER_25_1437 ();
 sg13g2_decap_8 FILLER_25_1458 ();
 sg13g2_decap_8 FILLER_25_1465 ();
 sg13g2_decap_8 FILLER_25_1472 ();
 sg13g2_decap_8 FILLER_25_1479 ();
 sg13g2_decap_8 FILLER_25_1486 ();
 sg13g2_decap_8 FILLER_25_1493 ();
 sg13g2_decap_8 FILLER_25_1500 ();
 sg13g2_decap_8 FILLER_25_1507 ();
 sg13g2_decap_8 FILLER_25_1514 ();
 sg13g2_decap_8 FILLER_25_1521 ();
 sg13g2_decap_4 FILLER_25_1528 ();
 sg13g2_decap_8 FILLER_25_1537 ();
 sg13g2_decap_4 FILLER_25_1544 ();
 sg13g2_fill_1 FILLER_25_1548 ();
 sg13g2_decap_4 FILLER_25_1554 ();
 sg13g2_fill_2 FILLER_25_1563 ();
 sg13g2_fill_1 FILLER_25_1565 ();
 sg13g2_fill_2 FILLER_25_1570 ();
 sg13g2_fill_2 FILLER_25_1577 ();
 sg13g2_fill_1 FILLER_25_1579 ();
 sg13g2_fill_1 FILLER_25_1584 ();
 sg13g2_decap_8 FILLER_25_1590 ();
 sg13g2_decap_8 FILLER_25_1597 ();
 sg13g2_decap_8 FILLER_25_1604 ();
 sg13g2_decap_8 FILLER_25_1611 ();
 sg13g2_decap_4 FILLER_25_1618 ();
 sg13g2_fill_1 FILLER_25_1622 ();
 sg13g2_decap_4 FILLER_25_1626 ();
 sg13g2_fill_1 FILLER_25_1630 ();
 sg13g2_decap_8 FILLER_25_1635 ();
 sg13g2_decap_8 FILLER_25_1642 ();
 sg13g2_decap_4 FILLER_25_1649 ();
 sg13g2_fill_2 FILLER_25_1653 ();
 sg13g2_fill_2 FILLER_25_1659 ();
 sg13g2_decap_8 FILLER_25_1676 ();
 sg13g2_decap_8 FILLER_25_1683 ();
 sg13g2_decap_4 FILLER_25_1690 ();
 sg13g2_fill_1 FILLER_25_1694 ();
 sg13g2_decap_8 FILLER_25_1701 ();
 sg13g2_decap_8 FILLER_25_1708 ();
 sg13g2_decap_8 FILLER_25_1715 ();
 sg13g2_decap_8 FILLER_25_1722 ();
 sg13g2_fill_2 FILLER_25_1734 ();
 sg13g2_fill_1 FILLER_25_1736 ();
 sg13g2_decap_8 FILLER_25_1740 ();
 sg13g2_decap_8 FILLER_25_1747 ();
 sg13g2_decap_8 FILLER_25_1754 ();
 sg13g2_decap_8 FILLER_25_1761 ();
 sg13g2_decap_8 FILLER_25_1768 ();
 sg13g2_decap_8 FILLER_25_1775 ();
 sg13g2_decap_8 FILLER_25_1782 ();
 sg13g2_decap_8 FILLER_25_1789 ();
 sg13g2_decap_8 FILLER_25_1796 ();
 sg13g2_decap_8 FILLER_25_1803 ();
 sg13g2_decap_8 FILLER_25_1810 ();
 sg13g2_decap_4 FILLER_25_1817 ();
 sg13g2_decap_8 FILLER_25_1826 ();
 sg13g2_decap_8 FILLER_25_1833 ();
 sg13g2_decap_8 FILLER_25_1840 ();
 sg13g2_decap_8 FILLER_25_1847 ();
 sg13g2_decap_8 FILLER_25_1854 ();
 sg13g2_decap_8 FILLER_25_1861 ();
 sg13g2_decap_8 FILLER_25_1868 ();
 sg13g2_decap_8 FILLER_25_1875 ();
 sg13g2_decap_8 FILLER_25_1882 ();
 sg13g2_fill_2 FILLER_25_1889 ();
 sg13g2_fill_1 FILLER_25_1891 ();
 sg13g2_decap_8 FILLER_25_1907 ();
 sg13g2_decap_8 FILLER_25_1914 ();
 sg13g2_decap_8 FILLER_25_1921 ();
 sg13g2_decap_8 FILLER_25_1928 ();
 sg13g2_decap_8 FILLER_25_1935 ();
 sg13g2_decap_8 FILLER_25_1942 ();
 sg13g2_decap_8 FILLER_25_1949 ();
 sg13g2_decap_8 FILLER_25_1956 ();
 sg13g2_decap_8 FILLER_25_1963 ();
 sg13g2_decap_8 FILLER_25_1970 ();
 sg13g2_decap_8 FILLER_25_1977 ();
 sg13g2_decap_8 FILLER_25_1984 ();
 sg13g2_decap_8 FILLER_25_1991 ();
 sg13g2_decap_8 FILLER_25_1998 ();
 sg13g2_decap_8 FILLER_25_2005 ();
 sg13g2_decap_8 FILLER_25_2012 ();
 sg13g2_decap_8 FILLER_25_2019 ();
 sg13g2_decap_8 FILLER_25_2026 ();
 sg13g2_decap_8 FILLER_25_2033 ();
 sg13g2_decap_8 FILLER_25_2040 ();
 sg13g2_decap_8 FILLER_25_2047 ();
 sg13g2_decap_8 FILLER_25_2054 ();
 sg13g2_decap_8 FILLER_25_2061 ();
 sg13g2_decap_8 FILLER_25_2068 ();
 sg13g2_decap_8 FILLER_25_2075 ();
 sg13g2_decap_8 FILLER_25_2082 ();
 sg13g2_decap_8 FILLER_25_2089 ();
 sg13g2_decap_8 FILLER_25_2096 ();
 sg13g2_decap_8 FILLER_25_2103 ();
 sg13g2_decap_8 FILLER_25_2110 ();
 sg13g2_decap_8 FILLER_25_2117 ();
 sg13g2_decap_8 FILLER_25_2124 ();
 sg13g2_decap_8 FILLER_25_2131 ();
 sg13g2_decap_8 FILLER_25_2138 ();
 sg13g2_decap_8 FILLER_25_2145 ();
 sg13g2_decap_8 FILLER_25_2152 ();
 sg13g2_decap_8 FILLER_25_2159 ();
 sg13g2_decap_8 FILLER_25_2166 ();
 sg13g2_decap_8 FILLER_25_2173 ();
 sg13g2_decap_8 FILLER_25_2180 ();
 sg13g2_decap_8 FILLER_25_2187 ();
 sg13g2_decap_8 FILLER_25_2194 ();
 sg13g2_decap_8 FILLER_25_2201 ();
 sg13g2_decap_8 FILLER_25_2208 ();
 sg13g2_decap_8 FILLER_25_2215 ();
 sg13g2_decap_8 FILLER_25_2222 ();
 sg13g2_decap_8 FILLER_25_2229 ();
 sg13g2_decap_8 FILLER_25_2236 ();
 sg13g2_decap_8 FILLER_25_2243 ();
 sg13g2_decap_8 FILLER_25_2250 ();
 sg13g2_decap_8 FILLER_25_2257 ();
 sg13g2_decap_8 FILLER_25_2264 ();
 sg13g2_decap_8 FILLER_25_2271 ();
 sg13g2_decap_8 FILLER_25_2278 ();
 sg13g2_decap_8 FILLER_25_2285 ();
 sg13g2_decap_8 FILLER_25_2292 ();
 sg13g2_decap_8 FILLER_25_2299 ();
 sg13g2_decap_8 FILLER_25_2306 ();
 sg13g2_decap_8 FILLER_25_2313 ();
 sg13g2_decap_8 FILLER_25_2320 ();
 sg13g2_decap_8 FILLER_25_2327 ();
 sg13g2_decap_8 FILLER_25_2334 ();
 sg13g2_decap_8 FILLER_25_2341 ();
 sg13g2_decap_8 FILLER_25_2348 ();
 sg13g2_decap_8 FILLER_25_2355 ();
 sg13g2_decap_8 FILLER_25_2362 ();
 sg13g2_decap_8 FILLER_25_2369 ();
 sg13g2_decap_8 FILLER_25_2376 ();
 sg13g2_decap_8 FILLER_25_2383 ();
 sg13g2_decap_8 FILLER_25_2390 ();
 sg13g2_decap_8 FILLER_25_2397 ();
 sg13g2_decap_8 FILLER_25_2404 ();
 sg13g2_decap_8 FILLER_25_2411 ();
 sg13g2_decap_8 FILLER_25_2418 ();
 sg13g2_decap_8 FILLER_25_2425 ();
 sg13g2_decap_8 FILLER_25_2432 ();
 sg13g2_decap_8 FILLER_25_2439 ();
 sg13g2_decap_8 FILLER_25_2446 ();
 sg13g2_decap_8 FILLER_25_2453 ();
 sg13g2_decap_8 FILLER_25_2460 ();
 sg13g2_decap_8 FILLER_25_2467 ();
 sg13g2_decap_8 FILLER_25_2474 ();
 sg13g2_decap_8 FILLER_25_2481 ();
 sg13g2_decap_8 FILLER_25_2488 ();
 sg13g2_decap_8 FILLER_25_2495 ();
 sg13g2_decap_8 FILLER_25_2502 ();
 sg13g2_decap_8 FILLER_25_2509 ();
 sg13g2_decap_8 FILLER_25_2516 ();
 sg13g2_decap_8 FILLER_25_2523 ();
 sg13g2_decap_8 FILLER_25_2530 ();
 sg13g2_decap_8 FILLER_25_2537 ();
 sg13g2_decap_8 FILLER_25_2544 ();
 sg13g2_decap_8 FILLER_25_2551 ();
 sg13g2_decap_8 FILLER_25_2558 ();
 sg13g2_decap_8 FILLER_25_2565 ();
 sg13g2_decap_8 FILLER_25_2572 ();
 sg13g2_decap_8 FILLER_25_2579 ();
 sg13g2_decap_8 FILLER_25_2586 ();
 sg13g2_decap_8 FILLER_25_2593 ();
 sg13g2_decap_8 FILLER_25_2600 ();
 sg13g2_decap_8 FILLER_25_2607 ();
 sg13g2_decap_8 FILLER_25_2614 ();
 sg13g2_decap_8 FILLER_25_2621 ();
 sg13g2_decap_8 FILLER_25_2628 ();
 sg13g2_decap_8 FILLER_25_2635 ();
 sg13g2_decap_8 FILLER_25_2642 ();
 sg13g2_decap_8 FILLER_25_2649 ();
 sg13g2_decap_8 FILLER_25_2656 ();
 sg13g2_decap_8 FILLER_25_2663 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_fill_2 FILLER_26_49 ();
 sg13g2_fill_1 FILLER_26_51 ();
 sg13g2_decap_8 FILLER_26_67 ();
 sg13g2_decap_8 FILLER_26_74 ();
 sg13g2_decap_8 FILLER_26_81 ();
 sg13g2_decap_8 FILLER_26_88 ();
 sg13g2_decap_8 FILLER_26_95 ();
 sg13g2_decap_4 FILLER_26_102 ();
 sg13g2_decap_8 FILLER_26_132 ();
 sg13g2_decap_8 FILLER_26_139 ();
 sg13g2_decap_8 FILLER_26_146 ();
 sg13g2_fill_2 FILLER_26_153 ();
 sg13g2_fill_1 FILLER_26_155 ();
 sg13g2_decap_8 FILLER_26_160 ();
 sg13g2_decap_8 FILLER_26_167 ();
 sg13g2_decap_8 FILLER_26_174 ();
 sg13g2_decap_8 FILLER_26_181 ();
 sg13g2_decap_8 FILLER_26_188 ();
 sg13g2_decap_8 FILLER_26_195 ();
 sg13g2_decap_8 FILLER_26_202 ();
 sg13g2_decap_8 FILLER_26_209 ();
 sg13g2_decap_8 FILLER_26_216 ();
 sg13g2_decap_8 FILLER_26_223 ();
 sg13g2_decap_8 FILLER_26_230 ();
 sg13g2_decap_8 FILLER_26_237 ();
 sg13g2_decap_8 FILLER_26_244 ();
 sg13g2_decap_8 FILLER_26_251 ();
 sg13g2_decap_8 FILLER_26_258 ();
 sg13g2_decap_8 FILLER_26_265 ();
 sg13g2_fill_2 FILLER_26_272 ();
 sg13g2_decap_8 FILLER_26_278 ();
 sg13g2_decap_8 FILLER_26_285 ();
 sg13g2_decap_8 FILLER_26_292 ();
 sg13g2_decap_8 FILLER_26_299 ();
 sg13g2_decap_4 FILLER_26_306 ();
 sg13g2_decap_8 FILLER_26_336 ();
 sg13g2_decap_8 FILLER_26_343 ();
 sg13g2_decap_8 FILLER_26_350 ();
 sg13g2_decap_8 FILLER_26_357 ();
 sg13g2_decap_8 FILLER_26_364 ();
 sg13g2_decap_8 FILLER_26_371 ();
 sg13g2_decap_8 FILLER_26_378 ();
 sg13g2_decap_8 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_4 FILLER_26_399 ();
 sg13g2_fill_1 FILLER_26_403 ();
 sg13g2_decap_8 FILLER_26_412 ();
 sg13g2_decap_8 FILLER_26_419 ();
 sg13g2_decap_8 FILLER_26_426 ();
 sg13g2_decap_8 FILLER_26_433 ();
 sg13g2_decap_8 FILLER_26_440 ();
 sg13g2_decap_8 FILLER_26_447 ();
 sg13g2_decap_8 FILLER_26_454 ();
 sg13g2_decap_8 FILLER_26_461 ();
 sg13g2_decap_8 FILLER_26_468 ();
 sg13g2_decap_8 FILLER_26_475 ();
 sg13g2_decap_8 FILLER_26_482 ();
 sg13g2_decap_8 FILLER_26_489 ();
 sg13g2_decap_8 FILLER_26_496 ();
 sg13g2_decap_8 FILLER_26_503 ();
 sg13g2_decap_8 FILLER_26_510 ();
 sg13g2_decap_8 FILLER_26_517 ();
 sg13g2_decap_8 FILLER_26_524 ();
 sg13g2_decap_8 FILLER_26_531 ();
 sg13g2_decap_8 FILLER_26_538 ();
 sg13g2_decap_8 FILLER_26_545 ();
 sg13g2_decap_8 FILLER_26_552 ();
 sg13g2_decap_8 FILLER_26_559 ();
 sg13g2_decap_8 FILLER_26_566 ();
 sg13g2_fill_1 FILLER_26_573 ();
 sg13g2_decap_8 FILLER_26_579 ();
 sg13g2_decap_8 FILLER_26_586 ();
 sg13g2_decap_8 FILLER_26_593 ();
 sg13g2_decap_8 FILLER_26_600 ();
 sg13g2_fill_2 FILLER_26_607 ();
 sg13g2_fill_2 FILLER_26_614 ();
 sg13g2_decap_8 FILLER_26_628 ();
 sg13g2_decap_8 FILLER_26_635 ();
 sg13g2_decap_8 FILLER_26_642 ();
 sg13g2_decap_8 FILLER_26_654 ();
 sg13g2_decap_8 FILLER_26_661 ();
 sg13g2_decap_8 FILLER_26_668 ();
 sg13g2_decap_8 FILLER_26_675 ();
 sg13g2_decap_8 FILLER_26_682 ();
 sg13g2_decap_8 FILLER_26_689 ();
 sg13g2_decap_8 FILLER_26_696 ();
 sg13g2_decap_8 FILLER_26_703 ();
 sg13g2_decap_8 FILLER_26_710 ();
 sg13g2_fill_2 FILLER_26_717 ();
 sg13g2_fill_1 FILLER_26_731 ();
 sg13g2_decap_4 FILLER_26_738 ();
 sg13g2_fill_2 FILLER_26_742 ();
 sg13g2_decap_8 FILLER_26_748 ();
 sg13g2_decap_8 FILLER_26_755 ();
 sg13g2_decap_8 FILLER_26_762 ();
 sg13g2_decap_4 FILLER_26_774 ();
 sg13g2_fill_2 FILLER_26_778 ();
 sg13g2_fill_2 FILLER_26_783 ();
 sg13g2_fill_1 FILLER_26_785 ();
 sg13g2_decap_8 FILLER_26_789 ();
 sg13g2_decap_8 FILLER_26_796 ();
 sg13g2_decap_8 FILLER_26_803 ();
 sg13g2_decap_8 FILLER_26_823 ();
 sg13g2_decap_8 FILLER_26_830 ();
 sg13g2_decap_8 FILLER_26_837 ();
 sg13g2_decap_8 FILLER_26_844 ();
 sg13g2_decap_8 FILLER_26_851 ();
 sg13g2_decap_8 FILLER_26_858 ();
 sg13g2_decap_8 FILLER_26_865 ();
 sg13g2_decap_8 FILLER_26_872 ();
 sg13g2_decap_8 FILLER_26_879 ();
 sg13g2_fill_1 FILLER_26_886 ();
 sg13g2_decap_8 FILLER_26_892 ();
 sg13g2_decap_8 FILLER_26_899 ();
 sg13g2_decap_8 FILLER_26_906 ();
 sg13g2_decap_8 FILLER_26_913 ();
 sg13g2_decap_8 FILLER_26_920 ();
 sg13g2_decap_8 FILLER_26_927 ();
 sg13g2_decap_8 FILLER_26_934 ();
 sg13g2_decap_8 FILLER_26_941 ();
 sg13g2_decap_8 FILLER_26_948 ();
 sg13g2_decap_8 FILLER_26_955 ();
 sg13g2_fill_2 FILLER_26_962 ();
 sg13g2_decap_8 FILLER_26_973 ();
 sg13g2_decap_8 FILLER_26_980 ();
 sg13g2_decap_8 FILLER_26_987 ();
 sg13g2_fill_1 FILLER_26_994 ();
 sg13g2_decap_8 FILLER_26_998 ();
 sg13g2_decap_8 FILLER_26_1005 ();
 sg13g2_decap_8 FILLER_26_1012 ();
 sg13g2_decap_8 FILLER_26_1019 ();
 sg13g2_decap_8 FILLER_26_1026 ();
 sg13g2_fill_1 FILLER_26_1033 ();
 sg13g2_decap_8 FILLER_26_1039 ();
 sg13g2_decap_8 FILLER_26_1046 ();
 sg13g2_decap_8 FILLER_26_1053 ();
 sg13g2_fill_1 FILLER_26_1060 ();
 sg13g2_decap_8 FILLER_26_1065 ();
 sg13g2_decap_8 FILLER_26_1072 ();
 sg13g2_decap_8 FILLER_26_1079 ();
 sg13g2_decap_8 FILLER_26_1086 ();
 sg13g2_decap_8 FILLER_26_1093 ();
 sg13g2_decap_8 FILLER_26_1100 ();
 sg13g2_decap_8 FILLER_26_1107 ();
 sg13g2_decap_8 FILLER_26_1114 ();
 sg13g2_decap_8 FILLER_26_1121 ();
 sg13g2_decap_4 FILLER_26_1128 ();
 sg13g2_decap_8 FILLER_26_1137 ();
 sg13g2_decap_8 FILLER_26_1144 ();
 sg13g2_decap_8 FILLER_26_1151 ();
 sg13g2_decap_8 FILLER_26_1158 ();
 sg13g2_decap_8 FILLER_26_1165 ();
 sg13g2_decap_8 FILLER_26_1172 ();
 sg13g2_decap_8 FILLER_26_1179 ();
 sg13g2_decap_4 FILLER_26_1186 ();
 sg13g2_fill_2 FILLER_26_1190 ();
 sg13g2_decap_8 FILLER_26_1196 ();
 sg13g2_decap_8 FILLER_26_1203 ();
 sg13g2_decap_8 FILLER_26_1210 ();
 sg13g2_decap_8 FILLER_26_1217 ();
 sg13g2_decap_8 FILLER_26_1224 ();
 sg13g2_decap_8 FILLER_26_1231 ();
 sg13g2_decap_8 FILLER_26_1238 ();
 sg13g2_decap_8 FILLER_26_1245 ();
 sg13g2_decap_8 FILLER_26_1252 ();
 sg13g2_decap_8 FILLER_26_1259 ();
 sg13g2_decap_8 FILLER_26_1266 ();
 sg13g2_decap_8 FILLER_26_1273 ();
 sg13g2_decap_8 FILLER_26_1280 ();
 sg13g2_decap_8 FILLER_26_1287 ();
 sg13g2_decap_8 FILLER_26_1294 ();
 sg13g2_decap_8 FILLER_26_1301 ();
 sg13g2_fill_2 FILLER_26_1308 ();
 sg13g2_decap_8 FILLER_26_1313 ();
 sg13g2_decap_8 FILLER_26_1320 ();
 sg13g2_decap_8 FILLER_26_1327 ();
 sg13g2_decap_8 FILLER_26_1338 ();
 sg13g2_decap_8 FILLER_26_1345 ();
 sg13g2_decap_8 FILLER_26_1352 ();
 sg13g2_decap_4 FILLER_26_1359 ();
 sg13g2_decap_8 FILLER_26_1366 ();
 sg13g2_decap_4 FILLER_26_1373 ();
 sg13g2_fill_1 FILLER_26_1377 ();
 sg13g2_decap_8 FILLER_26_1393 ();
 sg13g2_decap_8 FILLER_26_1400 ();
 sg13g2_decap_4 FILLER_26_1407 ();
 sg13g2_fill_1 FILLER_26_1411 ();
 sg13g2_decap_8 FILLER_26_1427 ();
 sg13g2_decap_4 FILLER_26_1434 ();
 sg13g2_decap_8 FILLER_26_1443 ();
 sg13g2_decap_8 FILLER_26_1450 ();
 sg13g2_decap_8 FILLER_26_1457 ();
 sg13g2_decap_8 FILLER_26_1464 ();
 sg13g2_decap_8 FILLER_26_1471 ();
 sg13g2_decap_8 FILLER_26_1478 ();
 sg13g2_decap_8 FILLER_26_1485 ();
 sg13g2_fill_1 FILLER_26_1492 ();
 sg13g2_decap_8 FILLER_26_1499 ();
 sg13g2_decap_8 FILLER_26_1506 ();
 sg13g2_decap_8 FILLER_26_1513 ();
 sg13g2_decap_8 FILLER_26_1520 ();
 sg13g2_decap_8 FILLER_26_1527 ();
 sg13g2_decap_8 FILLER_26_1534 ();
 sg13g2_decap_8 FILLER_26_1541 ();
 sg13g2_decap_8 FILLER_26_1548 ();
 sg13g2_decap_8 FILLER_26_1555 ();
 sg13g2_decap_8 FILLER_26_1562 ();
 sg13g2_decap_8 FILLER_26_1569 ();
 sg13g2_decap_8 FILLER_26_1576 ();
 sg13g2_decap_8 FILLER_26_1583 ();
 sg13g2_decap_8 FILLER_26_1590 ();
 sg13g2_decap_8 FILLER_26_1597 ();
 sg13g2_decap_8 FILLER_26_1604 ();
 sg13g2_decap_8 FILLER_26_1611 ();
 sg13g2_decap_8 FILLER_26_1618 ();
 sg13g2_decap_8 FILLER_26_1625 ();
 sg13g2_decap_8 FILLER_26_1632 ();
 sg13g2_decap_8 FILLER_26_1639 ();
 sg13g2_decap_8 FILLER_26_1646 ();
 sg13g2_decap_8 FILLER_26_1653 ();
 sg13g2_fill_1 FILLER_26_1660 ();
 sg13g2_decap_4 FILLER_26_1666 ();
 sg13g2_fill_1 FILLER_26_1670 ();
 sg13g2_decap_8 FILLER_26_1680 ();
 sg13g2_decap_8 FILLER_26_1687 ();
 sg13g2_fill_1 FILLER_26_1694 ();
 sg13g2_decap_4 FILLER_26_1699 ();
 sg13g2_decap_8 FILLER_26_1707 ();
 sg13g2_decap_8 FILLER_26_1714 ();
 sg13g2_decap_8 FILLER_26_1721 ();
 sg13g2_decap_8 FILLER_26_1728 ();
 sg13g2_decap_4 FILLER_26_1735 ();
 sg13g2_decap_8 FILLER_26_1748 ();
 sg13g2_decap_8 FILLER_26_1755 ();
 sg13g2_decap_8 FILLER_26_1762 ();
 sg13g2_decap_8 FILLER_26_1769 ();
 sg13g2_decap_8 FILLER_26_1776 ();
 sg13g2_decap_8 FILLER_26_1783 ();
 sg13g2_decap_8 FILLER_26_1790 ();
 sg13g2_decap_8 FILLER_26_1797 ();
 sg13g2_decap_8 FILLER_26_1804 ();
 sg13g2_decap_4 FILLER_26_1811 ();
 sg13g2_fill_2 FILLER_26_1815 ();
 sg13g2_decap_8 FILLER_26_1826 ();
 sg13g2_fill_1 FILLER_26_1833 ();
 sg13g2_decap_8 FILLER_26_1840 ();
 sg13g2_decap_8 FILLER_26_1847 ();
 sg13g2_decap_4 FILLER_26_1854 ();
 sg13g2_fill_1 FILLER_26_1858 ();
 sg13g2_decap_8 FILLER_26_1872 ();
 sg13g2_decap_8 FILLER_26_1879 ();
 sg13g2_decap_4 FILLER_26_1886 ();
 sg13g2_fill_2 FILLER_26_1890 ();
 sg13g2_decap_8 FILLER_26_1896 ();
 sg13g2_decap_8 FILLER_26_1903 ();
 sg13g2_decap_8 FILLER_26_1910 ();
 sg13g2_decap_8 FILLER_26_1917 ();
 sg13g2_decap_8 FILLER_26_1924 ();
 sg13g2_decap_8 FILLER_26_1931 ();
 sg13g2_decap_8 FILLER_26_1938 ();
 sg13g2_decap_8 FILLER_26_1945 ();
 sg13g2_decap_8 FILLER_26_1952 ();
 sg13g2_decap_8 FILLER_26_1959 ();
 sg13g2_decap_8 FILLER_26_1966 ();
 sg13g2_decap_8 FILLER_26_1973 ();
 sg13g2_decap_8 FILLER_26_1980 ();
 sg13g2_decap_8 FILLER_26_1987 ();
 sg13g2_decap_8 FILLER_26_1994 ();
 sg13g2_decap_8 FILLER_26_2001 ();
 sg13g2_decap_8 FILLER_26_2008 ();
 sg13g2_decap_8 FILLER_26_2015 ();
 sg13g2_decap_8 FILLER_26_2022 ();
 sg13g2_decap_8 FILLER_26_2029 ();
 sg13g2_decap_8 FILLER_26_2036 ();
 sg13g2_decap_8 FILLER_26_2043 ();
 sg13g2_decap_8 FILLER_26_2050 ();
 sg13g2_decap_8 FILLER_26_2057 ();
 sg13g2_decap_8 FILLER_26_2064 ();
 sg13g2_decap_8 FILLER_26_2071 ();
 sg13g2_decap_8 FILLER_26_2078 ();
 sg13g2_decap_8 FILLER_26_2085 ();
 sg13g2_decap_8 FILLER_26_2092 ();
 sg13g2_decap_8 FILLER_26_2099 ();
 sg13g2_decap_8 FILLER_26_2106 ();
 sg13g2_decap_8 FILLER_26_2113 ();
 sg13g2_decap_8 FILLER_26_2120 ();
 sg13g2_decap_8 FILLER_26_2127 ();
 sg13g2_decap_8 FILLER_26_2134 ();
 sg13g2_decap_8 FILLER_26_2141 ();
 sg13g2_decap_8 FILLER_26_2148 ();
 sg13g2_decap_8 FILLER_26_2155 ();
 sg13g2_decap_8 FILLER_26_2162 ();
 sg13g2_decap_8 FILLER_26_2169 ();
 sg13g2_decap_8 FILLER_26_2176 ();
 sg13g2_decap_8 FILLER_26_2183 ();
 sg13g2_decap_8 FILLER_26_2190 ();
 sg13g2_decap_8 FILLER_26_2197 ();
 sg13g2_decap_8 FILLER_26_2204 ();
 sg13g2_decap_8 FILLER_26_2211 ();
 sg13g2_decap_8 FILLER_26_2218 ();
 sg13g2_decap_8 FILLER_26_2225 ();
 sg13g2_decap_8 FILLER_26_2232 ();
 sg13g2_decap_8 FILLER_26_2239 ();
 sg13g2_decap_8 FILLER_26_2246 ();
 sg13g2_decap_8 FILLER_26_2253 ();
 sg13g2_decap_8 FILLER_26_2260 ();
 sg13g2_decap_8 FILLER_26_2267 ();
 sg13g2_decap_8 FILLER_26_2274 ();
 sg13g2_decap_8 FILLER_26_2281 ();
 sg13g2_decap_8 FILLER_26_2288 ();
 sg13g2_decap_8 FILLER_26_2295 ();
 sg13g2_decap_8 FILLER_26_2302 ();
 sg13g2_decap_8 FILLER_26_2309 ();
 sg13g2_decap_8 FILLER_26_2316 ();
 sg13g2_decap_8 FILLER_26_2323 ();
 sg13g2_decap_8 FILLER_26_2330 ();
 sg13g2_decap_8 FILLER_26_2337 ();
 sg13g2_decap_8 FILLER_26_2344 ();
 sg13g2_decap_8 FILLER_26_2351 ();
 sg13g2_decap_8 FILLER_26_2358 ();
 sg13g2_decap_8 FILLER_26_2365 ();
 sg13g2_decap_8 FILLER_26_2372 ();
 sg13g2_decap_8 FILLER_26_2379 ();
 sg13g2_decap_8 FILLER_26_2386 ();
 sg13g2_decap_8 FILLER_26_2393 ();
 sg13g2_decap_8 FILLER_26_2400 ();
 sg13g2_decap_8 FILLER_26_2407 ();
 sg13g2_decap_8 FILLER_26_2414 ();
 sg13g2_decap_8 FILLER_26_2421 ();
 sg13g2_decap_8 FILLER_26_2428 ();
 sg13g2_decap_8 FILLER_26_2435 ();
 sg13g2_decap_8 FILLER_26_2442 ();
 sg13g2_decap_8 FILLER_26_2449 ();
 sg13g2_decap_8 FILLER_26_2456 ();
 sg13g2_decap_8 FILLER_26_2463 ();
 sg13g2_decap_8 FILLER_26_2470 ();
 sg13g2_decap_8 FILLER_26_2477 ();
 sg13g2_decap_8 FILLER_26_2484 ();
 sg13g2_decap_8 FILLER_26_2491 ();
 sg13g2_decap_8 FILLER_26_2498 ();
 sg13g2_decap_8 FILLER_26_2505 ();
 sg13g2_decap_8 FILLER_26_2512 ();
 sg13g2_decap_8 FILLER_26_2519 ();
 sg13g2_decap_8 FILLER_26_2526 ();
 sg13g2_decap_8 FILLER_26_2533 ();
 sg13g2_decap_8 FILLER_26_2540 ();
 sg13g2_decap_8 FILLER_26_2547 ();
 sg13g2_decap_8 FILLER_26_2554 ();
 sg13g2_decap_8 FILLER_26_2561 ();
 sg13g2_decap_8 FILLER_26_2568 ();
 sg13g2_decap_8 FILLER_26_2575 ();
 sg13g2_decap_8 FILLER_26_2582 ();
 sg13g2_decap_8 FILLER_26_2589 ();
 sg13g2_decap_8 FILLER_26_2596 ();
 sg13g2_decap_8 FILLER_26_2603 ();
 sg13g2_decap_8 FILLER_26_2610 ();
 sg13g2_decap_8 FILLER_26_2617 ();
 sg13g2_decap_8 FILLER_26_2624 ();
 sg13g2_decap_8 FILLER_26_2631 ();
 sg13g2_decap_8 FILLER_26_2638 ();
 sg13g2_decap_8 FILLER_26_2645 ();
 sg13g2_decap_8 FILLER_26_2652 ();
 sg13g2_decap_8 FILLER_26_2659 ();
 sg13g2_decap_4 FILLER_26_2666 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_4 FILLER_27_49 ();
 sg13g2_fill_2 FILLER_27_53 ();
 sg13g2_decap_8 FILLER_27_81 ();
 sg13g2_decap_8 FILLER_27_88 ();
 sg13g2_decap_8 FILLER_27_95 ();
 sg13g2_decap_8 FILLER_27_102 ();
 sg13g2_fill_2 FILLER_27_109 ();
 sg13g2_decap_8 FILLER_27_115 ();
 sg13g2_decap_8 FILLER_27_122 ();
 sg13g2_decap_8 FILLER_27_129 ();
 sg13g2_decap_8 FILLER_27_136 ();
 sg13g2_decap_4 FILLER_27_143 ();
 sg13g2_fill_2 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_231 ();
 sg13g2_decap_8 FILLER_27_238 ();
 sg13g2_fill_1 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_255 ();
 sg13g2_decap_8 FILLER_27_262 ();
 sg13g2_decap_8 FILLER_27_269 ();
 sg13g2_decap_8 FILLER_27_276 ();
 sg13g2_decap_8 FILLER_27_283 ();
 sg13g2_decap_8 FILLER_27_290 ();
 sg13g2_decap_8 FILLER_27_297 ();
 sg13g2_decap_8 FILLER_27_304 ();
 sg13g2_decap_4 FILLER_27_311 ();
 sg13g2_decap_8 FILLER_27_319 ();
 sg13g2_decap_8 FILLER_27_326 ();
 sg13g2_decap_8 FILLER_27_333 ();
 sg13g2_decap_8 FILLER_27_340 ();
 sg13g2_decap_8 FILLER_27_347 ();
 sg13g2_decap_8 FILLER_27_354 ();
 sg13g2_decap_8 FILLER_27_361 ();
 sg13g2_decap_4 FILLER_27_368 ();
 sg13g2_fill_1 FILLER_27_372 ();
 sg13g2_decap_8 FILLER_27_377 ();
 sg13g2_decap_8 FILLER_27_384 ();
 sg13g2_decap_8 FILLER_27_391 ();
 sg13g2_decap_8 FILLER_27_398 ();
 sg13g2_decap_8 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_27_412 ();
 sg13g2_decap_8 FILLER_27_419 ();
 sg13g2_decap_8 FILLER_27_426 ();
 sg13g2_decap_8 FILLER_27_433 ();
 sg13g2_decap_8 FILLER_27_445 ();
 sg13g2_decap_8 FILLER_27_452 ();
 sg13g2_decap_8 FILLER_27_459 ();
 sg13g2_fill_1 FILLER_27_466 ();
 sg13g2_fill_2 FILLER_27_471 ();
 sg13g2_fill_1 FILLER_27_473 ();
 sg13g2_decap_8 FILLER_27_478 ();
 sg13g2_decap_8 FILLER_27_485 ();
 sg13g2_decap_8 FILLER_27_492 ();
 sg13g2_decap_8 FILLER_27_499 ();
 sg13g2_decap_8 FILLER_27_506 ();
 sg13g2_decap_8 FILLER_27_513 ();
 sg13g2_decap_8 FILLER_27_520 ();
 sg13g2_decap_8 FILLER_27_527 ();
 sg13g2_decap_8 FILLER_27_534 ();
 sg13g2_decap_8 FILLER_27_541 ();
 sg13g2_decap_8 FILLER_27_548 ();
 sg13g2_decap_8 FILLER_27_555 ();
 sg13g2_decap_4 FILLER_27_562 ();
 sg13g2_fill_1 FILLER_27_566 ();
 sg13g2_fill_1 FILLER_27_578 ();
 sg13g2_decap_8 FILLER_27_584 ();
 sg13g2_decap_8 FILLER_27_591 ();
 sg13g2_fill_1 FILLER_27_612 ();
 sg13g2_decap_8 FILLER_27_623 ();
 sg13g2_decap_8 FILLER_27_630 ();
 sg13g2_decap_8 FILLER_27_637 ();
 sg13g2_decap_8 FILLER_27_644 ();
 sg13g2_decap_8 FILLER_27_651 ();
 sg13g2_fill_2 FILLER_27_658 ();
 sg13g2_decap_4 FILLER_27_667 ();
 sg13g2_fill_2 FILLER_27_671 ();
 sg13g2_fill_1 FILLER_27_685 ();
 sg13g2_decap_4 FILLER_27_694 ();
 sg13g2_fill_2 FILLER_27_698 ();
 sg13g2_decap_8 FILLER_27_704 ();
 sg13g2_decap_8 FILLER_27_711 ();
 sg13g2_decap_8 FILLER_27_718 ();
 sg13g2_decap_8 FILLER_27_733 ();
 sg13g2_decap_8 FILLER_27_740 ();
 sg13g2_decap_8 FILLER_27_747 ();
 sg13g2_decap_8 FILLER_27_754 ();
 sg13g2_decap_8 FILLER_27_761 ();
 sg13g2_decap_8 FILLER_27_768 ();
 sg13g2_decap_4 FILLER_27_775 ();
 sg13g2_fill_1 FILLER_27_779 ();
 sg13g2_fill_1 FILLER_27_785 ();
 sg13g2_decap_8 FILLER_27_796 ();
 sg13g2_decap_4 FILLER_27_807 ();
 sg13g2_fill_1 FILLER_27_811 ();
 sg13g2_fill_2 FILLER_27_816 ();
 sg13g2_decap_8 FILLER_27_821 ();
 sg13g2_decap_8 FILLER_27_828 ();
 sg13g2_decap_8 FILLER_27_835 ();
 sg13g2_decap_8 FILLER_27_842 ();
 sg13g2_decap_8 FILLER_27_849 ();
 sg13g2_decap_8 FILLER_27_856 ();
 sg13g2_decap_8 FILLER_27_863 ();
 sg13g2_decap_8 FILLER_27_870 ();
 sg13g2_decap_8 FILLER_27_877 ();
 sg13g2_decap_8 FILLER_27_884 ();
 sg13g2_decap_8 FILLER_27_891 ();
 sg13g2_decap_8 FILLER_27_898 ();
 sg13g2_decap_8 FILLER_27_905 ();
 sg13g2_decap_8 FILLER_27_912 ();
 sg13g2_decap_4 FILLER_27_919 ();
 sg13g2_fill_2 FILLER_27_933 ();
 sg13g2_decap_4 FILLER_27_940 ();
 sg13g2_fill_1 FILLER_27_944 ();
 sg13g2_decap_4 FILLER_27_955 ();
 sg13g2_fill_2 FILLER_27_959 ();
 sg13g2_decap_4 FILLER_27_972 ();
 sg13g2_fill_1 FILLER_27_976 ();
 sg13g2_decap_8 FILLER_27_982 ();
 sg13g2_decap_8 FILLER_27_989 ();
 sg13g2_decap_8 FILLER_27_996 ();
 sg13g2_decap_8 FILLER_27_1003 ();
 sg13g2_decap_8 FILLER_27_1010 ();
 sg13g2_decap_8 FILLER_27_1017 ();
 sg13g2_fill_2 FILLER_27_1024 ();
 sg13g2_decap_8 FILLER_27_1029 ();
 sg13g2_decap_8 FILLER_27_1036 ();
 sg13g2_decap_8 FILLER_27_1043 ();
 sg13g2_decap_8 FILLER_27_1050 ();
 sg13g2_decap_8 FILLER_27_1057 ();
 sg13g2_decap_8 FILLER_27_1064 ();
 sg13g2_fill_2 FILLER_27_1071 ();
 sg13g2_decap_4 FILLER_27_1077 ();
 sg13g2_decap_8 FILLER_27_1085 ();
 sg13g2_fill_2 FILLER_27_1104 ();
 sg13g2_decap_8 FILLER_27_1112 ();
 sg13g2_decap_8 FILLER_27_1119 ();
 sg13g2_decap_8 FILLER_27_1126 ();
 sg13g2_decap_8 FILLER_27_1133 ();
 sg13g2_decap_4 FILLER_27_1140 ();
 sg13g2_fill_2 FILLER_27_1144 ();
 sg13g2_decap_8 FILLER_27_1150 ();
 sg13g2_decap_8 FILLER_27_1157 ();
 sg13g2_decap_8 FILLER_27_1164 ();
 sg13g2_decap_4 FILLER_27_1171 ();
 sg13g2_fill_1 FILLER_27_1175 ();
 sg13g2_decap_8 FILLER_27_1182 ();
 sg13g2_decap_8 FILLER_27_1189 ();
 sg13g2_decap_8 FILLER_27_1196 ();
 sg13g2_decap_8 FILLER_27_1203 ();
 sg13g2_decap_8 FILLER_27_1210 ();
 sg13g2_decap_8 FILLER_27_1217 ();
 sg13g2_decap_8 FILLER_27_1224 ();
 sg13g2_decap_8 FILLER_27_1231 ();
 sg13g2_decap_8 FILLER_27_1243 ();
 sg13g2_decap_8 FILLER_27_1250 ();
 sg13g2_decap_8 FILLER_27_1257 ();
 sg13g2_decap_8 FILLER_27_1264 ();
 sg13g2_decap_4 FILLER_27_1271 ();
 sg13g2_decap_8 FILLER_27_1290 ();
 sg13g2_decap_8 FILLER_27_1297 ();
 sg13g2_fill_2 FILLER_27_1304 ();
 sg13g2_fill_1 FILLER_27_1306 ();
 sg13g2_decap_8 FILLER_27_1314 ();
 sg13g2_decap_8 FILLER_27_1321 ();
 sg13g2_decap_8 FILLER_27_1328 ();
 sg13g2_decap_8 FILLER_27_1335 ();
 sg13g2_decap_8 FILLER_27_1342 ();
 sg13g2_decap_4 FILLER_27_1349 ();
 sg13g2_fill_2 FILLER_27_1353 ();
 sg13g2_decap_8 FILLER_27_1364 ();
 sg13g2_decap_8 FILLER_27_1371 ();
 sg13g2_decap_8 FILLER_27_1382 ();
 sg13g2_decap_8 FILLER_27_1389 ();
 sg13g2_decap_8 FILLER_27_1396 ();
 sg13g2_fill_1 FILLER_27_1406 ();
 sg13g2_fill_2 FILLER_27_1410 ();
 sg13g2_decap_8 FILLER_27_1427 ();
 sg13g2_decap_4 FILLER_27_1434 ();
 sg13g2_decap_8 FILLER_27_1441 ();
 sg13g2_decap_8 FILLER_27_1448 ();
 sg13g2_decap_8 FILLER_27_1455 ();
 sg13g2_decap_8 FILLER_27_1462 ();
 sg13g2_fill_1 FILLER_27_1469 ();
 sg13g2_decap_8 FILLER_27_1473 ();
 sg13g2_fill_2 FILLER_27_1480 ();
 sg13g2_decap_8 FILLER_27_1486 ();
 sg13g2_decap_4 FILLER_27_1493 ();
 sg13g2_fill_2 FILLER_27_1497 ();
 sg13g2_decap_8 FILLER_27_1504 ();
 sg13g2_decap_8 FILLER_27_1511 ();
 sg13g2_decap_4 FILLER_27_1518 ();
 sg13g2_fill_1 FILLER_27_1522 ();
 sg13g2_decap_8 FILLER_27_1529 ();
 sg13g2_decap_8 FILLER_27_1536 ();
 sg13g2_decap_8 FILLER_27_1543 ();
 sg13g2_decap_8 FILLER_27_1550 ();
 sg13g2_decap_8 FILLER_27_1557 ();
 sg13g2_decap_8 FILLER_27_1564 ();
 sg13g2_decap_4 FILLER_27_1571 ();
 sg13g2_fill_2 FILLER_27_1575 ();
 sg13g2_decap_8 FILLER_27_1592 ();
 sg13g2_decap_8 FILLER_27_1599 ();
 sg13g2_fill_1 FILLER_27_1606 ();
 sg13g2_decap_8 FILLER_27_1611 ();
 sg13g2_decap_8 FILLER_27_1618 ();
 sg13g2_decap_8 FILLER_27_1625 ();
 sg13g2_decap_8 FILLER_27_1632 ();
 sg13g2_fill_2 FILLER_27_1639 ();
 sg13g2_decap_8 FILLER_27_1649 ();
 sg13g2_decap_8 FILLER_27_1656 ();
 sg13g2_decap_8 FILLER_27_1663 ();
 sg13g2_decap_8 FILLER_27_1670 ();
 sg13g2_decap_8 FILLER_27_1677 ();
 sg13g2_decap_8 FILLER_27_1684 ();
 sg13g2_decap_8 FILLER_27_1691 ();
 sg13g2_decap_8 FILLER_27_1698 ();
 sg13g2_decap_8 FILLER_27_1705 ();
 sg13g2_decap_8 FILLER_27_1712 ();
 sg13g2_decap_8 FILLER_27_1719 ();
 sg13g2_decap_8 FILLER_27_1726 ();
 sg13g2_decap_8 FILLER_27_1733 ();
 sg13g2_decap_8 FILLER_27_1740 ();
 sg13g2_decap_8 FILLER_27_1747 ();
 sg13g2_decap_8 FILLER_27_1754 ();
 sg13g2_decap_8 FILLER_27_1761 ();
 sg13g2_decap_4 FILLER_27_1768 ();
 sg13g2_fill_2 FILLER_27_1772 ();
 sg13g2_fill_1 FILLER_27_1778 ();
 sg13g2_decap_8 FILLER_27_1783 ();
 sg13g2_decap_8 FILLER_27_1790 ();
 sg13g2_decap_8 FILLER_27_1797 ();
 sg13g2_decap_8 FILLER_27_1804 ();
 sg13g2_decap_8 FILLER_27_1811 ();
 sg13g2_decap_8 FILLER_27_1818 ();
 sg13g2_decap_8 FILLER_27_1825 ();
 sg13g2_decap_8 FILLER_27_1832 ();
 sg13g2_decap_8 FILLER_27_1839 ();
 sg13g2_decap_8 FILLER_27_1846 ();
 sg13g2_decap_8 FILLER_27_1853 ();
 sg13g2_decap_8 FILLER_27_1860 ();
 sg13g2_decap_8 FILLER_27_1867 ();
 sg13g2_decap_8 FILLER_27_1874 ();
 sg13g2_decap_8 FILLER_27_1881 ();
 sg13g2_decap_8 FILLER_27_1888 ();
 sg13g2_fill_2 FILLER_27_1895 ();
 sg13g2_decap_8 FILLER_27_1910 ();
 sg13g2_decap_8 FILLER_27_1917 ();
 sg13g2_decap_8 FILLER_27_1924 ();
 sg13g2_decap_8 FILLER_27_1931 ();
 sg13g2_decap_8 FILLER_27_1938 ();
 sg13g2_decap_8 FILLER_27_1945 ();
 sg13g2_decap_8 FILLER_27_1952 ();
 sg13g2_decap_8 FILLER_27_1959 ();
 sg13g2_decap_8 FILLER_27_1966 ();
 sg13g2_decap_8 FILLER_27_1973 ();
 sg13g2_decap_8 FILLER_27_1980 ();
 sg13g2_decap_8 FILLER_27_1987 ();
 sg13g2_decap_8 FILLER_27_1994 ();
 sg13g2_decap_8 FILLER_27_2001 ();
 sg13g2_decap_8 FILLER_27_2008 ();
 sg13g2_decap_8 FILLER_27_2015 ();
 sg13g2_decap_8 FILLER_27_2022 ();
 sg13g2_decap_8 FILLER_27_2029 ();
 sg13g2_decap_8 FILLER_27_2036 ();
 sg13g2_decap_8 FILLER_27_2043 ();
 sg13g2_decap_8 FILLER_27_2050 ();
 sg13g2_decap_8 FILLER_27_2057 ();
 sg13g2_decap_8 FILLER_27_2064 ();
 sg13g2_decap_8 FILLER_27_2071 ();
 sg13g2_decap_8 FILLER_27_2078 ();
 sg13g2_decap_8 FILLER_27_2085 ();
 sg13g2_decap_8 FILLER_27_2092 ();
 sg13g2_decap_8 FILLER_27_2099 ();
 sg13g2_decap_8 FILLER_27_2106 ();
 sg13g2_decap_8 FILLER_27_2113 ();
 sg13g2_decap_8 FILLER_27_2120 ();
 sg13g2_decap_8 FILLER_27_2127 ();
 sg13g2_decap_8 FILLER_27_2134 ();
 sg13g2_decap_8 FILLER_27_2141 ();
 sg13g2_decap_8 FILLER_27_2148 ();
 sg13g2_decap_8 FILLER_27_2155 ();
 sg13g2_decap_8 FILLER_27_2162 ();
 sg13g2_decap_8 FILLER_27_2169 ();
 sg13g2_decap_8 FILLER_27_2176 ();
 sg13g2_decap_8 FILLER_27_2183 ();
 sg13g2_decap_8 FILLER_27_2190 ();
 sg13g2_decap_8 FILLER_27_2197 ();
 sg13g2_decap_8 FILLER_27_2204 ();
 sg13g2_decap_8 FILLER_27_2211 ();
 sg13g2_decap_8 FILLER_27_2218 ();
 sg13g2_decap_8 FILLER_27_2225 ();
 sg13g2_decap_8 FILLER_27_2232 ();
 sg13g2_decap_8 FILLER_27_2239 ();
 sg13g2_decap_8 FILLER_27_2246 ();
 sg13g2_decap_8 FILLER_27_2253 ();
 sg13g2_decap_8 FILLER_27_2260 ();
 sg13g2_decap_8 FILLER_27_2267 ();
 sg13g2_decap_8 FILLER_27_2274 ();
 sg13g2_decap_8 FILLER_27_2281 ();
 sg13g2_decap_8 FILLER_27_2288 ();
 sg13g2_decap_8 FILLER_27_2295 ();
 sg13g2_decap_8 FILLER_27_2302 ();
 sg13g2_decap_8 FILLER_27_2309 ();
 sg13g2_decap_8 FILLER_27_2316 ();
 sg13g2_decap_8 FILLER_27_2323 ();
 sg13g2_decap_8 FILLER_27_2330 ();
 sg13g2_decap_8 FILLER_27_2337 ();
 sg13g2_decap_8 FILLER_27_2344 ();
 sg13g2_decap_8 FILLER_27_2351 ();
 sg13g2_decap_8 FILLER_27_2358 ();
 sg13g2_decap_8 FILLER_27_2365 ();
 sg13g2_decap_8 FILLER_27_2372 ();
 sg13g2_decap_8 FILLER_27_2379 ();
 sg13g2_decap_8 FILLER_27_2386 ();
 sg13g2_decap_8 FILLER_27_2393 ();
 sg13g2_decap_8 FILLER_27_2400 ();
 sg13g2_decap_8 FILLER_27_2407 ();
 sg13g2_decap_8 FILLER_27_2414 ();
 sg13g2_decap_8 FILLER_27_2421 ();
 sg13g2_decap_8 FILLER_27_2428 ();
 sg13g2_decap_8 FILLER_27_2435 ();
 sg13g2_decap_8 FILLER_27_2442 ();
 sg13g2_decap_8 FILLER_27_2449 ();
 sg13g2_decap_8 FILLER_27_2456 ();
 sg13g2_decap_8 FILLER_27_2463 ();
 sg13g2_decap_8 FILLER_27_2470 ();
 sg13g2_decap_8 FILLER_27_2477 ();
 sg13g2_decap_8 FILLER_27_2484 ();
 sg13g2_decap_8 FILLER_27_2491 ();
 sg13g2_decap_8 FILLER_27_2498 ();
 sg13g2_decap_8 FILLER_27_2505 ();
 sg13g2_decap_8 FILLER_27_2512 ();
 sg13g2_decap_8 FILLER_27_2519 ();
 sg13g2_decap_8 FILLER_27_2526 ();
 sg13g2_decap_8 FILLER_27_2533 ();
 sg13g2_decap_8 FILLER_27_2540 ();
 sg13g2_decap_8 FILLER_27_2547 ();
 sg13g2_decap_8 FILLER_27_2554 ();
 sg13g2_decap_8 FILLER_27_2561 ();
 sg13g2_decap_8 FILLER_27_2568 ();
 sg13g2_decap_8 FILLER_27_2575 ();
 sg13g2_decap_8 FILLER_27_2582 ();
 sg13g2_decap_8 FILLER_27_2589 ();
 sg13g2_decap_8 FILLER_27_2596 ();
 sg13g2_decap_8 FILLER_27_2603 ();
 sg13g2_decap_8 FILLER_27_2610 ();
 sg13g2_decap_8 FILLER_27_2617 ();
 sg13g2_decap_8 FILLER_27_2624 ();
 sg13g2_decap_8 FILLER_27_2631 ();
 sg13g2_decap_8 FILLER_27_2638 ();
 sg13g2_decap_8 FILLER_27_2645 ();
 sg13g2_decap_8 FILLER_27_2652 ();
 sg13g2_decap_8 FILLER_27_2659 ();
 sg13g2_decap_4 FILLER_27_2666 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_4 FILLER_28_49 ();
 sg13g2_fill_1 FILLER_28_53 ();
 sg13g2_fill_2 FILLER_28_58 ();
 sg13g2_decap_8 FILLER_28_64 ();
 sg13g2_decap_8 FILLER_28_71 ();
 sg13g2_decap_8 FILLER_28_78 ();
 sg13g2_decap_8 FILLER_28_85 ();
 sg13g2_decap_8 FILLER_28_92 ();
 sg13g2_decap_8 FILLER_28_99 ();
 sg13g2_decap_8 FILLER_28_106 ();
 sg13g2_decap_8 FILLER_28_113 ();
 sg13g2_decap_8 FILLER_28_120 ();
 sg13g2_decap_8 FILLER_28_127 ();
 sg13g2_decap_8 FILLER_28_134 ();
 sg13g2_decap_8 FILLER_28_141 ();
 sg13g2_decap_8 FILLER_28_148 ();
 sg13g2_decap_8 FILLER_28_155 ();
 sg13g2_decap_8 FILLER_28_162 ();
 sg13g2_decap_8 FILLER_28_169 ();
 sg13g2_decap_8 FILLER_28_176 ();
 sg13g2_decap_8 FILLER_28_183 ();
 sg13g2_decap_8 FILLER_28_190 ();
 sg13g2_decap_8 FILLER_28_197 ();
 sg13g2_decap_8 FILLER_28_204 ();
 sg13g2_decap_8 FILLER_28_211 ();
 sg13g2_decap_8 FILLER_28_218 ();
 sg13g2_decap_8 FILLER_28_225 ();
 sg13g2_decap_8 FILLER_28_232 ();
 sg13g2_decap_8 FILLER_28_239 ();
 sg13g2_decap_8 FILLER_28_246 ();
 sg13g2_decap_8 FILLER_28_253 ();
 sg13g2_decap_8 FILLER_28_260 ();
 sg13g2_decap_8 FILLER_28_267 ();
 sg13g2_decap_8 FILLER_28_274 ();
 sg13g2_decap_8 FILLER_28_281 ();
 sg13g2_decap_8 FILLER_28_288 ();
 sg13g2_decap_8 FILLER_28_295 ();
 sg13g2_decap_8 FILLER_28_302 ();
 sg13g2_decap_8 FILLER_28_309 ();
 sg13g2_decap_8 FILLER_28_316 ();
 sg13g2_decap_8 FILLER_28_323 ();
 sg13g2_decap_8 FILLER_28_330 ();
 sg13g2_decap_8 FILLER_28_337 ();
 sg13g2_decap_8 FILLER_28_344 ();
 sg13g2_decap_8 FILLER_28_351 ();
 sg13g2_decap_8 FILLER_28_358 ();
 sg13g2_decap_8 FILLER_28_365 ();
 sg13g2_decap_8 FILLER_28_372 ();
 sg13g2_decap_8 FILLER_28_379 ();
 sg13g2_decap_8 FILLER_28_386 ();
 sg13g2_decap_8 FILLER_28_393 ();
 sg13g2_decap_8 FILLER_28_400 ();
 sg13g2_decap_8 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_28_414 ();
 sg13g2_decap_8 FILLER_28_421 ();
 sg13g2_decap_4 FILLER_28_428 ();
 sg13g2_fill_1 FILLER_28_435 ();
 sg13g2_decap_4 FILLER_28_445 ();
 sg13g2_fill_1 FILLER_28_449 ();
 sg13g2_decap_8 FILLER_28_465 ();
 sg13g2_decap_8 FILLER_28_472 ();
 sg13g2_decap_8 FILLER_28_479 ();
 sg13g2_decap_8 FILLER_28_486 ();
 sg13g2_decap_4 FILLER_28_493 ();
 sg13g2_fill_1 FILLER_28_497 ();
 sg13g2_decap_8 FILLER_28_502 ();
 sg13g2_decap_4 FILLER_28_509 ();
 sg13g2_decap_8 FILLER_28_518 ();
 sg13g2_decap_8 FILLER_28_525 ();
 sg13g2_decap_8 FILLER_28_532 ();
 sg13g2_fill_2 FILLER_28_539 ();
 sg13g2_decap_8 FILLER_28_549 ();
 sg13g2_decap_8 FILLER_28_556 ();
 sg13g2_decap_8 FILLER_28_563 ();
 sg13g2_fill_1 FILLER_28_570 ();
 sg13g2_decap_8 FILLER_28_576 ();
 sg13g2_decap_8 FILLER_28_583 ();
 sg13g2_decap_8 FILLER_28_590 ();
 sg13g2_decap_8 FILLER_28_597 ();
 sg13g2_decap_8 FILLER_28_604 ();
 sg13g2_decap_8 FILLER_28_615 ();
 sg13g2_decap_8 FILLER_28_622 ();
 sg13g2_decap_8 FILLER_28_629 ();
 sg13g2_fill_2 FILLER_28_636 ();
 sg13g2_decap_8 FILLER_28_660 ();
 sg13g2_fill_2 FILLER_28_667 ();
 sg13g2_fill_1 FILLER_28_669 ();
 sg13g2_decap_8 FILLER_28_690 ();
 sg13g2_decap_8 FILLER_28_697 ();
 sg13g2_fill_1 FILLER_28_704 ();
 sg13g2_decap_8 FILLER_28_720 ();
 sg13g2_decap_4 FILLER_28_727 ();
 sg13g2_fill_1 FILLER_28_731 ();
 sg13g2_decap_8 FILLER_28_735 ();
 sg13g2_decap_8 FILLER_28_742 ();
 sg13g2_decap_8 FILLER_28_749 ();
 sg13g2_decap_8 FILLER_28_756 ();
 sg13g2_decap_8 FILLER_28_763 ();
 sg13g2_decap_8 FILLER_28_770 ();
 sg13g2_decap_8 FILLER_28_777 ();
 sg13g2_fill_2 FILLER_28_784 ();
 sg13g2_decap_8 FILLER_28_791 ();
 sg13g2_decap_8 FILLER_28_798 ();
 sg13g2_decap_8 FILLER_28_805 ();
 sg13g2_decap_8 FILLER_28_812 ();
 sg13g2_decap_8 FILLER_28_819 ();
 sg13g2_decap_8 FILLER_28_826 ();
 sg13g2_decap_8 FILLER_28_833 ();
 sg13g2_decap_4 FILLER_28_840 ();
 sg13g2_fill_1 FILLER_28_844 ();
 sg13g2_decap_8 FILLER_28_852 ();
 sg13g2_decap_8 FILLER_28_859 ();
 sg13g2_decap_8 FILLER_28_866 ();
 sg13g2_decap_8 FILLER_28_873 ();
 sg13g2_decap_8 FILLER_28_880 ();
 sg13g2_decap_8 FILLER_28_887 ();
 sg13g2_fill_2 FILLER_28_894 ();
 sg13g2_decap_8 FILLER_28_900 ();
 sg13g2_decap_8 FILLER_28_907 ();
 sg13g2_decap_8 FILLER_28_914 ();
 sg13g2_decap_8 FILLER_28_921 ();
 sg13g2_decap_8 FILLER_28_928 ();
 sg13g2_decap_8 FILLER_28_935 ();
 sg13g2_decap_4 FILLER_28_942 ();
 sg13g2_decap_8 FILLER_28_950 ();
 sg13g2_decap_8 FILLER_28_957 ();
 sg13g2_fill_2 FILLER_28_964 ();
 sg13g2_decap_8 FILLER_28_970 ();
 sg13g2_decap_8 FILLER_28_977 ();
 sg13g2_decap_8 FILLER_28_984 ();
 sg13g2_decap_8 FILLER_28_991 ();
 sg13g2_decap_8 FILLER_28_998 ();
 sg13g2_decap_8 FILLER_28_1005 ();
 sg13g2_decap_8 FILLER_28_1012 ();
 sg13g2_decap_8 FILLER_28_1019 ();
 sg13g2_decap_8 FILLER_28_1026 ();
 sg13g2_decap_8 FILLER_28_1033 ();
 sg13g2_decap_8 FILLER_28_1040 ();
 sg13g2_decap_8 FILLER_28_1047 ();
 sg13g2_decap_8 FILLER_28_1054 ();
 sg13g2_decap_8 FILLER_28_1061 ();
 sg13g2_decap_8 FILLER_28_1068 ();
 sg13g2_decap_8 FILLER_28_1075 ();
 sg13g2_decap_8 FILLER_28_1082 ();
 sg13g2_decap_4 FILLER_28_1089 ();
 sg13g2_fill_2 FILLER_28_1093 ();
 sg13g2_decap_8 FILLER_28_1109 ();
 sg13g2_decap_8 FILLER_28_1116 ();
 sg13g2_decap_8 FILLER_28_1123 ();
 sg13g2_decap_8 FILLER_28_1130 ();
 sg13g2_decap_8 FILLER_28_1137 ();
 sg13g2_decap_8 FILLER_28_1144 ();
 sg13g2_decap_8 FILLER_28_1151 ();
 sg13g2_decap_8 FILLER_28_1158 ();
 sg13g2_decap_8 FILLER_28_1165 ();
 sg13g2_decap_8 FILLER_28_1172 ();
 sg13g2_decap_8 FILLER_28_1185 ();
 sg13g2_decap_8 FILLER_28_1192 ();
 sg13g2_decap_8 FILLER_28_1199 ();
 sg13g2_decap_8 FILLER_28_1206 ();
 sg13g2_decap_8 FILLER_28_1213 ();
 sg13g2_decap_8 FILLER_28_1220 ();
 sg13g2_decap_8 FILLER_28_1227 ();
 sg13g2_decap_8 FILLER_28_1234 ();
 sg13g2_decap_8 FILLER_28_1241 ();
 sg13g2_decap_8 FILLER_28_1248 ();
 sg13g2_decap_8 FILLER_28_1255 ();
 sg13g2_decap_8 FILLER_28_1262 ();
 sg13g2_decap_8 FILLER_28_1285 ();
 sg13g2_decap_8 FILLER_28_1292 ();
 sg13g2_decap_8 FILLER_28_1299 ();
 sg13g2_fill_1 FILLER_28_1306 ();
 sg13g2_decap_8 FILLER_28_1312 ();
 sg13g2_decap_8 FILLER_28_1319 ();
 sg13g2_decap_8 FILLER_28_1326 ();
 sg13g2_decap_8 FILLER_28_1333 ();
 sg13g2_decap_8 FILLER_28_1340 ();
 sg13g2_fill_2 FILLER_28_1347 ();
 sg13g2_decap_8 FILLER_28_1362 ();
 sg13g2_decap_8 FILLER_28_1369 ();
 sg13g2_decap_8 FILLER_28_1376 ();
 sg13g2_decap_8 FILLER_28_1383 ();
 sg13g2_decap_8 FILLER_28_1390 ();
 sg13g2_decap_4 FILLER_28_1397 ();
 sg13g2_fill_2 FILLER_28_1410 ();
 sg13g2_decap_8 FILLER_28_1417 ();
 sg13g2_decap_8 FILLER_28_1424 ();
 sg13g2_decap_8 FILLER_28_1431 ();
 sg13g2_decap_8 FILLER_28_1438 ();
 sg13g2_decap_8 FILLER_28_1445 ();
 sg13g2_decap_4 FILLER_28_1452 ();
 sg13g2_decap_8 FILLER_28_1460 ();
 sg13g2_decap_8 FILLER_28_1475 ();
 sg13g2_decap_8 FILLER_28_1482 ();
 sg13g2_decap_4 FILLER_28_1489 ();
 sg13g2_fill_2 FILLER_28_1493 ();
 sg13g2_decap_8 FILLER_28_1511 ();
 sg13g2_decap_8 FILLER_28_1518 ();
 sg13g2_decap_8 FILLER_28_1525 ();
 sg13g2_decap_8 FILLER_28_1532 ();
 sg13g2_decap_8 FILLER_28_1539 ();
 sg13g2_decap_8 FILLER_28_1546 ();
 sg13g2_decap_8 FILLER_28_1553 ();
 sg13g2_fill_2 FILLER_28_1560 ();
 sg13g2_fill_1 FILLER_28_1562 ();
 sg13g2_decap_8 FILLER_28_1566 ();
 sg13g2_decap_8 FILLER_28_1582 ();
 sg13g2_decap_8 FILLER_28_1589 ();
 sg13g2_decap_4 FILLER_28_1596 ();
 sg13g2_decap_8 FILLER_28_1612 ();
 sg13g2_decap_8 FILLER_28_1619 ();
 sg13g2_fill_1 FILLER_28_1626 ();
 sg13g2_decap_8 FILLER_28_1636 ();
 sg13g2_decap_8 FILLER_28_1643 ();
 sg13g2_decap_8 FILLER_28_1650 ();
 sg13g2_decap_4 FILLER_28_1657 ();
 sg13g2_decap_8 FILLER_28_1667 ();
 sg13g2_fill_2 FILLER_28_1674 ();
 sg13g2_decap_8 FILLER_28_1684 ();
 sg13g2_decap_8 FILLER_28_1691 ();
 sg13g2_decap_8 FILLER_28_1698 ();
 sg13g2_decap_8 FILLER_28_1705 ();
 sg13g2_decap_8 FILLER_28_1712 ();
 sg13g2_decap_8 FILLER_28_1719 ();
 sg13g2_decap_8 FILLER_28_1726 ();
 sg13g2_decap_8 FILLER_28_1733 ();
 sg13g2_decap_8 FILLER_28_1740 ();
 sg13g2_decap_8 FILLER_28_1747 ();
 sg13g2_decap_8 FILLER_28_1754 ();
 sg13g2_decap_8 FILLER_28_1761 ();
 sg13g2_decap_8 FILLER_28_1768 ();
 sg13g2_decap_8 FILLER_28_1775 ();
 sg13g2_decap_8 FILLER_28_1782 ();
 sg13g2_decap_8 FILLER_28_1789 ();
 sg13g2_decap_8 FILLER_28_1796 ();
 sg13g2_decap_8 FILLER_28_1803 ();
 sg13g2_decap_8 FILLER_28_1810 ();
 sg13g2_decap_8 FILLER_28_1817 ();
 sg13g2_decap_8 FILLER_28_1824 ();
 sg13g2_decap_8 FILLER_28_1831 ();
 sg13g2_decap_8 FILLER_28_1838 ();
 sg13g2_decap_8 FILLER_28_1845 ();
 sg13g2_decap_8 FILLER_28_1852 ();
 sg13g2_decap_8 FILLER_28_1859 ();
 sg13g2_decap_8 FILLER_28_1866 ();
 sg13g2_decap_8 FILLER_28_1873 ();
 sg13g2_decap_8 FILLER_28_1880 ();
 sg13g2_decap_8 FILLER_28_1887 ();
 sg13g2_decap_8 FILLER_28_1894 ();
 sg13g2_decap_8 FILLER_28_1901 ();
 sg13g2_decap_8 FILLER_28_1908 ();
 sg13g2_decap_8 FILLER_28_1915 ();
 sg13g2_decap_8 FILLER_28_1922 ();
 sg13g2_decap_8 FILLER_28_1929 ();
 sg13g2_decap_8 FILLER_28_1936 ();
 sg13g2_decap_8 FILLER_28_1943 ();
 sg13g2_decap_8 FILLER_28_1950 ();
 sg13g2_decap_8 FILLER_28_1957 ();
 sg13g2_decap_8 FILLER_28_1964 ();
 sg13g2_decap_8 FILLER_28_1971 ();
 sg13g2_decap_8 FILLER_28_1978 ();
 sg13g2_decap_8 FILLER_28_1985 ();
 sg13g2_decap_8 FILLER_28_1992 ();
 sg13g2_decap_8 FILLER_28_1999 ();
 sg13g2_decap_8 FILLER_28_2006 ();
 sg13g2_decap_8 FILLER_28_2013 ();
 sg13g2_decap_8 FILLER_28_2020 ();
 sg13g2_decap_8 FILLER_28_2027 ();
 sg13g2_decap_8 FILLER_28_2034 ();
 sg13g2_decap_8 FILLER_28_2041 ();
 sg13g2_decap_8 FILLER_28_2048 ();
 sg13g2_decap_8 FILLER_28_2055 ();
 sg13g2_decap_8 FILLER_28_2062 ();
 sg13g2_decap_8 FILLER_28_2069 ();
 sg13g2_decap_8 FILLER_28_2076 ();
 sg13g2_decap_8 FILLER_28_2083 ();
 sg13g2_decap_8 FILLER_28_2090 ();
 sg13g2_decap_8 FILLER_28_2097 ();
 sg13g2_decap_8 FILLER_28_2104 ();
 sg13g2_decap_8 FILLER_28_2111 ();
 sg13g2_decap_8 FILLER_28_2118 ();
 sg13g2_decap_8 FILLER_28_2125 ();
 sg13g2_decap_8 FILLER_28_2132 ();
 sg13g2_decap_8 FILLER_28_2139 ();
 sg13g2_decap_8 FILLER_28_2146 ();
 sg13g2_decap_8 FILLER_28_2153 ();
 sg13g2_decap_8 FILLER_28_2160 ();
 sg13g2_decap_8 FILLER_28_2167 ();
 sg13g2_decap_8 FILLER_28_2174 ();
 sg13g2_decap_8 FILLER_28_2181 ();
 sg13g2_decap_8 FILLER_28_2188 ();
 sg13g2_decap_8 FILLER_28_2195 ();
 sg13g2_decap_8 FILLER_28_2202 ();
 sg13g2_decap_8 FILLER_28_2209 ();
 sg13g2_decap_8 FILLER_28_2216 ();
 sg13g2_decap_8 FILLER_28_2223 ();
 sg13g2_decap_8 FILLER_28_2230 ();
 sg13g2_decap_8 FILLER_28_2237 ();
 sg13g2_decap_8 FILLER_28_2244 ();
 sg13g2_decap_8 FILLER_28_2251 ();
 sg13g2_decap_8 FILLER_28_2258 ();
 sg13g2_decap_8 FILLER_28_2265 ();
 sg13g2_decap_8 FILLER_28_2272 ();
 sg13g2_decap_8 FILLER_28_2279 ();
 sg13g2_decap_8 FILLER_28_2286 ();
 sg13g2_decap_8 FILLER_28_2293 ();
 sg13g2_decap_8 FILLER_28_2300 ();
 sg13g2_decap_8 FILLER_28_2307 ();
 sg13g2_decap_8 FILLER_28_2314 ();
 sg13g2_decap_8 FILLER_28_2321 ();
 sg13g2_decap_8 FILLER_28_2328 ();
 sg13g2_decap_8 FILLER_28_2335 ();
 sg13g2_decap_8 FILLER_28_2342 ();
 sg13g2_decap_8 FILLER_28_2349 ();
 sg13g2_decap_8 FILLER_28_2356 ();
 sg13g2_decap_8 FILLER_28_2363 ();
 sg13g2_decap_8 FILLER_28_2370 ();
 sg13g2_decap_8 FILLER_28_2377 ();
 sg13g2_decap_8 FILLER_28_2384 ();
 sg13g2_decap_8 FILLER_28_2391 ();
 sg13g2_decap_8 FILLER_28_2398 ();
 sg13g2_decap_8 FILLER_28_2405 ();
 sg13g2_decap_8 FILLER_28_2412 ();
 sg13g2_decap_8 FILLER_28_2419 ();
 sg13g2_decap_8 FILLER_28_2426 ();
 sg13g2_decap_8 FILLER_28_2433 ();
 sg13g2_decap_8 FILLER_28_2440 ();
 sg13g2_decap_8 FILLER_28_2447 ();
 sg13g2_decap_8 FILLER_28_2454 ();
 sg13g2_decap_8 FILLER_28_2461 ();
 sg13g2_decap_8 FILLER_28_2468 ();
 sg13g2_decap_8 FILLER_28_2475 ();
 sg13g2_decap_8 FILLER_28_2482 ();
 sg13g2_decap_8 FILLER_28_2489 ();
 sg13g2_decap_8 FILLER_28_2496 ();
 sg13g2_decap_8 FILLER_28_2503 ();
 sg13g2_decap_8 FILLER_28_2510 ();
 sg13g2_decap_8 FILLER_28_2517 ();
 sg13g2_decap_8 FILLER_28_2524 ();
 sg13g2_decap_8 FILLER_28_2531 ();
 sg13g2_decap_8 FILLER_28_2538 ();
 sg13g2_decap_8 FILLER_28_2545 ();
 sg13g2_decap_8 FILLER_28_2552 ();
 sg13g2_decap_8 FILLER_28_2559 ();
 sg13g2_decap_8 FILLER_28_2566 ();
 sg13g2_decap_8 FILLER_28_2573 ();
 sg13g2_decap_8 FILLER_28_2580 ();
 sg13g2_decap_8 FILLER_28_2587 ();
 sg13g2_decap_8 FILLER_28_2594 ();
 sg13g2_decap_8 FILLER_28_2601 ();
 sg13g2_decap_8 FILLER_28_2608 ();
 sg13g2_decap_8 FILLER_28_2615 ();
 sg13g2_decap_8 FILLER_28_2622 ();
 sg13g2_decap_8 FILLER_28_2629 ();
 sg13g2_decap_8 FILLER_28_2636 ();
 sg13g2_decap_8 FILLER_28_2643 ();
 sg13g2_decap_8 FILLER_28_2650 ();
 sg13g2_decap_8 FILLER_28_2657 ();
 sg13g2_decap_4 FILLER_28_2664 ();
 sg13g2_fill_2 FILLER_28_2668 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_fill_1 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_76 ();
 sg13g2_decap_8 FILLER_29_83 ();
 sg13g2_decap_8 FILLER_29_90 ();
 sg13g2_decap_8 FILLER_29_97 ();
 sg13g2_decap_8 FILLER_29_104 ();
 sg13g2_decap_8 FILLER_29_111 ();
 sg13g2_decap_8 FILLER_29_118 ();
 sg13g2_decap_8 FILLER_29_125 ();
 sg13g2_decap_8 FILLER_29_132 ();
 sg13g2_decap_8 FILLER_29_139 ();
 sg13g2_fill_2 FILLER_29_146 ();
 sg13g2_fill_1 FILLER_29_148 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_decap_8 FILLER_29_182 ();
 sg13g2_decap_8 FILLER_29_189 ();
 sg13g2_fill_2 FILLER_29_196 ();
 sg13g2_fill_1 FILLER_29_198 ();
 sg13g2_decap_8 FILLER_29_225 ();
 sg13g2_decap_8 FILLER_29_232 ();
 sg13g2_decap_8 FILLER_29_239 ();
 sg13g2_decap_8 FILLER_29_246 ();
 sg13g2_decap_8 FILLER_29_253 ();
 sg13g2_decap_8 FILLER_29_260 ();
 sg13g2_decap_8 FILLER_29_267 ();
 sg13g2_decap_8 FILLER_29_274 ();
 sg13g2_decap_8 FILLER_29_281 ();
 sg13g2_decap_8 FILLER_29_288 ();
 sg13g2_decap_8 FILLER_29_295 ();
 sg13g2_decap_8 FILLER_29_302 ();
 sg13g2_decap_8 FILLER_29_309 ();
 sg13g2_decap_8 FILLER_29_316 ();
 sg13g2_decap_8 FILLER_29_323 ();
 sg13g2_decap_8 FILLER_29_330 ();
 sg13g2_decap_8 FILLER_29_337 ();
 sg13g2_decap_8 FILLER_29_344 ();
 sg13g2_decap_8 FILLER_29_351 ();
 sg13g2_decap_8 FILLER_29_358 ();
 sg13g2_decap_8 FILLER_29_365 ();
 sg13g2_decap_8 FILLER_29_372 ();
 sg13g2_decap_8 FILLER_29_379 ();
 sg13g2_decap_8 FILLER_29_386 ();
 sg13g2_decap_8 FILLER_29_393 ();
 sg13g2_fill_2 FILLER_29_400 ();
 sg13g2_fill_1 FILLER_29_402 ();
 sg13g2_decap_8 FILLER_29_412 ();
 sg13g2_decap_8 FILLER_29_419 ();
 sg13g2_decap_8 FILLER_29_426 ();
 sg13g2_decap_8 FILLER_29_433 ();
 sg13g2_decap_8 FILLER_29_440 ();
 sg13g2_decap_4 FILLER_29_447 ();
 sg13g2_fill_2 FILLER_29_451 ();
 sg13g2_decap_8 FILLER_29_458 ();
 sg13g2_decap_8 FILLER_29_465 ();
 sg13g2_decap_8 FILLER_29_472 ();
 sg13g2_decap_8 FILLER_29_479 ();
 sg13g2_decap_8 FILLER_29_486 ();
 sg13g2_decap_8 FILLER_29_493 ();
 sg13g2_decap_8 FILLER_29_500 ();
 sg13g2_decap_8 FILLER_29_507 ();
 sg13g2_decap_8 FILLER_29_514 ();
 sg13g2_decap_8 FILLER_29_521 ();
 sg13g2_decap_8 FILLER_29_528 ();
 sg13g2_fill_2 FILLER_29_535 ();
 sg13g2_decap_8 FILLER_29_540 ();
 sg13g2_decap_8 FILLER_29_547 ();
 sg13g2_decap_8 FILLER_29_554 ();
 sg13g2_decap_8 FILLER_29_561 ();
 sg13g2_decap_8 FILLER_29_568 ();
 sg13g2_decap_8 FILLER_29_575 ();
 sg13g2_decap_8 FILLER_29_582 ();
 sg13g2_decap_8 FILLER_29_589 ();
 sg13g2_decap_8 FILLER_29_596 ();
 sg13g2_fill_2 FILLER_29_603 ();
 sg13g2_fill_1 FILLER_29_605 ();
 sg13g2_decap_8 FILLER_29_610 ();
 sg13g2_decap_8 FILLER_29_617 ();
 sg13g2_decap_8 FILLER_29_624 ();
 sg13g2_decap_8 FILLER_29_631 ();
 sg13g2_decap_8 FILLER_29_638 ();
 sg13g2_fill_2 FILLER_29_645 ();
 sg13g2_fill_2 FILLER_29_651 ();
 sg13g2_decap_8 FILLER_29_657 ();
 sg13g2_decap_8 FILLER_29_664 ();
 sg13g2_decap_8 FILLER_29_671 ();
 sg13g2_decap_8 FILLER_29_678 ();
 sg13g2_decap_8 FILLER_29_685 ();
 sg13g2_decap_4 FILLER_29_692 ();
 sg13g2_decap_8 FILLER_29_716 ();
 sg13g2_decap_8 FILLER_29_723 ();
 sg13g2_decap_8 FILLER_29_730 ();
 sg13g2_decap_8 FILLER_29_737 ();
 sg13g2_decap_8 FILLER_29_744 ();
 sg13g2_decap_8 FILLER_29_751 ();
 sg13g2_decap_8 FILLER_29_758 ();
 sg13g2_decap_8 FILLER_29_765 ();
 sg13g2_decap_8 FILLER_29_772 ();
 sg13g2_decap_8 FILLER_29_779 ();
 sg13g2_fill_2 FILLER_29_786 ();
 sg13g2_decap_8 FILLER_29_816 ();
 sg13g2_decap_8 FILLER_29_823 ();
 sg13g2_decap_8 FILLER_29_830 ();
 sg13g2_decap_8 FILLER_29_837 ();
 sg13g2_decap_8 FILLER_29_844 ();
 sg13g2_decap_8 FILLER_29_851 ();
 sg13g2_decap_8 FILLER_29_858 ();
 sg13g2_decap_8 FILLER_29_865 ();
 sg13g2_decap_8 FILLER_29_872 ();
 sg13g2_decap_8 FILLER_29_879 ();
 sg13g2_decap_8 FILLER_29_886 ();
 sg13g2_decap_4 FILLER_29_893 ();
 sg13g2_fill_1 FILLER_29_897 ();
 sg13g2_decap_8 FILLER_29_922 ();
 sg13g2_decap_8 FILLER_29_929 ();
 sg13g2_decap_8 FILLER_29_936 ();
 sg13g2_decap_8 FILLER_29_943 ();
 sg13g2_decap_8 FILLER_29_950 ();
 sg13g2_decap_8 FILLER_29_957 ();
 sg13g2_decap_8 FILLER_29_964 ();
 sg13g2_decap_8 FILLER_29_971 ();
 sg13g2_decap_4 FILLER_29_978 ();
 sg13g2_fill_2 FILLER_29_982 ();
 sg13g2_decap_8 FILLER_29_988 ();
 sg13g2_decap_8 FILLER_29_995 ();
 sg13g2_decap_8 FILLER_29_1002 ();
 sg13g2_decap_8 FILLER_29_1009 ();
 sg13g2_decap_8 FILLER_29_1016 ();
 sg13g2_decap_4 FILLER_29_1023 ();
 sg13g2_fill_2 FILLER_29_1027 ();
 sg13g2_fill_1 FILLER_29_1044 ();
 sg13g2_decap_8 FILLER_29_1054 ();
 sg13g2_decap_4 FILLER_29_1061 ();
 sg13g2_decap_8 FILLER_29_1092 ();
 sg13g2_fill_2 FILLER_29_1099 ();
 sg13g2_decap_8 FILLER_29_1107 ();
 sg13g2_decap_8 FILLER_29_1114 ();
 sg13g2_decap_8 FILLER_29_1121 ();
 sg13g2_decap_8 FILLER_29_1128 ();
 sg13g2_decap_8 FILLER_29_1135 ();
 sg13g2_decap_8 FILLER_29_1142 ();
 sg13g2_decap_8 FILLER_29_1149 ();
 sg13g2_decap_8 FILLER_29_1156 ();
 sg13g2_decap_4 FILLER_29_1163 ();
 sg13g2_fill_1 FILLER_29_1167 ();
 sg13g2_decap_8 FILLER_29_1188 ();
 sg13g2_decap_8 FILLER_29_1195 ();
 sg13g2_decap_8 FILLER_29_1210 ();
 sg13g2_decap_8 FILLER_29_1217 ();
 sg13g2_decap_8 FILLER_29_1224 ();
 sg13g2_decap_8 FILLER_29_1231 ();
 sg13g2_decap_8 FILLER_29_1238 ();
 sg13g2_decap_8 FILLER_29_1245 ();
 sg13g2_decap_8 FILLER_29_1252 ();
 sg13g2_decap_8 FILLER_29_1259 ();
 sg13g2_decap_8 FILLER_29_1266 ();
 sg13g2_decap_4 FILLER_29_1273 ();
 sg13g2_decap_8 FILLER_29_1282 ();
 sg13g2_decap_8 FILLER_29_1289 ();
 sg13g2_decap_8 FILLER_29_1296 ();
 sg13g2_decap_4 FILLER_29_1303 ();
 sg13g2_decap_8 FILLER_29_1313 ();
 sg13g2_decap_8 FILLER_29_1320 ();
 sg13g2_decap_4 FILLER_29_1327 ();
 sg13g2_fill_2 FILLER_29_1331 ();
 sg13g2_decap_8 FILLER_29_1337 ();
 sg13g2_fill_1 FILLER_29_1344 ();
 sg13g2_decap_8 FILLER_29_1349 ();
 sg13g2_decap_8 FILLER_29_1356 ();
 sg13g2_decap_8 FILLER_29_1363 ();
 sg13g2_decap_8 FILLER_29_1370 ();
 sg13g2_decap_8 FILLER_29_1377 ();
 sg13g2_decap_8 FILLER_29_1384 ();
 sg13g2_decap_8 FILLER_29_1391 ();
 sg13g2_decap_4 FILLER_29_1398 ();
 sg13g2_fill_2 FILLER_29_1402 ();
 sg13g2_fill_2 FILLER_29_1409 ();
 sg13g2_fill_1 FILLER_29_1411 ();
 sg13g2_decap_8 FILLER_29_1432 ();
 sg13g2_decap_8 FILLER_29_1439 ();
 sg13g2_decap_8 FILLER_29_1446 ();
 sg13g2_decap_8 FILLER_29_1453 ();
 sg13g2_fill_1 FILLER_29_1460 ();
 sg13g2_decap_4 FILLER_29_1465 ();
 sg13g2_fill_1 FILLER_29_1469 ();
 sg13g2_decap_8 FILLER_29_1473 ();
 sg13g2_decap_8 FILLER_29_1480 ();
 sg13g2_decap_8 FILLER_29_1487 ();
 sg13g2_decap_4 FILLER_29_1494 ();
 sg13g2_fill_2 FILLER_29_1498 ();
 sg13g2_fill_1 FILLER_29_1503 ();
 sg13g2_decap_8 FILLER_29_1517 ();
 sg13g2_decap_8 FILLER_29_1524 ();
 sg13g2_decap_8 FILLER_29_1531 ();
 sg13g2_decap_8 FILLER_29_1538 ();
 sg13g2_decap_8 FILLER_29_1545 ();
 sg13g2_decap_4 FILLER_29_1552 ();
 sg13g2_fill_1 FILLER_29_1556 ();
 sg13g2_fill_1 FILLER_29_1573 ();
 sg13g2_decap_4 FILLER_29_1591 ();
 sg13g2_fill_1 FILLER_29_1595 ();
 sg13g2_fill_1 FILLER_29_1599 ();
 sg13g2_decap_8 FILLER_29_1607 ();
 sg13g2_decap_4 FILLER_29_1626 ();
 sg13g2_fill_2 FILLER_29_1640 ();
 sg13g2_fill_1 FILLER_29_1642 ();
 sg13g2_decap_8 FILLER_29_1648 ();
 sg13g2_decap_8 FILLER_29_1655 ();
 sg13g2_fill_1 FILLER_29_1662 ();
 sg13g2_decap_8 FILLER_29_1668 ();
 sg13g2_decap_8 FILLER_29_1675 ();
 sg13g2_decap_8 FILLER_29_1682 ();
 sg13g2_decap_8 FILLER_29_1689 ();
 sg13g2_fill_1 FILLER_29_1696 ();
 sg13g2_decap_8 FILLER_29_1707 ();
 sg13g2_decap_8 FILLER_29_1714 ();
 sg13g2_decap_8 FILLER_29_1721 ();
 sg13g2_decap_8 FILLER_29_1728 ();
 sg13g2_decap_8 FILLER_29_1735 ();
 sg13g2_decap_8 FILLER_29_1742 ();
 sg13g2_decap_8 FILLER_29_1749 ();
 sg13g2_decap_8 FILLER_29_1756 ();
 sg13g2_decap_8 FILLER_29_1763 ();
 sg13g2_fill_2 FILLER_29_1770 ();
 sg13g2_decap_4 FILLER_29_1776 ();
 sg13g2_decap_8 FILLER_29_1795 ();
 sg13g2_decap_8 FILLER_29_1802 ();
 sg13g2_decap_8 FILLER_29_1809 ();
 sg13g2_decap_8 FILLER_29_1816 ();
 sg13g2_decap_8 FILLER_29_1823 ();
 sg13g2_decap_8 FILLER_29_1830 ();
 sg13g2_decap_8 FILLER_29_1837 ();
 sg13g2_decap_8 FILLER_29_1844 ();
 sg13g2_decap_8 FILLER_29_1851 ();
 sg13g2_fill_2 FILLER_29_1858 ();
 sg13g2_fill_1 FILLER_29_1860 ();
 sg13g2_decap_8 FILLER_29_1876 ();
 sg13g2_decap_8 FILLER_29_1883 ();
 sg13g2_decap_8 FILLER_29_1890 ();
 sg13g2_decap_8 FILLER_29_1897 ();
 sg13g2_decap_8 FILLER_29_1904 ();
 sg13g2_decap_8 FILLER_29_1911 ();
 sg13g2_decap_8 FILLER_29_1918 ();
 sg13g2_decap_8 FILLER_29_1925 ();
 sg13g2_decap_8 FILLER_29_1932 ();
 sg13g2_decap_8 FILLER_29_1939 ();
 sg13g2_decap_8 FILLER_29_1946 ();
 sg13g2_decap_8 FILLER_29_1953 ();
 sg13g2_decap_8 FILLER_29_1960 ();
 sg13g2_decap_8 FILLER_29_1967 ();
 sg13g2_decap_8 FILLER_29_1974 ();
 sg13g2_decap_8 FILLER_29_1981 ();
 sg13g2_decap_8 FILLER_29_1988 ();
 sg13g2_decap_8 FILLER_29_1995 ();
 sg13g2_decap_8 FILLER_29_2002 ();
 sg13g2_decap_8 FILLER_29_2009 ();
 sg13g2_decap_8 FILLER_29_2016 ();
 sg13g2_decap_8 FILLER_29_2023 ();
 sg13g2_decap_8 FILLER_29_2030 ();
 sg13g2_decap_8 FILLER_29_2037 ();
 sg13g2_decap_8 FILLER_29_2044 ();
 sg13g2_decap_8 FILLER_29_2051 ();
 sg13g2_decap_8 FILLER_29_2058 ();
 sg13g2_decap_8 FILLER_29_2065 ();
 sg13g2_decap_8 FILLER_29_2072 ();
 sg13g2_decap_8 FILLER_29_2079 ();
 sg13g2_decap_8 FILLER_29_2086 ();
 sg13g2_decap_8 FILLER_29_2093 ();
 sg13g2_decap_8 FILLER_29_2100 ();
 sg13g2_decap_8 FILLER_29_2107 ();
 sg13g2_decap_8 FILLER_29_2114 ();
 sg13g2_decap_8 FILLER_29_2121 ();
 sg13g2_decap_8 FILLER_29_2128 ();
 sg13g2_decap_8 FILLER_29_2135 ();
 sg13g2_decap_8 FILLER_29_2142 ();
 sg13g2_decap_8 FILLER_29_2149 ();
 sg13g2_decap_8 FILLER_29_2156 ();
 sg13g2_decap_8 FILLER_29_2163 ();
 sg13g2_decap_8 FILLER_29_2170 ();
 sg13g2_decap_8 FILLER_29_2177 ();
 sg13g2_decap_8 FILLER_29_2184 ();
 sg13g2_decap_8 FILLER_29_2191 ();
 sg13g2_decap_8 FILLER_29_2198 ();
 sg13g2_decap_8 FILLER_29_2205 ();
 sg13g2_decap_8 FILLER_29_2212 ();
 sg13g2_decap_8 FILLER_29_2219 ();
 sg13g2_decap_8 FILLER_29_2226 ();
 sg13g2_decap_8 FILLER_29_2233 ();
 sg13g2_decap_8 FILLER_29_2240 ();
 sg13g2_decap_8 FILLER_29_2247 ();
 sg13g2_decap_8 FILLER_29_2254 ();
 sg13g2_decap_8 FILLER_29_2261 ();
 sg13g2_decap_8 FILLER_29_2268 ();
 sg13g2_decap_8 FILLER_29_2275 ();
 sg13g2_decap_8 FILLER_29_2282 ();
 sg13g2_decap_8 FILLER_29_2289 ();
 sg13g2_decap_8 FILLER_29_2296 ();
 sg13g2_decap_8 FILLER_29_2303 ();
 sg13g2_decap_8 FILLER_29_2310 ();
 sg13g2_decap_8 FILLER_29_2317 ();
 sg13g2_decap_8 FILLER_29_2324 ();
 sg13g2_decap_8 FILLER_29_2331 ();
 sg13g2_decap_8 FILLER_29_2338 ();
 sg13g2_decap_8 FILLER_29_2345 ();
 sg13g2_decap_8 FILLER_29_2352 ();
 sg13g2_decap_8 FILLER_29_2359 ();
 sg13g2_decap_8 FILLER_29_2366 ();
 sg13g2_decap_8 FILLER_29_2373 ();
 sg13g2_decap_8 FILLER_29_2380 ();
 sg13g2_decap_8 FILLER_29_2387 ();
 sg13g2_decap_8 FILLER_29_2394 ();
 sg13g2_decap_8 FILLER_29_2401 ();
 sg13g2_decap_8 FILLER_29_2408 ();
 sg13g2_decap_8 FILLER_29_2415 ();
 sg13g2_decap_8 FILLER_29_2422 ();
 sg13g2_decap_8 FILLER_29_2429 ();
 sg13g2_decap_8 FILLER_29_2436 ();
 sg13g2_decap_8 FILLER_29_2443 ();
 sg13g2_decap_8 FILLER_29_2450 ();
 sg13g2_decap_8 FILLER_29_2457 ();
 sg13g2_decap_8 FILLER_29_2464 ();
 sg13g2_decap_8 FILLER_29_2471 ();
 sg13g2_decap_8 FILLER_29_2478 ();
 sg13g2_decap_8 FILLER_29_2485 ();
 sg13g2_decap_8 FILLER_29_2492 ();
 sg13g2_decap_8 FILLER_29_2499 ();
 sg13g2_decap_8 FILLER_29_2506 ();
 sg13g2_decap_8 FILLER_29_2513 ();
 sg13g2_decap_8 FILLER_29_2520 ();
 sg13g2_decap_8 FILLER_29_2527 ();
 sg13g2_decap_8 FILLER_29_2534 ();
 sg13g2_decap_8 FILLER_29_2541 ();
 sg13g2_decap_8 FILLER_29_2548 ();
 sg13g2_decap_8 FILLER_29_2555 ();
 sg13g2_decap_8 FILLER_29_2562 ();
 sg13g2_decap_8 FILLER_29_2569 ();
 sg13g2_decap_8 FILLER_29_2576 ();
 sg13g2_decap_8 FILLER_29_2583 ();
 sg13g2_decap_8 FILLER_29_2590 ();
 sg13g2_decap_8 FILLER_29_2597 ();
 sg13g2_decap_8 FILLER_29_2604 ();
 sg13g2_decap_8 FILLER_29_2611 ();
 sg13g2_decap_8 FILLER_29_2618 ();
 sg13g2_decap_8 FILLER_29_2625 ();
 sg13g2_decap_8 FILLER_29_2632 ();
 sg13g2_decap_8 FILLER_29_2639 ();
 sg13g2_decap_8 FILLER_29_2646 ();
 sg13g2_decap_8 FILLER_29_2653 ();
 sg13g2_decap_8 FILLER_29_2660 ();
 sg13g2_fill_2 FILLER_29_2667 ();
 sg13g2_fill_1 FILLER_29_2669 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_fill_2 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_118 ();
 sg13g2_decap_8 FILLER_30_125 ();
 sg13g2_decap_8 FILLER_30_132 ();
 sg13g2_decap_8 FILLER_30_139 ();
 sg13g2_decap_8 FILLER_30_146 ();
 sg13g2_decap_4 FILLER_30_153 ();
 sg13g2_fill_1 FILLER_30_157 ();
 sg13g2_decap_8 FILLER_30_162 ();
 sg13g2_decap_8 FILLER_30_169 ();
 sg13g2_decap_8 FILLER_30_176 ();
 sg13g2_decap_8 FILLER_30_183 ();
 sg13g2_decap_8 FILLER_30_190 ();
 sg13g2_decap_8 FILLER_30_197 ();
 sg13g2_fill_1 FILLER_30_204 ();
 sg13g2_decap_8 FILLER_30_209 ();
 sg13g2_decap_8 FILLER_30_216 ();
 sg13g2_decap_8 FILLER_30_223 ();
 sg13g2_decap_8 FILLER_30_230 ();
 sg13g2_decap_8 FILLER_30_237 ();
 sg13g2_decap_8 FILLER_30_244 ();
 sg13g2_decap_8 FILLER_30_251 ();
 sg13g2_decap_8 FILLER_30_258 ();
 sg13g2_decap_8 FILLER_30_265 ();
 sg13g2_decap_8 FILLER_30_272 ();
 sg13g2_decap_8 FILLER_30_279 ();
 sg13g2_decap_8 FILLER_30_286 ();
 sg13g2_decap_8 FILLER_30_293 ();
 sg13g2_decap_8 FILLER_30_300 ();
 sg13g2_decap_8 FILLER_30_307 ();
 sg13g2_decap_8 FILLER_30_314 ();
 sg13g2_decap_8 FILLER_30_321 ();
 sg13g2_decap_8 FILLER_30_328 ();
 sg13g2_decap_8 FILLER_30_335 ();
 sg13g2_decap_8 FILLER_30_342 ();
 sg13g2_decap_8 FILLER_30_349 ();
 sg13g2_decap_8 FILLER_30_356 ();
 sg13g2_decap_8 FILLER_30_363 ();
 sg13g2_decap_8 FILLER_30_370 ();
 sg13g2_decap_8 FILLER_30_377 ();
 sg13g2_decap_8 FILLER_30_384 ();
 sg13g2_decap_8 FILLER_30_391 ();
 sg13g2_fill_1 FILLER_30_398 ();
 sg13g2_decap_8 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_30_414 ();
 sg13g2_decap_8 FILLER_30_421 ();
 sg13g2_decap_8 FILLER_30_428 ();
 sg13g2_decap_8 FILLER_30_435 ();
 sg13g2_decap_8 FILLER_30_442 ();
 sg13g2_decap_8 FILLER_30_449 ();
 sg13g2_decap_8 FILLER_30_456 ();
 sg13g2_decap_8 FILLER_30_463 ();
 sg13g2_decap_8 FILLER_30_470 ();
 sg13g2_decap_8 FILLER_30_477 ();
 sg13g2_decap_8 FILLER_30_484 ();
 sg13g2_decap_8 FILLER_30_496 ();
 sg13g2_decap_8 FILLER_30_503 ();
 sg13g2_decap_8 FILLER_30_510 ();
 sg13g2_decap_8 FILLER_30_517 ();
 sg13g2_decap_8 FILLER_30_524 ();
 sg13g2_decap_4 FILLER_30_531 ();
 sg13g2_fill_2 FILLER_30_535 ();
 sg13g2_decap_8 FILLER_30_542 ();
 sg13g2_decap_8 FILLER_30_549 ();
 sg13g2_decap_8 FILLER_30_556 ();
 sg13g2_decap_8 FILLER_30_563 ();
 sg13g2_decap_4 FILLER_30_570 ();
 sg13g2_decap_8 FILLER_30_589 ();
 sg13g2_decap_8 FILLER_30_596 ();
 sg13g2_decap_8 FILLER_30_603 ();
 sg13g2_decap_8 FILLER_30_610 ();
 sg13g2_decap_8 FILLER_30_617 ();
 sg13g2_decap_8 FILLER_30_624 ();
 sg13g2_decap_8 FILLER_30_631 ();
 sg13g2_decap_8 FILLER_30_638 ();
 sg13g2_decap_8 FILLER_30_645 ();
 sg13g2_decap_8 FILLER_30_652 ();
 sg13g2_decap_8 FILLER_30_659 ();
 sg13g2_decap_8 FILLER_30_666 ();
 sg13g2_fill_2 FILLER_30_673 ();
 sg13g2_decap_8 FILLER_30_681 ();
 sg13g2_decap_8 FILLER_30_688 ();
 sg13g2_decap_4 FILLER_30_695 ();
 sg13g2_fill_1 FILLER_30_699 ();
 sg13g2_decap_8 FILLER_30_704 ();
 sg13g2_decap_8 FILLER_30_711 ();
 sg13g2_decap_8 FILLER_30_718 ();
 sg13g2_decap_4 FILLER_30_725 ();
 sg13g2_fill_2 FILLER_30_729 ();
 sg13g2_decap_8 FILLER_30_736 ();
 sg13g2_decap_8 FILLER_30_743 ();
 sg13g2_decap_8 FILLER_30_750 ();
 sg13g2_decap_8 FILLER_30_757 ();
 sg13g2_decap_8 FILLER_30_764 ();
 sg13g2_decap_8 FILLER_30_771 ();
 sg13g2_decap_8 FILLER_30_778 ();
 sg13g2_decap_8 FILLER_30_785 ();
 sg13g2_decap_8 FILLER_30_792 ();
 sg13g2_decap_4 FILLER_30_799 ();
 sg13g2_fill_1 FILLER_30_803 ();
 sg13g2_decap_8 FILLER_30_807 ();
 sg13g2_decap_8 FILLER_30_814 ();
 sg13g2_fill_2 FILLER_30_821 ();
 sg13g2_decap_8 FILLER_30_827 ();
 sg13g2_decap_8 FILLER_30_834 ();
 sg13g2_decap_4 FILLER_30_841 ();
 sg13g2_fill_1 FILLER_30_845 ();
 sg13g2_decap_8 FILLER_30_850 ();
 sg13g2_decap_8 FILLER_30_860 ();
 sg13g2_decap_8 FILLER_30_867 ();
 sg13g2_decap_8 FILLER_30_874 ();
 sg13g2_decap_8 FILLER_30_881 ();
 sg13g2_decap_4 FILLER_30_888 ();
 sg13g2_fill_2 FILLER_30_892 ();
 sg13g2_fill_1 FILLER_30_901 ();
 sg13g2_fill_1 FILLER_30_906 ();
 sg13g2_decap_8 FILLER_30_920 ();
 sg13g2_decap_4 FILLER_30_927 ();
 sg13g2_fill_1 FILLER_30_931 ();
 sg13g2_decap_8 FILLER_30_935 ();
 sg13g2_decap_8 FILLER_30_942 ();
 sg13g2_fill_2 FILLER_30_949 ();
 sg13g2_decap_8 FILLER_30_958 ();
 sg13g2_decap_8 FILLER_30_965 ();
 sg13g2_decap_8 FILLER_30_972 ();
 sg13g2_decap_8 FILLER_30_979 ();
 sg13g2_decap_8 FILLER_30_986 ();
 sg13g2_decap_8 FILLER_30_993 ();
 sg13g2_decap_8 FILLER_30_1000 ();
 sg13g2_decap_8 FILLER_30_1007 ();
 sg13g2_decap_8 FILLER_30_1014 ();
 sg13g2_decap_8 FILLER_30_1021 ();
 sg13g2_decap_8 FILLER_30_1028 ();
 sg13g2_fill_2 FILLER_30_1035 ();
 sg13g2_fill_1 FILLER_30_1037 ();
 sg13g2_decap_8 FILLER_30_1049 ();
 sg13g2_decap_4 FILLER_30_1056 ();
 sg13g2_fill_2 FILLER_30_1060 ();
 sg13g2_fill_1 FILLER_30_1085 ();
 sg13g2_decap_8 FILLER_30_1098 ();
 sg13g2_decap_8 FILLER_30_1105 ();
 sg13g2_decap_8 FILLER_30_1112 ();
 sg13g2_decap_8 FILLER_30_1119 ();
 sg13g2_decap_8 FILLER_30_1126 ();
 sg13g2_decap_8 FILLER_30_1133 ();
 sg13g2_decap_8 FILLER_30_1140 ();
 sg13g2_decap_8 FILLER_30_1147 ();
 sg13g2_decap_8 FILLER_30_1154 ();
 sg13g2_decap_8 FILLER_30_1161 ();
 sg13g2_fill_2 FILLER_30_1168 ();
 sg13g2_fill_1 FILLER_30_1170 ();
 sg13g2_decap_8 FILLER_30_1185 ();
 sg13g2_decap_8 FILLER_30_1192 ();
 sg13g2_decap_8 FILLER_30_1199 ();
 sg13g2_decap_8 FILLER_30_1206 ();
 sg13g2_decap_8 FILLER_30_1213 ();
 sg13g2_decap_8 FILLER_30_1220 ();
 sg13g2_decap_8 FILLER_30_1227 ();
 sg13g2_fill_2 FILLER_30_1234 ();
 sg13g2_fill_1 FILLER_30_1236 ();
 sg13g2_decap_8 FILLER_30_1242 ();
 sg13g2_decap_8 FILLER_30_1249 ();
 sg13g2_decap_8 FILLER_30_1256 ();
 sg13g2_decap_8 FILLER_30_1263 ();
 sg13g2_decap_8 FILLER_30_1270 ();
 sg13g2_fill_1 FILLER_30_1277 ();
 sg13g2_decap_8 FILLER_30_1282 ();
 sg13g2_decap_8 FILLER_30_1289 ();
 sg13g2_decap_8 FILLER_30_1296 ();
 sg13g2_fill_2 FILLER_30_1303 ();
 sg13g2_fill_1 FILLER_30_1305 ();
 sg13g2_decap_8 FILLER_30_1315 ();
 sg13g2_decap_8 FILLER_30_1322 ();
 sg13g2_decap_8 FILLER_30_1329 ();
 sg13g2_decap_8 FILLER_30_1336 ();
 sg13g2_decap_4 FILLER_30_1343 ();
 sg13g2_decap_8 FILLER_30_1351 ();
 sg13g2_decap_8 FILLER_30_1358 ();
 sg13g2_decap_8 FILLER_30_1365 ();
 sg13g2_decap_8 FILLER_30_1372 ();
 sg13g2_decap_8 FILLER_30_1379 ();
 sg13g2_decap_8 FILLER_30_1386 ();
 sg13g2_decap_8 FILLER_30_1393 ();
 sg13g2_decap_8 FILLER_30_1400 ();
 sg13g2_decap_8 FILLER_30_1407 ();
 sg13g2_decap_8 FILLER_30_1414 ();
 sg13g2_decap_8 FILLER_30_1421 ();
 sg13g2_decap_8 FILLER_30_1428 ();
 sg13g2_decap_8 FILLER_30_1435 ();
 sg13g2_decap_8 FILLER_30_1442 ();
 sg13g2_decap_8 FILLER_30_1449 ();
 sg13g2_decap_8 FILLER_30_1456 ();
 sg13g2_decap_8 FILLER_30_1463 ();
 sg13g2_decap_8 FILLER_30_1470 ();
 sg13g2_decap_8 FILLER_30_1477 ();
 sg13g2_decap_8 FILLER_30_1484 ();
 sg13g2_decap_8 FILLER_30_1491 ();
 sg13g2_decap_8 FILLER_30_1498 ();
 sg13g2_decap_4 FILLER_30_1505 ();
 sg13g2_decap_8 FILLER_30_1513 ();
 sg13g2_decap_4 FILLER_30_1539 ();
 sg13g2_fill_2 FILLER_30_1543 ();
 sg13g2_decap_4 FILLER_30_1548 ();
 sg13g2_fill_2 FILLER_30_1552 ();
 sg13g2_fill_1 FILLER_30_1565 ();
 sg13g2_fill_1 FILLER_30_1595 ();
 sg13g2_decap_4 FILLER_30_1601 ();
 sg13g2_fill_2 FILLER_30_1605 ();
 sg13g2_decap_4 FILLER_30_1619 ();
 sg13g2_fill_1 FILLER_30_1623 ();
 sg13g2_decap_8 FILLER_30_1644 ();
 sg13g2_decap_4 FILLER_30_1651 ();
 sg13g2_decap_8 FILLER_30_1659 ();
 sg13g2_decap_8 FILLER_30_1666 ();
 sg13g2_decap_8 FILLER_30_1673 ();
 sg13g2_decap_8 FILLER_30_1680 ();
 sg13g2_decap_8 FILLER_30_1687 ();
 sg13g2_decap_8 FILLER_30_1694 ();
 sg13g2_decap_8 FILLER_30_1705 ();
 sg13g2_decap_8 FILLER_30_1712 ();
 sg13g2_fill_2 FILLER_30_1719 ();
 sg13g2_fill_1 FILLER_30_1721 ();
 sg13g2_decap_8 FILLER_30_1728 ();
 sg13g2_fill_1 FILLER_30_1735 ();
 sg13g2_fill_1 FILLER_30_1740 ();
 sg13g2_decap_8 FILLER_30_1746 ();
 sg13g2_decap_8 FILLER_30_1753 ();
 sg13g2_decap_8 FILLER_30_1760 ();
 sg13g2_decap_8 FILLER_30_1767 ();
 sg13g2_decap_4 FILLER_30_1774 ();
 sg13g2_fill_2 FILLER_30_1778 ();
 sg13g2_decap_8 FILLER_30_1786 ();
 sg13g2_decap_8 FILLER_30_1793 ();
 sg13g2_decap_8 FILLER_30_1800 ();
 sg13g2_decap_8 FILLER_30_1807 ();
 sg13g2_fill_1 FILLER_30_1814 ();
 sg13g2_fill_2 FILLER_30_1820 ();
 sg13g2_decap_8 FILLER_30_1826 ();
 sg13g2_decap_8 FILLER_30_1833 ();
 sg13g2_decap_8 FILLER_30_1840 ();
 sg13g2_decap_8 FILLER_30_1847 ();
 sg13g2_decap_8 FILLER_30_1854 ();
 sg13g2_decap_8 FILLER_30_1867 ();
 sg13g2_decap_8 FILLER_30_1874 ();
 sg13g2_decap_8 FILLER_30_1881 ();
 sg13g2_decap_8 FILLER_30_1888 ();
 sg13g2_decap_8 FILLER_30_1895 ();
 sg13g2_decap_8 FILLER_30_1902 ();
 sg13g2_decap_8 FILLER_30_1909 ();
 sg13g2_decap_8 FILLER_30_1916 ();
 sg13g2_decap_8 FILLER_30_1923 ();
 sg13g2_decap_8 FILLER_30_1930 ();
 sg13g2_decap_8 FILLER_30_1937 ();
 sg13g2_decap_8 FILLER_30_1944 ();
 sg13g2_decap_8 FILLER_30_1951 ();
 sg13g2_decap_8 FILLER_30_1958 ();
 sg13g2_decap_8 FILLER_30_1965 ();
 sg13g2_decap_8 FILLER_30_1972 ();
 sg13g2_decap_8 FILLER_30_1979 ();
 sg13g2_decap_8 FILLER_30_1986 ();
 sg13g2_decap_8 FILLER_30_1993 ();
 sg13g2_decap_8 FILLER_30_2000 ();
 sg13g2_decap_8 FILLER_30_2007 ();
 sg13g2_decap_8 FILLER_30_2014 ();
 sg13g2_decap_8 FILLER_30_2021 ();
 sg13g2_decap_8 FILLER_30_2028 ();
 sg13g2_decap_8 FILLER_30_2035 ();
 sg13g2_decap_8 FILLER_30_2042 ();
 sg13g2_decap_8 FILLER_30_2049 ();
 sg13g2_decap_8 FILLER_30_2056 ();
 sg13g2_decap_8 FILLER_30_2063 ();
 sg13g2_decap_8 FILLER_30_2070 ();
 sg13g2_decap_8 FILLER_30_2077 ();
 sg13g2_decap_8 FILLER_30_2084 ();
 sg13g2_decap_8 FILLER_30_2091 ();
 sg13g2_decap_8 FILLER_30_2098 ();
 sg13g2_decap_8 FILLER_30_2105 ();
 sg13g2_decap_8 FILLER_30_2112 ();
 sg13g2_decap_8 FILLER_30_2119 ();
 sg13g2_decap_8 FILLER_30_2126 ();
 sg13g2_decap_8 FILLER_30_2133 ();
 sg13g2_decap_8 FILLER_30_2140 ();
 sg13g2_decap_8 FILLER_30_2147 ();
 sg13g2_decap_8 FILLER_30_2154 ();
 sg13g2_decap_8 FILLER_30_2161 ();
 sg13g2_decap_8 FILLER_30_2168 ();
 sg13g2_decap_8 FILLER_30_2175 ();
 sg13g2_decap_8 FILLER_30_2182 ();
 sg13g2_decap_8 FILLER_30_2189 ();
 sg13g2_decap_8 FILLER_30_2196 ();
 sg13g2_decap_8 FILLER_30_2203 ();
 sg13g2_decap_8 FILLER_30_2210 ();
 sg13g2_decap_8 FILLER_30_2217 ();
 sg13g2_decap_8 FILLER_30_2224 ();
 sg13g2_decap_8 FILLER_30_2231 ();
 sg13g2_decap_8 FILLER_30_2238 ();
 sg13g2_decap_8 FILLER_30_2245 ();
 sg13g2_decap_8 FILLER_30_2252 ();
 sg13g2_decap_8 FILLER_30_2259 ();
 sg13g2_decap_8 FILLER_30_2266 ();
 sg13g2_decap_8 FILLER_30_2273 ();
 sg13g2_decap_8 FILLER_30_2280 ();
 sg13g2_decap_8 FILLER_30_2287 ();
 sg13g2_decap_8 FILLER_30_2294 ();
 sg13g2_decap_8 FILLER_30_2301 ();
 sg13g2_decap_8 FILLER_30_2308 ();
 sg13g2_decap_8 FILLER_30_2315 ();
 sg13g2_decap_8 FILLER_30_2322 ();
 sg13g2_decap_8 FILLER_30_2329 ();
 sg13g2_decap_8 FILLER_30_2336 ();
 sg13g2_decap_8 FILLER_30_2343 ();
 sg13g2_decap_8 FILLER_30_2350 ();
 sg13g2_decap_8 FILLER_30_2357 ();
 sg13g2_decap_8 FILLER_30_2364 ();
 sg13g2_decap_8 FILLER_30_2371 ();
 sg13g2_decap_8 FILLER_30_2378 ();
 sg13g2_decap_8 FILLER_30_2385 ();
 sg13g2_decap_8 FILLER_30_2392 ();
 sg13g2_decap_8 FILLER_30_2399 ();
 sg13g2_decap_8 FILLER_30_2406 ();
 sg13g2_decap_8 FILLER_30_2413 ();
 sg13g2_decap_8 FILLER_30_2420 ();
 sg13g2_decap_8 FILLER_30_2427 ();
 sg13g2_decap_8 FILLER_30_2434 ();
 sg13g2_decap_8 FILLER_30_2441 ();
 sg13g2_decap_8 FILLER_30_2448 ();
 sg13g2_decap_8 FILLER_30_2455 ();
 sg13g2_decap_8 FILLER_30_2462 ();
 sg13g2_decap_8 FILLER_30_2469 ();
 sg13g2_decap_8 FILLER_30_2476 ();
 sg13g2_decap_8 FILLER_30_2483 ();
 sg13g2_decap_8 FILLER_30_2490 ();
 sg13g2_decap_8 FILLER_30_2497 ();
 sg13g2_decap_8 FILLER_30_2504 ();
 sg13g2_decap_8 FILLER_30_2511 ();
 sg13g2_decap_8 FILLER_30_2518 ();
 sg13g2_decap_8 FILLER_30_2525 ();
 sg13g2_decap_8 FILLER_30_2532 ();
 sg13g2_decap_8 FILLER_30_2539 ();
 sg13g2_decap_8 FILLER_30_2546 ();
 sg13g2_decap_8 FILLER_30_2553 ();
 sg13g2_decap_8 FILLER_30_2560 ();
 sg13g2_decap_8 FILLER_30_2567 ();
 sg13g2_decap_8 FILLER_30_2574 ();
 sg13g2_decap_8 FILLER_30_2581 ();
 sg13g2_decap_8 FILLER_30_2588 ();
 sg13g2_decap_8 FILLER_30_2595 ();
 sg13g2_decap_8 FILLER_30_2602 ();
 sg13g2_decap_8 FILLER_30_2609 ();
 sg13g2_decap_8 FILLER_30_2616 ();
 sg13g2_decap_8 FILLER_30_2623 ();
 sg13g2_decap_8 FILLER_30_2630 ();
 sg13g2_decap_8 FILLER_30_2637 ();
 sg13g2_decap_8 FILLER_30_2644 ();
 sg13g2_decap_8 FILLER_30_2651 ();
 sg13g2_decap_8 FILLER_30_2658 ();
 sg13g2_decap_4 FILLER_30_2665 ();
 sg13g2_fill_1 FILLER_30_2669 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_fill_2 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_decap_8 FILLER_31_182 ();
 sg13g2_decap_8 FILLER_31_189 ();
 sg13g2_decap_8 FILLER_31_196 ();
 sg13g2_decap_8 FILLER_31_203 ();
 sg13g2_decap_8 FILLER_31_210 ();
 sg13g2_decap_8 FILLER_31_217 ();
 sg13g2_decap_8 FILLER_31_224 ();
 sg13g2_decap_8 FILLER_31_231 ();
 sg13g2_decap_8 FILLER_31_238 ();
 sg13g2_decap_8 FILLER_31_245 ();
 sg13g2_decap_8 FILLER_31_252 ();
 sg13g2_decap_8 FILLER_31_259 ();
 sg13g2_decap_8 FILLER_31_266 ();
 sg13g2_decap_8 FILLER_31_273 ();
 sg13g2_decap_8 FILLER_31_280 ();
 sg13g2_decap_4 FILLER_31_287 ();
 sg13g2_fill_1 FILLER_31_291 ();
 sg13g2_decap_8 FILLER_31_296 ();
 sg13g2_decap_8 FILLER_31_303 ();
 sg13g2_decap_8 FILLER_31_310 ();
 sg13g2_decap_8 FILLER_31_317 ();
 sg13g2_decap_8 FILLER_31_324 ();
 sg13g2_decap_8 FILLER_31_331 ();
 sg13g2_decap_8 FILLER_31_338 ();
 sg13g2_decap_8 FILLER_31_345 ();
 sg13g2_decap_8 FILLER_31_352 ();
 sg13g2_decap_8 FILLER_31_359 ();
 sg13g2_decap_8 FILLER_31_366 ();
 sg13g2_decap_8 FILLER_31_373 ();
 sg13g2_fill_2 FILLER_31_380 ();
 sg13g2_fill_1 FILLER_31_382 ();
 sg13g2_decap_8 FILLER_31_388 ();
 sg13g2_decap_8 FILLER_31_395 ();
 sg13g2_decap_8 FILLER_31_402 ();
 sg13g2_decap_8 FILLER_31_409 ();
 sg13g2_decap_8 FILLER_31_416 ();
 sg13g2_decap_8 FILLER_31_423 ();
 sg13g2_decap_8 FILLER_31_430 ();
 sg13g2_decap_8 FILLER_31_437 ();
 sg13g2_decap_8 FILLER_31_444 ();
 sg13g2_decap_8 FILLER_31_451 ();
 sg13g2_decap_8 FILLER_31_458 ();
 sg13g2_decap_8 FILLER_31_465 ();
 sg13g2_decap_8 FILLER_31_472 ();
 sg13g2_decap_4 FILLER_31_479 ();
 sg13g2_fill_2 FILLER_31_483 ();
 sg13g2_decap_8 FILLER_31_490 ();
 sg13g2_decap_8 FILLER_31_497 ();
 sg13g2_decap_8 FILLER_31_504 ();
 sg13g2_decap_8 FILLER_31_511 ();
 sg13g2_fill_1 FILLER_31_518 ();
 sg13g2_decap_8 FILLER_31_534 ();
 sg13g2_decap_8 FILLER_31_541 ();
 sg13g2_decap_8 FILLER_31_548 ();
 sg13g2_decap_8 FILLER_31_555 ();
 sg13g2_decap_8 FILLER_31_562 ();
 sg13g2_fill_2 FILLER_31_569 ();
 sg13g2_fill_1 FILLER_31_580 ();
 sg13g2_decap_8 FILLER_31_593 ();
 sg13g2_decap_4 FILLER_31_600 ();
 sg13g2_fill_2 FILLER_31_604 ();
 sg13g2_decap_8 FILLER_31_611 ();
 sg13g2_decap_8 FILLER_31_618 ();
 sg13g2_decap_8 FILLER_31_625 ();
 sg13g2_decap_8 FILLER_31_632 ();
 sg13g2_decap_4 FILLER_31_639 ();
 sg13g2_fill_2 FILLER_31_643 ();
 sg13g2_decap_8 FILLER_31_650 ();
 sg13g2_decap_8 FILLER_31_657 ();
 sg13g2_decap_4 FILLER_31_664 ();
 sg13g2_fill_1 FILLER_31_668 ();
 sg13g2_fill_1 FILLER_31_674 ();
 sg13g2_decap_8 FILLER_31_693 ();
 sg13g2_decap_8 FILLER_31_700 ();
 sg13g2_decap_4 FILLER_31_707 ();
 sg13g2_fill_1 FILLER_31_711 ();
 sg13g2_fill_2 FILLER_31_727 ();
 sg13g2_decap_8 FILLER_31_734 ();
 sg13g2_decap_8 FILLER_31_741 ();
 sg13g2_decap_8 FILLER_31_748 ();
 sg13g2_decap_8 FILLER_31_755 ();
 sg13g2_decap_8 FILLER_31_762 ();
 sg13g2_decap_8 FILLER_31_769 ();
 sg13g2_decap_8 FILLER_31_776 ();
 sg13g2_fill_1 FILLER_31_783 ();
 sg13g2_decap_8 FILLER_31_793 ();
 sg13g2_decap_4 FILLER_31_800 ();
 sg13g2_decap_8 FILLER_31_808 ();
 sg13g2_decap_8 FILLER_31_815 ();
 sg13g2_decap_8 FILLER_31_822 ();
 sg13g2_decap_8 FILLER_31_829 ();
 sg13g2_decap_8 FILLER_31_836 ();
 sg13g2_decap_8 FILLER_31_843 ();
 sg13g2_decap_8 FILLER_31_850 ();
 sg13g2_fill_2 FILLER_31_861 ();
 sg13g2_fill_1 FILLER_31_863 ();
 sg13g2_decap_8 FILLER_31_868 ();
 sg13g2_fill_2 FILLER_31_875 ();
 sg13g2_decap_8 FILLER_31_882 ();
 sg13g2_decap_8 FILLER_31_889 ();
 sg13g2_decap_8 FILLER_31_896 ();
 sg13g2_decap_8 FILLER_31_903 ();
 sg13g2_fill_1 FILLER_31_922 ();
 sg13g2_decap_8 FILLER_31_926 ();
 sg13g2_decap_8 FILLER_31_933 ();
 sg13g2_decap_8 FILLER_31_940 ();
 sg13g2_fill_1 FILLER_31_947 ();
 sg13g2_decap_8 FILLER_31_956 ();
 sg13g2_decap_8 FILLER_31_963 ();
 sg13g2_decap_8 FILLER_31_970 ();
 sg13g2_decap_4 FILLER_31_977 ();
 sg13g2_fill_1 FILLER_31_981 ();
 sg13g2_decap_8 FILLER_31_986 ();
 sg13g2_decap_8 FILLER_31_993 ();
 sg13g2_decap_8 FILLER_31_1000 ();
 sg13g2_decap_4 FILLER_31_1007 ();
 sg13g2_fill_1 FILLER_31_1011 ();
 sg13g2_decap_8 FILLER_31_1015 ();
 sg13g2_decap_8 FILLER_31_1022 ();
 sg13g2_decap_8 FILLER_31_1029 ();
 sg13g2_fill_1 FILLER_31_1036 ();
 sg13g2_fill_2 FILLER_31_1042 ();
 sg13g2_decap_8 FILLER_31_1050 ();
 sg13g2_decap_8 FILLER_31_1057 ();
 sg13g2_decap_8 FILLER_31_1064 ();
 sg13g2_decap_8 FILLER_31_1092 ();
 sg13g2_decap_8 FILLER_31_1099 ();
 sg13g2_decap_8 FILLER_31_1106 ();
 sg13g2_decap_8 FILLER_31_1113 ();
 sg13g2_decap_4 FILLER_31_1120 ();
 sg13g2_fill_1 FILLER_31_1124 ();
 sg13g2_fill_2 FILLER_31_1134 ();
 sg13g2_decap_8 FILLER_31_1149 ();
 sg13g2_fill_1 FILLER_31_1156 ();
 sg13g2_decap_8 FILLER_31_1163 ();
 sg13g2_decap_8 FILLER_31_1170 ();
 sg13g2_fill_2 FILLER_31_1180 ();
 sg13g2_fill_1 FILLER_31_1182 ();
 sg13g2_decap_8 FILLER_31_1198 ();
 sg13g2_decap_8 FILLER_31_1205 ();
 sg13g2_decap_8 FILLER_31_1212 ();
 sg13g2_decap_8 FILLER_31_1219 ();
 sg13g2_decap_4 FILLER_31_1226 ();
 sg13g2_fill_2 FILLER_31_1230 ();
 sg13g2_decap_8 FILLER_31_1241 ();
 sg13g2_decap_8 FILLER_31_1248 ();
 sg13g2_decap_8 FILLER_31_1255 ();
 sg13g2_decap_8 FILLER_31_1262 ();
 sg13g2_decap_8 FILLER_31_1269 ();
 sg13g2_decap_8 FILLER_31_1276 ();
 sg13g2_decap_8 FILLER_31_1283 ();
 sg13g2_decap_8 FILLER_31_1290 ();
 sg13g2_decap_8 FILLER_31_1297 ();
 sg13g2_decap_8 FILLER_31_1304 ();
 sg13g2_decap_8 FILLER_31_1311 ();
 sg13g2_decap_8 FILLER_31_1318 ();
 sg13g2_decap_8 FILLER_31_1325 ();
 sg13g2_decap_8 FILLER_31_1332 ();
 sg13g2_decap_8 FILLER_31_1339 ();
 sg13g2_decap_4 FILLER_31_1346 ();
 sg13g2_decap_8 FILLER_31_1356 ();
 sg13g2_decap_8 FILLER_31_1363 ();
 sg13g2_decap_8 FILLER_31_1370 ();
 sg13g2_decap_4 FILLER_31_1377 ();
 sg13g2_fill_1 FILLER_31_1381 ();
 sg13g2_decap_4 FILLER_31_1389 ();
 sg13g2_fill_1 FILLER_31_1393 ();
 sg13g2_decap_8 FILLER_31_1398 ();
 sg13g2_decap_8 FILLER_31_1405 ();
 sg13g2_decap_8 FILLER_31_1412 ();
 sg13g2_decap_8 FILLER_31_1419 ();
 sg13g2_fill_1 FILLER_31_1426 ();
 sg13g2_decap_8 FILLER_31_1431 ();
 sg13g2_fill_1 FILLER_31_1438 ();
 sg13g2_fill_1 FILLER_31_1443 ();
 sg13g2_decap_4 FILLER_31_1448 ();
 sg13g2_fill_2 FILLER_31_1452 ();
 sg13g2_decap_8 FILLER_31_1460 ();
 sg13g2_fill_2 FILLER_31_1467 ();
 sg13g2_decap_8 FILLER_31_1484 ();
 sg13g2_decap_8 FILLER_31_1491 ();
 sg13g2_decap_8 FILLER_31_1498 ();
 sg13g2_fill_1 FILLER_31_1505 ();
 sg13g2_decap_8 FILLER_31_1511 ();
 sg13g2_fill_2 FILLER_31_1518 ();
 sg13g2_decap_8 FILLER_31_1524 ();
 sg13g2_decap_8 FILLER_31_1531 ();
 sg13g2_fill_1 FILLER_31_1538 ();
 sg13g2_fill_2 FILLER_31_1559 ();
 sg13g2_fill_1 FILLER_31_1561 ();
 sg13g2_fill_2 FILLER_31_1574 ();
 sg13g2_fill_1 FILLER_31_1576 ();
 sg13g2_decap_8 FILLER_31_1589 ();
 sg13g2_decap_8 FILLER_31_1596 ();
 sg13g2_decap_8 FILLER_31_1603 ();
 sg13g2_decap_8 FILLER_31_1610 ();
 sg13g2_decap_8 FILLER_31_1617 ();
 sg13g2_decap_8 FILLER_31_1632 ();
 sg13g2_decap_8 FILLER_31_1639 ();
 sg13g2_decap_8 FILLER_31_1665 ();
 sg13g2_decap_8 FILLER_31_1672 ();
 sg13g2_decap_8 FILLER_31_1679 ();
 sg13g2_decap_8 FILLER_31_1686 ();
 sg13g2_decap_8 FILLER_31_1698 ();
 sg13g2_decap_8 FILLER_31_1705 ();
 sg13g2_decap_8 FILLER_31_1712 ();
 sg13g2_decap_8 FILLER_31_1719 ();
 sg13g2_fill_2 FILLER_31_1726 ();
 sg13g2_decap_8 FILLER_31_1736 ();
 sg13g2_decap_8 FILLER_31_1743 ();
 sg13g2_decap_8 FILLER_31_1750 ();
 sg13g2_decap_8 FILLER_31_1757 ();
 sg13g2_decap_8 FILLER_31_1764 ();
 sg13g2_decap_8 FILLER_31_1771 ();
 sg13g2_decap_8 FILLER_31_1778 ();
 sg13g2_decap_8 FILLER_31_1785 ();
 sg13g2_decap_8 FILLER_31_1792 ();
 sg13g2_decap_8 FILLER_31_1799 ();
 sg13g2_decap_8 FILLER_31_1806 ();
 sg13g2_decap_8 FILLER_31_1813 ();
 sg13g2_decap_8 FILLER_31_1820 ();
 sg13g2_decap_8 FILLER_31_1827 ();
 sg13g2_decap_8 FILLER_31_1834 ();
 sg13g2_decap_8 FILLER_31_1841 ();
 sg13g2_decap_8 FILLER_31_1848 ();
 sg13g2_decap_8 FILLER_31_1855 ();
 sg13g2_decap_8 FILLER_31_1862 ();
 sg13g2_decap_8 FILLER_31_1869 ();
 sg13g2_decap_8 FILLER_31_1876 ();
 sg13g2_decap_8 FILLER_31_1883 ();
 sg13g2_decap_8 FILLER_31_1890 ();
 sg13g2_decap_8 FILLER_31_1897 ();
 sg13g2_decap_8 FILLER_31_1904 ();
 sg13g2_decap_8 FILLER_31_1911 ();
 sg13g2_decap_8 FILLER_31_1918 ();
 sg13g2_decap_8 FILLER_31_1925 ();
 sg13g2_decap_8 FILLER_31_1932 ();
 sg13g2_decap_8 FILLER_31_1939 ();
 sg13g2_decap_8 FILLER_31_1946 ();
 sg13g2_decap_8 FILLER_31_1953 ();
 sg13g2_decap_8 FILLER_31_1960 ();
 sg13g2_decap_8 FILLER_31_1967 ();
 sg13g2_decap_8 FILLER_31_1974 ();
 sg13g2_decap_8 FILLER_31_1981 ();
 sg13g2_decap_8 FILLER_31_1988 ();
 sg13g2_decap_8 FILLER_31_1995 ();
 sg13g2_decap_8 FILLER_31_2002 ();
 sg13g2_decap_8 FILLER_31_2009 ();
 sg13g2_decap_8 FILLER_31_2016 ();
 sg13g2_decap_8 FILLER_31_2023 ();
 sg13g2_decap_8 FILLER_31_2030 ();
 sg13g2_decap_8 FILLER_31_2037 ();
 sg13g2_decap_8 FILLER_31_2044 ();
 sg13g2_decap_8 FILLER_31_2051 ();
 sg13g2_decap_8 FILLER_31_2058 ();
 sg13g2_decap_8 FILLER_31_2065 ();
 sg13g2_decap_8 FILLER_31_2072 ();
 sg13g2_decap_8 FILLER_31_2079 ();
 sg13g2_decap_8 FILLER_31_2086 ();
 sg13g2_decap_8 FILLER_31_2093 ();
 sg13g2_decap_8 FILLER_31_2100 ();
 sg13g2_decap_8 FILLER_31_2107 ();
 sg13g2_decap_8 FILLER_31_2114 ();
 sg13g2_decap_8 FILLER_31_2121 ();
 sg13g2_decap_8 FILLER_31_2128 ();
 sg13g2_decap_8 FILLER_31_2135 ();
 sg13g2_decap_8 FILLER_31_2142 ();
 sg13g2_decap_8 FILLER_31_2149 ();
 sg13g2_decap_8 FILLER_31_2156 ();
 sg13g2_decap_8 FILLER_31_2163 ();
 sg13g2_decap_8 FILLER_31_2170 ();
 sg13g2_decap_8 FILLER_31_2177 ();
 sg13g2_decap_8 FILLER_31_2184 ();
 sg13g2_decap_8 FILLER_31_2191 ();
 sg13g2_decap_8 FILLER_31_2198 ();
 sg13g2_decap_8 FILLER_31_2205 ();
 sg13g2_decap_8 FILLER_31_2212 ();
 sg13g2_decap_8 FILLER_31_2219 ();
 sg13g2_decap_8 FILLER_31_2226 ();
 sg13g2_decap_8 FILLER_31_2233 ();
 sg13g2_decap_8 FILLER_31_2240 ();
 sg13g2_decap_8 FILLER_31_2247 ();
 sg13g2_decap_8 FILLER_31_2254 ();
 sg13g2_decap_8 FILLER_31_2261 ();
 sg13g2_decap_8 FILLER_31_2268 ();
 sg13g2_decap_8 FILLER_31_2275 ();
 sg13g2_decap_8 FILLER_31_2282 ();
 sg13g2_decap_8 FILLER_31_2289 ();
 sg13g2_decap_8 FILLER_31_2296 ();
 sg13g2_decap_8 FILLER_31_2303 ();
 sg13g2_decap_8 FILLER_31_2310 ();
 sg13g2_decap_8 FILLER_31_2317 ();
 sg13g2_decap_8 FILLER_31_2324 ();
 sg13g2_decap_8 FILLER_31_2331 ();
 sg13g2_decap_8 FILLER_31_2338 ();
 sg13g2_decap_8 FILLER_31_2345 ();
 sg13g2_decap_8 FILLER_31_2352 ();
 sg13g2_decap_8 FILLER_31_2359 ();
 sg13g2_decap_8 FILLER_31_2366 ();
 sg13g2_decap_8 FILLER_31_2373 ();
 sg13g2_decap_8 FILLER_31_2380 ();
 sg13g2_decap_8 FILLER_31_2387 ();
 sg13g2_decap_8 FILLER_31_2394 ();
 sg13g2_decap_8 FILLER_31_2401 ();
 sg13g2_decap_8 FILLER_31_2408 ();
 sg13g2_decap_8 FILLER_31_2415 ();
 sg13g2_decap_8 FILLER_31_2422 ();
 sg13g2_decap_8 FILLER_31_2429 ();
 sg13g2_decap_8 FILLER_31_2436 ();
 sg13g2_decap_8 FILLER_31_2443 ();
 sg13g2_decap_8 FILLER_31_2450 ();
 sg13g2_decap_8 FILLER_31_2457 ();
 sg13g2_decap_8 FILLER_31_2464 ();
 sg13g2_decap_8 FILLER_31_2471 ();
 sg13g2_decap_8 FILLER_31_2478 ();
 sg13g2_decap_8 FILLER_31_2485 ();
 sg13g2_decap_8 FILLER_31_2492 ();
 sg13g2_decap_8 FILLER_31_2499 ();
 sg13g2_decap_8 FILLER_31_2506 ();
 sg13g2_decap_8 FILLER_31_2513 ();
 sg13g2_decap_8 FILLER_31_2520 ();
 sg13g2_decap_8 FILLER_31_2527 ();
 sg13g2_decap_8 FILLER_31_2534 ();
 sg13g2_decap_8 FILLER_31_2541 ();
 sg13g2_decap_8 FILLER_31_2548 ();
 sg13g2_decap_8 FILLER_31_2555 ();
 sg13g2_decap_8 FILLER_31_2562 ();
 sg13g2_decap_8 FILLER_31_2569 ();
 sg13g2_decap_8 FILLER_31_2576 ();
 sg13g2_decap_8 FILLER_31_2583 ();
 sg13g2_decap_8 FILLER_31_2590 ();
 sg13g2_decap_8 FILLER_31_2597 ();
 sg13g2_decap_8 FILLER_31_2604 ();
 sg13g2_decap_8 FILLER_31_2611 ();
 sg13g2_decap_8 FILLER_31_2618 ();
 sg13g2_decap_8 FILLER_31_2625 ();
 sg13g2_decap_8 FILLER_31_2632 ();
 sg13g2_decap_8 FILLER_31_2639 ();
 sg13g2_decap_8 FILLER_31_2646 ();
 sg13g2_decap_8 FILLER_31_2653 ();
 sg13g2_decap_8 FILLER_31_2660 ();
 sg13g2_fill_2 FILLER_31_2667 ();
 sg13g2_fill_1 FILLER_31_2669 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_103 ();
 sg13g2_decap_8 FILLER_32_110 ();
 sg13g2_decap_8 FILLER_32_117 ();
 sg13g2_decap_8 FILLER_32_124 ();
 sg13g2_decap_8 FILLER_32_131 ();
 sg13g2_decap_8 FILLER_32_138 ();
 sg13g2_decap_8 FILLER_32_145 ();
 sg13g2_decap_8 FILLER_32_152 ();
 sg13g2_decap_8 FILLER_32_159 ();
 sg13g2_decap_8 FILLER_32_166 ();
 sg13g2_decap_8 FILLER_32_173 ();
 sg13g2_decap_8 FILLER_32_180 ();
 sg13g2_decap_8 FILLER_32_187 ();
 sg13g2_decap_8 FILLER_32_194 ();
 sg13g2_decap_8 FILLER_32_201 ();
 sg13g2_decap_8 FILLER_32_208 ();
 sg13g2_decap_8 FILLER_32_215 ();
 sg13g2_decap_8 FILLER_32_222 ();
 sg13g2_decap_8 FILLER_32_229 ();
 sg13g2_decap_8 FILLER_32_236 ();
 sg13g2_decap_8 FILLER_32_243 ();
 sg13g2_decap_8 FILLER_32_250 ();
 sg13g2_decap_8 FILLER_32_257 ();
 sg13g2_decap_4 FILLER_32_264 ();
 sg13g2_fill_1 FILLER_32_268 ();
 sg13g2_decap_8 FILLER_32_274 ();
 sg13g2_decap_4 FILLER_32_281 ();
 sg13g2_decap_8 FILLER_32_311 ();
 sg13g2_decap_8 FILLER_32_318 ();
 sg13g2_decap_8 FILLER_32_325 ();
 sg13g2_decap_8 FILLER_32_332 ();
 sg13g2_decap_8 FILLER_32_339 ();
 sg13g2_decap_8 FILLER_32_346 ();
 sg13g2_decap_4 FILLER_32_353 ();
 sg13g2_decap_8 FILLER_32_365 ();
 sg13g2_decap_8 FILLER_32_372 ();
 sg13g2_decap_8 FILLER_32_379 ();
 sg13g2_decap_8 FILLER_32_386 ();
 sg13g2_fill_1 FILLER_32_393 ();
 sg13g2_decap_8 FILLER_32_402 ();
 sg13g2_decap_8 FILLER_32_409 ();
 sg13g2_decap_8 FILLER_32_416 ();
 sg13g2_decap_8 FILLER_32_423 ();
 sg13g2_decap_8 FILLER_32_430 ();
 sg13g2_decap_8 FILLER_32_437 ();
 sg13g2_decap_8 FILLER_32_444 ();
 sg13g2_decap_8 FILLER_32_451 ();
 sg13g2_decap_8 FILLER_32_458 ();
 sg13g2_decap_8 FILLER_32_465 ();
 sg13g2_decap_8 FILLER_32_472 ();
 sg13g2_decap_8 FILLER_32_479 ();
 sg13g2_decap_8 FILLER_32_486 ();
 sg13g2_decap_8 FILLER_32_493 ();
 sg13g2_fill_2 FILLER_32_500 ();
 sg13g2_fill_1 FILLER_32_502 ();
 sg13g2_decap_8 FILLER_32_507 ();
 sg13g2_decap_8 FILLER_32_514 ();
 sg13g2_fill_1 FILLER_32_521 ();
 sg13g2_decap_4 FILLER_32_526 ();
 sg13g2_fill_2 FILLER_32_530 ();
 sg13g2_decap_8 FILLER_32_542 ();
 sg13g2_decap_8 FILLER_32_549 ();
 sg13g2_decap_8 FILLER_32_556 ();
 sg13g2_decap_8 FILLER_32_563 ();
 sg13g2_decap_4 FILLER_32_586 ();
 sg13g2_fill_1 FILLER_32_590 ();
 sg13g2_decap_8 FILLER_32_596 ();
 sg13g2_decap_8 FILLER_32_603 ();
 sg13g2_decap_8 FILLER_32_610 ();
 sg13g2_decap_8 FILLER_32_617 ();
 sg13g2_decap_8 FILLER_32_624 ();
 sg13g2_fill_1 FILLER_32_631 ();
 sg13g2_decap_8 FILLER_32_636 ();
 sg13g2_decap_8 FILLER_32_643 ();
 sg13g2_decap_8 FILLER_32_650 ();
 sg13g2_decap_8 FILLER_32_657 ();
 sg13g2_decap_8 FILLER_32_664 ();
 sg13g2_fill_2 FILLER_32_671 ();
 sg13g2_decap_8 FILLER_32_695 ();
 sg13g2_decap_8 FILLER_32_702 ();
 sg13g2_decap_8 FILLER_32_709 ();
 sg13g2_decap_8 FILLER_32_716 ();
 sg13g2_fill_1 FILLER_32_723 ();
 sg13g2_fill_2 FILLER_32_728 ();
 sg13g2_fill_2 FILLER_32_733 ();
 sg13g2_fill_1 FILLER_32_735 ();
 sg13g2_decap_8 FILLER_32_751 ();
 sg13g2_decap_8 FILLER_32_758 ();
 sg13g2_decap_8 FILLER_32_765 ();
 sg13g2_decap_4 FILLER_32_772 ();
 sg13g2_fill_2 FILLER_32_776 ();
 sg13g2_decap_8 FILLER_32_791 ();
 sg13g2_decap_8 FILLER_32_798 ();
 sg13g2_decap_8 FILLER_32_805 ();
 sg13g2_decap_8 FILLER_32_812 ();
 sg13g2_decap_8 FILLER_32_819 ();
 sg13g2_decap_8 FILLER_32_826 ();
 sg13g2_decap_8 FILLER_32_833 ();
 sg13g2_decap_8 FILLER_32_840 ();
 sg13g2_fill_2 FILLER_32_847 ();
 sg13g2_decap_8 FILLER_32_852 ();
 sg13g2_decap_8 FILLER_32_859 ();
 sg13g2_decap_8 FILLER_32_866 ();
 sg13g2_decap_8 FILLER_32_873 ();
 sg13g2_decap_8 FILLER_32_880 ();
 sg13g2_decap_4 FILLER_32_887 ();
 sg13g2_fill_2 FILLER_32_891 ();
 sg13g2_decap_8 FILLER_32_905 ();
 sg13g2_decap_4 FILLER_32_912 ();
 sg13g2_fill_2 FILLER_32_916 ();
 sg13g2_fill_2 FILLER_32_921 ();
 sg13g2_fill_1 FILLER_32_923 ();
 sg13g2_decap_8 FILLER_32_927 ();
 sg13g2_decap_8 FILLER_32_934 ();
 sg13g2_decap_8 FILLER_32_941 ();
 sg13g2_decap_8 FILLER_32_948 ();
 sg13g2_decap_8 FILLER_32_955 ();
 sg13g2_fill_2 FILLER_32_962 ();
 sg13g2_fill_1 FILLER_32_964 ();
 sg13g2_decap_4 FILLER_32_970 ();
 sg13g2_fill_1 FILLER_32_974 ();
 sg13g2_fill_2 FILLER_32_987 ();
 sg13g2_fill_1 FILLER_32_989 ();
 sg13g2_fill_1 FILLER_32_1005 ();
 sg13g2_decap_8 FILLER_32_1013 ();
 sg13g2_decap_8 FILLER_32_1020 ();
 sg13g2_fill_2 FILLER_32_1027 ();
 sg13g2_decap_4 FILLER_32_1035 ();
 sg13g2_fill_2 FILLER_32_1039 ();
 sg13g2_decap_8 FILLER_32_1056 ();
 sg13g2_decap_8 FILLER_32_1063 ();
 sg13g2_decap_8 FILLER_32_1070 ();
 sg13g2_decap_8 FILLER_32_1077 ();
 sg13g2_decap_8 FILLER_32_1084 ();
 sg13g2_decap_8 FILLER_32_1091 ();
 sg13g2_decap_8 FILLER_32_1098 ();
 sg13g2_decap_8 FILLER_32_1105 ();
 sg13g2_decap_8 FILLER_32_1112 ();
 sg13g2_decap_4 FILLER_32_1119 ();
 sg13g2_fill_2 FILLER_32_1123 ();
 sg13g2_decap_8 FILLER_32_1140 ();
 sg13g2_decap_4 FILLER_32_1147 ();
 sg13g2_decap_8 FILLER_32_1168 ();
 sg13g2_decap_4 FILLER_32_1175 ();
 sg13g2_fill_2 FILLER_32_1183 ();
 sg13g2_fill_1 FILLER_32_1185 ();
 sg13g2_decap_8 FILLER_32_1191 ();
 sg13g2_decap_8 FILLER_32_1198 ();
 sg13g2_decap_8 FILLER_32_1205 ();
 sg13g2_decap_8 FILLER_32_1212 ();
 sg13g2_decap_8 FILLER_32_1219 ();
 sg13g2_decap_8 FILLER_32_1226 ();
 sg13g2_decap_8 FILLER_32_1233 ();
 sg13g2_decap_4 FILLER_32_1240 ();
 sg13g2_decap_8 FILLER_32_1248 ();
 sg13g2_decap_8 FILLER_32_1255 ();
 sg13g2_decap_8 FILLER_32_1262 ();
 sg13g2_decap_8 FILLER_32_1269 ();
 sg13g2_fill_2 FILLER_32_1276 ();
 sg13g2_fill_2 FILLER_32_1281 ();
 sg13g2_decap_8 FILLER_32_1289 ();
 sg13g2_decap_8 FILLER_32_1296 ();
 sg13g2_decap_8 FILLER_32_1303 ();
 sg13g2_decap_8 FILLER_32_1310 ();
 sg13g2_decap_8 FILLER_32_1317 ();
 sg13g2_decap_8 FILLER_32_1324 ();
 sg13g2_fill_2 FILLER_32_1331 ();
 sg13g2_decap_8 FILLER_32_1339 ();
 sg13g2_decap_4 FILLER_32_1346 ();
 sg13g2_decap_8 FILLER_32_1355 ();
 sg13g2_decap_4 FILLER_32_1362 ();
 sg13g2_fill_1 FILLER_32_1366 ();
 sg13g2_decap_8 FILLER_32_1373 ();
 sg13g2_decap_8 FILLER_32_1380 ();
 sg13g2_decap_8 FILLER_32_1387 ();
 sg13g2_decap_8 FILLER_32_1394 ();
 sg13g2_decap_8 FILLER_32_1401 ();
 sg13g2_decap_8 FILLER_32_1408 ();
 sg13g2_decap_8 FILLER_32_1415 ();
 sg13g2_decap_8 FILLER_32_1422 ();
 sg13g2_decap_8 FILLER_32_1429 ();
 sg13g2_decap_8 FILLER_32_1436 ();
 sg13g2_fill_2 FILLER_32_1443 ();
 sg13g2_fill_1 FILLER_32_1445 ();
 sg13g2_decap_8 FILLER_32_1450 ();
 sg13g2_decap_8 FILLER_32_1457 ();
 sg13g2_decap_4 FILLER_32_1464 ();
 sg13g2_fill_1 FILLER_32_1468 ();
 sg13g2_decap_8 FILLER_32_1473 ();
 sg13g2_decap_8 FILLER_32_1480 ();
 sg13g2_decap_8 FILLER_32_1487 ();
 sg13g2_decap_8 FILLER_32_1494 ();
 sg13g2_decap_8 FILLER_32_1501 ();
 sg13g2_decap_8 FILLER_32_1508 ();
 sg13g2_decap_8 FILLER_32_1515 ();
 sg13g2_decap_8 FILLER_32_1522 ();
 sg13g2_decap_8 FILLER_32_1529 ();
 sg13g2_fill_2 FILLER_32_1536 ();
 sg13g2_fill_1 FILLER_32_1538 ();
 sg13g2_decap_8 FILLER_32_1544 ();
 sg13g2_decap_8 FILLER_32_1551 ();
 sg13g2_decap_4 FILLER_32_1558 ();
 sg13g2_decap_4 FILLER_32_1592 ();
 sg13g2_fill_1 FILLER_32_1596 ();
 sg13g2_decap_8 FILLER_32_1602 ();
 sg13g2_decap_8 FILLER_32_1609 ();
 sg13g2_decap_8 FILLER_32_1616 ();
 sg13g2_decap_8 FILLER_32_1623 ();
 sg13g2_fill_2 FILLER_32_1630 ();
 sg13g2_fill_1 FILLER_32_1632 ();
 sg13g2_decap_8 FILLER_32_1638 ();
 sg13g2_fill_1 FILLER_32_1645 ();
 sg13g2_decap_8 FILLER_32_1650 ();
 sg13g2_decap_8 FILLER_32_1657 ();
 sg13g2_decap_8 FILLER_32_1664 ();
 sg13g2_fill_2 FILLER_32_1671 ();
 sg13g2_fill_1 FILLER_32_1673 ();
 sg13g2_decap_4 FILLER_32_1679 ();
 sg13g2_fill_1 FILLER_32_1683 ();
 sg13g2_decap_8 FILLER_32_1690 ();
 sg13g2_decap_8 FILLER_32_1697 ();
 sg13g2_decap_8 FILLER_32_1704 ();
 sg13g2_decap_8 FILLER_32_1711 ();
 sg13g2_decap_8 FILLER_32_1718 ();
 sg13g2_decap_8 FILLER_32_1725 ();
 sg13g2_decap_8 FILLER_32_1732 ();
 sg13g2_decap_8 FILLER_32_1739 ();
 sg13g2_decap_8 FILLER_32_1746 ();
 sg13g2_decap_8 FILLER_32_1753 ();
 sg13g2_decap_8 FILLER_32_1760 ();
 sg13g2_decap_4 FILLER_32_1767 ();
 sg13g2_fill_2 FILLER_32_1771 ();
 sg13g2_decap_4 FILLER_32_1778 ();
 sg13g2_fill_1 FILLER_32_1782 ();
 sg13g2_decap_8 FILLER_32_1787 ();
 sg13g2_decap_8 FILLER_32_1794 ();
 sg13g2_decap_8 FILLER_32_1801 ();
 sg13g2_decap_8 FILLER_32_1808 ();
 sg13g2_fill_2 FILLER_32_1815 ();
 sg13g2_fill_1 FILLER_32_1817 ();
 sg13g2_decap_8 FILLER_32_1833 ();
 sg13g2_decap_8 FILLER_32_1840 ();
 sg13g2_decap_8 FILLER_32_1847 ();
 sg13g2_decap_8 FILLER_32_1866 ();
 sg13g2_decap_8 FILLER_32_1873 ();
 sg13g2_decap_8 FILLER_32_1880 ();
 sg13g2_fill_2 FILLER_32_1887 ();
 sg13g2_decap_8 FILLER_32_1904 ();
 sg13g2_decap_8 FILLER_32_1911 ();
 sg13g2_decap_8 FILLER_32_1918 ();
 sg13g2_decap_8 FILLER_32_1925 ();
 sg13g2_decap_8 FILLER_32_1932 ();
 sg13g2_decap_8 FILLER_32_1939 ();
 sg13g2_decap_8 FILLER_32_1946 ();
 sg13g2_decap_8 FILLER_32_1953 ();
 sg13g2_decap_8 FILLER_32_1960 ();
 sg13g2_decap_8 FILLER_32_1967 ();
 sg13g2_decap_8 FILLER_32_1974 ();
 sg13g2_decap_8 FILLER_32_1981 ();
 sg13g2_decap_8 FILLER_32_1988 ();
 sg13g2_decap_8 FILLER_32_1995 ();
 sg13g2_decap_8 FILLER_32_2002 ();
 sg13g2_decap_8 FILLER_32_2009 ();
 sg13g2_decap_8 FILLER_32_2016 ();
 sg13g2_decap_8 FILLER_32_2023 ();
 sg13g2_decap_8 FILLER_32_2030 ();
 sg13g2_decap_8 FILLER_32_2037 ();
 sg13g2_decap_8 FILLER_32_2044 ();
 sg13g2_decap_8 FILLER_32_2051 ();
 sg13g2_decap_8 FILLER_32_2058 ();
 sg13g2_decap_8 FILLER_32_2065 ();
 sg13g2_decap_8 FILLER_32_2072 ();
 sg13g2_decap_8 FILLER_32_2079 ();
 sg13g2_decap_8 FILLER_32_2086 ();
 sg13g2_decap_8 FILLER_32_2093 ();
 sg13g2_decap_8 FILLER_32_2100 ();
 sg13g2_decap_8 FILLER_32_2107 ();
 sg13g2_decap_8 FILLER_32_2114 ();
 sg13g2_decap_8 FILLER_32_2121 ();
 sg13g2_decap_8 FILLER_32_2128 ();
 sg13g2_decap_8 FILLER_32_2135 ();
 sg13g2_decap_8 FILLER_32_2142 ();
 sg13g2_decap_8 FILLER_32_2149 ();
 sg13g2_decap_8 FILLER_32_2156 ();
 sg13g2_decap_8 FILLER_32_2163 ();
 sg13g2_decap_8 FILLER_32_2170 ();
 sg13g2_decap_8 FILLER_32_2177 ();
 sg13g2_decap_8 FILLER_32_2184 ();
 sg13g2_decap_8 FILLER_32_2191 ();
 sg13g2_decap_8 FILLER_32_2198 ();
 sg13g2_decap_8 FILLER_32_2205 ();
 sg13g2_decap_8 FILLER_32_2212 ();
 sg13g2_decap_8 FILLER_32_2219 ();
 sg13g2_decap_8 FILLER_32_2226 ();
 sg13g2_decap_8 FILLER_32_2233 ();
 sg13g2_decap_8 FILLER_32_2240 ();
 sg13g2_decap_8 FILLER_32_2247 ();
 sg13g2_decap_8 FILLER_32_2254 ();
 sg13g2_decap_8 FILLER_32_2261 ();
 sg13g2_decap_8 FILLER_32_2268 ();
 sg13g2_decap_8 FILLER_32_2275 ();
 sg13g2_decap_8 FILLER_32_2282 ();
 sg13g2_decap_8 FILLER_32_2289 ();
 sg13g2_decap_8 FILLER_32_2296 ();
 sg13g2_decap_8 FILLER_32_2303 ();
 sg13g2_decap_8 FILLER_32_2310 ();
 sg13g2_decap_8 FILLER_32_2317 ();
 sg13g2_decap_8 FILLER_32_2324 ();
 sg13g2_decap_8 FILLER_32_2331 ();
 sg13g2_decap_8 FILLER_32_2338 ();
 sg13g2_decap_8 FILLER_32_2345 ();
 sg13g2_decap_8 FILLER_32_2352 ();
 sg13g2_decap_8 FILLER_32_2359 ();
 sg13g2_decap_8 FILLER_32_2366 ();
 sg13g2_decap_8 FILLER_32_2373 ();
 sg13g2_decap_8 FILLER_32_2380 ();
 sg13g2_decap_8 FILLER_32_2387 ();
 sg13g2_decap_8 FILLER_32_2394 ();
 sg13g2_decap_8 FILLER_32_2401 ();
 sg13g2_decap_8 FILLER_32_2408 ();
 sg13g2_decap_8 FILLER_32_2415 ();
 sg13g2_decap_8 FILLER_32_2422 ();
 sg13g2_decap_8 FILLER_32_2429 ();
 sg13g2_decap_8 FILLER_32_2436 ();
 sg13g2_decap_8 FILLER_32_2443 ();
 sg13g2_decap_8 FILLER_32_2450 ();
 sg13g2_decap_8 FILLER_32_2457 ();
 sg13g2_decap_8 FILLER_32_2464 ();
 sg13g2_decap_8 FILLER_32_2471 ();
 sg13g2_decap_8 FILLER_32_2478 ();
 sg13g2_decap_8 FILLER_32_2485 ();
 sg13g2_decap_8 FILLER_32_2492 ();
 sg13g2_decap_8 FILLER_32_2499 ();
 sg13g2_decap_8 FILLER_32_2506 ();
 sg13g2_decap_8 FILLER_32_2513 ();
 sg13g2_decap_8 FILLER_32_2520 ();
 sg13g2_decap_8 FILLER_32_2527 ();
 sg13g2_decap_8 FILLER_32_2534 ();
 sg13g2_decap_8 FILLER_32_2541 ();
 sg13g2_decap_8 FILLER_32_2548 ();
 sg13g2_decap_8 FILLER_32_2555 ();
 sg13g2_decap_8 FILLER_32_2562 ();
 sg13g2_decap_8 FILLER_32_2569 ();
 sg13g2_decap_8 FILLER_32_2576 ();
 sg13g2_decap_8 FILLER_32_2583 ();
 sg13g2_decap_8 FILLER_32_2590 ();
 sg13g2_decap_8 FILLER_32_2597 ();
 sg13g2_decap_8 FILLER_32_2604 ();
 sg13g2_decap_8 FILLER_32_2611 ();
 sg13g2_decap_8 FILLER_32_2618 ();
 sg13g2_decap_8 FILLER_32_2625 ();
 sg13g2_decap_8 FILLER_32_2632 ();
 sg13g2_decap_8 FILLER_32_2639 ();
 sg13g2_decap_8 FILLER_32_2646 ();
 sg13g2_decap_8 FILLER_32_2653 ();
 sg13g2_decap_8 FILLER_32_2660 ();
 sg13g2_fill_2 FILLER_32_2667 ();
 sg13g2_fill_1 FILLER_32_2669 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_4 FILLER_33_77 ();
 sg13g2_fill_1 FILLER_33_81 ();
 sg13g2_decap_8 FILLER_33_86 ();
 sg13g2_decap_8 FILLER_33_93 ();
 sg13g2_decap_8 FILLER_33_100 ();
 sg13g2_decap_8 FILLER_33_107 ();
 sg13g2_decap_8 FILLER_33_114 ();
 sg13g2_decap_8 FILLER_33_121 ();
 sg13g2_decap_8 FILLER_33_128 ();
 sg13g2_decap_8 FILLER_33_135 ();
 sg13g2_decap_8 FILLER_33_142 ();
 sg13g2_decap_8 FILLER_33_149 ();
 sg13g2_decap_8 FILLER_33_156 ();
 sg13g2_decap_8 FILLER_33_163 ();
 sg13g2_decap_8 FILLER_33_170 ();
 sg13g2_decap_8 FILLER_33_177 ();
 sg13g2_decap_8 FILLER_33_184 ();
 sg13g2_decap_8 FILLER_33_191 ();
 sg13g2_decap_8 FILLER_33_198 ();
 sg13g2_decap_8 FILLER_33_205 ();
 sg13g2_decap_8 FILLER_33_212 ();
 sg13g2_decap_8 FILLER_33_219 ();
 sg13g2_decap_8 FILLER_33_226 ();
 sg13g2_decap_8 FILLER_33_233 ();
 sg13g2_decap_8 FILLER_33_240 ();
 sg13g2_decap_8 FILLER_33_247 ();
 sg13g2_decap_8 FILLER_33_254 ();
 sg13g2_decap_8 FILLER_33_261 ();
 sg13g2_decap_8 FILLER_33_268 ();
 sg13g2_decap_8 FILLER_33_275 ();
 sg13g2_decap_8 FILLER_33_282 ();
 sg13g2_decap_8 FILLER_33_289 ();
 sg13g2_decap_8 FILLER_33_296 ();
 sg13g2_decap_8 FILLER_33_303 ();
 sg13g2_decap_8 FILLER_33_310 ();
 sg13g2_decap_8 FILLER_33_317 ();
 sg13g2_decap_8 FILLER_33_324 ();
 sg13g2_decap_8 FILLER_33_331 ();
 sg13g2_decap_8 FILLER_33_338 ();
 sg13g2_decap_8 FILLER_33_345 ();
 sg13g2_decap_8 FILLER_33_352 ();
 sg13g2_decap_8 FILLER_33_359 ();
 sg13g2_decap_8 FILLER_33_366 ();
 sg13g2_decap_8 FILLER_33_373 ();
 sg13g2_decap_8 FILLER_33_380 ();
 sg13g2_decap_8 FILLER_33_387 ();
 sg13g2_decap_8 FILLER_33_394 ();
 sg13g2_decap_8 FILLER_33_401 ();
 sg13g2_decap_8 FILLER_33_408 ();
 sg13g2_fill_1 FILLER_33_415 ();
 sg13g2_decap_8 FILLER_33_422 ();
 sg13g2_decap_8 FILLER_33_429 ();
 sg13g2_fill_2 FILLER_33_436 ();
 sg13g2_decap_4 FILLER_33_442 ();
 sg13g2_fill_2 FILLER_33_446 ();
 sg13g2_decap_4 FILLER_33_453 ();
 sg13g2_decap_8 FILLER_33_466 ();
 sg13g2_decap_8 FILLER_33_473 ();
 sg13g2_decap_8 FILLER_33_480 ();
 sg13g2_decap_8 FILLER_33_487 ();
 sg13g2_decap_8 FILLER_33_494 ();
 sg13g2_decap_8 FILLER_33_501 ();
 sg13g2_decap_4 FILLER_33_508 ();
 sg13g2_fill_1 FILLER_33_512 ();
 sg13g2_decap_8 FILLER_33_539 ();
 sg13g2_fill_2 FILLER_33_546 ();
 sg13g2_decap_8 FILLER_33_563 ();
 sg13g2_decap_8 FILLER_33_570 ();
 sg13g2_decap_4 FILLER_33_577 ();
 sg13g2_fill_1 FILLER_33_581 ();
 sg13g2_decap_8 FILLER_33_586 ();
 sg13g2_decap_8 FILLER_33_593 ();
 sg13g2_decap_8 FILLER_33_600 ();
 sg13g2_decap_8 FILLER_33_607 ();
 sg13g2_decap_8 FILLER_33_614 ();
 sg13g2_decap_8 FILLER_33_621 ();
 sg13g2_decap_4 FILLER_33_628 ();
 sg13g2_fill_2 FILLER_33_632 ();
 sg13g2_decap_8 FILLER_33_638 ();
 sg13g2_decap_8 FILLER_33_645 ();
 sg13g2_decap_8 FILLER_33_652 ();
 sg13g2_decap_8 FILLER_33_659 ();
 sg13g2_decap_8 FILLER_33_666 ();
 sg13g2_decap_8 FILLER_33_673 ();
 sg13g2_decap_8 FILLER_33_680 ();
 sg13g2_decap_8 FILLER_33_687 ();
 sg13g2_decap_8 FILLER_33_694 ();
 sg13g2_decap_8 FILLER_33_701 ();
 sg13g2_decap_8 FILLER_33_708 ();
 sg13g2_decap_8 FILLER_33_715 ();
 sg13g2_fill_1 FILLER_33_729 ();
 sg13g2_decap_8 FILLER_33_746 ();
 sg13g2_decap_8 FILLER_33_753 ();
 sg13g2_decap_8 FILLER_33_760 ();
 sg13g2_decap_4 FILLER_33_767 ();
 sg13g2_fill_2 FILLER_33_771 ();
 sg13g2_decap_8 FILLER_33_777 ();
 sg13g2_fill_2 FILLER_33_784 ();
 sg13g2_fill_1 FILLER_33_786 ();
 sg13g2_fill_2 FILLER_33_799 ();
 sg13g2_decap_8 FILLER_33_805 ();
 sg13g2_decap_8 FILLER_33_812 ();
 sg13g2_decap_8 FILLER_33_819 ();
 sg13g2_decap_8 FILLER_33_826 ();
 sg13g2_decap_4 FILLER_33_833 ();
 sg13g2_fill_2 FILLER_33_837 ();
 sg13g2_fill_2 FILLER_33_842 ();
 sg13g2_fill_1 FILLER_33_844 ();
 sg13g2_decap_8 FILLER_33_857 ();
 sg13g2_decap_8 FILLER_33_864 ();
 sg13g2_decap_8 FILLER_33_871 ();
 sg13g2_decap_8 FILLER_33_878 ();
 sg13g2_decap_4 FILLER_33_885 ();
 sg13g2_fill_1 FILLER_33_889 ();
 sg13g2_decap_8 FILLER_33_898 ();
 sg13g2_decap_8 FILLER_33_905 ();
 sg13g2_decap_4 FILLER_33_912 ();
 sg13g2_fill_2 FILLER_33_916 ();
 sg13g2_decap_8 FILLER_33_923 ();
 sg13g2_decap_8 FILLER_33_930 ();
 sg13g2_decap_8 FILLER_33_937 ();
 sg13g2_decap_8 FILLER_33_944 ();
 sg13g2_decap_8 FILLER_33_951 ();
 sg13g2_decap_8 FILLER_33_958 ();
 sg13g2_fill_2 FILLER_33_965 ();
 sg13g2_fill_1 FILLER_33_971 ();
 sg13g2_decap_8 FILLER_33_984 ();
 sg13g2_fill_2 FILLER_33_991 ();
 sg13g2_decap_8 FILLER_33_998 ();
 sg13g2_decap_4 FILLER_33_1005 ();
 sg13g2_decap_8 FILLER_33_1016 ();
 sg13g2_decap_4 FILLER_33_1023 ();
 sg13g2_fill_2 FILLER_33_1027 ();
 sg13g2_decap_8 FILLER_33_1037 ();
 sg13g2_decap_8 FILLER_33_1044 ();
 sg13g2_decap_8 FILLER_33_1051 ();
 sg13g2_decap_8 FILLER_33_1058 ();
 sg13g2_decap_8 FILLER_33_1065 ();
 sg13g2_decap_8 FILLER_33_1072 ();
 sg13g2_decap_4 FILLER_33_1079 ();
 sg13g2_fill_1 FILLER_33_1083 ();
 sg13g2_decap_8 FILLER_33_1093 ();
 sg13g2_decap_8 FILLER_33_1100 ();
 sg13g2_decap_8 FILLER_33_1107 ();
 sg13g2_fill_2 FILLER_33_1114 ();
 sg13g2_decap_8 FILLER_33_1133 ();
 sg13g2_decap_8 FILLER_33_1140 ();
 sg13g2_decap_8 FILLER_33_1147 ();
 sg13g2_decap_8 FILLER_33_1154 ();
 sg13g2_fill_2 FILLER_33_1161 ();
 sg13g2_fill_1 FILLER_33_1163 ();
 sg13g2_decap_8 FILLER_33_1178 ();
 sg13g2_decap_4 FILLER_33_1185 ();
 sg13g2_decap_8 FILLER_33_1193 ();
 sg13g2_decap_8 FILLER_33_1200 ();
 sg13g2_decap_8 FILLER_33_1207 ();
 sg13g2_decap_8 FILLER_33_1214 ();
 sg13g2_decap_8 FILLER_33_1221 ();
 sg13g2_decap_4 FILLER_33_1228 ();
 sg13g2_decap_8 FILLER_33_1236 ();
 sg13g2_decap_8 FILLER_33_1243 ();
 sg13g2_decap_8 FILLER_33_1250 ();
 sg13g2_decap_8 FILLER_33_1257 ();
 sg13g2_decap_8 FILLER_33_1264 ();
 sg13g2_decap_8 FILLER_33_1271 ();
 sg13g2_decap_8 FILLER_33_1287 ();
 sg13g2_decap_8 FILLER_33_1294 ();
 sg13g2_decap_4 FILLER_33_1301 ();
 sg13g2_fill_1 FILLER_33_1305 ();
 sg13g2_fill_1 FILLER_33_1332 ();
 sg13g2_fill_2 FILLER_33_1339 ();
 sg13g2_decap_8 FILLER_33_1346 ();
 sg13g2_decap_4 FILLER_33_1353 ();
 sg13g2_fill_1 FILLER_33_1357 ();
 sg13g2_fill_2 FILLER_33_1370 ();
 sg13g2_fill_2 FILLER_33_1378 ();
 sg13g2_fill_1 FILLER_33_1380 ();
 sg13g2_decap_8 FILLER_33_1386 ();
 sg13g2_decap_8 FILLER_33_1393 ();
 sg13g2_decap_8 FILLER_33_1400 ();
 sg13g2_decap_8 FILLER_33_1407 ();
 sg13g2_decap_8 FILLER_33_1414 ();
 sg13g2_decap_8 FILLER_33_1421 ();
 sg13g2_decap_8 FILLER_33_1428 ();
 sg13g2_decap_8 FILLER_33_1435 ();
 sg13g2_decap_8 FILLER_33_1442 ();
 sg13g2_decap_8 FILLER_33_1457 ();
 sg13g2_decap_8 FILLER_33_1464 ();
 sg13g2_decap_8 FILLER_33_1471 ();
 sg13g2_decap_8 FILLER_33_1478 ();
 sg13g2_decap_8 FILLER_33_1485 ();
 sg13g2_decap_8 FILLER_33_1492 ();
 sg13g2_fill_2 FILLER_33_1499 ();
 sg13g2_decap_8 FILLER_33_1505 ();
 sg13g2_decap_8 FILLER_33_1512 ();
 sg13g2_decap_8 FILLER_33_1519 ();
 sg13g2_decap_8 FILLER_33_1526 ();
 sg13g2_decap_8 FILLER_33_1533 ();
 sg13g2_fill_1 FILLER_33_1540 ();
 sg13g2_fill_2 FILLER_33_1545 ();
 sg13g2_fill_1 FILLER_33_1547 ();
 sg13g2_decap_8 FILLER_33_1553 ();
 sg13g2_decap_8 FILLER_33_1560 ();
 sg13g2_decap_8 FILLER_33_1567 ();
 sg13g2_decap_8 FILLER_33_1574 ();
 sg13g2_decap_8 FILLER_33_1581 ();
 sg13g2_decap_8 FILLER_33_1588 ();
 sg13g2_decap_8 FILLER_33_1595 ();
 sg13g2_decap_8 FILLER_33_1602 ();
 sg13g2_fill_1 FILLER_33_1609 ();
 sg13g2_decap_8 FILLER_33_1616 ();
 sg13g2_decap_8 FILLER_33_1623 ();
 sg13g2_decap_8 FILLER_33_1630 ();
 sg13g2_decap_8 FILLER_33_1637 ();
 sg13g2_fill_2 FILLER_33_1644 ();
 sg13g2_fill_2 FILLER_33_1649 ();
 sg13g2_decap_8 FILLER_33_1669 ();
 sg13g2_decap_8 FILLER_33_1676 ();
 sg13g2_decap_8 FILLER_33_1683 ();
 sg13g2_decap_8 FILLER_33_1690 ();
 sg13g2_decap_8 FILLER_33_1697 ();
 sg13g2_decap_8 FILLER_33_1704 ();
 sg13g2_decap_8 FILLER_33_1711 ();
 sg13g2_fill_2 FILLER_33_1718 ();
 sg13g2_fill_1 FILLER_33_1720 ();
 sg13g2_decap_8 FILLER_33_1732 ();
 sg13g2_decap_8 FILLER_33_1739 ();
 sg13g2_decap_8 FILLER_33_1746 ();
 sg13g2_decap_8 FILLER_33_1753 ();
 sg13g2_decap_8 FILLER_33_1760 ();
 sg13g2_decap_8 FILLER_33_1767 ();
 sg13g2_decap_8 FILLER_33_1774 ();
 sg13g2_decap_8 FILLER_33_1781 ();
 sg13g2_decap_8 FILLER_33_1788 ();
 sg13g2_decap_8 FILLER_33_1795 ();
 sg13g2_decap_8 FILLER_33_1802 ();
 sg13g2_decap_8 FILLER_33_1809 ();
 sg13g2_fill_2 FILLER_33_1816 ();
 sg13g2_decap_8 FILLER_33_1822 ();
 sg13g2_decap_8 FILLER_33_1829 ();
 sg13g2_decap_8 FILLER_33_1836 ();
 sg13g2_decap_8 FILLER_33_1843 ();
 sg13g2_decap_8 FILLER_33_1850 ();
 sg13g2_decap_4 FILLER_33_1857 ();
 sg13g2_decap_8 FILLER_33_1870 ();
 sg13g2_decap_8 FILLER_33_1877 ();
 sg13g2_decap_4 FILLER_33_1884 ();
 sg13g2_fill_1 FILLER_33_1888 ();
 sg13g2_decap_8 FILLER_33_1902 ();
 sg13g2_decap_8 FILLER_33_1909 ();
 sg13g2_decap_8 FILLER_33_1916 ();
 sg13g2_decap_8 FILLER_33_1923 ();
 sg13g2_decap_8 FILLER_33_1930 ();
 sg13g2_decap_8 FILLER_33_1937 ();
 sg13g2_decap_8 FILLER_33_1944 ();
 sg13g2_decap_8 FILLER_33_1951 ();
 sg13g2_decap_8 FILLER_33_1958 ();
 sg13g2_decap_8 FILLER_33_1965 ();
 sg13g2_decap_8 FILLER_33_1972 ();
 sg13g2_decap_8 FILLER_33_1979 ();
 sg13g2_decap_8 FILLER_33_1986 ();
 sg13g2_decap_8 FILLER_33_1993 ();
 sg13g2_decap_8 FILLER_33_2000 ();
 sg13g2_decap_8 FILLER_33_2007 ();
 sg13g2_decap_8 FILLER_33_2014 ();
 sg13g2_decap_8 FILLER_33_2021 ();
 sg13g2_decap_8 FILLER_33_2028 ();
 sg13g2_decap_8 FILLER_33_2035 ();
 sg13g2_decap_8 FILLER_33_2042 ();
 sg13g2_decap_8 FILLER_33_2049 ();
 sg13g2_decap_8 FILLER_33_2056 ();
 sg13g2_decap_8 FILLER_33_2063 ();
 sg13g2_decap_8 FILLER_33_2070 ();
 sg13g2_decap_8 FILLER_33_2077 ();
 sg13g2_decap_8 FILLER_33_2084 ();
 sg13g2_decap_8 FILLER_33_2091 ();
 sg13g2_decap_8 FILLER_33_2098 ();
 sg13g2_decap_8 FILLER_33_2105 ();
 sg13g2_decap_8 FILLER_33_2112 ();
 sg13g2_decap_8 FILLER_33_2119 ();
 sg13g2_decap_8 FILLER_33_2126 ();
 sg13g2_decap_8 FILLER_33_2133 ();
 sg13g2_decap_8 FILLER_33_2140 ();
 sg13g2_decap_8 FILLER_33_2147 ();
 sg13g2_decap_8 FILLER_33_2154 ();
 sg13g2_decap_8 FILLER_33_2161 ();
 sg13g2_decap_8 FILLER_33_2168 ();
 sg13g2_decap_8 FILLER_33_2175 ();
 sg13g2_decap_8 FILLER_33_2182 ();
 sg13g2_decap_8 FILLER_33_2189 ();
 sg13g2_decap_8 FILLER_33_2196 ();
 sg13g2_decap_8 FILLER_33_2203 ();
 sg13g2_decap_8 FILLER_33_2210 ();
 sg13g2_decap_8 FILLER_33_2217 ();
 sg13g2_decap_8 FILLER_33_2224 ();
 sg13g2_decap_8 FILLER_33_2231 ();
 sg13g2_decap_8 FILLER_33_2238 ();
 sg13g2_decap_8 FILLER_33_2245 ();
 sg13g2_decap_8 FILLER_33_2252 ();
 sg13g2_decap_8 FILLER_33_2259 ();
 sg13g2_decap_8 FILLER_33_2266 ();
 sg13g2_decap_8 FILLER_33_2273 ();
 sg13g2_decap_8 FILLER_33_2280 ();
 sg13g2_decap_8 FILLER_33_2287 ();
 sg13g2_decap_8 FILLER_33_2294 ();
 sg13g2_decap_8 FILLER_33_2301 ();
 sg13g2_decap_8 FILLER_33_2308 ();
 sg13g2_decap_8 FILLER_33_2315 ();
 sg13g2_decap_8 FILLER_33_2322 ();
 sg13g2_decap_8 FILLER_33_2329 ();
 sg13g2_decap_8 FILLER_33_2336 ();
 sg13g2_decap_8 FILLER_33_2343 ();
 sg13g2_decap_8 FILLER_33_2350 ();
 sg13g2_decap_8 FILLER_33_2357 ();
 sg13g2_decap_8 FILLER_33_2364 ();
 sg13g2_decap_8 FILLER_33_2371 ();
 sg13g2_decap_8 FILLER_33_2378 ();
 sg13g2_decap_8 FILLER_33_2385 ();
 sg13g2_decap_8 FILLER_33_2392 ();
 sg13g2_decap_8 FILLER_33_2399 ();
 sg13g2_decap_8 FILLER_33_2406 ();
 sg13g2_decap_8 FILLER_33_2413 ();
 sg13g2_decap_8 FILLER_33_2420 ();
 sg13g2_decap_8 FILLER_33_2427 ();
 sg13g2_decap_8 FILLER_33_2434 ();
 sg13g2_decap_8 FILLER_33_2441 ();
 sg13g2_decap_8 FILLER_33_2448 ();
 sg13g2_decap_8 FILLER_33_2455 ();
 sg13g2_decap_8 FILLER_33_2462 ();
 sg13g2_decap_8 FILLER_33_2469 ();
 sg13g2_decap_8 FILLER_33_2476 ();
 sg13g2_decap_8 FILLER_33_2483 ();
 sg13g2_decap_8 FILLER_33_2490 ();
 sg13g2_decap_8 FILLER_33_2497 ();
 sg13g2_decap_8 FILLER_33_2504 ();
 sg13g2_decap_8 FILLER_33_2511 ();
 sg13g2_decap_8 FILLER_33_2518 ();
 sg13g2_decap_8 FILLER_33_2525 ();
 sg13g2_decap_8 FILLER_33_2532 ();
 sg13g2_decap_8 FILLER_33_2539 ();
 sg13g2_decap_8 FILLER_33_2546 ();
 sg13g2_decap_8 FILLER_33_2553 ();
 sg13g2_decap_8 FILLER_33_2560 ();
 sg13g2_decap_8 FILLER_33_2567 ();
 sg13g2_decap_8 FILLER_33_2574 ();
 sg13g2_decap_8 FILLER_33_2581 ();
 sg13g2_decap_8 FILLER_33_2588 ();
 sg13g2_decap_8 FILLER_33_2595 ();
 sg13g2_decap_8 FILLER_33_2602 ();
 sg13g2_decap_8 FILLER_33_2609 ();
 sg13g2_decap_8 FILLER_33_2616 ();
 sg13g2_decap_8 FILLER_33_2623 ();
 sg13g2_decap_8 FILLER_33_2630 ();
 sg13g2_decap_8 FILLER_33_2637 ();
 sg13g2_decap_8 FILLER_33_2644 ();
 sg13g2_decap_8 FILLER_33_2651 ();
 sg13g2_decap_8 FILLER_33_2658 ();
 sg13g2_decap_4 FILLER_33_2665 ();
 sg13g2_fill_1 FILLER_33_2669 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_4 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_134 ();
 sg13g2_decap_8 FILLER_34_141 ();
 sg13g2_decap_8 FILLER_34_148 ();
 sg13g2_decap_8 FILLER_34_155 ();
 sg13g2_decap_8 FILLER_34_162 ();
 sg13g2_decap_8 FILLER_34_169 ();
 sg13g2_decap_8 FILLER_34_176 ();
 sg13g2_decap_8 FILLER_34_183 ();
 sg13g2_decap_8 FILLER_34_190 ();
 sg13g2_decap_4 FILLER_34_197 ();
 sg13g2_fill_1 FILLER_34_201 ();
 sg13g2_decap_8 FILLER_34_206 ();
 sg13g2_decap_8 FILLER_34_213 ();
 sg13g2_decap_8 FILLER_34_220 ();
 sg13g2_decap_8 FILLER_34_227 ();
 sg13g2_decap_8 FILLER_34_234 ();
 sg13g2_decap_8 FILLER_34_241 ();
 sg13g2_decap_8 FILLER_34_248 ();
 sg13g2_decap_8 FILLER_34_255 ();
 sg13g2_decap_8 FILLER_34_262 ();
 sg13g2_decap_8 FILLER_34_269 ();
 sg13g2_decap_8 FILLER_34_276 ();
 sg13g2_decap_8 FILLER_34_283 ();
 sg13g2_decap_4 FILLER_34_290 ();
 sg13g2_fill_1 FILLER_34_294 ();
 sg13g2_decap_8 FILLER_34_299 ();
 sg13g2_decap_8 FILLER_34_306 ();
 sg13g2_decap_8 FILLER_34_313 ();
 sg13g2_decap_8 FILLER_34_320 ();
 sg13g2_decap_8 FILLER_34_327 ();
 sg13g2_decap_8 FILLER_34_334 ();
 sg13g2_decap_8 FILLER_34_341 ();
 sg13g2_decap_8 FILLER_34_348 ();
 sg13g2_decap_8 FILLER_34_355 ();
 sg13g2_decap_8 FILLER_34_362 ();
 sg13g2_decap_8 FILLER_34_369 ();
 sg13g2_decap_8 FILLER_34_376 ();
 sg13g2_fill_2 FILLER_34_383 ();
 sg13g2_fill_1 FILLER_34_385 ();
 sg13g2_fill_1 FILLER_34_401 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_fill_1 FILLER_34_409 ();
 sg13g2_decap_8 FILLER_34_423 ();
 sg13g2_decap_4 FILLER_34_430 ();
 sg13g2_fill_1 FILLER_34_434 ();
 sg13g2_decap_8 FILLER_34_439 ();
 sg13g2_decap_8 FILLER_34_446 ();
 sg13g2_decap_8 FILLER_34_453 ();
 sg13g2_decap_8 FILLER_34_460 ();
 sg13g2_decap_8 FILLER_34_467 ();
 sg13g2_decap_8 FILLER_34_474 ();
 sg13g2_decap_4 FILLER_34_481 ();
 sg13g2_fill_1 FILLER_34_485 ();
 sg13g2_decap_8 FILLER_34_490 ();
 sg13g2_decap_8 FILLER_34_502 ();
 sg13g2_decap_8 FILLER_34_509 ();
 sg13g2_decap_8 FILLER_34_516 ();
 sg13g2_fill_2 FILLER_34_523 ();
 sg13g2_decap_8 FILLER_34_528 ();
 sg13g2_fill_1 FILLER_34_535 ();
 sg13g2_decap_8 FILLER_34_541 ();
 sg13g2_fill_2 FILLER_34_548 ();
 sg13g2_fill_1 FILLER_34_550 ();
 sg13g2_decap_8 FILLER_34_555 ();
 sg13g2_decap_4 FILLER_34_562 ();
 sg13g2_fill_2 FILLER_34_566 ();
 sg13g2_decap_4 FILLER_34_576 ();
 sg13g2_fill_2 FILLER_34_584 ();
 sg13g2_fill_1 FILLER_34_586 ();
 sg13g2_fill_1 FILLER_34_597 ();
 sg13g2_decap_8 FILLER_34_602 ();
 sg13g2_decap_8 FILLER_34_609 ();
 sg13g2_decap_8 FILLER_34_616 ();
 sg13g2_decap_8 FILLER_34_623 ();
 sg13g2_decap_8 FILLER_34_630 ();
 sg13g2_decap_8 FILLER_34_637 ();
 sg13g2_decap_8 FILLER_34_644 ();
 sg13g2_decap_8 FILLER_34_651 ();
 sg13g2_decap_8 FILLER_34_658 ();
 sg13g2_decap_8 FILLER_34_665 ();
 sg13g2_decap_4 FILLER_34_672 ();
 sg13g2_fill_1 FILLER_34_676 ();
 sg13g2_decap_8 FILLER_34_692 ();
 sg13g2_decap_8 FILLER_34_699 ();
 sg13g2_decap_8 FILLER_34_706 ();
 sg13g2_decap_8 FILLER_34_713 ();
 sg13g2_decap_4 FILLER_34_720 ();
 sg13g2_fill_1 FILLER_34_724 ();
 sg13g2_decap_8 FILLER_34_728 ();
 sg13g2_decap_8 FILLER_34_735 ();
 sg13g2_decap_8 FILLER_34_742 ();
 sg13g2_decap_8 FILLER_34_749 ();
 sg13g2_decap_8 FILLER_34_756 ();
 sg13g2_decap_8 FILLER_34_763 ();
 sg13g2_decap_8 FILLER_34_770 ();
 sg13g2_decap_4 FILLER_34_777 ();
 sg13g2_fill_2 FILLER_34_795 ();
 sg13g2_fill_1 FILLER_34_797 ();
 sg13g2_decap_8 FILLER_34_813 ();
 sg13g2_fill_1 FILLER_34_820 ();
 sg13g2_decap_8 FILLER_34_825 ();
 sg13g2_decap_8 FILLER_34_832 ();
 sg13g2_decap_8 FILLER_34_845 ();
 sg13g2_decap_8 FILLER_34_852 ();
 sg13g2_decap_8 FILLER_34_859 ();
 sg13g2_decap_8 FILLER_34_866 ();
 sg13g2_decap_8 FILLER_34_873 ();
 sg13g2_decap_8 FILLER_34_880 ();
 sg13g2_decap_8 FILLER_34_887 ();
 sg13g2_decap_8 FILLER_34_894 ();
 sg13g2_decap_8 FILLER_34_901 ();
 sg13g2_decap_8 FILLER_34_908 ();
 sg13g2_fill_2 FILLER_34_915 ();
 sg13g2_decap_8 FILLER_34_922 ();
 sg13g2_decap_8 FILLER_34_929 ();
 sg13g2_decap_8 FILLER_34_936 ();
 sg13g2_decap_8 FILLER_34_943 ();
 sg13g2_decap_8 FILLER_34_950 ();
 sg13g2_decap_8 FILLER_34_957 ();
 sg13g2_decap_8 FILLER_34_964 ();
 sg13g2_decap_8 FILLER_34_971 ();
 sg13g2_decap_8 FILLER_34_978 ();
 sg13g2_decap_8 FILLER_34_985 ();
 sg13g2_decap_8 FILLER_34_992 ();
 sg13g2_decap_8 FILLER_34_999 ();
 sg13g2_decap_4 FILLER_34_1006 ();
 sg13g2_fill_2 FILLER_34_1010 ();
 sg13g2_decap_8 FILLER_34_1019 ();
 sg13g2_fill_1 FILLER_34_1026 ();
 sg13g2_decap_8 FILLER_34_1035 ();
 sg13g2_decap_8 FILLER_34_1042 ();
 sg13g2_decap_4 FILLER_34_1049 ();
 sg13g2_fill_2 FILLER_34_1053 ();
 sg13g2_decap_8 FILLER_34_1064 ();
 sg13g2_decap_8 FILLER_34_1071 ();
 sg13g2_fill_1 FILLER_34_1078 ();
 sg13g2_decap_8 FILLER_34_1095 ();
 sg13g2_decap_8 FILLER_34_1102 ();
 sg13g2_decap_8 FILLER_34_1109 ();
 sg13g2_decap_4 FILLER_34_1116 ();
 sg13g2_fill_1 FILLER_34_1120 ();
 sg13g2_fill_2 FILLER_34_1125 ();
 sg13g2_fill_1 FILLER_34_1127 ();
 sg13g2_decap_8 FILLER_34_1139 ();
 sg13g2_decap_8 FILLER_34_1146 ();
 sg13g2_decap_8 FILLER_34_1153 ();
 sg13g2_decap_8 FILLER_34_1160 ();
 sg13g2_decap_8 FILLER_34_1172 ();
 sg13g2_decap_8 FILLER_34_1179 ();
 sg13g2_decap_8 FILLER_34_1186 ();
 sg13g2_decap_8 FILLER_34_1193 ();
 sg13g2_decap_8 FILLER_34_1200 ();
 sg13g2_decap_8 FILLER_34_1207 ();
 sg13g2_decap_8 FILLER_34_1218 ();
 sg13g2_decap_8 FILLER_34_1225 ();
 sg13g2_decap_8 FILLER_34_1232 ();
 sg13g2_decap_8 FILLER_34_1239 ();
 sg13g2_decap_8 FILLER_34_1246 ();
 sg13g2_decap_8 FILLER_34_1253 ();
 sg13g2_decap_4 FILLER_34_1260 ();
 sg13g2_fill_2 FILLER_34_1264 ();
 sg13g2_decap_8 FILLER_34_1278 ();
 sg13g2_decap_8 FILLER_34_1285 ();
 sg13g2_decap_8 FILLER_34_1292 ();
 sg13g2_decap_8 FILLER_34_1299 ();
 sg13g2_decap_8 FILLER_34_1306 ();
 sg13g2_decap_4 FILLER_34_1313 ();
 sg13g2_fill_1 FILLER_34_1317 ();
 sg13g2_fill_1 FILLER_34_1324 ();
 sg13g2_fill_2 FILLER_34_1330 ();
 sg13g2_fill_1 FILLER_34_1332 ();
 sg13g2_decap_8 FILLER_34_1345 ();
 sg13g2_fill_2 FILLER_34_1352 ();
 sg13g2_fill_1 FILLER_34_1354 ();
 sg13g2_decap_8 FILLER_34_1367 ();
 sg13g2_decap_8 FILLER_34_1374 ();
 sg13g2_decap_8 FILLER_34_1381 ();
 sg13g2_decap_8 FILLER_34_1388 ();
 sg13g2_decap_8 FILLER_34_1395 ();
 sg13g2_fill_2 FILLER_34_1402 ();
 sg13g2_decap_8 FILLER_34_1412 ();
 sg13g2_decap_8 FILLER_34_1419 ();
 sg13g2_decap_8 FILLER_34_1426 ();
 sg13g2_decap_8 FILLER_34_1433 ();
 sg13g2_decap_8 FILLER_34_1440 ();
 sg13g2_fill_2 FILLER_34_1447 ();
 sg13g2_fill_1 FILLER_34_1449 ();
 sg13g2_fill_2 FILLER_34_1456 ();
 sg13g2_fill_2 FILLER_34_1471 ();
 sg13g2_fill_1 FILLER_34_1473 ();
 sg13g2_decap_8 FILLER_34_1478 ();
 sg13g2_decap_8 FILLER_34_1485 ();
 sg13g2_decap_8 FILLER_34_1492 ();
 sg13g2_fill_2 FILLER_34_1499 ();
 sg13g2_decap_8 FILLER_34_1521 ();
 sg13g2_decap_8 FILLER_34_1528 ();
 sg13g2_decap_8 FILLER_34_1535 ();
 sg13g2_decap_8 FILLER_34_1542 ();
 sg13g2_decap_8 FILLER_34_1549 ();
 sg13g2_decap_8 FILLER_34_1556 ();
 sg13g2_decap_8 FILLER_34_1563 ();
 sg13g2_decap_8 FILLER_34_1570 ();
 sg13g2_decap_8 FILLER_34_1577 ();
 sg13g2_decap_8 FILLER_34_1584 ();
 sg13g2_decap_8 FILLER_34_1591 ();
 sg13g2_fill_2 FILLER_34_1598 ();
 sg13g2_fill_1 FILLER_34_1600 ();
 sg13g2_decap_8 FILLER_34_1606 ();
 sg13g2_decap_8 FILLER_34_1613 ();
 sg13g2_decap_8 FILLER_34_1620 ();
 sg13g2_decap_8 FILLER_34_1627 ();
 sg13g2_decap_8 FILLER_34_1634 ();
 sg13g2_decap_8 FILLER_34_1641 ();
 sg13g2_fill_2 FILLER_34_1648 ();
 sg13g2_fill_1 FILLER_34_1650 ();
 sg13g2_decap_8 FILLER_34_1657 ();
 sg13g2_decap_4 FILLER_34_1664 ();
 sg13g2_fill_1 FILLER_34_1668 ();
 sg13g2_decap_8 FILLER_34_1674 ();
 sg13g2_decap_8 FILLER_34_1681 ();
 sg13g2_decap_8 FILLER_34_1688 ();
 sg13g2_decap_8 FILLER_34_1695 ();
 sg13g2_fill_1 FILLER_34_1702 ();
 sg13g2_decap_8 FILLER_34_1715 ();
 sg13g2_decap_8 FILLER_34_1722 ();
 sg13g2_decap_8 FILLER_34_1729 ();
 sg13g2_fill_1 FILLER_34_1736 ();
 sg13g2_decap_8 FILLER_34_1747 ();
 sg13g2_decap_8 FILLER_34_1754 ();
 sg13g2_decap_8 FILLER_34_1761 ();
 sg13g2_fill_2 FILLER_34_1768 ();
 sg13g2_fill_1 FILLER_34_1770 ();
 sg13g2_decap_8 FILLER_34_1775 ();
 sg13g2_decap_8 FILLER_34_1782 ();
 sg13g2_decap_8 FILLER_34_1789 ();
 sg13g2_decap_8 FILLER_34_1796 ();
 sg13g2_decap_8 FILLER_34_1803 ();
 sg13g2_decap_8 FILLER_34_1810 ();
 sg13g2_decap_8 FILLER_34_1817 ();
 sg13g2_fill_2 FILLER_34_1837 ();
 sg13g2_decap_8 FILLER_34_1844 ();
 sg13g2_decap_8 FILLER_34_1851 ();
 sg13g2_decap_8 FILLER_34_1858 ();
 sg13g2_decap_8 FILLER_34_1865 ();
 sg13g2_decap_8 FILLER_34_1872 ();
 sg13g2_decap_8 FILLER_34_1879 ();
 sg13g2_decap_8 FILLER_34_1886 ();
 sg13g2_decap_8 FILLER_34_1893 ();
 sg13g2_decap_8 FILLER_34_1900 ();
 sg13g2_decap_8 FILLER_34_1907 ();
 sg13g2_decap_8 FILLER_34_1914 ();
 sg13g2_decap_8 FILLER_34_1921 ();
 sg13g2_decap_8 FILLER_34_1928 ();
 sg13g2_decap_8 FILLER_34_1935 ();
 sg13g2_decap_8 FILLER_34_1942 ();
 sg13g2_decap_8 FILLER_34_1949 ();
 sg13g2_decap_8 FILLER_34_1956 ();
 sg13g2_decap_8 FILLER_34_1963 ();
 sg13g2_decap_8 FILLER_34_1970 ();
 sg13g2_decap_8 FILLER_34_1977 ();
 sg13g2_decap_8 FILLER_34_1984 ();
 sg13g2_decap_8 FILLER_34_1991 ();
 sg13g2_decap_8 FILLER_34_1998 ();
 sg13g2_decap_8 FILLER_34_2005 ();
 sg13g2_decap_8 FILLER_34_2012 ();
 sg13g2_decap_8 FILLER_34_2019 ();
 sg13g2_decap_8 FILLER_34_2026 ();
 sg13g2_decap_8 FILLER_34_2033 ();
 sg13g2_decap_8 FILLER_34_2040 ();
 sg13g2_decap_8 FILLER_34_2047 ();
 sg13g2_decap_8 FILLER_34_2054 ();
 sg13g2_decap_8 FILLER_34_2061 ();
 sg13g2_decap_8 FILLER_34_2068 ();
 sg13g2_decap_8 FILLER_34_2075 ();
 sg13g2_decap_8 FILLER_34_2082 ();
 sg13g2_decap_8 FILLER_34_2089 ();
 sg13g2_decap_8 FILLER_34_2096 ();
 sg13g2_decap_8 FILLER_34_2103 ();
 sg13g2_decap_8 FILLER_34_2110 ();
 sg13g2_decap_8 FILLER_34_2117 ();
 sg13g2_decap_8 FILLER_34_2124 ();
 sg13g2_decap_8 FILLER_34_2131 ();
 sg13g2_decap_8 FILLER_34_2138 ();
 sg13g2_decap_8 FILLER_34_2145 ();
 sg13g2_decap_8 FILLER_34_2152 ();
 sg13g2_decap_8 FILLER_34_2159 ();
 sg13g2_decap_8 FILLER_34_2166 ();
 sg13g2_decap_8 FILLER_34_2173 ();
 sg13g2_decap_8 FILLER_34_2180 ();
 sg13g2_decap_8 FILLER_34_2187 ();
 sg13g2_decap_8 FILLER_34_2194 ();
 sg13g2_decap_8 FILLER_34_2201 ();
 sg13g2_decap_8 FILLER_34_2208 ();
 sg13g2_decap_8 FILLER_34_2215 ();
 sg13g2_decap_8 FILLER_34_2222 ();
 sg13g2_decap_8 FILLER_34_2229 ();
 sg13g2_decap_8 FILLER_34_2236 ();
 sg13g2_decap_8 FILLER_34_2243 ();
 sg13g2_decap_8 FILLER_34_2250 ();
 sg13g2_decap_8 FILLER_34_2257 ();
 sg13g2_decap_8 FILLER_34_2264 ();
 sg13g2_decap_8 FILLER_34_2271 ();
 sg13g2_decap_8 FILLER_34_2278 ();
 sg13g2_decap_8 FILLER_34_2285 ();
 sg13g2_decap_8 FILLER_34_2292 ();
 sg13g2_decap_8 FILLER_34_2299 ();
 sg13g2_decap_8 FILLER_34_2306 ();
 sg13g2_decap_8 FILLER_34_2313 ();
 sg13g2_decap_8 FILLER_34_2320 ();
 sg13g2_decap_8 FILLER_34_2327 ();
 sg13g2_decap_8 FILLER_34_2334 ();
 sg13g2_decap_8 FILLER_34_2341 ();
 sg13g2_decap_8 FILLER_34_2348 ();
 sg13g2_decap_8 FILLER_34_2355 ();
 sg13g2_decap_8 FILLER_34_2362 ();
 sg13g2_decap_8 FILLER_34_2369 ();
 sg13g2_decap_8 FILLER_34_2376 ();
 sg13g2_decap_8 FILLER_34_2383 ();
 sg13g2_decap_8 FILLER_34_2390 ();
 sg13g2_decap_8 FILLER_34_2397 ();
 sg13g2_decap_8 FILLER_34_2404 ();
 sg13g2_decap_8 FILLER_34_2411 ();
 sg13g2_decap_8 FILLER_34_2418 ();
 sg13g2_decap_8 FILLER_34_2425 ();
 sg13g2_decap_8 FILLER_34_2432 ();
 sg13g2_decap_8 FILLER_34_2439 ();
 sg13g2_decap_8 FILLER_34_2446 ();
 sg13g2_decap_8 FILLER_34_2453 ();
 sg13g2_decap_8 FILLER_34_2460 ();
 sg13g2_decap_8 FILLER_34_2467 ();
 sg13g2_decap_8 FILLER_34_2474 ();
 sg13g2_decap_8 FILLER_34_2481 ();
 sg13g2_decap_8 FILLER_34_2488 ();
 sg13g2_decap_8 FILLER_34_2495 ();
 sg13g2_decap_8 FILLER_34_2502 ();
 sg13g2_decap_8 FILLER_34_2509 ();
 sg13g2_decap_8 FILLER_34_2516 ();
 sg13g2_decap_8 FILLER_34_2523 ();
 sg13g2_decap_8 FILLER_34_2530 ();
 sg13g2_decap_8 FILLER_34_2537 ();
 sg13g2_decap_8 FILLER_34_2544 ();
 sg13g2_decap_8 FILLER_34_2551 ();
 sg13g2_decap_8 FILLER_34_2558 ();
 sg13g2_decap_8 FILLER_34_2565 ();
 sg13g2_decap_8 FILLER_34_2572 ();
 sg13g2_decap_8 FILLER_34_2579 ();
 sg13g2_decap_8 FILLER_34_2586 ();
 sg13g2_decap_8 FILLER_34_2593 ();
 sg13g2_decap_8 FILLER_34_2600 ();
 sg13g2_decap_8 FILLER_34_2607 ();
 sg13g2_decap_8 FILLER_34_2614 ();
 sg13g2_decap_8 FILLER_34_2621 ();
 sg13g2_decap_8 FILLER_34_2628 ();
 sg13g2_decap_8 FILLER_34_2635 ();
 sg13g2_decap_8 FILLER_34_2642 ();
 sg13g2_decap_8 FILLER_34_2649 ();
 sg13g2_decap_8 FILLER_34_2656 ();
 sg13g2_decap_8 FILLER_34_2663 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_65 ();
 sg13g2_decap_8 FILLER_35_72 ();
 sg13g2_decap_8 FILLER_35_79 ();
 sg13g2_decap_8 FILLER_35_86 ();
 sg13g2_decap_8 FILLER_35_93 ();
 sg13g2_decap_8 FILLER_35_100 ();
 sg13g2_decap_8 FILLER_35_107 ();
 sg13g2_decap_8 FILLER_35_114 ();
 sg13g2_decap_8 FILLER_35_121 ();
 sg13g2_decap_8 FILLER_35_128 ();
 sg13g2_decap_8 FILLER_35_135 ();
 sg13g2_decap_8 FILLER_35_142 ();
 sg13g2_decap_8 FILLER_35_149 ();
 sg13g2_decap_8 FILLER_35_156 ();
 sg13g2_decap_8 FILLER_35_163 ();
 sg13g2_decap_8 FILLER_35_170 ();
 sg13g2_decap_8 FILLER_35_177 ();
 sg13g2_decap_8 FILLER_35_184 ();
 sg13g2_decap_4 FILLER_35_191 ();
 sg13g2_decap_8 FILLER_35_221 ();
 sg13g2_decap_8 FILLER_35_228 ();
 sg13g2_decap_8 FILLER_35_235 ();
 sg13g2_decap_8 FILLER_35_242 ();
 sg13g2_decap_8 FILLER_35_249 ();
 sg13g2_decap_8 FILLER_35_256 ();
 sg13g2_decap_8 FILLER_35_263 ();
 sg13g2_decap_4 FILLER_35_270 ();
 sg13g2_decap_8 FILLER_35_280 ();
 sg13g2_decap_8 FILLER_35_287 ();
 sg13g2_decap_8 FILLER_35_294 ();
 sg13g2_decap_8 FILLER_35_301 ();
 sg13g2_decap_8 FILLER_35_308 ();
 sg13g2_decap_8 FILLER_35_315 ();
 sg13g2_decap_8 FILLER_35_322 ();
 sg13g2_decap_8 FILLER_35_329 ();
 sg13g2_decap_8 FILLER_35_336 ();
 sg13g2_decap_8 FILLER_35_343 ();
 sg13g2_decap_8 FILLER_35_350 ();
 sg13g2_decap_8 FILLER_35_357 ();
 sg13g2_decap_8 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_371 ();
 sg13g2_decap_4 FILLER_35_378 ();
 sg13g2_fill_1 FILLER_35_382 ();
 sg13g2_fill_2 FILLER_35_393 ();
 sg13g2_decap_8 FILLER_35_399 ();
 sg13g2_decap_8 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_413 ();
 sg13g2_decap_8 FILLER_35_429 ();
 sg13g2_decap_8 FILLER_35_436 ();
 sg13g2_decap_8 FILLER_35_443 ();
 sg13g2_decap_8 FILLER_35_450 ();
 sg13g2_decap_8 FILLER_35_457 ();
 sg13g2_decap_8 FILLER_35_464 ();
 sg13g2_decap_8 FILLER_35_471 ();
 sg13g2_decap_4 FILLER_35_478 ();
 sg13g2_decap_8 FILLER_35_486 ();
 sg13g2_decap_8 FILLER_35_493 ();
 sg13g2_decap_8 FILLER_35_500 ();
 sg13g2_decap_8 FILLER_35_507 ();
 sg13g2_decap_4 FILLER_35_514 ();
 sg13g2_fill_2 FILLER_35_518 ();
 sg13g2_fill_1 FILLER_35_535 ();
 sg13g2_decap_8 FILLER_35_539 ();
 sg13g2_decap_4 FILLER_35_546 ();
 sg13g2_fill_1 FILLER_35_550 ();
 sg13g2_decap_8 FILLER_35_554 ();
 sg13g2_fill_2 FILLER_35_561 ();
 sg13g2_fill_1 FILLER_35_563 ();
 sg13g2_decap_8 FILLER_35_569 ();
 sg13g2_decap_8 FILLER_35_576 ();
 sg13g2_decap_8 FILLER_35_583 ();
 sg13g2_decap_8 FILLER_35_590 ();
 sg13g2_decap_8 FILLER_35_597 ();
 sg13g2_decap_8 FILLER_35_604 ();
 sg13g2_decap_8 FILLER_35_611 ();
 sg13g2_decap_8 FILLER_35_618 ();
 sg13g2_decap_8 FILLER_35_625 ();
 sg13g2_decap_8 FILLER_35_632 ();
 sg13g2_decap_8 FILLER_35_639 ();
 sg13g2_decap_8 FILLER_35_646 ();
 sg13g2_decap_8 FILLER_35_653 ();
 sg13g2_decap_8 FILLER_35_660 ();
 sg13g2_fill_2 FILLER_35_667 ();
 sg13g2_fill_1 FILLER_35_669 ();
 sg13g2_decap_8 FILLER_35_673 ();
 sg13g2_decap_8 FILLER_35_684 ();
 sg13g2_decap_8 FILLER_35_691 ();
 sg13g2_decap_8 FILLER_35_698 ();
 sg13g2_decap_8 FILLER_35_705 ();
 sg13g2_decap_4 FILLER_35_712 ();
 sg13g2_fill_1 FILLER_35_716 ();
 sg13g2_decap_8 FILLER_35_720 ();
 sg13g2_decap_4 FILLER_35_727 ();
 sg13g2_fill_1 FILLER_35_731 ();
 sg13g2_decap_8 FILLER_35_736 ();
 sg13g2_decap_8 FILLER_35_743 ();
 sg13g2_decap_8 FILLER_35_750 ();
 sg13g2_decap_8 FILLER_35_757 ();
 sg13g2_decap_8 FILLER_35_764 ();
 sg13g2_decap_4 FILLER_35_771 ();
 sg13g2_fill_2 FILLER_35_775 ();
 sg13g2_fill_1 FILLER_35_785 ();
 sg13g2_decap_8 FILLER_35_809 ();
 sg13g2_decap_8 FILLER_35_816 ();
 sg13g2_fill_2 FILLER_35_823 ();
 sg13g2_fill_1 FILLER_35_825 ();
 sg13g2_fill_2 FILLER_35_831 ();
 sg13g2_fill_1 FILLER_35_838 ();
 sg13g2_fill_2 FILLER_35_844 ();
 sg13g2_decap_8 FILLER_35_851 ();
 sg13g2_decap_8 FILLER_35_858 ();
 sg13g2_decap_8 FILLER_35_865 ();
 sg13g2_decap_8 FILLER_35_872 ();
 sg13g2_decap_8 FILLER_35_879 ();
 sg13g2_decap_8 FILLER_35_886 ();
 sg13g2_decap_8 FILLER_35_893 ();
 sg13g2_decap_8 FILLER_35_900 ();
 sg13g2_decap_8 FILLER_35_907 ();
 sg13g2_decap_8 FILLER_35_914 ();
 sg13g2_decap_8 FILLER_35_921 ();
 sg13g2_decap_8 FILLER_35_928 ();
 sg13g2_decap_8 FILLER_35_935 ();
 sg13g2_decap_8 FILLER_35_942 ();
 sg13g2_decap_8 FILLER_35_949 ();
 sg13g2_decap_8 FILLER_35_956 ();
 sg13g2_decap_8 FILLER_35_963 ();
 sg13g2_decap_8 FILLER_35_970 ();
 sg13g2_decap_8 FILLER_35_977 ();
 sg13g2_decap_8 FILLER_35_984 ();
 sg13g2_fill_1 FILLER_35_991 ();
 sg13g2_decap_8 FILLER_35_1001 ();
 sg13g2_decap_8 FILLER_35_1008 ();
 sg13g2_decap_8 FILLER_35_1015 ();
 sg13g2_decap_8 FILLER_35_1022 ();
 sg13g2_decap_8 FILLER_35_1029 ();
 sg13g2_decap_8 FILLER_35_1036 ();
 sg13g2_decap_4 FILLER_35_1043 ();
 sg13g2_fill_2 FILLER_35_1047 ();
 sg13g2_decap_8 FILLER_35_1063 ();
 sg13g2_decap_8 FILLER_35_1070 ();
 sg13g2_decap_8 FILLER_35_1077 ();
 sg13g2_decap_8 FILLER_35_1084 ();
 sg13g2_decap_8 FILLER_35_1091 ();
 sg13g2_decap_8 FILLER_35_1098 ();
 sg13g2_decap_8 FILLER_35_1105 ();
 sg13g2_decap_8 FILLER_35_1112 ();
 sg13g2_fill_2 FILLER_35_1119 ();
 sg13g2_decap_8 FILLER_35_1154 ();
 sg13g2_decap_8 FILLER_35_1161 ();
 sg13g2_decap_4 FILLER_35_1168 ();
 sg13g2_decap_8 FILLER_35_1177 ();
 sg13g2_decap_8 FILLER_35_1184 ();
 sg13g2_decap_8 FILLER_35_1191 ();
 sg13g2_decap_8 FILLER_35_1198 ();
 sg13g2_decap_8 FILLER_35_1205 ();
 sg13g2_fill_2 FILLER_35_1212 ();
 sg13g2_fill_1 FILLER_35_1218 ();
 sg13g2_decap_8 FILLER_35_1234 ();
 sg13g2_decap_8 FILLER_35_1241 ();
 sg13g2_decap_8 FILLER_35_1248 ();
 sg13g2_decap_4 FILLER_35_1255 ();
 sg13g2_fill_1 FILLER_35_1259 ();
 sg13g2_fill_1 FILLER_35_1270 ();
 sg13g2_decap_8 FILLER_35_1277 ();
 sg13g2_decap_8 FILLER_35_1284 ();
 sg13g2_decap_8 FILLER_35_1291 ();
 sg13g2_decap_8 FILLER_35_1298 ();
 sg13g2_decap_8 FILLER_35_1305 ();
 sg13g2_decap_4 FILLER_35_1312 ();
 sg13g2_fill_2 FILLER_35_1316 ();
 sg13g2_decap_8 FILLER_35_1321 ();
 sg13g2_decap_8 FILLER_35_1328 ();
 sg13g2_decap_8 FILLER_35_1335 ();
 sg13g2_decap_8 FILLER_35_1342 ();
 sg13g2_decap_8 FILLER_35_1349 ();
 sg13g2_decap_8 FILLER_35_1356 ();
 sg13g2_decap_8 FILLER_35_1363 ();
 sg13g2_decap_8 FILLER_35_1370 ();
 sg13g2_decap_8 FILLER_35_1377 ();
 sg13g2_decap_8 FILLER_35_1384 ();
 sg13g2_decap_8 FILLER_35_1391 ();
 sg13g2_decap_8 FILLER_35_1405 ();
 sg13g2_decap_8 FILLER_35_1412 ();
 sg13g2_decap_8 FILLER_35_1419 ();
 sg13g2_decap_8 FILLER_35_1426 ();
 sg13g2_decap_8 FILLER_35_1433 ();
 sg13g2_decap_8 FILLER_35_1440 ();
 sg13g2_decap_8 FILLER_35_1466 ();
 sg13g2_decap_8 FILLER_35_1473 ();
 sg13g2_decap_8 FILLER_35_1480 ();
 sg13g2_decap_4 FILLER_35_1487 ();
 sg13g2_fill_2 FILLER_35_1491 ();
 sg13g2_decap_8 FILLER_35_1504 ();
 sg13g2_decap_8 FILLER_35_1511 ();
 sg13g2_decap_8 FILLER_35_1518 ();
 sg13g2_decap_8 FILLER_35_1525 ();
 sg13g2_decap_8 FILLER_35_1532 ();
 sg13g2_decap_8 FILLER_35_1539 ();
 sg13g2_decap_8 FILLER_35_1549 ();
 sg13g2_decap_8 FILLER_35_1556 ();
 sg13g2_decap_8 FILLER_35_1563 ();
 sg13g2_decap_8 FILLER_35_1570 ();
 sg13g2_decap_8 FILLER_35_1581 ();
 sg13g2_decap_8 FILLER_35_1588 ();
 sg13g2_decap_8 FILLER_35_1595 ();
 sg13g2_fill_1 FILLER_35_1602 ();
 sg13g2_decap_8 FILLER_35_1607 ();
 sg13g2_decap_8 FILLER_35_1614 ();
 sg13g2_decap_4 FILLER_35_1621 ();
 sg13g2_fill_1 FILLER_35_1625 ();
 sg13g2_decap_8 FILLER_35_1630 ();
 sg13g2_decap_8 FILLER_35_1637 ();
 sg13g2_decap_8 FILLER_35_1644 ();
 sg13g2_decap_8 FILLER_35_1651 ();
 sg13g2_decap_8 FILLER_35_1658 ();
 sg13g2_decap_8 FILLER_35_1665 ();
 sg13g2_decap_8 FILLER_35_1672 ();
 sg13g2_decap_8 FILLER_35_1679 ();
 sg13g2_decap_8 FILLER_35_1686 ();
 sg13g2_decap_8 FILLER_35_1693 ();
 sg13g2_decap_8 FILLER_35_1700 ();
 sg13g2_decap_8 FILLER_35_1707 ();
 sg13g2_decap_8 FILLER_35_1714 ();
 sg13g2_decap_8 FILLER_35_1721 ();
 sg13g2_decap_8 FILLER_35_1728 ();
 sg13g2_decap_8 FILLER_35_1735 ();
 sg13g2_decap_8 FILLER_35_1742 ();
 sg13g2_fill_1 FILLER_35_1749 ();
 sg13g2_decap_8 FILLER_35_1754 ();
 sg13g2_decap_8 FILLER_35_1761 ();
 sg13g2_decap_8 FILLER_35_1768 ();
 sg13g2_decap_8 FILLER_35_1775 ();
 sg13g2_decap_8 FILLER_35_1782 ();
 sg13g2_decap_8 FILLER_35_1789 ();
 sg13g2_decap_8 FILLER_35_1796 ();
 sg13g2_decap_8 FILLER_35_1803 ();
 sg13g2_decap_8 FILLER_35_1810 ();
 sg13g2_decap_8 FILLER_35_1817 ();
 sg13g2_decap_8 FILLER_35_1824 ();
 sg13g2_decap_8 FILLER_35_1831 ();
 sg13g2_decap_8 FILLER_35_1838 ();
 sg13g2_decap_8 FILLER_35_1845 ();
 sg13g2_decap_4 FILLER_35_1852 ();
 sg13g2_fill_2 FILLER_35_1856 ();
 sg13g2_decap_8 FILLER_35_1875 ();
 sg13g2_decap_8 FILLER_35_1882 ();
 sg13g2_decap_8 FILLER_35_1889 ();
 sg13g2_decap_8 FILLER_35_1896 ();
 sg13g2_decap_8 FILLER_35_1903 ();
 sg13g2_decap_8 FILLER_35_1910 ();
 sg13g2_decap_8 FILLER_35_1917 ();
 sg13g2_decap_8 FILLER_35_1924 ();
 sg13g2_decap_8 FILLER_35_1931 ();
 sg13g2_decap_8 FILLER_35_1938 ();
 sg13g2_decap_8 FILLER_35_1945 ();
 sg13g2_decap_8 FILLER_35_1952 ();
 sg13g2_decap_8 FILLER_35_1959 ();
 sg13g2_decap_8 FILLER_35_1966 ();
 sg13g2_decap_8 FILLER_35_1973 ();
 sg13g2_decap_8 FILLER_35_1980 ();
 sg13g2_decap_8 FILLER_35_1987 ();
 sg13g2_decap_8 FILLER_35_1994 ();
 sg13g2_decap_8 FILLER_35_2001 ();
 sg13g2_decap_8 FILLER_35_2008 ();
 sg13g2_decap_8 FILLER_35_2015 ();
 sg13g2_decap_8 FILLER_35_2022 ();
 sg13g2_decap_8 FILLER_35_2029 ();
 sg13g2_decap_8 FILLER_35_2036 ();
 sg13g2_decap_8 FILLER_35_2043 ();
 sg13g2_decap_8 FILLER_35_2050 ();
 sg13g2_decap_8 FILLER_35_2057 ();
 sg13g2_decap_8 FILLER_35_2064 ();
 sg13g2_decap_8 FILLER_35_2071 ();
 sg13g2_decap_8 FILLER_35_2078 ();
 sg13g2_decap_8 FILLER_35_2085 ();
 sg13g2_decap_8 FILLER_35_2092 ();
 sg13g2_decap_8 FILLER_35_2099 ();
 sg13g2_decap_8 FILLER_35_2106 ();
 sg13g2_decap_8 FILLER_35_2113 ();
 sg13g2_decap_8 FILLER_35_2120 ();
 sg13g2_decap_8 FILLER_35_2127 ();
 sg13g2_decap_8 FILLER_35_2134 ();
 sg13g2_decap_8 FILLER_35_2141 ();
 sg13g2_decap_8 FILLER_35_2148 ();
 sg13g2_decap_8 FILLER_35_2155 ();
 sg13g2_decap_8 FILLER_35_2162 ();
 sg13g2_decap_8 FILLER_35_2169 ();
 sg13g2_decap_8 FILLER_35_2176 ();
 sg13g2_decap_8 FILLER_35_2183 ();
 sg13g2_decap_8 FILLER_35_2190 ();
 sg13g2_decap_8 FILLER_35_2197 ();
 sg13g2_decap_8 FILLER_35_2204 ();
 sg13g2_decap_8 FILLER_35_2211 ();
 sg13g2_decap_8 FILLER_35_2218 ();
 sg13g2_decap_8 FILLER_35_2225 ();
 sg13g2_decap_8 FILLER_35_2232 ();
 sg13g2_decap_8 FILLER_35_2239 ();
 sg13g2_decap_8 FILLER_35_2246 ();
 sg13g2_decap_8 FILLER_35_2253 ();
 sg13g2_decap_8 FILLER_35_2260 ();
 sg13g2_decap_8 FILLER_35_2267 ();
 sg13g2_decap_8 FILLER_35_2274 ();
 sg13g2_decap_8 FILLER_35_2281 ();
 sg13g2_decap_8 FILLER_35_2288 ();
 sg13g2_decap_8 FILLER_35_2295 ();
 sg13g2_decap_8 FILLER_35_2302 ();
 sg13g2_decap_8 FILLER_35_2309 ();
 sg13g2_decap_8 FILLER_35_2316 ();
 sg13g2_decap_8 FILLER_35_2323 ();
 sg13g2_decap_8 FILLER_35_2330 ();
 sg13g2_decap_8 FILLER_35_2337 ();
 sg13g2_decap_8 FILLER_35_2344 ();
 sg13g2_decap_8 FILLER_35_2351 ();
 sg13g2_decap_8 FILLER_35_2358 ();
 sg13g2_decap_8 FILLER_35_2365 ();
 sg13g2_decap_8 FILLER_35_2372 ();
 sg13g2_decap_8 FILLER_35_2379 ();
 sg13g2_decap_8 FILLER_35_2386 ();
 sg13g2_decap_8 FILLER_35_2393 ();
 sg13g2_decap_8 FILLER_35_2400 ();
 sg13g2_decap_8 FILLER_35_2407 ();
 sg13g2_decap_8 FILLER_35_2414 ();
 sg13g2_decap_8 FILLER_35_2421 ();
 sg13g2_decap_8 FILLER_35_2428 ();
 sg13g2_decap_8 FILLER_35_2435 ();
 sg13g2_decap_8 FILLER_35_2442 ();
 sg13g2_decap_8 FILLER_35_2449 ();
 sg13g2_decap_8 FILLER_35_2456 ();
 sg13g2_decap_8 FILLER_35_2463 ();
 sg13g2_decap_8 FILLER_35_2470 ();
 sg13g2_decap_8 FILLER_35_2477 ();
 sg13g2_decap_8 FILLER_35_2484 ();
 sg13g2_decap_8 FILLER_35_2491 ();
 sg13g2_decap_8 FILLER_35_2498 ();
 sg13g2_decap_8 FILLER_35_2505 ();
 sg13g2_decap_8 FILLER_35_2512 ();
 sg13g2_decap_8 FILLER_35_2519 ();
 sg13g2_decap_8 FILLER_35_2526 ();
 sg13g2_decap_8 FILLER_35_2533 ();
 sg13g2_decap_8 FILLER_35_2540 ();
 sg13g2_decap_8 FILLER_35_2547 ();
 sg13g2_decap_8 FILLER_35_2554 ();
 sg13g2_decap_8 FILLER_35_2561 ();
 sg13g2_decap_8 FILLER_35_2568 ();
 sg13g2_decap_8 FILLER_35_2575 ();
 sg13g2_decap_8 FILLER_35_2582 ();
 sg13g2_decap_8 FILLER_35_2589 ();
 sg13g2_decap_8 FILLER_35_2596 ();
 sg13g2_decap_8 FILLER_35_2603 ();
 sg13g2_decap_8 FILLER_35_2610 ();
 sg13g2_decap_8 FILLER_35_2617 ();
 sg13g2_decap_8 FILLER_35_2624 ();
 sg13g2_decap_8 FILLER_35_2631 ();
 sg13g2_decap_8 FILLER_35_2638 ();
 sg13g2_decap_8 FILLER_35_2645 ();
 sg13g2_decap_8 FILLER_35_2652 ();
 sg13g2_decap_8 FILLER_35_2659 ();
 sg13g2_decap_4 FILLER_35_2666 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_fill_2 FILLER_36_119 ();
 sg13g2_fill_1 FILLER_36_121 ();
 sg13g2_decap_8 FILLER_36_127 ();
 sg13g2_decap_8 FILLER_36_134 ();
 sg13g2_decap_4 FILLER_36_141 ();
 sg13g2_fill_2 FILLER_36_145 ();
 sg13g2_decap_8 FILLER_36_151 ();
 sg13g2_decap_8 FILLER_36_158 ();
 sg13g2_decap_8 FILLER_36_165 ();
 sg13g2_decap_8 FILLER_36_172 ();
 sg13g2_decap_8 FILLER_36_179 ();
 sg13g2_decap_8 FILLER_36_186 ();
 sg13g2_decap_8 FILLER_36_193 ();
 sg13g2_decap_8 FILLER_36_200 ();
 sg13g2_decap_8 FILLER_36_207 ();
 sg13g2_decap_8 FILLER_36_214 ();
 sg13g2_decap_8 FILLER_36_221 ();
 sg13g2_decap_8 FILLER_36_228 ();
 sg13g2_decap_8 FILLER_36_235 ();
 sg13g2_decap_8 FILLER_36_242 ();
 sg13g2_decap_8 FILLER_36_249 ();
 sg13g2_decap_8 FILLER_36_256 ();
 sg13g2_decap_8 FILLER_36_263 ();
 sg13g2_fill_1 FILLER_36_276 ();
 sg13g2_decap_8 FILLER_36_287 ();
 sg13g2_decap_8 FILLER_36_294 ();
 sg13g2_decap_8 FILLER_36_301 ();
 sg13g2_decap_8 FILLER_36_308 ();
 sg13g2_decap_8 FILLER_36_315 ();
 sg13g2_fill_1 FILLER_36_322 ();
 sg13g2_decap_8 FILLER_36_327 ();
 sg13g2_decap_8 FILLER_36_334 ();
 sg13g2_fill_2 FILLER_36_341 ();
 sg13g2_fill_1 FILLER_36_343 ();
 sg13g2_fill_2 FILLER_36_351 ();
 sg13g2_fill_1 FILLER_36_353 ();
 sg13g2_fill_1 FILLER_36_377 ();
 sg13g2_decap_8 FILLER_36_387 ();
 sg13g2_decap_8 FILLER_36_394 ();
 sg13g2_fill_1 FILLER_36_401 ();
 sg13g2_decap_8 FILLER_36_425 ();
 sg13g2_fill_2 FILLER_36_436 ();
 sg13g2_fill_1 FILLER_36_438 ();
 sg13g2_decap_8 FILLER_36_465 ();
 sg13g2_decap_8 FILLER_36_472 ();
 sg13g2_decap_8 FILLER_36_479 ();
 sg13g2_decap_8 FILLER_36_486 ();
 sg13g2_decap_8 FILLER_36_493 ();
 sg13g2_decap_8 FILLER_36_500 ();
 sg13g2_decap_8 FILLER_36_507 ();
 sg13g2_decap_8 FILLER_36_514 ();
 sg13g2_decap_4 FILLER_36_521 ();
 sg13g2_fill_1 FILLER_36_525 ();
 sg13g2_fill_2 FILLER_36_530 ();
 sg13g2_fill_1 FILLER_36_532 ();
 sg13g2_decap_8 FILLER_36_537 ();
 sg13g2_decap_8 FILLER_36_544 ();
 sg13g2_decap_8 FILLER_36_551 ();
 sg13g2_decap_8 FILLER_36_558 ();
 sg13g2_decap_8 FILLER_36_565 ();
 sg13g2_decap_8 FILLER_36_572 ();
 sg13g2_decap_8 FILLER_36_579 ();
 sg13g2_decap_8 FILLER_36_586 ();
 sg13g2_decap_8 FILLER_36_593 ();
 sg13g2_decap_8 FILLER_36_600 ();
 sg13g2_decap_8 FILLER_36_607 ();
 sg13g2_fill_1 FILLER_36_614 ();
 sg13g2_decap_4 FILLER_36_620 ();
 sg13g2_fill_2 FILLER_36_624 ();
 sg13g2_decap_4 FILLER_36_631 ();
 sg13g2_fill_1 FILLER_36_635 ();
 sg13g2_decap_8 FILLER_36_641 ();
 sg13g2_decap_8 FILLER_36_648 ();
 sg13g2_fill_2 FILLER_36_655 ();
 sg13g2_fill_1 FILLER_36_657 ();
 sg13g2_fill_1 FILLER_36_667 ();
 sg13g2_fill_1 FILLER_36_683 ();
 sg13g2_decap_8 FILLER_36_702 ();
 sg13g2_fill_2 FILLER_36_709 ();
 sg13g2_fill_1 FILLER_36_711 ();
 sg13g2_decap_8 FILLER_36_733 ();
 sg13g2_decap_8 FILLER_36_740 ();
 sg13g2_decap_8 FILLER_36_747 ();
 sg13g2_decap_8 FILLER_36_754 ();
 sg13g2_decap_8 FILLER_36_761 ();
 sg13g2_decap_8 FILLER_36_768 ();
 sg13g2_decap_4 FILLER_36_775 ();
 sg13g2_fill_1 FILLER_36_779 ();
 sg13g2_decap_4 FILLER_36_783 ();
 sg13g2_decap_4 FILLER_36_790 ();
 sg13g2_fill_1 FILLER_36_794 ();
 sg13g2_decap_8 FILLER_36_803 ();
 sg13g2_decap_8 FILLER_36_810 ();
 sg13g2_decap_8 FILLER_36_817 ();
 sg13g2_decap_4 FILLER_36_824 ();
 sg13g2_fill_2 FILLER_36_828 ();
 sg13g2_fill_1 FILLER_36_838 ();
 sg13g2_fill_1 FILLER_36_845 ();
 sg13g2_decap_8 FILLER_36_849 ();
 sg13g2_decap_8 FILLER_36_856 ();
 sg13g2_decap_8 FILLER_36_863 ();
 sg13g2_decap_8 FILLER_36_870 ();
 sg13g2_decap_8 FILLER_36_877 ();
 sg13g2_decap_8 FILLER_36_884 ();
 sg13g2_decap_8 FILLER_36_891 ();
 sg13g2_decap_8 FILLER_36_898 ();
 sg13g2_decap_4 FILLER_36_905 ();
 sg13g2_fill_1 FILLER_36_909 ();
 sg13g2_decap_8 FILLER_36_913 ();
 sg13g2_fill_1 FILLER_36_920 ();
 sg13g2_decap_8 FILLER_36_928 ();
 sg13g2_decap_8 FILLER_36_935 ();
 sg13g2_fill_2 FILLER_36_942 ();
 sg13g2_fill_1 FILLER_36_944 ();
 sg13g2_decap_8 FILLER_36_949 ();
 sg13g2_decap_8 FILLER_36_956 ();
 sg13g2_decap_8 FILLER_36_963 ();
 sg13g2_decap_8 FILLER_36_970 ();
 sg13g2_decap_8 FILLER_36_977 ();
 sg13g2_decap_4 FILLER_36_984 ();
 sg13g2_fill_2 FILLER_36_988 ();
 sg13g2_decap_8 FILLER_36_994 ();
 sg13g2_decap_8 FILLER_36_1001 ();
 sg13g2_decap_8 FILLER_36_1008 ();
 sg13g2_decap_8 FILLER_36_1015 ();
 sg13g2_decap_8 FILLER_36_1022 ();
 sg13g2_decap_4 FILLER_36_1029 ();
 sg13g2_fill_1 FILLER_36_1033 ();
 sg13g2_decap_4 FILLER_36_1046 ();
 sg13g2_fill_1 FILLER_36_1050 ();
 sg13g2_decap_8 FILLER_36_1076 ();
 sg13g2_fill_2 FILLER_36_1083 ();
 sg13g2_fill_1 FILLER_36_1085 ();
 sg13g2_decap_8 FILLER_36_1091 ();
 sg13g2_decap_8 FILLER_36_1098 ();
 sg13g2_decap_8 FILLER_36_1105 ();
 sg13g2_decap_8 FILLER_36_1112 ();
 sg13g2_fill_2 FILLER_36_1119 ();
 sg13g2_fill_1 FILLER_36_1121 ();
 sg13g2_fill_2 FILLER_36_1137 ();
 sg13g2_decap_8 FILLER_36_1149 ();
 sg13g2_decap_8 FILLER_36_1156 ();
 sg13g2_decap_8 FILLER_36_1163 ();
 sg13g2_decap_8 FILLER_36_1170 ();
 sg13g2_decap_8 FILLER_36_1177 ();
 sg13g2_decap_8 FILLER_36_1184 ();
 sg13g2_decap_8 FILLER_36_1191 ();
 sg13g2_decap_8 FILLER_36_1198 ();
 sg13g2_decap_8 FILLER_36_1205 ();
 sg13g2_decap_4 FILLER_36_1212 ();
 sg13g2_fill_1 FILLER_36_1216 ();
 sg13g2_fill_2 FILLER_36_1228 ();
 sg13g2_decap_8 FILLER_36_1234 ();
 sg13g2_decap_8 FILLER_36_1241 ();
 sg13g2_decap_8 FILLER_36_1248 ();
 sg13g2_fill_2 FILLER_36_1264 ();
 sg13g2_decap_8 FILLER_36_1273 ();
 sg13g2_decap_8 FILLER_36_1280 ();
 sg13g2_decap_8 FILLER_36_1287 ();
 sg13g2_decap_8 FILLER_36_1294 ();
 sg13g2_decap_8 FILLER_36_1301 ();
 sg13g2_decap_8 FILLER_36_1308 ();
 sg13g2_decap_8 FILLER_36_1315 ();
 sg13g2_decap_8 FILLER_36_1322 ();
 sg13g2_decap_8 FILLER_36_1329 ();
 sg13g2_decap_8 FILLER_36_1336 ();
 sg13g2_decap_8 FILLER_36_1343 ();
 sg13g2_decap_8 FILLER_36_1350 ();
 sg13g2_decap_4 FILLER_36_1357 ();
 sg13g2_fill_1 FILLER_36_1361 ();
 sg13g2_decap_8 FILLER_36_1366 ();
 sg13g2_decap_8 FILLER_36_1373 ();
 sg13g2_decap_8 FILLER_36_1380 ();
 sg13g2_decap_4 FILLER_36_1387 ();
 sg13g2_decap_8 FILLER_36_1403 ();
 sg13g2_decap_8 FILLER_36_1410 ();
 sg13g2_decap_8 FILLER_36_1417 ();
 sg13g2_decap_8 FILLER_36_1424 ();
 sg13g2_decap_8 FILLER_36_1431 ();
 sg13g2_decap_8 FILLER_36_1438 ();
 sg13g2_fill_2 FILLER_36_1445 ();
 sg13g2_fill_1 FILLER_36_1456 ();
 sg13g2_fill_2 FILLER_36_1460 ();
 sg13g2_fill_1 FILLER_36_1470 ();
 sg13g2_decap_8 FILLER_36_1475 ();
 sg13g2_decap_8 FILLER_36_1482 ();
 sg13g2_decap_8 FILLER_36_1489 ();
 sg13g2_decap_4 FILLER_36_1496 ();
 sg13g2_fill_1 FILLER_36_1500 ();
 sg13g2_decap_8 FILLER_36_1505 ();
 sg13g2_decap_8 FILLER_36_1512 ();
 sg13g2_decap_8 FILLER_36_1519 ();
 sg13g2_decap_8 FILLER_36_1526 ();
 sg13g2_decap_8 FILLER_36_1533 ();
 sg13g2_decap_4 FILLER_36_1540 ();
 sg13g2_fill_1 FILLER_36_1544 ();
 sg13g2_fill_1 FILLER_36_1560 ();
 sg13g2_decap_8 FILLER_36_1565 ();
 sg13g2_decap_8 FILLER_36_1572 ();
 sg13g2_decap_8 FILLER_36_1579 ();
 sg13g2_decap_8 FILLER_36_1586 ();
 sg13g2_decap_4 FILLER_36_1593 ();
 sg13g2_fill_2 FILLER_36_1597 ();
 sg13g2_decap_8 FILLER_36_1615 ();
 sg13g2_decap_8 FILLER_36_1622 ();
 sg13g2_decap_8 FILLER_36_1629 ();
 sg13g2_decap_8 FILLER_36_1636 ();
 sg13g2_decap_8 FILLER_36_1643 ();
 sg13g2_decap_4 FILLER_36_1650 ();
 sg13g2_fill_1 FILLER_36_1654 ();
 sg13g2_decap_8 FILLER_36_1659 ();
 sg13g2_decap_8 FILLER_36_1670 ();
 sg13g2_decap_8 FILLER_36_1677 ();
 sg13g2_decap_8 FILLER_36_1684 ();
 sg13g2_decap_8 FILLER_36_1691 ();
 sg13g2_decap_4 FILLER_36_1698 ();
 sg13g2_fill_2 FILLER_36_1702 ();
 sg13g2_decap_8 FILLER_36_1710 ();
 sg13g2_decap_8 FILLER_36_1717 ();
 sg13g2_decap_8 FILLER_36_1724 ();
 sg13g2_decap_4 FILLER_36_1731 ();
 sg13g2_decap_8 FILLER_36_1745 ();
 sg13g2_decap_8 FILLER_36_1752 ();
 sg13g2_decap_8 FILLER_36_1759 ();
 sg13g2_decap_8 FILLER_36_1766 ();
 sg13g2_decap_8 FILLER_36_1773 ();
 sg13g2_decap_8 FILLER_36_1780 ();
 sg13g2_fill_2 FILLER_36_1787 ();
 sg13g2_decap_8 FILLER_36_1794 ();
 sg13g2_decap_8 FILLER_36_1801 ();
 sg13g2_decap_8 FILLER_36_1808 ();
 sg13g2_decap_4 FILLER_36_1815 ();
 sg13g2_fill_2 FILLER_36_1819 ();
 sg13g2_decap_8 FILLER_36_1826 ();
 sg13g2_decap_8 FILLER_36_1833 ();
 sg13g2_decap_8 FILLER_36_1840 ();
 sg13g2_decap_8 FILLER_36_1847 ();
 sg13g2_decap_8 FILLER_36_1854 ();
 sg13g2_decap_8 FILLER_36_1861 ();
 sg13g2_decap_8 FILLER_36_1868 ();
 sg13g2_decap_8 FILLER_36_1875 ();
 sg13g2_decap_8 FILLER_36_1882 ();
 sg13g2_decap_8 FILLER_36_1889 ();
 sg13g2_decap_8 FILLER_36_1896 ();
 sg13g2_decap_8 FILLER_36_1903 ();
 sg13g2_decap_8 FILLER_36_1910 ();
 sg13g2_decap_8 FILLER_36_1917 ();
 sg13g2_decap_8 FILLER_36_1924 ();
 sg13g2_decap_8 FILLER_36_1931 ();
 sg13g2_decap_8 FILLER_36_1938 ();
 sg13g2_decap_8 FILLER_36_1945 ();
 sg13g2_decap_8 FILLER_36_1952 ();
 sg13g2_decap_8 FILLER_36_1959 ();
 sg13g2_decap_8 FILLER_36_1966 ();
 sg13g2_decap_8 FILLER_36_1973 ();
 sg13g2_decap_8 FILLER_36_1980 ();
 sg13g2_decap_8 FILLER_36_1987 ();
 sg13g2_decap_8 FILLER_36_1994 ();
 sg13g2_decap_8 FILLER_36_2001 ();
 sg13g2_decap_8 FILLER_36_2008 ();
 sg13g2_decap_8 FILLER_36_2015 ();
 sg13g2_decap_8 FILLER_36_2022 ();
 sg13g2_decap_8 FILLER_36_2029 ();
 sg13g2_decap_8 FILLER_36_2036 ();
 sg13g2_decap_8 FILLER_36_2043 ();
 sg13g2_decap_8 FILLER_36_2050 ();
 sg13g2_decap_8 FILLER_36_2057 ();
 sg13g2_decap_8 FILLER_36_2064 ();
 sg13g2_decap_8 FILLER_36_2071 ();
 sg13g2_decap_8 FILLER_36_2078 ();
 sg13g2_decap_8 FILLER_36_2085 ();
 sg13g2_decap_8 FILLER_36_2092 ();
 sg13g2_decap_8 FILLER_36_2099 ();
 sg13g2_decap_8 FILLER_36_2106 ();
 sg13g2_decap_8 FILLER_36_2113 ();
 sg13g2_decap_8 FILLER_36_2120 ();
 sg13g2_decap_8 FILLER_36_2127 ();
 sg13g2_decap_8 FILLER_36_2134 ();
 sg13g2_decap_8 FILLER_36_2141 ();
 sg13g2_decap_8 FILLER_36_2148 ();
 sg13g2_decap_8 FILLER_36_2155 ();
 sg13g2_decap_8 FILLER_36_2162 ();
 sg13g2_decap_8 FILLER_36_2169 ();
 sg13g2_decap_8 FILLER_36_2176 ();
 sg13g2_decap_8 FILLER_36_2183 ();
 sg13g2_decap_8 FILLER_36_2190 ();
 sg13g2_decap_8 FILLER_36_2197 ();
 sg13g2_decap_8 FILLER_36_2204 ();
 sg13g2_decap_8 FILLER_36_2211 ();
 sg13g2_decap_8 FILLER_36_2218 ();
 sg13g2_decap_8 FILLER_36_2225 ();
 sg13g2_decap_8 FILLER_36_2232 ();
 sg13g2_decap_8 FILLER_36_2239 ();
 sg13g2_decap_8 FILLER_36_2246 ();
 sg13g2_decap_8 FILLER_36_2253 ();
 sg13g2_decap_8 FILLER_36_2260 ();
 sg13g2_decap_8 FILLER_36_2267 ();
 sg13g2_decap_8 FILLER_36_2274 ();
 sg13g2_decap_8 FILLER_36_2281 ();
 sg13g2_decap_8 FILLER_36_2288 ();
 sg13g2_decap_8 FILLER_36_2295 ();
 sg13g2_decap_8 FILLER_36_2302 ();
 sg13g2_decap_8 FILLER_36_2309 ();
 sg13g2_decap_8 FILLER_36_2316 ();
 sg13g2_decap_8 FILLER_36_2323 ();
 sg13g2_decap_8 FILLER_36_2330 ();
 sg13g2_decap_8 FILLER_36_2337 ();
 sg13g2_decap_8 FILLER_36_2344 ();
 sg13g2_decap_8 FILLER_36_2351 ();
 sg13g2_decap_8 FILLER_36_2358 ();
 sg13g2_decap_8 FILLER_36_2365 ();
 sg13g2_decap_8 FILLER_36_2372 ();
 sg13g2_decap_8 FILLER_36_2379 ();
 sg13g2_decap_8 FILLER_36_2386 ();
 sg13g2_decap_8 FILLER_36_2393 ();
 sg13g2_decap_8 FILLER_36_2400 ();
 sg13g2_decap_8 FILLER_36_2407 ();
 sg13g2_decap_8 FILLER_36_2414 ();
 sg13g2_decap_8 FILLER_36_2421 ();
 sg13g2_decap_8 FILLER_36_2428 ();
 sg13g2_decap_8 FILLER_36_2435 ();
 sg13g2_decap_8 FILLER_36_2442 ();
 sg13g2_decap_8 FILLER_36_2449 ();
 sg13g2_decap_8 FILLER_36_2456 ();
 sg13g2_decap_8 FILLER_36_2463 ();
 sg13g2_decap_8 FILLER_36_2470 ();
 sg13g2_decap_8 FILLER_36_2477 ();
 sg13g2_decap_8 FILLER_36_2484 ();
 sg13g2_decap_8 FILLER_36_2491 ();
 sg13g2_decap_8 FILLER_36_2498 ();
 sg13g2_decap_8 FILLER_36_2505 ();
 sg13g2_decap_8 FILLER_36_2512 ();
 sg13g2_decap_8 FILLER_36_2519 ();
 sg13g2_decap_8 FILLER_36_2526 ();
 sg13g2_decap_8 FILLER_36_2533 ();
 sg13g2_decap_8 FILLER_36_2540 ();
 sg13g2_decap_8 FILLER_36_2547 ();
 sg13g2_decap_8 FILLER_36_2554 ();
 sg13g2_decap_8 FILLER_36_2561 ();
 sg13g2_decap_8 FILLER_36_2568 ();
 sg13g2_decap_8 FILLER_36_2575 ();
 sg13g2_decap_8 FILLER_36_2582 ();
 sg13g2_decap_8 FILLER_36_2589 ();
 sg13g2_decap_8 FILLER_36_2596 ();
 sg13g2_decap_8 FILLER_36_2603 ();
 sg13g2_decap_8 FILLER_36_2610 ();
 sg13g2_decap_8 FILLER_36_2617 ();
 sg13g2_decap_8 FILLER_36_2624 ();
 sg13g2_decap_8 FILLER_36_2631 ();
 sg13g2_decap_8 FILLER_36_2638 ();
 sg13g2_decap_8 FILLER_36_2645 ();
 sg13g2_decap_8 FILLER_36_2652 ();
 sg13g2_decap_8 FILLER_36_2659 ();
 sg13g2_decap_4 FILLER_36_2666 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_fill_2 FILLER_37_84 ();
 sg13g2_fill_1 FILLER_37_86 ();
 sg13g2_decap_8 FILLER_37_90 ();
 sg13g2_decap_4 FILLER_37_97 ();
 sg13g2_fill_2 FILLER_37_101 ();
 sg13g2_decap_4 FILLER_37_113 ();
 sg13g2_fill_1 FILLER_37_117 ();
 sg13g2_decap_8 FILLER_37_123 ();
 sg13g2_fill_2 FILLER_37_130 ();
 sg13g2_decap_8 FILLER_37_137 ();
 sg13g2_decap_8 FILLER_37_144 ();
 sg13g2_decap_8 FILLER_37_151 ();
 sg13g2_decap_8 FILLER_37_158 ();
 sg13g2_decap_8 FILLER_37_165 ();
 sg13g2_decap_8 FILLER_37_172 ();
 sg13g2_decap_8 FILLER_37_179 ();
 sg13g2_decap_8 FILLER_37_186 ();
 sg13g2_decap_8 FILLER_37_193 ();
 sg13g2_decap_8 FILLER_37_200 ();
 sg13g2_decap_8 FILLER_37_207 ();
 sg13g2_decap_8 FILLER_37_214 ();
 sg13g2_decap_8 FILLER_37_221 ();
 sg13g2_decap_8 FILLER_37_228 ();
 sg13g2_decap_8 FILLER_37_235 ();
 sg13g2_decap_8 FILLER_37_242 ();
 sg13g2_decap_8 FILLER_37_249 ();
 sg13g2_decap_8 FILLER_37_256 ();
 sg13g2_decap_8 FILLER_37_263 ();
 sg13g2_decap_8 FILLER_37_270 ();
 sg13g2_decap_8 FILLER_37_277 ();
 sg13g2_decap_8 FILLER_37_284 ();
 sg13g2_decap_8 FILLER_37_291 ();
 sg13g2_decap_8 FILLER_37_298 ();
 sg13g2_decap_8 FILLER_37_305 ();
 sg13g2_decap_8 FILLER_37_312 ();
 sg13g2_decap_4 FILLER_37_319 ();
 sg13g2_fill_2 FILLER_37_323 ();
 sg13g2_decap_8 FILLER_37_330 ();
 sg13g2_decap_8 FILLER_37_337 ();
 sg13g2_decap_8 FILLER_37_344 ();
 sg13g2_decap_8 FILLER_37_351 ();
 sg13g2_decap_8 FILLER_37_358 ();
 sg13g2_decap_8 FILLER_37_365 ();
 sg13g2_decap_8 FILLER_37_372 ();
 sg13g2_decap_8 FILLER_37_379 ();
 sg13g2_decap_8 FILLER_37_386 ();
 sg13g2_decap_8 FILLER_37_393 ();
 sg13g2_decap_8 FILLER_37_400 ();
 sg13g2_decap_8 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_37_414 ();
 sg13g2_decap_8 FILLER_37_421 ();
 sg13g2_decap_8 FILLER_37_428 ();
 sg13g2_decap_8 FILLER_37_435 ();
 sg13g2_decap_8 FILLER_37_468 ();
 sg13g2_decap_8 FILLER_37_475 ();
 sg13g2_decap_8 FILLER_37_482 ();
 sg13g2_decap_8 FILLER_37_489 ();
 sg13g2_decap_8 FILLER_37_496 ();
 sg13g2_decap_8 FILLER_37_503 ();
 sg13g2_decap_8 FILLER_37_510 ();
 sg13g2_decap_4 FILLER_37_517 ();
 sg13g2_fill_1 FILLER_37_521 ();
 sg13g2_decap_4 FILLER_37_527 ();
 sg13g2_decap_8 FILLER_37_535 ();
 sg13g2_decap_8 FILLER_37_542 ();
 sg13g2_decap_4 FILLER_37_549 ();
 sg13g2_fill_1 FILLER_37_553 ();
 sg13g2_decap_8 FILLER_37_569 ();
 sg13g2_decap_8 FILLER_37_576 ();
 sg13g2_decap_8 FILLER_37_583 ();
 sg13g2_decap_8 FILLER_37_590 ();
 sg13g2_decap_4 FILLER_37_597 ();
 sg13g2_fill_1 FILLER_37_601 ();
 sg13g2_decap_8 FILLER_37_617 ();
 sg13g2_decap_8 FILLER_37_624 ();
 sg13g2_decap_8 FILLER_37_631 ();
 sg13g2_decap_8 FILLER_37_638 ();
 sg13g2_decap_8 FILLER_37_645 ();
 sg13g2_decap_8 FILLER_37_671 ();
 sg13g2_decap_8 FILLER_37_678 ();
 sg13g2_fill_2 FILLER_37_685 ();
 sg13g2_decap_8 FILLER_37_694 ();
 sg13g2_decap_8 FILLER_37_701 ();
 sg13g2_decap_8 FILLER_37_733 ();
 sg13g2_decap_8 FILLER_37_740 ();
 sg13g2_decap_8 FILLER_37_747 ();
 sg13g2_decap_8 FILLER_37_754 ();
 sg13g2_decap_8 FILLER_37_761 ();
 sg13g2_fill_1 FILLER_37_768 ();
 sg13g2_decap_8 FILLER_37_772 ();
 sg13g2_decap_8 FILLER_37_779 ();
 sg13g2_decap_8 FILLER_37_786 ();
 sg13g2_decap_8 FILLER_37_793 ();
 sg13g2_decap_8 FILLER_37_800 ();
 sg13g2_decap_8 FILLER_37_807 ();
 sg13g2_decap_8 FILLER_37_814 ();
 sg13g2_decap_8 FILLER_37_821 ();
 sg13g2_decap_8 FILLER_37_828 ();
 sg13g2_decap_8 FILLER_37_835 ();
 sg13g2_fill_1 FILLER_37_842 ();
 sg13g2_decap_8 FILLER_37_853 ();
 sg13g2_decap_8 FILLER_37_860 ();
 sg13g2_decap_8 FILLER_37_867 ();
 sg13g2_decap_8 FILLER_37_874 ();
 sg13g2_decap_8 FILLER_37_881 ();
 sg13g2_decap_8 FILLER_37_888 ();
 sg13g2_decap_4 FILLER_37_895 ();
 sg13g2_fill_2 FILLER_37_899 ();
 sg13g2_decap_8 FILLER_37_917 ();
 sg13g2_fill_1 FILLER_37_924 ();
 sg13g2_decap_8 FILLER_37_929 ();
 sg13g2_decap_4 FILLER_37_936 ();
 sg13g2_fill_1 FILLER_37_940 ();
 sg13g2_decap_8 FILLER_37_946 ();
 sg13g2_decap_8 FILLER_37_953 ();
 sg13g2_decap_8 FILLER_37_960 ();
 sg13g2_decap_8 FILLER_37_967 ();
 sg13g2_decap_8 FILLER_37_974 ();
 sg13g2_decap_8 FILLER_37_981 ();
 sg13g2_decap_4 FILLER_37_988 ();
 sg13g2_decap_8 FILLER_37_1002 ();
 sg13g2_decap_8 FILLER_37_1009 ();
 sg13g2_decap_8 FILLER_37_1016 ();
 sg13g2_decap_8 FILLER_37_1023 ();
 sg13g2_fill_1 FILLER_37_1030 ();
 sg13g2_decap_8 FILLER_37_1039 ();
 sg13g2_decap_8 FILLER_37_1046 ();
 sg13g2_decap_8 FILLER_37_1053 ();
 sg13g2_decap_4 FILLER_37_1060 ();
 sg13g2_fill_2 FILLER_37_1064 ();
 sg13g2_decap_8 FILLER_37_1071 ();
 sg13g2_decap_8 FILLER_37_1078 ();
 sg13g2_decap_8 FILLER_37_1085 ();
 sg13g2_decap_8 FILLER_37_1092 ();
 sg13g2_decap_8 FILLER_37_1099 ();
 sg13g2_decap_8 FILLER_37_1106 ();
 sg13g2_decap_8 FILLER_37_1113 ();
 sg13g2_decap_8 FILLER_37_1120 ();
 sg13g2_fill_2 FILLER_37_1127 ();
 sg13g2_fill_1 FILLER_37_1129 ();
 sg13g2_decap_8 FILLER_37_1139 ();
 sg13g2_decap_8 FILLER_37_1146 ();
 sg13g2_decap_8 FILLER_37_1153 ();
 sg13g2_decap_8 FILLER_37_1160 ();
 sg13g2_decap_8 FILLER_37_1167 ();
 sg13g2_decap_8 FILLER_37_1174 ();
 sg13g2_decap_8 FILLER_37_1181 ();
 sg13g2_decap_8 FILLER_37_1188 ();
 sg13g2_decap_8 FILLER_37_1195 ();
 sg13g2_decap_8 FILLER_37_1202 ();
 sg13g2_decap_8 FILLER_37_1209 ();
 sg13g2_decap_8 FILLER_37_1216 ();
 sg13g2_decap_8 FILLER_37_1223 ();
 sg13g2_fill_2 FILLER_37_1230 ();
 sg13g2_decap_8 FILLER_37_1236 ();
 sg13g2_decap_8 FILLER_37_1243 ();
 sg13g2_fill_2 FILLER_37_1250 ();
 sg13g2_decap_8 FILLER_37_1262 ();
 sg13g2_decap_8 FILLER_37_1269 ();
 sg13g2_decap_8 FILLER_37_1282 ();
 sg13g2_decap_8 FILLER_37_1289 ();
 sg13g2_decap_8 FILLER_37_1296 ();
 sg13g2_fill_2 FILLER_37_1303 ();
 sg13g2_fill_1 FILLER_37_1305 ();
 sg13g2_decap_8 FILLER_37_1310 ();
 sg13g2_decap_8 FILLER_37_1317 ();
 sg13g2_decap_8 FILLER_37_1324 ();
 sg13g2_decap_8 FILLER_37_1331 ();
 sg13g2_decap_8 FILLER_37_1338 ();
 sg13g2_decap_8 FILLER_37_1345 ();
 sg13g2_decap_8 FILLER_37_1352 ();
 sg13g2_decap_8 FILLER_37_1359 ();
 sg13g2_decap_8 FILLER_37_1366 ();
 sg13g2_decap_8 FILLER_37_1373 ();
 sg13g2_decap_8 FILLER_37_1380 ();
 sg13g2_decap_4 FILLER_37_1387 ();
 sg13g2_fill_1 FILLER_37_1391 ();
 sg13g2_decap_8 FILLER_37_1398 ();
 sg13g2_decap_8 FILLER_37_1405 ();
 sg13g2_decap_8 FILLER_37_1412 ();
 sg13g2_decap_8 FILLER_37_1419 ();
 sg13g2_decap_8 FILLER_37_1426 ();
 sg13g2_decap_4 FILLER_37_1433 ();
 sg13g2_fill_2 FILLER_37_1458 ();
 sg13g2_decap_4 FILLER_37_1469 ();
 sg13g2_decap_8 FILLER_37_1493 ();
 sg13g2_decap_8 FILLER_37_1500 ();
 sg13g2_decap_8 FILLER_37_1507 ();
 sg13g2_decap_8 FILLER_37_1514 ();
 sg13g2_decap_8 FILLER_37_1521 ();
 sg13g2_decap_8 FILLER_37_1528 ();
 sg13g2_decap_8 FILLER_37_1535 ();
 sg13g2_fill_2 FILLER_37_1542 ();
 sg13g2_fill_1 FILLER_37_1544 ();
 sg13g2_decap_4 FILLER_37_1550 ();
 sg13g2_decap_8 FILLER_37_1558 ();
 sg13g2_decap_8 FILLER_37_1565 ();
 sg13g2_decap_4 FILLER_37_1572 ();
 sg13g2_fill_2 FILLER_37_1576 ();
 sg13g2_decap_8 FILLER_37_1583 ();
 sg13g2_decap_8 FILLER_37_1590 ();
 sg13g2_fill_2 FILLER_37_1597 ();
 sg13g2_decap_8 FILLER_37_1604 ();
 sg13g2_fill_2 FILLER_37_1611 ();
 sg13g2_decap_8 FILLER_37_1616 ();
 sg13g2_decap_4 FILLER_37_1623 ();
 sg13g2_decap_8 FILLER_37_1631 ();
 sg13g2_decap_8 FILLER_37_1638 ();
 sg13g2_decap_8 FILLER_37_1645 ();
 sg13g2_decap_8 FILLER_37_1652 ();
 sg13g2_decap_8 FILLER_37_1659 ();
 sg13g2_decap_8 FILLER_37_1666 ();
 sg13g2_decap_8 FILLER_37_1673 ();
 sg13g2_decap_8 FILLER_37_1680 ();
 sg13g2_decap_8 FILLER_37_1687 ();
 sg13g2_decap_8 FILLER_37_1694 ();
 sg13g2_decap_8 FILLER_37_1701 ();
 sg13g2_decap_8 FILLER_37_1708 ();
 sg13g2_decap_8 FILLER_37_1715 ();
 sg13g2_decap_8 FILLER_37_1722 ();
 sg13g2_decap_8 FILLER_37_1729 ();
 sg13g2_fill_1 FILLER_37_1736 ();
 sg13g2_decap_8 FILLER_37_1742 ();
 sg13g2_decap_8 FILLER_37_1749 ();
 sg13g2_decap_8 FILLER_37_1756 ();
 sg13g2_decap_8 FILLER_37_1763 ();
 sg13g2_decap_8 FILLER_37_1770 ();
 sg13g2_decap_8 FILLER_37_1777 ();
 sg13g2_decap_4 FILLER_37_1784 ();
 sg13g2_decap_8 FILLER_37_1793 ();
 sg13g2_decap_8 FILLER_37_1800 ();
 sg13g2_decap_8 FILLER_37_1807 ();
 sg13g2_decap_8 FILLER_37_1814 ();
 sg13g2_decap_8 FILLER_37_1821 ();
 sg13g2_decap_8 FILLER_37_1828 ();
 sg13g2_decap_8 FILLER_37_1835 ();
 sg13g2_decap_8 FILLER_37_1842 ();
 sg13g2_decap_8 FILLER_37_1849 ();
 sg13g2_decap_8 FILLER_37_1856 ();
 sg13g2_decap_8 FILLER_37_1863 ();
 sg13g2_decap_8 FILLER_37_1870 ();
 sg13g2_decap_8 FILLER_37_1877 ();
 sg13g2_decap_8 FILLER_37_1884 ();
 sg13g2_decap_8 FILLER_37_1891 ();
 sg13g2_decap_8 FILLER_37_1898 ();
 sg13g2_decap_8 FILLER_37_1905 ();
 sg13g2_decap_8 FILLER_37_1912 ();
 sg13g2_decap_8 FILLER_37_1919 ();
 sg13g2_decap_8 FILLER_37_1926 ();
 sg13g2_decap_8 FILLER_37_1933 ();
 sg13g2_decap_8 FILLER_37_1940 ();
 sg13g2_decap_8 FILLER_37_1947 ();
 sg13g2_decap_8 FILLER_37_1954 ();
 sg13g2_decap_8 FILLER_37_1961 ();
 sg13g2_decap_8 FILLER_37_1968 ();
 sg13g2_decap_8 FILLER_37_1975 ();
 sg13g2_decap_8 FILLER_37_1982 ();
 sg13g2_decap_8 FILLER_37_1989 ();
 sg13g2_decap_8 FILLER_37_1996 ();
 sg13g2_decap_8 FILLER_37_2003 ();
 sg13g2_decap_8 FILLER_37_2010 ();
 sg13g2_decap_8 FILLER_37_2017 ();
 sg13g2_decap_8 FILLER_37_2024 ();
 sg13g2_decap_8 FILLER_37_2031 ();
 sg13g2_decap_8 FILLER_37_2038 ();
 sg13g2_decap_8 FILLER_37_2045 ();
 sg13g2_decap_8 FILLER_37_2052 ();
 sg13g2_decap_8 FILLER_37_2059 ();
 sg13g2_decap_8 FILLER_37_2066 ();
 sg13g2_decap_8 FILLER_37_2073 ();
 sg13g2_decap_8 FILLER_37_2080 ();
 sg13g2_decap_8 FILLER_37_2087 ();
 sg13g2_decap_8 FILLER_37_2094 ();
 sg13g2_decap_8 FILLER_37_2101 ();
 sg13g2_decap_8 FILLER_37_2108 ();
 sg13g2_decap_8 FILLER_37_2115 ();
 sg13g2_decap_8 FILLER_37_2122 ();
 sg13g2_decap_8 FILLER_37_2129 ();
 sg13g2_decap_8 FILLER_37_2136 ();
 sg13g2_decap_8 FILLER_37_2143 ();
 sg13g2_decap_8 FILLER_37_2150 ();
 sg13g2_decap_8 FILLER_37_2157 ();
 sg13g2_decap_8 FILLER_37_2164 ();
 sg13g2_decap_8 FILLER_37_2171 ();
 sg13g2_decap_8 FILLER_37_2178 ();
 sg13g2_decap_8 FILLER_37_2185 ();
 sg13g2_decap_8 FILLER_37_2192 ();
 sg13g2_decap_8 FILLER_37_2199 ();
 sg13g2_decap_8 FILLER_37_2206 ();
 sg13g2_decap_8 FILLER_37_2213 ();
 sg13g2_decap_8 FILLER_37_2220 ();
 sg13g2_decap_8 FILLER_37_2227 ();
 sg13g2_decap_8 FILLER_37_2234 ();
 sg13g2_decap_8 FILLER_37_2241 ();
 sg13g2_decap_8 FILLER_37_2248 ();
 sg13g2_decap_8 FILLER_37_2255 ();
 sg13g2_decap_8 FILLER_37_2262 ();
 sg13g2_decap_8 FILLER_37_2269 ();
 sg13g2_decap_8 FILLER_37_2276 ();
 sg13g2_decap_8 FILLER_37_2283 ();
 sg13g2_decap_8 FILLER_37_2290 ();
 sg13g2_decap_8 FILLER_37_2297 ();
 sg13g2_decap_8 FILLER_37_2304 ();
 sg13g2_decap_8 FILLER_37_2311 ();
 sg13g2_decap_8 FILLER_37_2318 ();
 sg13g2_decap_8 FILLER_37_2325 ();
 sg13g2_decap_8 FILLER_37_2332 ();
 sg13g2_decap_8 FILLER_37_2339 ();
 sg13g2_decap_8 FILLER_37_2346 ();
 sg13g2_decap_8 FILLER_37_2353 ();
 sg13g2_decap_8 FILLER_37_2360 ();
 sg13g2_decap_8 FILLER_37_2367 ();
 sg13g2_decap_8 FILLER_37_2374 ();
 sg13g2_decap_8 FILLER_37_2381 ();
 sg13g2_decap_8 FILLER_37_2388 ();
 sg13g2_decap_8 FILLER_37_2395 ();
 sg13g2_decap_8 FILLER_37_2402 ();
 sg13g2_decap_8 FILLER_37_2409 ();
 sg13g2_decap_8 FILLER_37_2416 ();
 sg13g2_decap_8 FILLER_37_2423 ();
 sg13g2_decap_8 FILLER_37_2430 ();
 sg13g2_decap_8 FILLER_37_2437 ();
 sg13g2_decap_8 FILLER_37_2444 ();
 sg13g2_decap_8 FILLER_37_2451 ();
 sg13g2_decap_8 FILLER_37_2458 ();
 sg13g2_decap_8 FILLER_37_2465 ();
 sg13g2_decap_8 FILLER_37_2472 ();
 sg13g2_decap_8 FILLER_37_2479 ();
 sg13g2_decap_8 FILLER_37_2486 ();
 sg13g2_decap_8 FILLER_37_2493 ();
 sg13g2_decap_8 FILLER_37_2500 ();
 sg13g2_decap_8 FILLER_37_2507 ();
 sg13g2_decap_8 FILLER_37_2514 ();
 sg13g2_decap_8 FILLER_37_2521 ();
 sg13g2_decap_8 FILLER_37_2528 ();
 sg13g2_decap_8 FILLER_37_2535 ();
 sg13g2_decap_8 FILLER_37_2542 ();
 sg13g2_decap_8 FILLER_37_2549 ();
 sg13g2_decap_8 FILLER_37_2556 ();
 sg13g2_decap_8 FILLER_37_2563 ();
 sg13g2_decap_8 FILLER_37_2570 ();
 sg13g2_decap_8 FILLER_37_2577 ();
 sg13g2_decap_8 FILLER_37_2584 ();
 sg13g2_decap_8 FILLER_37_2591 ();
 sg13g2_decap_8 FILLER_37_2598 ();
 sg13g2_decap_8 FILLER_37_2605 ();
 sg13g2_decap_8 FILLER_37_2612 ();
 sg13g2_decap_8 FILLER_37_2619 ();
 sg13g2_decap_8 FILLER_37_2626 ();
 sg13g2_decap_8 FILLER_37_2633 ();
 sg13g2_decap_8 FILLER_37_2640 ();
 sg13g2_decap_8 FILLER_37_2647 ();
 sg13g2_decap_8 FILLER_37_2654 ();
 sg13g2_decap_8 FILLER_37_2661 ();
 sg13g2_fill_2 FILLER_37_2668 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_4 FILLER_38_119 ();
 sg13g2_decap_8 FILLER_38_128 ();
 sg13g2_decap_8 FILLER_38_135 ();
 sg13g2_decap_8 FILLER_38_142 ();
 sg13g2_decap_8 FILLER_38_149 ();
 sg13g2_decap_8 FILLER_38_156 ();
 sg13g2_decap_8 FILLER_38_163 ();
 sg13g2_decap_8 FILLER_38_170 ();
 sg13g2_decap_8 FILLER_38_177 ();
 sg13g2_decap_8 FILLER_38_184 ();
 sg13g2_decap_8 FILLER_38_191 ();
 sg13g2_decap_8 FILLER_38_198 ();
 sg13g2_decap_8 FILLER_38_205 ();
 sg13g2_decap_8 FILLER_38_212 ();
 sg13g2_decap_8 FILLER_38_219 ();
 sg13g2_decap_8 FILLER_38_226 ();
 sg13g2_decap_8 FILLER_38_233 ();
 sg13g2_decap_8 FILLER_38_240 ();
 sg13g2_decap_8 FILLER_38_247 ();
 sg13g2_decap_8 FILLER_38_254 ();
 sg13g2_decap_8 FILLER_38_261 ();
 sg13g2_decap_8 FILLER_38_268 ();
 sg13g2_decap_8 FILLER_38_275 ();
 sg13g2_decap_8 FILLER_38_282 ();
 sg13g2_decap_8 FILLER_38_289 ();
 sg13g2_decap_8 FILLER_38_296 ();
 sg13g2_decap_8 FILLER_38_303 ();
 sg13g2_decap_8 FILLER_38_310 ();
 sg13g2_decap_8 FILLER_38_317 ();
 sg13g2_decap_8 FILLER_38_324 ();
 sg13g2_decap_8 FILLER_38_331 ();
 sg13g2_decap_8 FILLER_38_338 ();
 sg13g2_decap_8 FILLER_38_345 ();
 sg13g2_decap_8 FILLER_38_352 ();
 sg13g2_decap_8 FILLER_38_359 ();
 sg13g2_decap_8 FILLER_38_366 ();
 sg13g2_decap_8 FILLER_38_373 ();
 sg13g2_decap_8 FILLER_38_380 ();
 sg13g2_decap_8 FILLER_38_387 ();
 sg13g2_decap_8 FILLER_38_394 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_decap_8 FILLER_38_408 ();
 sg13g2_decap_8 FILLER_38_415 ();
 sg13g2_decap_8 FILLER_38_422 ();
 sg13g2_decap_8 FILLER_38_429 ();
 sg13g2_fill_1 FILLER_38_451 ();
 sg13g2_decap_8 FILLER_38_461 ();
 sg13g2_decap_8 FILLER_38_468 ();
 sg13g2_decap_8 FILLER_38_475 ();
 sg13g2_decap_8 FILLER_38_482 ();
 sg13g2_decap_8 FILLER_38_489 ();
 sg13g2_decap_8 FILLER_38_496 ();
 sg13g2_decap_8 FILLER_38_503 ();
 sg13g2_decap_8 FILLER_38_510 ();
 sg13g2_decap_8 FILLER_38_517 ();
 sg13g2_decap_8 FILLER_38_524 ();
 sg13g2_decap_8 FILLER_38_531 ();
 sg13g2_decap_8 FILLER_38_538 ();
 sg13g2_decap_8 FILLER_38_564 ();
 sg13g2_decap_8 FILLER_38_571 ();
 sg13g2_decap_8 FILLER_38_578 ();
 sg13g2_decap_8 FILLER_38_585 ();
 sg13g2_fill_1 FILLER_38_597 ();
 sg13g2_fill_2 FILLER_38_603 ();
 sg13g2_decap_8 FILLER_38_610 ();
 sg13g2_decap_8 FILLER_38_617 ();
 sg13g2_decap_8 FILLER_38_624 ();
 sg13g2_decap_8 FILLER_38_631 ();
 sg13g2_decap_8 FILLER_38_638 ();
 sg13g2_decap_8 FILLER_38_645 ();
 sg13g2_decap_8 FILLER_38_652 ();
 sg13g2_decap_4 FILLER_38_659 ();
 sg13g2_decap_4 FILLER_38_668 ();
 sg13g2_fill_2 FILLER_38_672 ();
 sg13g2_fill_1 FILLER_38_683 ();
 sg13g2_decap_8 FILLER_38_702 ();
 sg13g2_fill_2 FILLER_38_709 ();
 sg13g2_decap_8 FILLER_38_726 ();
 sg13g2_decap_8 FILLER_38_733 ();
 sg13g2_decap_8 FILLER_38_740 ();
 sg13g2_decap_8 FILLER_38_747 ();
 sg13g2_decap_8 FILLER_38_754 ();
 sg13g2_decap_4 FILLER_38_761 ();
 sg13g2_decap_8 FILLER_38_773 ();
 sg13g2_decap_8 FILLER_38_780 ();
 sg13g2_decap_8 FILLER_38_787 ();
 sg13g2_decap_8 FILLER_38_794 ();
 sg13g2_decap_8 FILLER_38_801 ();
 sg13g2_decap_8 FILLER_38_808 ();
 sg13g2_decap_8 FILLER_38_815 ();
 sg13g2_decap_8 FILLER_38_822 ();
 sg13g2_decap_8 FILLER_38_829 ();
 sg13g2_decap_8 FILLER_38_836 ();
 sg13g2_decap_8 FILLER_38_843 ();
 sg13g2_decap_8 FILLER_38_850 ();
 sg13g2_decap_8 FILLER_38_857 ();
 sg13g2_fill_1 FILLER_38_864 ();
 sg13g2_decap_8 FILLER_38_880 ();
 sg13g2_decap_8 FILLER_38_887 ();
 sg13g2_decap_8 FILLER_38_894 ();
 sg13g2_decap_8 FILLER_38_901 ();
 sg13g2_decap_8 FILLER_38_908 ();
 sg13g2_decap_8 FILLER_38_915 ();
 sg13g2_fill_2 FILLER_38_922 ();
 sg13g2_fill_1 FILLER_38_924 ();
 sg13g2_decap_8 FILLER_38_928 ();
 sg13g2_decap_8 FILLER_38_935 ();
 sg13g2_decap_8 FILLER_38_942 ();
 sg13g2_decap_8 FILLER_38_949 ();
 sg13g2_decap_8 FILLER_38_956 ();
 sg13g2_decap_8 FILLER_38_963 ();
 sg13g2_decap_8 FILLER_38_970 ();
 sg13g2_decap_8 FILLER_38_977 ();
 sg13g2_decap_8 FILLER_38_984 ();
 sg13g2_decap_8 FILLER_38_991 ();
 sg13g2_fill_2 FILLER_38_998 ();
 sg13g2_decap_8 FILLER_38_1003 ();
 sg13g2_decap_8 FILLER_38_1010 ();
 sg13g2_decap_8 FILLER_38_1017 ();
 sg13g2_decap_4 FILLER_38_1024 ();
 sg13g2_decap_8 FILLER_38_1033 ();
 sg13g2_decap_8 FILLER_38_1040 ();
 sg13g2_decap_8 FILLER_38_1047 ();
 sg13g2_decap_8 FILLER_38_1054 ();
 sg13g2_decap_8 FILLER_38_1061 ();
 sg13g2_decap_8 FILLER_38_1068 ();
 sg13g2_decap_8 FILLER_38_1075 ();
 sg13g2_decap_8 FILLER_38_1082 ();
 sg13g2_decap_8 FILLER_38_1089 ();
 sg13g2_decap_8 FILLER_38_1096 ();
 sg13g2_decap_8 FILLER_38_1103 ();
 sg13g2_decap_8 FILLER_38_1110 ();
 sg13g2_decap_8 FILLER_38_1117 ();
 sg13g2_fill_1 FILLER_38_1124 ();
 sg13g2_decap_8 FILLER_38_1130 ();
 sg13g2_decap_8 FILLER_38_1137 ();
 sg13g2_decap_8 FILLER_38_1144 ();
 sg13g2_decap_8 FILLER_38_1151 ();
 sg13g2_decap_8 FILLER_38_1158 ();
 sg13g2_fill_1 FILLER_38_1165 ();
 sg13g2_decap_8 FILLER_38_1173 ();
 sg13g2_decap_8 FILLER_38_1180 ();
 sg13g2_decap_8 FILLER_38_1199 ();
 sg13g2_decap_8 FILLER_38_1206 ();
 sg13g2_decap_8 FILLER_38_1213 ();
 sg13g2_decap_8 FILLER_38_1220 ();
 sg13g2_decap_8 FILLER_38_1227 ();
 sg13g2_fill_2 FILLER_38_1234 ();
 sg13g2_fill_1 FILLER_38_1236 ();
 sg13g2_decap_8 FILLER_38_1240 ();
 sg13g2_decap_8 FILLER_38_1247 ();
 sg13g2_decap_8 FILLER_38_1254 ();
 sg13g2_decap_8 FILLER_38_1261 ();
 sg13g2_decap_4 FILLER_38_1268 ();
 sg13g2_fill_1 FILLER_38_1272 ();
 sg13g2_fill_1 FILLER_38_1277 ();
 sg13g2_decap_8 FILLER_38_1282 ();
 sg13g2_decap_8 FILLER_38_1289 ();
 sg13g2_decap_8 FILLER_38_1296 ();
 sg13g2_decap_8 FILLER_38_1303 ();
 sg13g2_decap_8 FILLER_38_1310 ();
 sg13g2_decap_8 FILLER_38_1317 ();
 sg13g2_decap_8 FILLER_38_1324 ();
 sg13g2_decap_4 FILLER_38_1331 ();
 sg13g2_decap_8 FILLER_38_1339 ();
 sg13g2_decap_8 FILLER_38_1346 ();
 sg13g2_decap_8 FILLER_38_1353 ();
 sg13g2_fill_2 FILLER_38_1360 ();
 sg13g2_fill_1 FILLER_38_1362 ();
 sg13g2_decap_8 FILLER_38_1372 ();
 sg13g2_decap_8 FILLER_38_1379 ();
 sg13g2_decap_8 FILLER_38_1386 ();
 sg13g2_fill_2 FILLER_38_1393 ();
 sg13g2_fill_1 FILLER_38_1395 ();
 sg13g2_decap_8 FILLER_38_1400 ();
 sg13g2_decap_8 FILLER_38_1407 ();
 sg13g2_decap_8 FILLER_38_1414 ();
 sg13g2_decap_8 FILLER_38_1421 ();
 sg13g2_decap_8 FILLER_38_1428 ();
 sg13g2_fill_2 FILLER_38_1435 ();
 sg13g2_decap_8 FILLER_38_1441 ();
 sg13g2_fill_2 FILLER_38_1470 ();
 sg13g2_fill_1 FILLER_38_1472 ();
 sg13g2_decap_8 FILLER_38_1477 ();
 sg13g2_decap_8 FILLER_38_1484 ();
 sg13g2_decap_8 FILLER_38_1491 ();
 sg13g2_fill_2 FILLER_38_1498 ();
 sg13g2_fill_1 FILLER_38_1500 ();
 sg13g2_decap_8 FILLER_38_1516 ();
 sg13g2_decap_8 FILLER_38_1523 ();
 sg13g2_decap_8 FILLER_38_1530 ();
 sg13g2_decap_8 FILLER_38_1537 ();
 sg13g2_fill_1 FILLER_38_1544 ();
 sg13g2_decap_8 FILLER_38_1556 ();
 sg13g2_decap_8 FILLER_38_1563 ();
 sg13g2_decap_8 FILLER_38_1570 ();
 sg13g2_decap_8 FILLER_38_1577 ();
 sg13g2_decap_8 FILLER_38_1584 ();
 sg13g2_decap_8 FILLER_38_1591 ();
 sg13g2_decap_8 FILLER_38_1598 ();
 sg13g2_decap_8 FILLER_38_1605 ();
 sg13g2_fill_2 FILLER_38_1612 ();
 sg13g2_decap_8 FILLER_38_1620 ();
 sg13g2_decap_8 FILLER_38_1627 ();
 sg13g2_decap_8 FILLER_38_1634 ();
 sg13g2_decap_8 FILLER_38_1641 ();
 sg13g2_decap_8 FILLER_38_1648 ();
 sg13g2_decap_8 FILLER_38_1655 ();
 sg13g2_fill_2 FILLER_38_1662 ();
 sg13g2_fill_1 FILLER_38_1664 ();
 sg13g2_decap_8 FILLER_38_1669 ();
 sg13g2_decap_8 FILLER_38_1676 ();
 sg13g2_decap_8 FILLER_38_1683 ();
 sg13g2_decap_8 FILLER_38_1690 ();
 sg13g2_decap_8 FILLER_38_1697 ();
 sg13g2_decap_8 FILLER_38_1704 ();
 sg13g2_decap_8 FILLER_38_1711 ();
 sg13g2_decap_8 FILLER_38_1718 ();
 sg13g2_decap_8 FILLER_38_1725 ();
 sg13g2_decap_8 FILLER_38_1732 ();
 sg13g2_decap_8 FILLER_38_1739 ();
 sg13g2_decap_8 FILLER_38_1746 ();
 sg13g2_decap_8 FILLER_38_1753 ();
 sg13g2_decap_8 FILLER_38_1760 ();
 sg13g2_decap_4 FILLER_38_1767 ();
 sg13g2_fill_2 FILLER_38_1771 ();
 sg13g2_decap_8 FILLER_38_1782 ();
 sg13g2_decap_8 FILLER_38_1789 ();
 sg13g2_decap_8 FILLER_38_1796 ();
 sg13g2_decap_8 FILLER_38_1803 ();
 sg13g2_decap_8 FILLER_38_1810 ();
 sg13g2_decap_8 FILLER_38_1817 ();
 sg13g2_decap_8 FILLER_38_1824 ();
 sg13g2_decap_8 FILLER_38_1831 ();
 sg13g2_decap_8 FILLER_38_1838 ();
 sg13g2_decap_8 FILLER_38_1845 ();
 sg13g2_decap_8 FILLER_38_1852 ();
 sg13g2_decap_8 FILLER_38_1859 ();
 sg13g2_decap_8 FILLER_38_1866 ();
 sg13g2_decap_8 FILLER_38_1873 ();
 sg13g2_decap_8 FILLER_38_1880 ();
 sg13g2_decap_8 FILLER_38_1887 ();
 sg13g2_decap_8 FILLER_38_1894 ();
 sg13g2_decap_8 FILLER_38_1901 ();
 sg13g2_decap_8 FILLER_38_1908 ();
 sg13g2_decap_8 FILLER_38_1915 ();
 sg13g2_decap_8 FILLER_38_1922 ();
 sg13g2_decap_8 FILLER_38_1929 ();
 sg13g2_decap_8 FILLER_38_1936 ();
 sg13g2_decap_8 FILLER_38_1943 ();
 sg13g2_decap_8 FILLER_38_1950 ();
 sg13g2_decap_8 FILLER_38_1957 ();
 sg13g2_decap_8 FILLER_38_1964 ();
 sg13g2_decap_8 FILLER_38_1971 ();
 sg13g2_decap_8 FILLER_38_1978 ();
 sg13g2_decap_8 FILLER_38_1985 ();
 sg13g2_decap_8 FILLER_38_1992 ();
 sg13g2_decap_8 FILLER_38_1999 ();
 sg13g2_decap_8 FILLER_38_2006 ();
 sg13g2_decap_8 FILLER_38_2013 ();
 sg13g2_decap_8 FILLER_38_2020 ();
 sg13g2_decap_8 FILLER_38_2027 ();
 sg13g2_decap_8 FILLER_38_2034 ();
 sg13g2_decap_8 FILLER_38_2041 ();
 sg13g2_decap_8 FILLER_38_2048 ();
 sg13g2_decap_8 FILLER_38_2055 ();
 sg13g2_decap_8 FILLER_38_2062 ();
 sg13g2_decap_8 FILLER_38_2069 ();
 sg13g2_decap_8 FILLER_38_2076 ();
 sg13g2_decap_8 FILLER_38_2083 ();
 sg13g2_decap_8 FILLER_38_2090 ();
 sg13g2_decap_8 FILLER_38_2097 ();
 sg13g2_decap_8 FILLER_38_2104 ();
 sg13g2_decap_8 FILLER_38_2111 ();
 sg13g2_decap_8 FILLER_38_2118 ();
 sg13g2_decap_8 FILLER_38_2125 ();
 sg13g2_decap_8 FILLER_38_2132 ();
 sg13g2_decap_8 FILLER_38_2139 ();
 sg13g2_decap_8 FILLER_38_2146 ();
 sg13g2_decap_8 FILLER_38_2153 ();
 sg13g2_decap_8 FILLER_38_2160 ();
 sg13g2_decap_8 FILLER_38_2167 ();
 sg13g2_decap_8 FILLER_38_2174 ();
 sg13g2_decap_8 FILLER_38_2181 ();
 sg13g2_decap_8 FILLER_38_2188 ();
 sg13g2_decap_8 FILLER_38_2195 ();
 sg13g2_decap_8 FILLER_38_2202 ();
 sg13g2_decap_8 FILLER_38_2209 ();
 sg13g2_decap_8 FILLER_38_2216 ();
 sg13g2_decap_8 FILLER_38_2223 ();
 sg13g2_decap_8 FILLER_38_2230 ();
 sg13g2_decap_8 FILLER_38_2237 ();
 sg13g2_decap_8 FILLER_38_2244 ();
 sg13g2_decap_8 FILLER_38_2251 ();
 sg13g2_decap_8 FILLER_38_2258 ();
 sg13g2_decap_8 FILLER_38_2265 ();
 sg13g2_decap_8 FILLER_38_2272 ();
 sg13g2_decap_8 FILLER_38_2279 ();
 sg13g2_decap_8 FILLER_38_2286 ();
 sg13g2_decap_8 FILLER_38_2293 ();
 sg13g2_decap_8 FILLER_38_2300 ();
 sg13g2_decap_8 FILLER_38_2307 ();
 sg13g2_decap_8 FILLER_38_2314 ();
 sg13g2_decap_8 FILLER_38_2321 ();
 sg13g2_decap_8 FILLER_38_2328 ();
 sg13g2_decap_8 FILLER_38_2335 ();
 sg13g2_decap_8 FILLER_38_2342 ();
 sg13g2_decap_8 FILLER_38_2349 ();
 sg13g2_decap_8 FILLER_38_2356 ();
 sg13g2_decap_8 FILLER_38_2363 ();
 sg13g2_decap_8 FILLER_38_2370 ();
 sg13g2_decap_8 FILLER_38_2377 ();
 sg13g2_decap_8 FILLER_38_2384 ();
 sg13g2_decap_8 FILLER_38_2391 ();
 sg13g2_decap_8 FILLER_38_2398 ();
 sg13g2_decap_8 FILLER_38_2405 ();
 sg13g2_decap_8 FILLER_38_2412 ();
 sg13g2_decap_8 FILLER_38_2419 ();
 sg13g2_decap_8 FILLER_38_2426 ();
 sg13g2_decap_8 FILLER_38_2433 ();
 sg13g2_decap_8 FILLER_38_2440 ();
 sg13g2_decap_8 FILLER_38_2447 ();
 sg13g2_decap_8 FILLER_38_2454 ();
 sg13g2_decap_8 FILLER_38_2461 ();
 sg13g2_decap_8 FILLER_38_2468 ();
 sg13g2_decap_8 FILLER_38_2475 ();
 sg13g2_decap_8 FILLER_38_2482 ();
 sg13g2_decap_8 FILLER_38_2489 ();
 sg13g2_decap_8 FILLER_38_2496 ();
 sg13g2_decap_8 FILLER_38_2503 ();
 sg13g2_decap_8 FILLER_38_2510 ();
 sg13g2_decap_8 FILLER_38_2517 ();
 sg13g2_decap_8 FILLER_38_2524 ();
 sg13g2_decap_8 FILLER_38_2531 ();
 sg13g2_decap_8 FILLER_38_2538 ();
 sg13g2_decap_8 FILLER_38_2545 ();
 sg13g2_decap_8 FILLER_38_2552 ();
 sg13g2_decap_8 FILLER_38_2559 ();
 sg13g2_decap_8 FILLER_38_2566 ();
 sg13g2_decap_8 FILLER_38_2573 ();
 sg13g2_decap_8 FILLER_38_2580 ();
 sg13g2_decap_8 FILLER_38_2587 ();
 sg13g2_decap_8 FILLER_38_2594 ();
 sg13g2_decap_8 FILLER_38_2601 ();
 sg13g2_decap_8 FILLER_38_2608 ();
 sg13g2_decap_8 FILLER_38_2615 ();
 sg13g2_decap_8 FILLER_38_2622 ();
 sg13g2_decap_8 FILLER_38_2629 ();
 sg13g2_decap_8 FILLER_38_2636 ();
 sg13g2_decap_8 FILLER_38_2643 ();
 sg13g2_decap_8 FILLER_38_2650 ();
 sg13g2_decap_8 FILLER_38_2657 ();
 sg13g2_decap_4 FILLER_38_2664 ();
 sg13g2_fill_2 FILLER_38_2668 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_fill_2 FILLER_39_70 ();
 sg13g2_fill_1 FILLER_39_72 ();
 sg13g2_fill_2 FILLER_39_83 ();
 sg13g2_decap_8 FILLER_39_88 ();
 sg13g2_decap_8 FILLER_39_95 ();
 sg13g2_decap_4 FILLER_39_102 ();
 sg13g2_fill_2 FILLER_39_106 ();
 sg13g2_decap_8 FILLER_39_113 ();
 sg13g2_decap_8 FILLER_39_120 ();
 sg13g2_decap_8 FILLER_39_127 ();
 sg13g2_decap_8 FILLER_39_134 ();
 sg13g2_decap_8 FILLER_39_141 ();
 sg13g2_decap_8 FILLER_39_148 ();
 sg13g2_decap_8 FILLER_39_155 ();
 sg13g2_decap_8 FILLER_39_162 ();
 sg13g2_decap_8 FILLER_39_169 ();
 sg13g2_decap_4 FILLER_39_176 ();
 sg13g2_fill_1 FILLER_39_180 ();
 sg13g2_fill_1 FILLER_39_184 ();
 sg13g2_decap_8 FILLER_39_190 ();
 sg13g2_decap_8 FILLER_39_197 ();
 sg13g2_decap_8 FILLER_39_204 ();
 sg13g2_decap_8 FILLER_39_211 ();
 sg13g2_decap_8 FILLER_39_218 ();
 sg13g2_decap_8 FILLER_39_225 ();
 sg13g2_fill_2 FILLER_39_232 ();
 sg13g2_fill_1 FILLER_39_234 ();
 sg13g2_decap_8 FILLER_39_261 ();
 sg13g2_decap_8 FILLER_39_268 ();
 sg13g2_decap_8 FILLER_39_275 ();
 sg13g2_decap_8 FILLER_39_282 ();
 sg13g2_decap_8 FILLER_39_289 ();
 sg13g2_decap_8 FILLER_39_296 ();
 sg13g2_decap_8 FILLER_39_303 ();
 sg13g2_decap_8 FILLER_39_310 ();
 sg13g2_decap_8 FILLER_39_317 ();
 sg13g2_decap_8 FILLER_39_324 ();
 sg13g2_decap_8 FILLER_39_331 ();
 sg13g2_decap_8 FILLER_39_338 ();
 sg13g2_decap_8 FILLER_39_345 ();
 sg13g2_decap_8 FILLER_39_352 ();
 sg13g2_decap_4 FILLER_39_359 ();
 sg13g2_fill_1 FILLER_39_363 ();
 sg13g2_decap_8 FILLER_39_372 ();
 sg13g2_decap_8 FILLER_39_379 ();
 sg13g2_decap_8 FILLER_39_386 ();
 sg13g2_decap_8 FILLER_39_393 ();
 sg13g2_decap_8 FILLER_39_400 ();
 sg13g2_decap_8 FILLER_39_407 ();
 sg13g2_decap_8 FILLER_39_414 ();
 sg13g2_decap_8 FILLER_39_421 ();
 sg13g2_decap_8 FILLER_39_428 ();
 sg13g2_decap_8 FILLER_39_435 ();
 sg13g2_decap_8 FILLER_39_446 ();
 sg13g2_decap_8 FILLER_39_453 ();
 sg13g2_decap_8 FILLER_39_460 ();
 sg13g2_decap_8 FILLER_39_467 ();
 sg13g2_decap_8 FILLER_39_474 ();
 sg13g2_decap_8 FILLER_39_481 ();
 sg13g2_decap_8 FILLER_39_488 ();
 sg13g2_decap_8 FILLER_39_495 ();
 sg13g2_decap_8 FILLER_39_502 ();
 sg13g2_decap_8 FILLER_39_509 ();
 sg13g2_decap_8 FILLER_39_516 ();
 sg13g2_decap_8 FILLER_39_523 ();
 sg13g2_decap_8 FILLER_39_530 ();
 sg13g2_decap_8 FILLER_39_537 ();
 sg13g2_decap_8 FILLER_39_544 ();
 sg13g2_decap_8 FILLER_39_551 ();
 sg13g2_decap_8 FILLER_39_558 ();
 sg13g2_decap_8 FILLER_39_565 ();
 sg13g2_fill_1 FILLER_39_572 ();
 sg13g2_decap_8 FILLER_39_588 ();
 sg13g2_decap_8 FILLER_39_595 ();
 sg13g2_decap_8 FILLER_39_602 ();
 sg13g2_decap_8 FILLER_39_609 ();
 sg13g2_decap_8 FILLER_39_616 ();
 sg13g2_decap_8 FILLER_39_623 ();
 sg13g2_decap_8 FILLER_39_630 ();
 sg13g2_decap_4 FILLER_39_637 ();
 sg13g2_fill_1 FILLER_39_641 ();
 sg13g2_decap_8 FILLER_39_657 ();
 sg13g2_decap_8 FILLER_39_664 ();
 sg13g2_fill_2 FILLER_39_671 ();
 sg13g2_fill_1 FILLER_39_673 ();
 sg13g2_decap_8 FILLER_39_692 ();
 sg13g2_decap_8 FILLER_39_699 ();
 sg13g2_decap_8 FILLER_39_706 ();
 sg13g2_decap_8 FILLER_39_713 ();
 sg13g2_decap_8 FILLER_39_720 ();
 sg13g2_decap_8 FILLER_39_727 ();
 sg13g2_decap_8 FILLER_39_734 ();
 sg13g2_decap_8 FILLER_39_741 ();
 sg13g2_fill_1 FILLER_39_748 ();
 sg13g2_decap_8 FILLER_39_776 ();
 sg13g2_decap_8 FILLER_39_783 ();
 sg13g2_decap_8 FILLER_39_790 ();
 sg13g2_fill_1 FILLER_39_797 ();
 sg13g2_decap_8 FILLER_39_813 ();
 sg13g2_decap_8 FILLER_39_820 ();
 sg13g2_fill_2 FILLER_39_827 ();
 sg13g2_decap_8 FILLER_39_832 ();
 sg13g2_fill_1 FILLER_39_839 ();
 sg13g2_decap_8 FILLER_39_844 ();
 sg13g2_decap_8 FILLER_39_851 ();
 sg13g2_decap_8 FILLER_39_858 ();
 sg13g2_fill_2 FILLER_39_865 ();
 sg13g2_fill_1 FILLER_39_867 ();
 sg13g2_decap_8 FILLER_39_873 ();
 sg13g2_decap_8 FILLER_39_880 ();
 sg13g2_decap_8 FILLER_39_887 ();
 sg13g2_fill_2 FILLER_39_894 ();
 sg13g2_decap_8 FILLER_39_900 ();
 sg13g2_decap_8 FILLER_39_907 ();
 sg13g2_decap_8 FILLER_39_914 ();
 sg13g2_decap_8 FILLER_39_921 ();
 sg13g2_decap_4 FILLER_39_932 ();
 sg13g2_decap_8 FILLER_39_944 ();
 sg13g2_decap_8 FILLER_39_951 ();
 sg13g2_decap_8 FILLER_39_958 ();
 sg13g2_decap_8 FILLER_39_965 ();
 sg13g2_decap_8 FILLER_39_972 ();
 sg13g2_decap_8 FILLER_39_979 ();
 sg13g2_decap_8 FILLER_39_986 ();
 sg13g2_decap_4 FILLER_39_993 ();
 sg13g2_decap_8 FILLER_39_1001 ();
 sg13g2_decap_8 FILLER_39_1008 ();
 sg13g2_decap_8 FILLER_39_1020 ();
 sg13g2_fill_2 FILLER_39_1027 ();
 sg13g2_decap_8 FILLER_39_1033 ();
 sg13g2_decap_8 FILLER_39_1040 ();
 sg13g2_decap_8 FILLER_39_1047 ();
 sg13g2_decap_8 FILLER_39_1054 ();
 sg13g2_decap_8 FILLER_39_1061 ();
 sg13g2_decap_8 FILLER_39_1068 ();
 sg13g2_decap_8 FILLER_39_1075 ();
 sg13g2_decap_8 FILLER_39_1082 ();
 sg13g2_decap_8 FILLER_39_1089 ();
 sg13g2_decap_8 FILLER_39_1096 ();
 sg13g2_decap_8 FILLER_39_1103 ();
 sg13g2_decap_8 FILLER_39_1110 ();
 sg13g2_decap_4 FILLER_39_1117 ();
 sg13g2_fill_1 FILLER_39_1121 ();
 sg13g2_decap_8 FILLER_39_1128 ();
 sg13g2_decap_8 FILLER_39_1135 ();
 sg13g2_decap_8 FILLER_39_1142 ();
 sg13g2_decap_8 FILLER_39_1149 ();
 sg13g2_decap_8 FILLER_39_1156 ();
 sg13g2_decap_4 FILLER_39_1163 ();
 sg13g2_fill_2 FILLER_39_1167 ();
 sg13g2_decap_8 FILLER_39_1172 ();
 sg13g2_decap_8 FILLER_39_1179 ();
 sg13g2_decap_8 FILLER_39_1186 ();
 sg13g2_decap_8 FILLER_39_1193 ();
 sg13g2_decap_8 FILLER_39_1200 ();
 sg13g2_decap_8 FILLER_39_1207 ();
 sg13g2_decap_8 FILLER_39_1214 ();
 sg13g2_decap_8 FILLER_39_1221 ();
 sg13g2_fill_2 FILLER_39_1228 ();
 sg13g2_fill_1 FILLER_39_1230 ();
 sg13g2_decap_8 FILLER_39_1249 ();
 sg13g2_decap_4 FILLER_39_1265 ();
 sg13g2_fill_2 FILLER_39_1269 ();
 sg13g2_decap_8 FILLER_39_1286 ();
 sg13g2_decap_8 FILLER_39_1293 ();
 sg13g2_decap_8 FILLER_39_1300 ();
 sg13g2_decap_8 FILLER_39_1307 ();
 sg13g2_decap_8 FILLER_39_1314 ();
 sg13g2_fill_2 FILLER_39_1321 ();
 sg13g2_decap_8 FILLER_39_1347 ();
 sg13g2_decap_8 FILLER_39_1354 ();
 sg13g2_fill_2 FILLER_39_1361 ();
 sg13g2_decap_8 FILLER_39_1368 ();
 sg13g2_decap_8 FILLER_39_1375 ();
 sg13g2_decap_8 FILLER_39_1382 ();
 sg13g2_decap_8 FILLER_39_1389 ();
 sg13g2_decap_8 FILLER_39_1396 ();
 sg13g2_decap_8 FILLER_39_1403 ();
 sg13g2_decap_8 FILLER_39_1410 ();
 sg13g2_decap_8 FILLER_39_1417 ();
 sg13g2_decap_8 FILLER_39_1424 ();
 sg13g2_decap_4 FILLER_39_1431 ();
 sg13g2_fill_2 FILLER_39_1435 ();
 sg13g2_decap_4 FILLER_39_1440 ();
 sg13g2_fill_1 FILLER_39_1444 ();
 sg13g2_decap_8 FILLER_39_1460 ();
 sg13g2_decap_8 FILLER_39_1467 ();
 sg13g2_decap_8 FILLER_39_1474 ();
 sg13g2_decap_8 FILLER_39_1481 ();
 sg13g2_decap_8 FILLER_39_1488 ();
 sg13g2_decap_4 FILLER_39_1495 ();
 sg13g2_fill_2 FILLER_39_1499 ();
 sg13g2_decap_4 FILLER_39_1511 ();
 sg13g2_decap_8 FILLER_39_1521 ();
 sg13g2_decap_8 FILLER_39_1528 ();
 sg13g2_decap_8 FILLER_39_1535 ();
 sg13g2_decap_8 FILLER_39_1542 ();
 sg13g2_decap_8 FILLER_39_1549 ();
 sg13g2_decap_8 FILLER_39_1556 ();
 sg13g2_decap_8 FILLER_39_1563 ();
 sg13g2_decap_8 FILLER_39_1570 ();
 sg13g2_decap_8 FILLER_39_1577 ();
 sg13g2_decap_8 FILLER_39_1584 ();
 sg13g2_decap_8 FILLER_39_1591 ();
 sg13g2_decap_8 FILLER_39_1598 ();
 sg13g2_decap_8 FILLER_39_1605 ();
 sg13g2_decap_8 FILLER_39_1612 ();
 sg13g2_fill_2 FILLER_39_1619 ();
 sg13g2_fill_1 FILLER_39_1621 ();
 sg13g2_decap_8 FILLER_39_1630 ();
 sg13g2_decap_8 FILLER_39_1640 ();
 sg13g2_decap_8 FILLER_39_1647 ();
 sg13g2_decap_8 FILLER_39_1654 ();
 sg13g2_decap_4 FILLER_39_1661 ();
 sg13g2_decap_8 FILLER_39_1671 ();
 sg13g2_decap_8 FILLER_39_1678 ();
 sg13g2_decap_8 FILLER_39_1685 ();
 sg13g2_decap_8 FILLER_39_1692 ();
 sg13g2_fill_2 FILLER_39_1699 ();
 sg13g2_fill_1 FILLER_39_1701 ();
 sg13g2_decap_8 FILLER_39_1708 ();
 sg13g2_decap_8 FILLER_39_1715 ();
 sg13g2_decap_8 FILLER_39_1722 ();
 sg13g2_decap_8 FILLER_39_1729 ();
 sg13g2_decap_8 FILLER_39_1736 ();
 sg13g2_fill_2 FILLER_39_1743 ();
 sg13g2_fill_1 FILLER_39_1745 ();
 sg13g2_decap_8 FILLER_39_1762 ();
 sg13g2_decap_8 FILLER_39_1769 ();
 sg13g2_decap_8 FILLER_39_1776 ();
 sg13g2_decap_8 FILLER_39_1783 ();
 sg13g2_decap_8 FILLER_39_1790 ();
 sg13g2_decap_8 FILLER_39_1797 ();
 sg13g2_decap_8 FILLER_39_1804 ();
 sg13g2_decap_8 FILLER_39_1811 ();
 sg13g2_decap_8 FILLER_39_1818 ();
 sg13g2_decap_8 FILLER_39_1825 ();
 sg13g2_decap_8 FILLER_39_1832 ();
 sg13g2_decap_8 FILLER_39_1839 ();
 sg13g2_decap_8 FILLER_39_1846 ();
 sg13g2_decap_8 FILLER_39_1853 ();
 sg13g2_decap_8 FILLER_39_1860 ();
 sg13g2_decap_8 FILLER_39_1867 ();
 sg13g2_decap_8 FILLER_39_1874 ();
 sg13g2_decap_8 FILLER_39_1881 ();
 sg13g2_decap_8 FILLER_39_1888 ();
 sg13g2_decap_8 FILLER_39_1895 ();
 sg13g2_decap_8 FILLER_39_1902 ();
 sg13g2_decap_8 FILLER_39_1909 ();
 sg13g2_decap_8 FILLER_39_1916 ();
 sg13g2_decap_8 FILLER_39_1923 ();
 sg13g2_decap_8 FILLER_39_1930 ();
 sg13g2_decap_8 FILLER_39_1937 ();
 sg13g2_decap_8 FILLER_39_1944 ();
 sg13g2_decap_8 FILLER_39_1951 ();
 sg13g2_decap_8 FILLER_39_1958 ();
 sg13g2_decap_8 FILLER_39_1965 ();
 sg13g2_decap_8 FILLER_39_1972 ();
 sg13g2_decap_8 FILLER_39_1979 ();
 sg13g2_fill_2 FILLER_39_1986 ();
 sg13g2_fill_1 FILLER_39_1988 ();
 sg13g2_decap_8 FILLER_39_1993 ();
 sg13g2_decap_8 FILLER_39_2000 ();
 sg13g2_decap_8 FILLER_39_2007 ();
 sg13g2_decap_8 FILLER_39_2014 ();
 sg13g2_decap_8 FILLER_39_2021 ();
 sg13g2_decap_8 FILLER_39_2028 ();
 sg13g2_decap_8 FILLER_39_2035 ();
 sg13g2_decap_8 FILLER_39_2042 ();
 sg13g2_decap_8 FILLER_39_2049 ();
 sg13g2_decap_8 FILLER_39_2056 ();
 sg13g2_decap_8 FILLER_39_2063 ();
 sg13g2_decap_8 FILLER_39_2070 ();
 sg13g2_decap_8 FILLER_39_2077 ();
 sg13g2_decap_8 FILLER_39_2084 ();
 sg13g2_decap_8 FILLER_39_2091 ();
 sg13g2_decap_8 FILLER_39_2098 ();
 sg13g2_decap_8 FILLER_39_2105 ();
 sg13g2_decap_8 FILLER_39_2112 ();
 sg13g2_decap_8 FILLER_39_2119 ();
 sg13g2_decap_8 FILLER_39_2126 ();
 sg13g2_decap_8 FILLER_39_2133 ();
 sg13g2_decap_8 FILLER_39_2140 ();
 sg13g2_decap_8 FILLER_39_2147 ();
 sg13g2_decap_8 FILLER_39_2154 ();
 sg13g2_decap_8 FILLER_39_2161 ();
 sg13g2_decap_8 FILLER_39_2168 ();
 sg13g2_decap_8 FILLER_39_2175 ();
 sg13g2_decap_8 FILLER_39_2182 ();
 sg13g2_decap_8 FILLER_39_2189 ();
 sg13g2_decap_8 FILLER_39_2196 ();
 sg13g2_decap_8 FILLER_39_2203 ();
 sg13g2_decap_8 FILLER_39_2210 ();
 sg13g2_decap_8 FILLER_39_2217 ();
 sg13g2_decap_8 FILLER_39_2224 ();
 sg13g2_decap_8 FILLER_39_2231 ();
 sg13g2_decap_8 FILLER_39_2238 ();
 sg13g2_decap_8 FILLER_39_2245 ();
 sg13g2_decap_8 FILLER_39_2252 ();
 sg13g2_decap_8 FILLER_39_2259 ();
 sg13g2_decap_8 FILLER_39_2266 ();
 sg13g2_decap_8 FILLER_39_2273 ();
 sg13g2_decap_8 FILLER_39_2280 ();
 sg13g2_decap_8 FILLER_39_2287 ();
 sg13g2_decap_8 FILLER_39_2294 ();
 sg13g2_decap_8 FILLER_39_2301 ();
 sg13g2_decap_8 FILLER_39_2308 ();
 sg13g2_decap_8 FILLER_39_2315 ();
 sg13g2_decap_8 FILLER_39_2322 ();
 sg13g2_decap_8 FILLER_39_2329 ();
 sg13g2_decap_8 FILLER_39_2336 ();
 sg13g2_decap_8 FILLER_39_2343 ();
 sg13g2_decap_8 FILLER_39_2350 ();
 sg13g2_decap_8 FILLER_39_2357 ();
 sg13g2_decap_8 FILLER_39_2364 ();
 sg13g2_decap_8 FILLER_39_2371 ();
 sg13g2_decap_8 FILLER_39_2378 ();
 sg13g2_decap_8 FILLER_39_2385 ();
 sg13g2_decap_8 FILLER_39_2392 ();
 sg13g2_decap_8 FILLER_39_2399 ();
 sg13g2_decap_8 FILLER_39_2406 ();
 sg13g2_decap_8 FILLER_39_2413 ();
 sg13g2_decap_8 FILLER_39_2420 ();
 sg13g2_decap_8 FILLER_39_2427 ();
 sg13g2_decap_8 FILLER_39_2434 ();
 sg13g2_decap_8 FILLER_39_2441 ();
 sg13g2_decap_8 FILLER_39_2448 ();
 sg13g2_decap_8 FILLER_39_2455 ();
 sg13g2_decap_8 FILLER_39_2462 ();
 sg13g2_decap_8 FILLER_39_2469 ();
 sg13g2_decap_8 FILLER_39_2476 ();
 sg13g2_decap_8 FILLER_39_2483 ();
 sg13g2_decap_8 FILLER_39_2490 ();
 sg13g2_decap_8 FILLER_39_2497 ();
 sg13g2_decap_8 FILLER_39_2504 ();
 sg13g2_decap_8 FILLER_39_2511 ();
 sg13g2_decap_8 FILLER_39_2518 ();
 sg13g2_decap_8 FILLER_39_2525 ();
 sg13g2_decap_8 FILLER_39_2532 ();
 sg13g2_decap_8 FILLER_39_2539 ();
 sg13g2_decap_8 FILLER_39_2546 ();
 sg13g2_decap_8 FILLER_39_2553 ();
 sg13g2_decap_8 FILLER_39_2560 ();
 sg13g2_decap_8 FILLER_39_2567 ();
 sg13g2_decap_8 FILLER_39_2574 ();
 sg13g2_decap_8 FILLER_39_2581 ();
 sg13g2_decap_8 FILLER_39_2588 ();
 sg13g2_decap_8 FILLER_39_2595 ();
 sg13g2_decap_8 FILLER_39_2602 ();
 sg13g2_decap_8 FILLER_39_2609 ();
 sg13g2_decap_8 FILLER_39_2616 ();
 sg13g2_decap_8 FILLER_39_2623 ();
 sg13g2_decap_8 FILLER_39_2630 ();
 sg13g2_decap_8 FILLER_39_2637 ();
 sg13g2_decap_8 FILLER_39_2644 ();
 sg13g2_decap_8 FILLER_39_2651 ();
 sg13g2_decap_8 FILLER_39_2658 ();
 sg13g2_decap_4 FILLER_39_2665 ();
 sg13g2_fill_1 FILLER_39_2669 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_4 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_50 ();
 sg13g2_fill_1 FILLER_40_57 ();
 sg13g2_decap_4 FILLER_40_62 ();
 sg13g2_fill_2 FILLER_40_66 ();
 sg13g2_decap_8 FILLER_40_73 ();
 sg13g2_decap_8 FILLER_40_80 ();
 sg13g2_fill_2 FILLER_40_87 ();
 sg13g2_fill_1 FILLER_40_89 ();
 sg13g2_decap_8 FILLER_40_94 ();
 sg13g2_decap_8 FILLER_40_101 ();
 sg13g2_decap_8 FILLER_40_108 ();
 sg13g2_decap_8 FILLER_40_115 ();
 sg13g2_decap_8 FILLER_40_122 ();
 sg13g2_decap_8 FILLER_40_129 ();
 sg13g2_decap_8 FILLER_40_136 ();
 sg13g2_decap_8 FILLER_40_143 ();
 sg13g2_fill_2 FILLER_40_150 ();
 sg13g2_fill_1 FILLER_40_152 ();
 sg13g2_decap_8 FILLER_40_156 ();
 sg13g2_decap_8 FILLER_40_163 ();
 sg13g2_decap_8 FILLER_40_170 ();
 sg13g2_fill_2 FILLER_40_177 ();
 sg13g2_decap_4 FILLER_40_184 ();
 sg13g2_fill_1 FILLER_40_188 ();
 sg13g2_decap_8 FILLER_40_194 ();
 sg13g2_decap_8 FILLER_40_201 ();
 sg13g2_decap_8 FILLER_40_216 ();
 sg13g2_decap_8 FILLER_40_223 ();
 sg13g2_decap_8 FILLER_40_230 ();
 sg13g2_decap_4 FILLER_40_237 ();
 sg13g2_decap_8 FILLER_40_245 ();
 sg13g2_decap_8 FILLER_40_252 ();
 sg13g2_decap_8 FILLER_40_259 ();
 sg13g2_decap_8 FILLER_40_266 ();
 sg13g2_decap_8 FILLER_40_273 ();
 sg13g2_decap_8 FILLER_40_280 ();
 sg13g2_decap_8 FILLER_40_287 ();
 sg13g2_decap_8 FILLER_40_294 ();
 sg13g2_decap_8 FILLER_40_301 ();
 sg13g2_decap_8 FILLER_40_308 ();
 sg13g2_decap_8 FILLER_40_315 ();
 sg13g2_fill_1 FILLER_40_322 ();
 sg13g2_decap_8 FILLER_40_331 ();
 sg13g2_fill_1 FILLER_40_338 ();
 sg13g2_decap_8 FILLER_40_343 ();
 sg13g2_decap_8 FILLER_40_350 ();
 sg13g2_decap_8 FILLER_40_357 ();
 sg13g2_decap_8 FILLER_40_364 ();
 sg13g2_decap_8 FILLER_40_371 ();
 sg13g2_decap_8 FILLER_40_378 ();
 sg13g2_decap_8 FILLER_40_385 ();
 sg13g2_decap_8 FILLER_40_392 ();
 sg13g2_decap_8 FILLER_40_399 ();
 sg13g2_decap_8 FILLER_40_406 ();
 sg13g2_decap_8 FILLER_40_413 ();
 sg13g2_decap_8 FILLER_40_420 ();
 sg13g2_decap_8 FILLER_40_427 ();
 sg13g2_decap_8 FILLER_40_434 ();
 sg13g2_decap_8 FILLER_40_441 ();
 sg13g2_decap_8 FILLER_40_448 ();
 sg13g2_decap_8 FILLER_40_455 ();
 sg13g2_decap_8 FILLER_40_462 ();
 sg13g2_decap_8 FILLER_40_469 ();
 sg13g2_decap_8 FILLER_40_476 ();
 sg13g2_decap_8 FILLER_40_483 ();
 sg13g2_decap_8 FILLER_40_490 ();
 sg13g2_decap_8 FILLER_40_497 ();
 sg13g2_decap_8 FILLER_40_504 ();
 sg13g2_decap_8 FILLER_40_511 ();
 sg13g2_decap_8 FILLER_40_518 ();
 sg13g2_decap_8 FILLER_40_525 ();
 sg13g2_decap_8 FILLER_40_532 ();
 sg13g2_decap_8 FILLER_40_539 ();
 sg13g2_decap_8 FILLER_40_546 ();
 sg13g2_decap_8 FILLER_40_553 ();
 sg13g2_decap_8 FILLER_40_560 ();
 sg13g2_decap_4 FILLER_40_567 ();
 sg13g2_fill_2 FILLER_40_571 ();
 sg13g2_decap_8 FILLER_40_581 ();
 sg13g2_decap_8 FILLER_40_588 ();
 sg13g2_decap_8 FILLER_40_595 ();
 sg13g2_decap_8 FILLER_40_602 ();
 sg13g2_decap_4 FILLER_40_609 ();
 sg13g2_fill_2 FILLER_40_617 ();
 sg13g2_decap_8 FILLER_40_623 ();
 sg13g2_decap_8 FILLER_40_630 ();
 sg13g2_decap_8 FILLER_40_637 ();
 sg13g2_fill_1 FILLER_40_644 ();
 sg13g2_decap_4 FILLER_40_650 ();
 sg13g2_fill_2 FILLER_40_654 ();
 sg13g2_fill_2 FILLER_40_675 ();
 sg13g2_decap_8 FILLER_40_688 ();
 sg13g2_decap_8 FILLER_40_695 ();
 sg13g2_decap_8 FILLER_40_702 ();
 sg13g2_decap_8 FILLER_40_709 ();
 sg13g2_decap_8 FILLER_40_716 ();
 sg13g2_decap_8 FILLER_40_723 ();
 sg13g2_decap_8 FILLER_40_730 ();
 sg13g2_decap_8 FILLER_40_737 ();
 sg13g2_decap_8 FILLER_40_744 ();
 sg13g2_fill_1 FILLER_40_751 ();
 sg13g2_decap_8 FILLER_40_769 ();
 sg13g2_decap_4 FILLER_40_776 ();
 sg13g2_decap_4 FILLER_40_784 ();
 sg13g2_fill_1 FILLER_40_792 ();
 sg13g2_decap_8 FILLER_40_806 ();
 sg13g2_decap_8 FILLER_40_813 ();
 sg13g2_decap_8 FILLER_40_820 ();
 sg13g2_fill_2 FILLER_40_827 ();
 sg13g2_decap_8 FILLER_40_834 ();
 sg13g2_decap_8 FILLER_40_841 ();
 sg13g2_decap_8 FILLER_40_848 ();
 sg13g2_decap_8 FILLER_40_855 ();
 sg13g2_fill_2 FILLER_40_862 ();
 sg13g2_fill_1 FILLER_40_864 ();
 sg13g2_decap_8 FILLER_40_880 ();
 sg13g2_fill_2 FILLER_40_891 ();
 sg13g2_fill_1 FILLER_40_893 ();
 sg13g2_decap_8 FILLER_40_904 ();
 sg13g2_decap_8 FILLER_40_911 ();
 sg13g2_decap_8 FILLER_40_918 ();
 sg13g2_decap_8 FILLER_40_925 ();
 sg13g2_decap_8 FILLER_40_932 ();
 sg13g2_decap_8 FILLER_40_939 ();
 sg13g2_decap_8 FILLER_40_946 ();
 sg13g2_fill_2 FILLER_40_953 ();
 sg13g2_fill_1 FILLER_40_955 ();
 sg13g2_decap_8 FILLER_40_960 ();
 sg13g2_decap_8 FILLER_40_967 ();
 sg13g2_decap_8 FILLER_40_974 ();
 sg13g2_decap_8 FILLER_40_981 ();
 sg13g2_decap_8 FILLER_40_988 ();
 sg13g2_fill_2 FILLER_40_995 ();
 sg13g2_decap_8 FILLER_40_1005 ();
 sg13g2_decap_8 FILLER_40_1012 ();
 sg13g2_decap_8 FILLER_40_1019 ();
 sg13g2_decap_8 FILLER_40_1026 ();
 sg13g2_decap_8 FILLER_40_1033 ();
 sg13g2_decap_8 FILLER_40_1040 ();
 sg13g2_decap_8 FILLER_40_1047 ();
 sg13g2_decap_8 FILLER_40_1054 ();
 sg13g2_decap_4 FILLER_40_1061 ();
 sg13g2_fill_1 FILLER_40_1065 ();
 sg13g2_decap_4 FILLER_40_1071 ();
 sg13g2_fill_2 FILLER_40_1075 ();
 sg13g2_decap_8 FILLER_40_1085 ();
 sg13g2_decap_8 FILLER_40_1092 ();
 sg13g2_decap_8 FILLER_40_1099 ();
 sg13g2_decap_8 FILLER_40_1106 ();
 sg13g2_decap_8 FILLER_40_1113 ();
 sg13g2_decap_8 FILLER_40_1120 ();
 sg13g2_decap_8 FILLER_40_1127 ();
 sg13g2_decap_8 FILLER_40_1134 ();
 sg13g2_fill_2 FILLER_40_1141 ();
 sg13g2_fill_2 FILLER_40_1155 ();
 sg13g2_decap_8 FILLER_40_1163 ();
 sg13g2_decap_8 FILLER_40_1170 ();
 sg13g2_decap_8 FILLER_40_1177 ();
 sg13g2_decap_8 FILLER_40_1184 ();
 sg13g2_decap_8 FILLER_40_1191 ();
 sg13g2_decap_8 FILLER_40_1198 ();
 sg13g2_decap_8 FILLER_40_1205 ();
 sg13g2_decap_8 FILLER_40_1212 ();
 sg13g2_decap_8 FILLER_40_1219 ();
 sg13g2_fill_2 FILLER_40_1226 ();
 sg13g2_decap_8 FILLER_40_1249 ();
 sg13g2_fill_1 FILLER_40_1261 ();
 sg13g2_decap_8 FILLER_40_1282 ();
 sg13g2_decap_8 FILLER_40_1289 ();
 sg13g2_decap_8 FILLER_40_1296 ();
 sg13g2_fill_1 FILLER_40_1303 ();
 sg13g2_decap_8 FILLER_40_1308 ();
 sg13g2_decap_8 FILLER_40_1315 ();
 sg13g2_decap_8 FILLER_40_1322 ();
 sg13g2_decap_4 FILLER_40_1329 ();
 sg13g2_fill_2 FILLER_40_1333 ();
 sg13g2_decap_4 FILLER_40_1340 ();
 sg13g2_decap_8 FILLER_40_1347 ();
 sg13g2_decap_8 FILLER_40_1354 ();
 sg13g2_decap_8 FILLER_40_1361 ();
 sg13g2_decap_8 FILLER_40_1368 ();
 sg13g2_decap_8 FILLER_40_1375 ();
 sg13g2_decap_8 FILLER_40_1382 ();
 sg13g2_decap_8 FILLER_40_1389 ();
 sg13g2_fill_1 FILLER_40_1396 ();
 sg13g2_decap_8 FILLER_40_1402 ();
 sg13g2_decap_8 FILLER_40_1409 ();
 sg13g2_decap_8 FILLER_40_1416 ();
 sg13g2_decap_8 FILLER_40_1423 ();
 sg13g2_decap_8 FILLER_40_1430 ();
 sg13g2_decap_8 FILLER_40_1437 ();
 sg13g2_fill_1 FILLER_40_1444 ();
 sg13g2_decap_8 FILLER_40_1450 ();
 sg13g2_decap_8 FILLER_40_1457 ();
 sg13g2_decap_8 FILLER_40_1464 ();
 sg13g2_fill_2 FILLER_40_1471 ();
 sg13g2_fill_1 FILLER_40_1473 ();
 sg13g2_decap_8 FILLER_40_1477 ();
 sg13g2_decap_8 FILLER_40_1484 ();
 sg13g2_decap_8 FILLER_40_1491 ();
 sg13g2_decap_8 FILLER_40_1498 ();
 sg13g2_decap_8 FILLER_40_1505 ();
 sg13g2_decap_8 FILLER_40_1512 ();
 sg13g2_decap_8 FILLER_40_1519 ();
 sg13g2_decap_8 FILLER_40_1526 ();
 sg13g2_decap_8 FILLER_40_1533 ();
 sg13g2_decap_8 FILLER_40_1540 ();
 sg13g2_decap_4 FILLER_40_1552 ();
 sg13g2_decap_8 FILLER_40_1562 ();
 sg13g2_decap_8 FILLER_40_1569 ();
 sg13g2_decap_8 FILLER_40_1576 ();
 sg13g2_decap_8 FILLER_40_1583 ();
 sg13g2_decap_8 FILLER_40_1590 ();
 sg13g2_fill_2 FILLER_40_1597 ();
 sg13g2_decap_8 FILLER_40_1603 ();
 sg13g2_decap_8 FILLER_40_1610 ();
 sg13g2_decap_4 FILLER_40_1617 ();
 sg13g2_fill_2 FILLER_40_1621 ();
 sg13g2_decap_4 FILLER_40_1629 ();
 sg13g2_fill_1 FILLER_40_1633 ();
 sg13g2_decap_8 FILLER_40_1644 ();
 sg13g2_decap_8 FILLER_40_1651 ();
 sg13g2_fill_2 FILLER_40_1658 ();
 sg13g2_fill_1 FILLER_40_1660 ();
 sg13g2_decap_8 FILLER_40_1673 ();
 sg13g2_decap_8 FILLER_40_1680 ();
 sg13g2_decap_4 FILLER_40_1687 ();
 sg13g2_fill_1 FILLER_40_1691 ();
 sg13g2_decap_8 FILLER_40_1698 ();
 sg13g2_decap_8 FILLER_40_1705 ();
 sg13g2_decap_8 FILLER_40_1712 ();
 sg13g2_decap_8 FILLER_40_1719 ();
 sg13g2_decap_8 FILLER_40_1726 ();
 sg13g2_decap_8 FILLER_40_1733 ();
 sg13g2_decap_8 FILLER_40_1740 ();
 sg13g2_decap_8 FILLER_40_1747 ();
 sg13g2_decap_8 FILLER_40_1754 ();
 sg13g2_fill_1 FILLER_40_1761 ();
 sg13g2_decap_8 FILLER_40_1765 ();
 sg13g2_decap_8 FILLER_40_1772 ();
 sg13g2_decap_8 FILLER_40_1779 ();
 sg13g2_decap_8 FILLER_40_1786 ();
 sg13g2_decap_8 FILLER_40_1793 ();
 sg13g2_decap_8 FILLER_40_1800 ();
 sg13g2_decap_4 FILLER_40_1807 ();
 sg13g2_fill_2 FILLER_40_1811 ();
 sg13g2_decap_8 FILLER_40_1826 ();
 sg13g2_decap_8 FILLER_40_1833 ();
 sg13g2_decap_8 FILLER_40_1840 ();
 sg13g2_decap_8 FILLER_40_1847 ();
 sg13g2_fill_2 FILLER_40_1854 ();
 sg13g2_decap_8 FILLER_40_1864 ();
 sg13g2_decap_8 FILLER_40_1871 ();
 sg13g2_decap_8 FILLER_40_1878 ();
 sg13g2_decap_8 FILLER_40_1885 ();
 sg13g2_decap_8 FILLER_40_1892 ();
 sg13g2_decap_8 FILLER_40_1899 ();
 sg13g2_decap_8 FILLER_40_1906 ();
 sg13g2_decap_8 FILLER_40_1913 ();
 sg13g2_decap_8 FILLER_40_1920 ();
 sg13g2_decap_8 FILLER_40_1927 ();
 sg13g2_decap_8 FILLER_40_1934 ();
 sg13g2_decap_4 FILLER_40_1941 ();
 sg13g2_decap_8 FILLER_40_1949 ();
 sg13g2_decap_8 FILLER_40_1956 ();
 sg13g2_decap_8 FILLER_40_1963 ();
 sg13g2_decap_4 FILLER_40_1970 ();
 sg13g2_decap_4 FILLER_40_1978 ();
 sg13g2_fill_1 FILLER_40_1982 ();
 sg13g2_decap_8 FILLER_40_2009 ();
 sg13g2_decap_8 FILLER_40_2016 ();
 sg13g2_decap_8 FILLER_40_2023 ();
 sg13g2_decap_8 FILLER_40_2030 ();
 sg13g2_decap_8 FILLER_40_2037 ();
 sg13g2_decap_8 FILLER_40_2044 ();
 sg13g2_decap_8 FILLER_40_2051 ();
 sg13g2_decap_8 FILLER_40_2058 ();
 sg13g2_decap_8 FILLER_40_2065 ();
 sg13g2_decap_8 FILLER_40_2072 ();
 sg13g2_decap_8 FILLER_40_2079 ();
 sg13g2_decap_8 FILLER_40_2086 ();
 sg13g2_decap_8 FILLER_40_2093 ();
 sg13g2_decap_8 FILLER_40_2100 ();
 sg13g2_decap_8 FILLER_40_2107 ();
 sg13g2_decap_8 FILLER_40_2114 ();
 sg13g2_decap_8 FILLER_40_2121 ();
 sg13g2_decap_8 FILLER_40_2128 ();
 sg13g2_decap_8 FILLER_40_2135 ();
 sg13g2_decap_8 FILLER_40_2142 ();
 sg13g2_decap_8 FILLER_40_2149 ();
 sg13g2_decap_8 FILLER_40_2156 ();
 sg13g2_decap_8 FILLER_40_2163 ();
 sg13g2_decap_8 FILLER_40_2170 ();
 sg13g2_decap_8 FILLER_40_2177 ();
 sg13g2_decap_8 FILLER_40_2184 ();
 sg13g2_decap_8 FILLER_40_2191 ();
 sg13g2_decap_8 FILLER_40_2198 ();
 sg13g2_decap_8 FILLER_40_2205 ();
 sg13g2_decap_8 FILLER_40_2212 ();
 sg13g2_decap_8 FILLER_40_2219 ();
 sg13g2_decap_8 FILLER_40_2226 ();
 sg13g2_decap_8 FILLER_40_2233 ();
 sg13g2_decap_8 FILLER_40_2240 ();
 sg13g2_decap_8 FILLER_40_2247 ();
 sg13g2_decap_8 FILLER_40_2254 ();
 sg13g2_decap_8 FILLER_40_2261 ();
 sg13g2_decap_8 FILLER_40_2268 ();
 sg13g2_decap_8 FILLER_40_2275 ();
 sg13g2_decap_8 FILLER_40_2282 ();
 sg13g2_decap_8 FILLER_40_2289 ();
 sg13g2_decap_8 FILLER_40_2296 ();
 sg13g2_decap_8 FILLER_40_2303 ();
 sg13g2_decap_8 FILLER_40_2310 ();
 sg13g2_decap_8 FILLER_40_2317 ();
 sg13g2_decap_8 FILLER_40_2324 ();
 sg13g2_decap_8 FILLER_40_2331 ();
 sg13g2_decap_8 FILLER_40_2338 ();
 sg13g2_decap_8 FILLER_40_2345 ();
 sg13g2_decap_8 FILLER_40_2352 ();
 sg13g2_decap_8 FILLER_40_2359 ();
 sg13g2_decap_8 FILLER_40_2366 ();
 sg13g2_decap_8 FILLER_40_2373 ();
 sg13g2_decap_8 FILLER_40_2380 ();
 sg13g2_decap_8 FILLER_40_2387 ();
 sg13g2_decap_8 FILLER_40_2394 ();
 sg13g2_decap_8 FILLER_40_2401 ();
 sg13g2_decap_8 FILLER_40_2408 ();
 sg13g2_decap_8 FILLER_40_2415 ();
 sg13g2_decap_8 FILLER_40_2422 ();
 sg13g2_decap_8 FILLER_40_2429 ();
 sg13g2_decap_8 FILLER_40_2436 ();
 sg13g2_decap_8 FILLER_40_2443 ();
 sg13g2_decap_8 FILLER_40_2450 ();
 sg13g2_decap_8 FILLER_40_2457 ();
 sg13g2_decap_8 FILLER_40_2464 ();
 sg13g2_decap_8 FILLER_40_2471 ();
 sg13g2_decap_8 FILLER_40_2478 ();
 sg13g2_decap_8 FILLER_40_2485 ();
 sg13g2_decap_8 FILLER_40_2492 ();
 sg13g2_decap_8 FILLER_40_2499 ();
 sg13g2_decap_8 FILLER_40_2506 ();
 sg13g2_decap_8 FILLER_40_2513 ();
 sg13g2_decap_8 FILLER_40_2520 ();
 sg13g2_decap_8 FILLER_40_2527 ();
 sg13g2_decap_8 FILLER_40_2534 ();
 sg13g2_decap_8 FILLER_40_2541 ();
 sg13g2_decap_8 FILLER_40_2548 ();
 sg13g2_decap_8 FILLER_40_2555 ();
 sg13g2_decap_8 FILLER_40_2562 ();
 sg13g2_decap_8 FILLER_40_2569 ();
 sg13g2_decap_8 FILLER_40_2576 ();
 sg13g2_decap_8 FILLER_40_2583 ();
 sg13g2_decap_8 FILLER_40_2590 ();
 sg13g2_decap_8 FILLER_40_2597 ();
 sg13g2_decap_8 FILLER_40_2604 ();
 sg13g2_decap_8 FILLER_40_2611 ();
 sg13g2_decap_8 FILLER_40_2618 ();
 sg13g2_decap_8 FILLER_40_2625 ();
 sg13g2_decap_8 FILLER_40_2632 ();
 sg13g2_decap_8 FILLER_40_2639 ();
 sg13g2_decap_8 FILLER_40_2646 ();
 sg13g2_decap_8 FILLER_40_2653 ();
 sg13g2_decap_8 FILLER_40_2660 ();
 sg13g2_fill_2 FILLER_40_2667 ();
 sg13g2_fill_1 FILLER_40_2669 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_fill_2 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_64 ();
 sg13g2_decap_8 FILLER_41_71 ();
 sg13g2_decap_8 FILLER_41_78 ();
 sg13g2_decap_8 FILLER_41_85 ();
 sg13g2_decap_8 FILLER_41_92 ();
 sg13g2_decap_4 FILLER_41_99 ();
 sg13g2_fill_2 FILLER_41_103 ();
 sg13g2_fill_2 FILLER_41_109 ();
 sg13g2_decap_8 FILLER_41_123 ();
 sg13g2_decap_8 FILLER_41_135 ();
 sg13g2_decap_8 FILLER_41_142 ();
 sg13g2_decap_8 FILLER_41_149 ();
 sg13g2_decap_4 FILLER_41_156 ();
 sg13g2_fill_2 FILLER_41_160 ();
 sg13g2_decap_8 FILLER_41_167 ();
 sg13g2_decap_8 FILLER_41_174 ();
 sg13g2_decap_8 FILLER_41_181 ();
 sg13g2_decap_8 FILLER_41_188 ();
 sg13g2_decap_8 FILLER_41_195 ();
 sg13g2_decap_8 FILLER_41_202 ();
 sg13g2_decap_8 FILLER_41_209 ();
 sg13g2_decap_8 FILLER_41_216 ();
 sg13g2_decap_8 FILLER_41_223 ();
 sg13g2_decap_8 FILLER_41_230 ();
 sg13g2_decap_8 FILLER_41_237 ();
 sg13g2_decap_8 FILLER_41_244 ();
 sg13g2_decap_8 FILLER_41_251 ();
 sg13g2_decap_8 FILLER_41_258 ();
 sg13g2_fill_1 FILLER_41_265 ();
 sg13g2_decap_4 FILLER_41_271 ();
 sg13g2_decap_8 FILLER_41_279 ();
 sg13g2_decap_8 FILLER_41_286 ();
 sg13g2_decap_8 FILLER_41_293 ();
 sg13g2_decap_8 FILLER_41_300 ();
 sg13g2_decap_8 FILLER_41_307 ();
 sg13g2_decap_8 FILLER_41_314 ();
 sg13g2_fill_2 FILLER_41_321 ();
 sg13g2_decap_8 FILLER_41_328 ();
 sg13g2_fill_2 FILLER_41_335 ();
 sg13g2_fill_1 FILLER_41_337 ();
 sg13g2_decap_8 FILLER_41_343 ();
 sg13g2_decap_8 FILLER_41_350 ();
 sg13g2_decap_8 FILLER_41_357 ();
 sg13g2_decap_8 FILLER_41_364 ();
 sg13g2_decap_8 FILLER_41_371 ();
 sg13g2_decap_8 FILLER_41_378 ();
 sg13g2_decap_8 FILLER_41_385 ();
 sg13g2_decap_8 FILLER_41_392 ();
 sg13g2_decap_8 FILLER_41_399 ();
 sg13g2_decap_8 FILLER_41_406 ();
 sg13g2_decap_8 FILLER_41_413 ();
 sg13g2_fill_2 FILLER_41_420 ();
 sg13g2_decap_8 FILLER_41_426 ();
 sg13g2_decap_8 FILLER_41_433 ();
 sg13g2_decap_8 FILLER_41_440 ();
 sg13g2_decap_8 FILLER_41_447 ();
 sg13g2_decap_8 FILLER_41_454 ();
 sg13g2_decap_8 FILLER_41_461 ();
 sg13g2_decap_8 FILLER_41_468 ();
 sg13g2_decap_4 FILLER_41_475 ();
 sg13g2_fill_1 FILLER_41_479 ();
 sg13g2_decap_8 FILLER_41_493 ();
 sg13g2_decap_8 FILLER_41_500 ();
 sg13g2_decap_8 FILLER_41_507 ();
 sg13g2_decap_8 FILLER_41_514 ();
 sg13g2_decap_8 FILLER_41_521 ();
 sg13g2_decap_8 FILLER_41_528 ();
 sg13g2_decap_8 FILLER_41_535 ();
 sg13g2_decap_8 FILLER_41_542 ();
 sg13g2_decap_8 FILLER_41_549 ();
 sg13g2_decap_8 FILLER_41_556 ();
 sg13g2_decap_4 FILLER_41_563 ();
 sg13g2_decap_8 FILLER_41_591 ();
 sg13g2_decap_8 FILLER_41_598 ();
 sg13g2_fill_1 FILLER_41_605 ();
 sg13g2_decap_8 FILLER_41_635 ();
 sg13g2_decap_8 FILLER_41_642 ();
 sg13g2_decap_8 FILLER_41_649 ();
 sg13g2_decap_4 FILLER_41_656 ();
 sg13g2_decap_4 FILLER_41_667 ();
 sg13g2_fill_1 FILLER_41_671 ();
 sg13g2_decap_8 FILLER_41_691 ();
 sg13g2_decap_8 FILLER_41_698 ();
 sg13g2_decap_8 FILLER_41_705 ();
 sg13g2_decap_8 FILLER_41_712 ();
 sg13g2_decap_8 FILLER_41_719 ();
 sg13g2_decap_8 FILLER_41_726 ();
 sg13g2_decap_8 FILLER_41_733 ();
 sg13g2_decap_8 FILLER_41_740 ();
 sg13g2_decap_8 FILLER_41_747 ();
 sg13g2_decap_8 FILLER_41_754 ();
 sg13g2_decap_8 FILLER_41_761 ();
 sg13g2_decap_8 FILLER_41_774 ();
 sg13g2_decap_8 FILLER_41_781 ();
 sg13g2_decap_8 FILLER_41_788 ();
 sg13g2_decap_8 FILLER_41_795 ();
 sg13g2_decap_8 FILLER_41_802 ();
 sg13g2_decap_8 FILLER_41_809 ();
 sg13g2_decap_8 FILLER_41_816 ();
 sg13g2_decap_4 FILLER_41_823 ();
 sg13g2_fill_2 FILLER_41_827 ();
 sg13g2_decap_8 FILLER_41_844 ();
 sg13g2_decap_8 FILLER_41_851 ();
 sg13g2_decap_8 FILLER_41_858 ();
 sg13g2_decap_8 FILLER_41_865 ();
 sg13g2_decap_8 FILLER_41_872 ();
 sg13g2_decap_8 FILLER_41_879 ();
 sg13g2_decap_4 FILLER_41_886 ();
 sg13g2_fill_2 FILLER_41_890 ();
 sg13g2_decap_8 FILLER_41_907 ();
 sg13g2_decap_8 FILLER_41_914 ();
 sg13g2_decap_8 FILLER_41_921 ();
 sg13g2_decap_4 FILLER_41_928 ();
 sg13g2_fill_1 FILLER_41_932 ();
 sg13g2_fill_2 FILLER_41_945 ();
 sg13g2_fill_1 FILLER_41_947 ();
 sg13g2_decap_8 FILLER_41_964 ();
 sg13g2_decap_8 FILLER_41_971 ();
 sg13g2_decap_8 FILLER_41_978 ();
 sg13g2_decap_8 FILLER_41_985 ();
 sg13g2_decap_8 FILLER_41_992 ();
 sg13g2_decap_8 FILLER_41_999 ();
 sg13g2_decap_8 FILLER_41_1006 ();
 sg13g2_decap_8 FILLER_41_1013 ();
 sg13g2_decap_8 FILLER_41_1020 ();
 sg13g2_decap_8 FILLER_41_1027 ();
 sg13g2_decap_8 FILLER_41_1034 ();
 sg13g2_decap_4 FILLER_41_1041 ();
 sg13g2_fill_1 FILLER_41_1045 ();
 sg13g2_decap_8 FILLER_41_1061 ();
 sg13g2_decap_8 FILLER_41_1068 ();
 sg13g2_decap_8 FILLER_41_1075 ();
 sg13g2_decap_8 FILLER_41_1082 ();
 sg13g2_decap_8 FILLER_41_1089 ();
 sg13g2_decap_8 FILLER_41_1096 ();
 sg13g2_decap_8 FILLER_41_1103 ();
 sg13g2_decap_8 FILLER_41_1110 ();
 sg13g2_decap_8 FILLER_41_1117 ();
 sg13g2_decap_8 FILLER_41_1124 ();
 sg13g2_fill_1 FILLER_41_1131 ();
 sg13g2_decap_8 FILLER_41_1135 ();
 sg13g2_decap_8 FILLER_41_1142 ();
 sg13g2_decap_8 FILLER_41_1149 ();
 sg13g2_fill_1 FILLER_41_1156 ();
 sg13g2_decap_8 FILLER_41_1162 ();
 sg13g2_decap_8 FILLER_41_1169 ();
 sg13g2_decap_8 FILLER_41_1176 ();
 sg13g2_decap_8 FILLER_41_1183 ();
 sg13g2_decap_8 FILLER_41_1190 ();
 sg13g2_decap_8 FILLER_41_1197 ();
 sg13g2_decap_8 FILLER_41_1204 ();
 sg13g2_decap_8 FILLER_41_1211 ();
 sg13g2_decap_8 FILLER_41_1218 ();
 sg13g2_decap_8 FILLER_41_1225 ();
 sg13g2_decap_8 FILLER_41_1240 ();
 sg13g2_decap_8 FILLER_41_1247 ();
 sg13g2_decap_8 FILLER_41_1254 ();
 sg13g2_decap_8 FILLER_41_1261 ();
 sg13g2_fill_1 FILLER_41_1268 ();
 sg13g2_decap_8 FILLER_41_1278 ();
 sg13g2_decap_8 FILLER_41_1285 ();
 sg13g2_decap_8 FILLER_41_1292 ();
 sg13g2_decap_8 FILLER_41_1299 ();
 sg13g2_decap_8 FILLER_41_1306 ();
 sg13g2_decap_8 FILLER_41_1313 ();
 sg13g2_decap_8 FILLER_41_1320 ();
 sg13g2_decap_8 FILLER_41_1327 ();
 sg13g2_decap_8 FILLER_41_1334 ();
 sg13g2_fill_2 FILLER_41_1341 ();
 sg13g2_fill_1 FILLER_41_1343 ();
 sg13g2_decap_8 FILLER_41_1362 ();
 sg13g2_decap_8 FILLER_41_1369 ();
 sg13g2_decap_8 FILLER_41_1376 ();
 sg13g2_fill_2 FILLER_41_1383 ();
 sg13g2_decap_8 FILLER_41_1388 ();
 sg13g2_decap_8 FILLER_41_1395 ();
 sg13g2_fill_2 FILLER_41_1402 ();
 sg13g2_fill_1 FILLER_41_1404 ();
 sg13g2_decap_8 FILLER_41_1415 ();
 sg13g2_decap_8 FILLER_41_1427 ();
 sg13g2_decap_8 FILLER_41_1434 ();
 sg13g2_decap_8 FILLER_41_1441 ();
 sg13g2_decap_8 FILLER_41_1448 ();
 sg13g2_decap_8 FILLER_41_1455 ();
 sg13g2_decap_8 FILLER_41_1462 ();
 sg13g2_decap_4 FILLER_41_1469 ();
 sg13g2_fill_1 FILLER_41_1473 ();
 sg13g2_decap_8 FILLER_41_1478 ();
 sg13g2_decap_8 FILLER_41_1485 ();
 sg13g2_decap_4 FILLER_41_1492 ();
 sg13g2_decap_8 FILLER_41_1500 ();
 sg13g2_decap_8 FILLER_41_1507 ();
 sg13g2_decap_8 FILLER_41_1514 ();
 sg13g2_decap_4 FILLER_41_1521 ();
 sg13g2_decap_8 FILLER_41_1530 ();
 sg13g2_fill_2 FILLER_41_1537 ();
 sg13g2_fill_1 FILLER_41_1539 ();
 sg13g2_decap_4 FILLER_41_1545 ();
 sg13g2_fill_1 FILLER_41_1549 ();
 sg13g2_decap_8 FILLER_41_1567 ();
 sg13g2_decap_8 FILLER_41_1574 ();
 sg13g2_decap_4 FILLER_41_1581 ();
 sg13g2_fill_1 FILLER_41_1585 ();
 sg13g2_decap_8 FILLER_41_1590 ();
 sg13g2_decap_8 FILLER_41_1597 ();
 sg13g2_fill_2 FILLER_41_1604 ();
 sg13g2_decap_8 FILLER_41_1616 ();
 sg13g2_decap_4 FILLER_41_1623 ();
 sg13g2_fill_2 FILLER_41_1627 ();
 sg13g2_decap_8 FILLER_41_1635 ();
 sg13g2_decap_8 FILLER_41_1642 ();
 sg13g2_decap_4 FILLER_41_1649 ();
 sg13g2_fill_1 FILLER_41_1665 ();
 sg13g2_decap_8 FILLER_41_1675 ();
 sg13g2_decap_8 FILLER_41_1682 ();
 sg13g2_decap_8 FILLER_41_1689 ();
 sg13g2_decap_8 FILLER_41_1696 ();
 sg13g2_decap_8 FILLER_41_1703 ();
 sg13g2_decap_8 FILLER_41_1710 ();
 sg13g2_decap_8 FILLER_41_1717 ();
 sg13g2_decap_8 FILLER_41_1724 ();
 sg13g2_decap_8 FILLER_41_1731 ();
 sg13g2_decap_8 FILLER_41_1738 ();
 sg13g2_decap_8 FILLER_41_1754 ();
 sg13g2_fill_1 FILLER_41_1761 ();
 sg13g2_decap_4 FILLER_41_1766 ();
 sg13g2_fill_1 FILLER_41_1770 ();
 sg13g2_fill_2 FILLER_41_1777 ();
 sg13g2_decap_8 FILLER_41_1782 ();
 sg13g2_decap_8 FILLER_41_1789 ();
 sg13g2_decap_8 FILLER_41_1796 ();
 sg13g2_decap_8 FILLER_41_1803 ();
 sg13g2_decap_8 FILLER_41_1810 ();
 sg13g2_decap_4 FILLER_41_1817 ();
 sg13g2_decap_8 FILLER_41_1825 ();
 sg13g2_decap_8 FILLER_41_1832 ();
 sg13g2_decap_8 FILLER_41_1839 ();
 sg13g2_decap_8 FILLER_41_1846 ();
 sg13g2_fill_2 FILLER_41_1853 ();
 sg13g2_fill_1 FILLER_41_1855 ();
 sg13g2_fill_2 FILLER_41_1861 ();
 sg13g2_decap_8 FILLER_41_1868 ();
 sg13g2_decap_8 FILLER_41_1875 ();
 sg13g2_decap_8 FILLER_41_1882 ();
 sg13g2_decap_8 FILLER_41_1889 ();
 sg13g2_decap_8 FILLER_41_1896 ();
 sg13g2_decap_8 FILLER_41_1903 ();
 sg13g2_decap_8 FILLER_41_1910 ();
 sg13g2_decap_8 FILLER_41_1917 ();
 sg13g2_decap_8 FILLER_41_1924 ();
 sg13g2_decap_8 FILLER_41_1931 ();
 sg13g2_decap_4 FILLER_41_1938 ();
 sg13g2_fill_1 FILLER_41_1942 ();
 sg13g2_decap_4 FILLER_41_1969 ();
 sg13g2_decap_8 FILLER_41_1982 ();
 sg13g2_decap_8 FILLER_41_1989 ();
 sg13g2_decap_8 FILLER_41_1996 ();
 sg13g2_decap_8 FILLER_41_2003 ();
 sg13g2_decap_8 FILLER_41_2010 ();
 sg13g2_decap_8 FILLER_41_2017 ();
 sg13g2_decap_8 FILLER_41_2024 ();
 sg13g2_decap_8 FILLER_41_2031 ();
 sg13g2_decap_8 FILLER_41_2038 ();
 sg13g2_decap_8 FILLER_41_2045 ();
 sg13g2_decap_8 FILLER_41_2052 ();
 sg13g2_decap_8 FILLER_41_2059 ();
 sg13g2_decap_8 FILLER_41_2066 ();
 sg13g2_decap_4 FILLER_41_2073 ();
 sg13g2_fill_1 FILLER_41_2077 ();
 sg13g2_decap_8 FILLER_41_2108 ();
 sg13g2_decap_8 FILLER_41_2115 ();
 sg13g2_decap_8 FILLER_41_2122 ();
 sg13g2_decap_8 FILLER_41_2129 ();
 sg13g2_decap_8 FILLER_41_2140 ();
 sg13g2_decap_8 FILLER_41_2147 ();
 sg13g2_decap_8 FILLER_41_2154 ();
 sg13g2_decap_8 FILLER_41_2161 ();
 sg13g2_decap_8 FILLER_41_2168 ();
 sg13g2_decap_8 FILLER_41_2175 ();
 sg13g2_decap_8 FILLER_41_2182 ();
 sg13g2_decap_8 FILLER_41_2189 ();
 sg13g2_decap_8 FILLER_41_2196 ();
 sg13g2_decap_8 FILLER_41_2203 ();
 sg13g2_decap_8 FILLER_41_2210 ();
 sg13g2_decap_8 FILLER_41_2217 ();
 sg13g2_decap_8 FILLER_41_2224 ();
 sg13g2_decap_8 FILLER_41_2231 ();
 sg13g2_decap_8 FILLER_41_2238 ();
 sg13g2_decap_8 FILLER_41_2245 ();
 sg13g2_decap_8 FILLER_41_2252 ();
 sg13g2_decap_8 FILLER_41_2259 ();
 sg13g2_decap_8 FILLER_41_2266 ();
 sg13g2_decap_8 FILLER_41_2273 ();
 sg13g2_decap_8 FILLER_41_2280 ();
 sg13g2_decap_8 FILLER_41_2287 ();
 sg13g2_decap_8 FILLER_41_2294 ();
 sg13g2_decap_8 FILLER_41_2301 ();
 sg13g2_decap_8 FILLER_41_2308 ();
 sg13g2_decap_8 FILLER_41_2315 ();
 sg13g2_decap_8 FILLER_41_2322 ();
 sg13g2_decap_8 FILLER_41_2329 ();
 sg13g2_decap_8 FILLER_41_2336 ();
 sg13g2_decap_8 FILLER_41_2343 ();
 sg13g2_decap_8 FILLER_41_2350 ();
 sg13g2_decap_8 FILLER_41_2357 ();
 sg13g2_decap_8 FILLER_41_2364 ();
 sg13g2_decap_8 FILLER_41_2371 ();
 sg13g2_decap_8 FILLER_41_2378 ();
 sg13g2_decap_8 FILLER_41_2385 ();
 sg13g2_decap_8 FILLER_41_2392 ();
 sg13g2_decap_8 FILLER_41_2399 ();
 sg13g2_decap_8 FILLER_41_2406 ();
 sg13g2_decap_8 FILLER_41_2413 ();
 sg13g2_decap_8 FILLER_41_2420 ();
 sg13g2_decap_8 FILLER_41_2427 ();
 sg13g2_decap_8 FILLER_41_2434 ();
 sg13g2_decap_8 FILLER_41_2441 ();
 sg13g2_decap_8 FILLER_41_2448 ();
 sg13g2_decap_8 FILLER_41_2455 ();
 sg13g2_decap_8 FILLER_41_2462 ();
 sg13g2_decap_8 FILLER_41_2469 ();
 sg13g2_decap_8 FILLER_41_2476 ();
 sg13g2_decap_8 FILLER_41_2483 ();
 sg13g2_decap_8 FILLER_41_2490 ();
 sg13g2_decap_8 FILLER_41_2497 ();
 sg13g2_decap_8 FILLER_41_2504 ();
 sg13g2_decap_8 FILLER_41_2511 ();
 sg13g2_decap_8 FILLER_41_2518 ();
 sg13g2_decap_8 FILLER_41_2525 ();
 sg13g2_decap_8 FILLER_41_2532 ();
 sg13g2_decap_8 FILLER_41_2539 ();
 sg13g2_decap_8 FILLER_41_2546 ();
 sg13g2_decap_8 FILLER_41_2553 ();
 sg13g2_decap_8 FILLER_41_2560 ();
 sg13g2_decap_8 FILLER_41_2567 ();
 sg13g2_decap_8 FILLER_41_2574 ();
 sg13g2_decap_8 FILLER_41_2581 ();
 sg13g2_decap_8 FILLER_41_2588 ();
 sg13g2_decap_8 FILLER_41_2595 ();
 sg13g2_decap_8 FILLER_41_2602 ();
 sg13g2_decap_8 FILLER_41_2609 ();
 sg13g2_decap_8 FILLER_41_2616 ();
 sg13g2_decap_8 FILLER_41_2623 ();
 sg13g2_decap_8 FILLER_41_2630 ();
 sg13g2_decap_8 FILLER_41_2637 ();
 sg13g2_decap_8 FILLER_41_2644 ();
 sg13g2_decap_8 FILLER_41_2651 ();
 sg13g2_decap_8 FILLER_41_2658 ();
 sg13g2_decap_4 FILLER_41_2665 ();
 sg13g2_fill_1 FILLER_41_2669 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_fill_2 FILLER_42_98 ();
 sg13g2_fill_1 FILLER_42_100 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_fill_1 FILLER_42_112 ();
 sg13g2_fill_2 FILLER_42_116 ();
 sg13g2_decap_8 FILLER_42_122 ();
 sg13g2_decap_8 FILLER_42_129 ();
 sg13g2_decap_8 FILLER_42_136 ();
 sg13g2_decap_8 FILLER_42_143 ();
 sg13g2_decap_8 FILLER_42_150 ();
 sg13g2_decap_8 FILLER_42_157 ();
 sg13g2_decap_8 FILLER_42_164 ();
 sg13g2_decap_8 FILLER_42_171 ();
 sg13g2_fill_1 FILLER_42_178 ();
 sg13g2_decap_4 FILLER_42_182 ();
 sg13g2_decap_8 FILLER_42_190 ();
 sg13g2_decap_8 FILLER_42_197 ();
 sg13g2_decap_8 FILLER_42_204 ();
 sg13g2_decap_8 FILLER_42_211 ();
 sg13g2_decap_8 FILLER_42_218 ();
 sg13g2_decap_8 FILLER_42_225 ();
 sg13g2_decap_8 FILLER_42_232 ();
 sg13g2_decap_8 FILLER_42_239 ();
 sg13g2_decap_8 FILLER_42_246 ();
 sg13g2_decap_8 FILLER_42_253 ();
 sg13g2_decap_4 FILLER_42_260 ();
 sg13g2_fill_1 FILLER_42_264 ();
 sg13g2_decap_8 FILLER_42_275 ();
 sg13g2_decap_8 FILLER_42_282 ();
 sg13g2_decap_8 FILLER_42_289 ();
 sg13g2_decap_8 FILLER_42_296 ();
 sg13g2_decap_8 FILLER_42_303 ();
 sg13g2_decap_8 FILLER_42_310 ();
 sg13g2_decap_8 FILLER_42_317 ();
 sg13g2_decap_8 FILLER_42_328 ();
 sg13g2_decap_8 FILLER_42_335 ();
 sg13g2_decap_8 FILLER_42_342 ();
 sg13g2_decap_8 FILLER_42_349 ();
 sg13g2_decap_8 FILLER_42_356 ();
 sg13g2_decap_8 FILLER_42_363 ();
 sg13g2_decap_8 FILLER_42_370 ();
 sg13g2_decap_8 FILLER_42_377 ();
 sg13g2_decap_8 FILLER_42_384 ();
 sg13g2_decap_8 FILLER_42_391 ();
 sg13g2_decap_8 FILLER_42_398 ();
 sg13g2_decap_8 FILLER_42_405 ();
 sg13g2_decap_8 FILLER_42_412 ();
 sg13g2_decap_8 FILLER_42_419 ();
 sg13g2_decap_8 FILLER_42_426 ();
 sg13g2_decap_8 FILLER_42_433 ();
 sg13g2_decap_8 FILLER_42_440 ();
 sg13g2_fill_1 FILLER_42_447 ();
 sg13g2_decap_8 FILLER_42_453 ();
 sg13g2_decap_8 FILLER_42_460 ();
 sg13g2_decap_8 FILLER_42_467 ();
 sg13g2_decap_8 FILLER_42_474 ();
 sg13g2_fill_2 FILLER_42_481 ();
 sg13g2_fill_1 FILLER_42_483 ();
 sg13g2_fill_1 FILLER_42_489 ();
 sg13g2_decap_8 FILLER_42_495 ();
 sg13g2_decap_4 FILLER_42_502 ();
 sg13g2_fill_1 FILLER_42_506 ();
 sg13g2_decap_8 FILLER_42_516 ();
 sg13g2_decap_8 FILLER_42_523 ();
 sg13g2_decap_8 FILLER_42_530 ();
 sg13g2_decap_8 FILLER_42_537 ();
 sg13g2_decap_8 FILLER_42_544 ();
 sg13g2_decap_8 FILLER_42_551 ();
 sg13g2_decap_8 FILLER_42_558 ();
 sg13g2_decap_8 FILLER_42_565 ();
 sg13g2_decap_8 FILLER_42_572 ();
 sg13g2_decap_8 FILLER_42_579 ();
 sg13g2_decap_8 FILLER_42_586 ();
 sg13g2_fill_1 FILLER_42_617 ();
 sg13g2_fill_2 FILLER_42_633 ();
 sg13g2_decap_8 FILLER_42_638 ();
 sg13g2_decap_8 FILLER_42_645 ();
 sg13g2_decap_8 FILLER_42_652 ();
 sg13g2_decap_8 FILLER_42_659 ();
 sg13g2_decap_8 FILLER_42_666 ();
 sg13g2_decap_8 FILLER_42_673 ();
 sg13g2_decap_8 FILLER_42_680 ();
 sg13g2_decap_8 FILLER_42_687 ();
 sg13g2_decap_8 FILLER_42_694 ();
 sg13g2_decap_8 FILLER_42_701 ();
 sg13g2_decap_4 FILLER_42_708 ();
 sg13g2_fill_1 FILLER_42_712 ();
 sg13g2_decap_8 FILLER_42_722 ();
 sg13g2_decap_4 FILLER_42_729 ();
 sg13g2_fill_2 FILLER_42_733 ();
 sg13g2_decap_8 FILLER_42_739 ();
 sg13g2_decap_8 FILLER_42_761 ();
 sg13g2_decap_8 FILLER_42_768 ();
 sg13g2_decap_8 FILLER_42_775 ();
 sg13g2_decap_8 FILLER_42_782 ();
 sg13g2_decap_8 FILLER_42_789 ();
 sg13g2_fill_1 FILLER_42_796 ();
 sg13g2_fill_1 FILLER_42_801 ();
 sg13g2_decap_8 FILLER_42_840 ();
 sg13g2_decap_8 FILLER_42_847 ();
 sg13g2_decap_8 FILLER_42_854 ();
 sg13g2_decap_8 FILLER_42_861 ();
 sg13g2_decap_8 FILLER_42_868 ();
 sg13g2_decap_8 FILLER_42_875 ();
 sg13g2_decap_8 FILLER_42_882 ();
 sg13g2_fill_2 FILLER_42_889 ();
 sg13g2_fill_1 FILLER_42_891 ();
 sg13g2_decap_8 FILLER_42_900 ();
 sg13g2_decap_8 FILLER_42_907 ();
 sg13g2_decap_8 FILLER_42_914 ();
 sg13g2_decap_8 FILLER_42_921 ();
 sg13g2_decap_4 FILLER_42_928 ();
 sg13g2_fill_1 FILLER_42_932 ();
 sg13g2_decap_8 FILLER_42_938 ();
 sg13g2_decap_8 FILLER_42_945 ();
 sg13g2_fill_2 FILLER_42_952 ();
 sg13g2_decap_8 FILLER_42_958 ();
 sg13g2_decap_8 FILLER_42_965 ();
 sg13g2_decap_8 FILLER_42_972 ();
 sg13g2_decap_8 FILLER_42_979 ();
 sg13g2_decap_8 FILLER_42_986 ();
 sg13g2_decap_8 FILLER_42_1001 ();
 sg13g2_decap_8 FILLER_42_1008 ();
 sg13g2_decap_8 FILLER_42_1015 ();
 sg13g2_decap_8 FILLER_42_1022 ();
 sg13g2_decap_4 FILLER_42_1029 ();
 sg13g2_fill_1 FILLER_42_1033 ();
 sg13g2_decap_8 FILLER_42_1042 ();
 sg13g2_decap_8 FILLER_42_1055 ();
 sg13g2_decap_8 FILLER_42_1062 ();
 sg13g2_decap_4 FILLER_42_1069 ();
 sg13g2_decap_8 FILLER_42_1077 ();
 sg13g2_decap_8 FILLER_42_1084 ();
 sg13g2_decap_8 FILLER_42_1091 ();
 sg13g2_fill_2 FILLER_42_1098 ();
 sg13g2_fill_1 FILLER_42_1100 ();
 sg13g2_decap_8 FILLER_42_1119 ();
 sg13g2_decap_8 FILLER_42_1126 ();
 sg13g2_decap_8 FILLER_42_1133 ();
 sg13g2_decap_8 FILLER_42_1140 ();
 sg13g2_decap_8 FILLER_42_1147 ();
 sg13g2_decap_8 FILLER_42_1154 ();
 sg13g2_decap_8 FILLER_42_1161 ();
 sg13g2_decap_8 FILLER_42_1168 ();
 sg13g2_decap_8 FILLER_42_1175 ();
 sg13g2_decap_8 FILLER_42_1182 ();
 sg13g2_decap_8 FILLER_42_1198 ();
 sg13g2_decap_8 FILLER_42_1205 ();
 sg13g2_decap_8 FILLER_42_1212 ();
 sg13g2_decap_8 FILLER_42_1219 ();
 sg13g2_decap_8 FILLER_42_1226 ();
 sg13g2_decap_8 FILLER_42_1233 ();
 sg13g2_decap_8 FILLER_42_1240 ();
 sg13g2_decap_8 FILLER_42_1247 ();
 sg13g2_decap_8 FILLER_42_1254 ();
 sg13g2_decap_4 FILLER_42_1261 ();
 sg13g2_fill_1 FILLER_42_1265 ();
 sg13g2_decap_4 FILLER_42_1281 ();
 sg13g2_fill_2 FILLER_42_1285 ();
 sg13g2_decap_8 FILLER_42_1291 ();
 sg13g2_decap_8 FILLER_42_1298 ();
 sg13g2_decap_8 FILLER_42_1305 ();
 sg13g2_decap_8 FILLER_42_1312 ();
 sg13g2_decap_4 FILLER_42_1319 ();
 sg13g2_fill_2 FILLER_42_1338 ();
 sg13g2_fill_1 FILLER_42_1343 ();
 sg13g2_decap_4 FILLER_42_1349 ();
 sg13g2_decap_8 FILLER_42_1358 ();
 sg13g2_decap_8 FILLER_42_1365 ();
 sg13g2_decap_8 FILLER_42_1372 ();
 sg13g2_decap_4 FILLER_42_1379 ();
 sg13g2_fill_2 FILLER_42_1383 ();
 sg13g2_decap_8 FILLER_42_1390 ();
 sg13g2_decap_8 FILLER_42_1397 ();
 sg13g2_decap_8 FILLER_42_1404 ();
 sg13g2_decap_4 FILLER_42_1411 ();
 sg13g2_fill_1 FILLER_42_1415 ();
 sg13g2_decap_8 FILLER_42_1421 ();
 sg13g2_decap_8 FILLER_42_1428 ();
 sg13g2_decap_8 FILLER_42_1435 ();
 sg13g2_decap_8 FILLER_42_1442 ();
 sg13g2_decap_8 FILLER_42_1449 ();
 sg13g2_decap_4 FILLER_42_1456 ();
 sg13g2_decap_8 FILLER_42_1465 ();
 sg13g2_decap_8 FILLER_42_1472 ();
 sg13g2_decap_8 FILLER_42_1479 ();
 sg13g2_decap_8 FILLER_42_1486 ();
 sg13g2_fill_2 FILLER_42_1493 ();
 sg13g2_fill_1 FILLER_42_1495 ();
 sg13g2_decap_8 FILLER_42_1500 ();
 sg13g2_decap_8 FILLER_42_1507 ();
 sg13g2_decap_8 FILLER_42_1514 ();
 sg13g2_decap_4 FILLER_42_1521 ();
 sg13g2_fill_2 FILLER_42_1525 ();
 sg13g2_decap_8 FILLER_42_1535 ();
 sg13g2_decap_4 FILLER_42_1542 ();
 sg13g2_decap_4 FILLER_42_1555 ();
 sg13g2_fill_1 FILLER_42_1559 ();
 sg13g2_decap_8 FILLER_42_1563 ();
 sg13g2_decap_4 FILLER_42_1570 ();
 sg13g2_fill_1 FILLER_42_1574 ();
 sg13g2_decap_4 FILLER_42_1579 ();
 sg13g2_fill_2 FILLER_42_1583 ();
 sg13g2_decap_8 FILLER_42_1589 ();
 sg13g2_decap_8 FILLER_42_1596 ();
 sg13g2_decap_8 FILLER_42_1603 ();
 sg13g2_decap_8 FILLER_42_1610 ();
 sg13g2_decap_8 FILLER_42_1617 ();
 sg13g2_decap_8 FILLER_42_1624 ();
 sg13g2_decap_8 FILLER_42_1631 ();
 sg13g2_decap_8 FILLER_42_1638 ();
 sg13g2_decap_8 FILLER_42_1645 ();
 sg13g2_decap_8 FILLER_42_1652 ();
 sg13g2_decap_8 FILLER_42_1668 ();
 sg13g2_decap_8 FILLER_42_1675 ();
 sg13g2_fill_2 FILLER_42_1682 ();
 sg13g2_fill_1 FILLER_42_1684 ();
 sg13g2_decap_8 FILLER_42_1688 ();
 sg13g2_fill_2 FILLER_42_1695 ();
 sg13g2_decap_8 FILLER_42_1706 ();
 sg13g2_decap_8 FILLER_42_1713 ();
 sg13g2_decap_8 FILLER_42_1720 ();
 sg13g2_decap_8 FILLER_42_1727 ();
 sg13g2_decap_8 FILLER_42_1734 ();
 sg13g2_decap_8 FILLER_42_1741 ();
 sg13g2_decap_8 FILLER_42_1748 ();
 sg13g2_decap_8 FILLER_42_1755 ();
 sg13g2_decap_8 FILLER_42_1762 ();
 sg13g2_decap_8 FILLER_42_1769 ();
 sg13g2_fill_2 FILLER_42_1776 ();
 sg13g2_fill_1 FILLER_42_1778 ();
 sg13g2_decap_8 FILLER_42_1792 ();
 sg13g2_decap_8 FILLER_42_1799 ();
 sg13g2_decap_8 FILLER_42_1806 ();
 sg13g2_decap_8 FILLER_42_1813 ();
 sg13g2_decap_8 FILLER_42_1820 ();
 sg13g2_decap_8 FILLER_42_1827 ();
 sg13g2_decap_8 FILLER_42_1834 ();
 sg13g2_decap_8 FILLER_42_1841 ();
 sg13g2_decap_8 FILLER_42_1848 ();
 sg13g2_decap_8 FILLER_42_1855 ();
 sg13g2_decap_8 FILLER_42_1862 ();
 sg13g2_decap_8 FILLER_42_1869 ();
 sg13g2_decap_8 FILLER_42_1876 ();
 sg13g2_decap_8 FILLER_42_1883 ();
 sg13g2_decap_8 FILLER_42_1890 ();
 sg13g2_decap_8 FILLER_42_1897 ();
 sg13g2_decap_8 FILLER_42_1904 ();
 sg13g2_decap_8 FILLER_42_1911 ();
 sg13g2_decap_8 FILLER_42_1918 ();
 sg13g2_decap_8 FILLER_42_1925 ();
 sg13g2_decap_8 FILLER_42_1932 ();
 sg13g2_decap_8 FILLER_42_1939 ();
 sg13g2_decap_8 FILLER_42_1946 ();
 sg13g2_decap_8 FILLER_42_1953 ();
 sg13g2_decap_4 FILLER_42_1960 ();
 sg13g2_fill_1 FILLER_42_1964 ();
 sg13g2_decap_4 FILLER_42_1970 ();
 sg13g2_fill_1 FILLER_42_1974 ();
 sg13g2_decap_8 FILLER_42_1978 ();
 sg13g2_decap_8 FILLER_42_1985 ();
 sg13g2_decap_8 FILLER_42_1992 ();
 sg13g2_decap_8 FILLER_42_1999 ();
 sg13g2_decap_8 FILLER_42_2006 ();
 sg13g2_decap_8 FILLER_42_2013 ();
 sg13g2_decap_8 FILLER_42_2020 ();
 sg13g2_decap_8 FILLER_42_2027 ();
 sg13g2_decap_8 FILLER_42_2034 ();
 sg13g2_decap_8 FILLER_42_2041 ();
 sg13g2_decap_8 FILLER_42_2048 ();
 sg13g2_decap_8 FILLER_42_2055 ();
 sg13g2_decap_8 FILLER_42_2062 ();
 sg13g2_decap_8 FILLER_42_2069 ();
 sg13g2_fill_2 FILLER_42_2076 ();
 sg13g2_fill_1 FILLER_42_2078 ();
 sg13g2_decap_8 FILLER_42_2083 ();
 sg13g2_decap_8 FILLER_42_2090 ();
 sg13g2_decap_8 FILLER_42_2097 ();
 sg13g2_decap_8 FILLER_42_2104 ();
 sg13g2_decap_8 FILLER_42_2111 ();
 sg13g2_decap_8 FILLER_42_2118 ();
 sg13g2_decap_8 FILLER_42_2155 ();
 sg13g2_decap_8 FILLER_42_2162 ();
 sg13g2_decap_8 FILLER_42_2169 ();
 sg13g2_decap_8 FILLER_42_2176 ();
 sg13g2_decap_8 FILLER_42_2183 ();
 sg13g2_decap_8 FILLER_42_2190 ();
 sg13g2_decap_8 FILLER_42_2197 ();
 sg13g2_decap_8 FILLER_42_2204 ();
 sg13g2_decap_8 FILLER_42_2211 ();
 sg13g2_decap_8 FILLER_42_2218 ();
 sg13g2_decap_8 FILLER_42_2225 ();
 sg13g2_decap_8 FILLER_42_2232 ();
 sg13g2_decap_8 FILLER_42_2239 ();
 sg13g2_decap_8 FILLER_42_2246 ();
 sg13g2_decap_8 FILLER_42_2253 ();
 sg13g2_decap_8 FILLER_42_2260 ();
 sg13g2_decap_8 FILLER_42_2267 ();
 sg13g2_decap_8 FILLER_42_2274 ();
 sg13g2_decap_8 FILLER_42_2281 ();
 sg13g2_decap_8 FILLER_42_2288 ();
 sg13g2_decap_8 FILLER_42_2295 ();
 sg13g2_decap_8 FILLER_42_2302 ();
 sg13g2_decap_8 FILLER_42_2309 ();
 sg13g2_decap_8 FILLER_42_2316 ();
 sg13g2_decap_8 FILLER_42_2323 ();
 sg13g2_decap_8 FILLER_42_2330 ();
 sg13g2_decap_8 FILLER_42_2337 ();
 sg13g2_decap_8 FILLER_42_2344 ();
 sg13g2_decap_8 FILLER_42_2351 ();
 sg13g2_decap_8 FILLER_42_2358 ();
 sg13g2_decap_8 FILLER_42_2365 ();
 sg13g2_decap_8 FILLER_42_2372 ();
 sg13g2_decap_8 FILLER_42_2379 ();
 sg13g2_decap_8 FILLER_42_2386 ();
 sg13g2_decap_8 FILLER_42_2393 ();
 sg13g2_decap_8 FILLER_42_2400 ();
 sg13g2_decap_8 FILLER_42_2407 ();
 sg13g2_decap_8 FILLER_42_2414 ();
 sg13g2_decap_8 FILLER_42_2421 ();
 sg13g2_decap_8 FILLER_42_2428 ();
 sg13g2_decap_8 FILLER_42_2435 ();
 sg13g2_decap_8 FILLER_42_2442 ();
 sg13g2_decap_8 FILLER_42_2449 ();
 sg13g2_decap_8 FILLER_42_2456 ();
 sg13g2_decap_8 FILLER_42_2463 ();
 sg13g2_decap_8 FILLER_42_2470 ();
 sg13g2_decap_8 FILLER_42_2477 ();
 sg13g2_decap_8 FILLER_42_2484 ();
 sg13g2_decap_8 FILLER_42_2491 ();
 sg13g2_decap_8 FILLER_42_2498 ();
 sg13g2_decap_8 FILLER_42_2505 ();
 sg13g2_decap_8 FILLER_42_2512 ();
 sg13g2_decap_8 FILLER_42_2519 ();
 sg13g2_decap_8 FILLER_42_2526 ();
 sg13g2_decap_8 FILLER_42_2533 ();
 sg13g2_decap_8 FILLER_42_2540 ();
 sg13g2_decap_8 FILLER_42_2547 ();
 sg13g2_decap_8 FILLER_42_2554 ();
 sg13g2_decap_8 FILLER_42_2561 ();
 sg13g2_decap_8 FILLER_42_2568 ();
 sg13g2_decap_8 FILLER_42_2575 ();
 sg13g2_decap_8 FILLER_42_2582 ();
 sg13g2_decap_8 FILLER_42_2589 ();
 sg13g2_decap_8 FILLER_42_2596 ();
 sg13g2_decap_8 FILLER_42_2603 ();
 sg13g2_decap_8 FILLER_42_2610 ();
 sg13g2_decap_8 FILLER_42_2617 ();
 sg13g2_decap_8 FILLER_42_2624 ();
 sg13g2_decap_8 FILLER_42_2631 ();
 sg13g2_decap_8 FILLER_42_2638 ();
 sg13g2_decap_8 FILLER_42_2645 ();
 sg13g2_decap_8 FILLER_42_2652 ();
 sg13g2_decap_8 FILLER_42_2659 ();
 sg13g2_decap_4 FILLER_42_2666 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_106 ();
 sg13g2_decap_8 FILLER_43_113 ();
 sg13g2_decap_8 FILLER_43_120 ();
 sg13g2_decap_8 FILLER_43_127 ();
 sg13g2_decap_8 FILLER_43_134 ();
 sg13g2_decap_8 FILLER_43_141 ();
 sg13g2_decap_8 FILLER_43_148 ();
 sg13g2_decap_8 FILLER_43_155 ();
 sg13g2_decap_8 FILLER_43_162 ();
 sg13g2_decap_8 FILLER_43_169 ();
 sg13g2_decap_4 FILLER_43_176 ();
 sg13g2_fill_2 FILLER_43_185 ();
 sg13g2_fill_1 FILLER_43_187 ();
 sg13g2_decap_8 FILLER_43_193 ();
 sg13g2_decap_8 FILLER_43_200 ();
 sg13g2_decap_8 FILLER_43_207 ();
 sg13g2_decap_8 FILLER_43_214 ();
 sg13g2_decap_8 FILLER_43_221 ();
 sg13g2_decap_8 FILLER_43_228 ();
 sg13g2_decap_8 FILLER_43_235 ();
 sg13g2_decap_8 FILLER_43_242 ();
 sg13g2_decap_8 FILLER_43_249 ();
 sg13g2_decap_8 FILLER_43_256 ();
 sg13g2_decap_8 FILLER_43_263 ();
 sg13g2_decap_8 FILLER_43_270 ();
 sg13g2_decap_8 FILLER_43_277 ();
 sg13g2_decap_8 FILLER_43_284 ();
 sg13g2_decap_8 FILLER_43_291 ();
 sg13g2_decap_8 FILLER_43_298 ();
 sg13g2_decap_8 FILLER_43_305 ();
 sg13g2_decap_4 FILLER_43_312 ();
 sg13g2_fill_1 FILLER_43_316 ();
 sg13g2_decap_8 FILLER_43_322 ();
 sg13g2_fill_1 FILLER_43_329 ();
 sg13g2_decap_8 FILLER_43_334 ();
 sg13g2_decap_8 FILLER_43_341 ();
 sg13g2_decap_8 FILLER_43_348 ();
 sg13g2_decap_8 FILLER_43_355 ();
 sg13g2_decap_8 FILLER_43_362 ();
 sg13g2_decap_8 FILLER_43_369 ();
 sg13g2_decap_8 FILLER_43_376 ();
 sg13g2_decap_8 FILLER_43_383 ();
 sg13g2_decap_8 FILLER_43_390 ();
 sg13g2_decap_8 FILLER_43_397 ();
 sg13g2_decap_8 FILLER_43_404 ();
 sg13g2_decap_8 FILLER_43_411 ();
 sg13g2_fill_2 FILLER_43_418 ();
 sg13g2_fill_1 FILLER_43_420 ();
 sg13g2_decap_8 FILLER_43_426 ();
 sg13g2_decap_8 FILLER_43_433 ();
 sg13g2_decap_8 FILLER_43_440 ();
 sg13g2_decap_8 FILLER_43_447 ();
 sg13g2_decap_8 FILLER_43_458 ();
 sg13g2_fill_2 FILLER_43_465 ();
 sg13g2_fill_1 FILLER_43_467 ();
 sg13g2_decap_8 FILLER_43_474 ();
 sg13g2_decap_8 FILLER_43_481 ();
 sg13g2_decap_8 FILLER_43_488 ();
 sg13g2_decap_8 FILLER_43_495 ();
 sg13g2_decap_8 FILLER_43_502 ();
 sg13g2_decap_4 FILLER_43_509 ();
 sg13g2_fill_1 FILLER_43_513 ();
 sg13g2_decap_4 FILLER_43_519 ();
 sg13g2_fill_2 FILLER_43_523 ();
 sg13g2_decap_8 FILLER_43_530 ();
 sg13g2_decap_8 FILLER_43_537 ();
 sg13g2_decap_8 FILLER_43_544 ();
 sg13g2_decap_8 FILLER_43_551 ();
 sg13g2_decap_8 FILLER_43_558 ();
 sg13g2_decap_8 FILLER_43_565 ();
 sg13g2_decap_4 FILLER_43_572 ();
 sg13g2_fill_1 FILLER_43_576 ();
 sg13g2_decap_8 FILLER_43_592 ();
 sg13g2_decap_4 FILLER_43_599 ();
 sg13g2_decap_4 FILLER_43_631 ();
 sg13g2_decap_4 FILLER_43_639 ();
 sg13g2_fill_1 FILLER_43_643 ();
 sg13g2_decap_8 FILLER_43_659 ();
 sg13g2_decap_8 FILLER_43_666 ();
 sg13g2_decap_8 FILLER_43_673 ();
 sg13g2_decap_8 FILLER_43_680 ();
 sg13g2_decap_8 FILLER_43_687 ();
 sg13g2_decap_8 FILLER_43_694 ();
 sg13g2_decap_8 FILLER_43_701 ();
 sg13g2_decap_8 FILLER_43_708 ();
 sg13g2_decap_8 FILLER_43_715 ();
 sg13g2_decap_8 FILLER_43_722 ();
 sg13g2_decap_8 FILLER_43_729 ();
 sg13g2_fill_1 FILLER_43_736 ();
 sg13g2_decap_8 FILLER_43_756 ();
 sg13g2_decap_8 FILLER_43_763 ();
 sg13g2_decap_8 FILLER_43_770 ();
 sg13g2_decap_8 FILLER_43_777 ();
 sg13g2_decap_8 FILLER_43_784 ();
 sg13g2_decap_8 FILLER_43_791 ();
 sg13g2_decap_8 FILLER_43_798 ();
 sg13g2_decap_8 FILLER_43_805 ();
 sg13g2_decap_4 FILLER_43_816 ();
 sg13g2_fill_2 FILLER_43_820 ();
 sg13g2_fill_2 FILLER_43_830 ();
 sg13g2_fill_1 FILLER_43_835 ();
 sg13g2_decap_8 FILLER_43_840 ();
 sg13g2_decap_8 FILLER_43_847 ();
 sg13g2_decap_8 FILLER_43_854 ();
 sg13g2_decap_8 FILLER_43_861 ();
 sg13g2_decap_8 FILLER_43_868 ();
 sg13g2_decap_8 FILLER_43_875 ();
 sg13g2_decap_8 FILLER_43_882 ();
 sg13g2_decap_8 FILLER_43_889 ();
 sg13g2_decap_8 FILLER_43_896 ();
 sg13g2_decap_8 FILLER_43_903 ();
 sg13g2_decap_4 FILLER_43_910 ();
 sg13g2_decap_4 FILLER_43_926 ();
 sg13g2_fill_2 FILLER_43_930 ();
 sg13g2_decap_8 FILLER_43_938 ();
 sg13g2_decap_8 FILLER_43_945 ();
 sg13g2_decap_8 FILLER_43_952 ();
 sg13g2_fill_2 FILLER_43_959 ();
 sg13g2_decap_8 FILLER_43_973 ();
 sg13g2_decap_8 FILLER_43_980 ();
 sg13g2_decap_4 FILLER_43_987 ();
 sg13g2_fill_1 FILLER_43_991 ();
 sg13g2_decap_8 FILLER_43_995 ();
 sg13g2_decap_8 FILLER_43_1002 ();
 sg13g2_decap_8 FILLER_43_1009 ();
 sg13g2_decap_8 FILLER_43_1016 ();
 sg13g2_decap_8 FILLER_43_1023 ();
 sg13g2_decap_8 FILLER_43_1030 ();
 sg13g2_decap_8 FILLER_43_1037 ();
 sg13g2_decap_8 FILLER_43_1044 ();
 sg13g2_decap_8 FILLER_43_1051 ();
 sg13g2_decap_8 FILLER_43_1058 ();
 sg13g2_decap_8 FILLER_43_1065 ();
 sg13g2_fill_2 FILLER_43_1072 ();
 sg13g2_decap_8 FILLER_43_1094 ();
 sg13g2_decap_8 FILLER_43_1101 ();
 sg13g2_decap_8 FILLER_43_1108 ();
 sg13g2_decap_8 FILLER_43_1115 ();
 sg13g2_decap_8 FILLER_43_1122 ();
 sg13g2_decap_8 FILLER_43_1129 ();
 sg13g2_decap_8 FILLER_43_1136 ();
 sg13g2_fill_2 FILLER_43_1143 ();
 sg13g2_decap_8 FILLER_43_1151 ();
 sg13g2_decap_8 FILLER_43_1158 ();
 sg13g2_decap_8 FILLER_43_1165 ();
 sg13g2_decap_8 FILLER_43_1172 ();
 sg13g2_decap_8 FILLER_43_1179 ();
 sg13g2_decap_8 FILLER_43_1186 ();
 sg13g2_fill_1 FILLER_43_1193 ();
 sg13g2_decap_8 FILLER_43_1198 ();
 sg13g2_decap_8 FILLER_43_1205 ();
 sg13g2_fill_2 FILLER_43_1212 ();
 sg13g2_fill_1 FILLER_43_1214 ();
 sg13g2_decap_8 FILLER_43_1230 ();
 sg13g2_fill_1 FILLER_43_1237 ();
 sg13g2_decap_8 FILLER_43_1243 ();
 sg13g2_decap_8 FILLER_43_1250 ();
 sg13g2_decap_8 FILLER_43_1257 ();
 sg13g2_decap_4 FILLER_43_1264 ();
 sg13g2_fill_2 FILLER_43_1268 ();
 sg13g2_decap_4 FILLER_43_1273 ();
 sg13g2_fill_1 FILLER_43_1277 ();
 sg13g2_decap_8 FILLER_43_1283 ();
 sg13g2_decap_8 FILLER_43_1290 ();
 sg13g2_decap_8 FILLER_43_1297 ();
 sg13g2_decap_8 FILLER_43_1304 ();
 sg13g2_decap_8 FILLER_43_1311 ();
 sg13g2_decap_4 FILLER_43_1318 ();
 sg13g2_fill_2 FILLER_43_1322 ();
 sg13g2_fill_2 FILLER_43_1332 ();
 sg13g2_fill_1 FILLER_43_1334 ();
 sg13g2_decap_8 FILLER_43_1353 ();
 sg13g2_decap_8 FILLER_43_1360 ();
 sg13g2_decap_8 FILLER_43_1367 ();
 sg13g2_decap_8 FILLER_43_1374 ();
 sg13g2_decap_8 FILLER_43_1381 ();
 sg13g2_decap_8 FILLER_43_1388 ();
 sg13g2_decap_4 FILLER_43_1395 ();
 sg13g2_decap_8 FILLER_43_1414 ();
 sg13g2_decap_8 FILLER_43_1421 ();
 sg13g2_decap_8 FILLER_43_1428 ();
 sg13g2_decap_8 FILLER_43_1435 ();
 sg13g2_fill_2 FILLER_43_1442 ();
 sg13g2_decap_8 FILLER_43_1448 ();
 sg13g2_decap_8 FILLER_43_1455 ();
 sg13g2_decap_8 FILLER_43_1462 ();
 sg13g2_decap_8 FILLER_43_1469 ();
 sg13g2_decap_8 FILLER_43_1476 ();
 sg13g2_decap_8 FILLER_43_1483 ();
 sg13g2_decap_8 FILLER_43_1490 ();
 sg13g2_decap_8 FILLER_43_1497 ();
 sg13g2_decap_8 FILLER_43_1504 ();
 sg13g2_decap_8 FILLER_43_1511 ();
 sg13g2_decap_8 FILLER_43_1518 ();
 sg13g2_decap_4 FILLER_43_1525 ();
 sg13g2_fill_1 FILLER_43_1529 ();
 sg13g2_decap_8 FILLER_43_1534 ();
 sg13g2_decap_8 FILLER_43_1541 ();
 sg13g2_decap_8 FILLER_43_1548 ();
 sg13g2_decap_8 FILLER_43_1555 ();
 sg13g2_decap_8 FILLER_43_1562 ();
 sg13g2_decap_4 FILLER_43_1569 ();
 sg13g2_fill_1 FILLER_43_1573 ();
 sg13g2_decap_8 FILLER_43_1578 ();
 sg13g2_decap_8 FILLER_43_1585 ();
 sg13g2_decap_8 FILLER_43_1592 ();
 sg13g2_decap_8 FILLER_43_1599 ();
 sg13g2_decap_8 FILLER_43_1606 ();
 sg13g2_decap_8 FILLER_43_1613 ();
 sg13g2_decap_8 FILLER_43_1620 ();
 sg13g2_fill_2 FILLER_43_1627 ();
 sg13g2_decap_8 FILLER_43_1644 ();
 sg13g2_decap_8 FILLER_43_1651 ();
 sg13g2_decap_8 FILLER_43_1658 ();
 sg13g2_decap_8 FILLER_43_1665 ();
 sg13g2_decap_8 FILLER_43_1672 ();
 sg13g2_fill_2 FILLER_43_1703 ();
 sg13g2_decap_8 FILLER_43_1719 ();
 sg13g2_decap_8 FILLER_43_1726 ();
 sg13g2_decap_8 FILLER_43_1733 ();
 sg13g2_decap_8 FILLER_43_1740 ();
 sg13g2_decap_8 FILLER_43_1747 ();
 sg13g2_decap_8 FILLER_43_1754 ();
 sg13g2_decap_8 FILLER_43_1761 ();
 sg13g2_decap_8 FILLER_43_1768 ();
 sg13g2_decap_4 FILLER_43_1775 ();
 sg13g2_decap_8 FILLER_43_1787 ();
 sg13g2_decap_8 FILLER_43_1794 ();
 sg13g2_decap_8 FILLER_43_1801 ();
 sg13g2_decap_8 FILLER_43_1808 ();
 sg13g2_decap_8 FILLER_43_1815 ();
 sg13g2_decap_8 FILLER_43_1822 ();
 sg13g2_decap_8 FILLER_43_1829 ();
 sg13g2_decap_8 FILLER_43_1836 ();
 sg13g2_decap_8 FILLER_43_1843 ();
 sg13g2_decap_8 FILLER_43_1850 ();
 sg13g2_decap_8 FILLER_43_1857 ();
 sg13g2_decap_8 FILLER_43_1864 ();
 sg13g2_decap_8 FILLER_43_1871 ();
 sg13g2_decap_8 FILLER_43_1878 ();
 sg13g2_decap_8 FILLER_43_1885 ();
 sg13g2_decap_8 FILLER_43_1892 ();
 sg13g2_decap_8 FILLER_43_1899 ();
 sg13g2_decap_8 FILLER_43_1906 ();
 sg13g2_decap_8 FILLER_43_1913 ();
 sg13g2_decap_8 FILLER_43_1920 ();
 sg13g2_decap_8 FILLER_43_1927 ();
 sg13g2_decap_8 FILLER_43_1934 ();
 sg13g2_decap_8 FILLER_43_1941 ();
 sg13g2_decap_8 FILLER_43_1948 ();
 sg13g2_decap_8 FILLER_43_1955 ();
 sg13g2_decap_8 FILLER_43_1962 ();
 sg13g2_decap_8 FILLER_43_1969 ();
 sg13g2_decap_8 FILLER_43_1976 ();
 sg13g2_decap_8 FILLER_43_1983 ();
 sg13g2_decap_8 FILLER_43_1990 ();
 sg13g2_decap_8 FILLER_43_1997 ();
 sg13g2_decap_8 FILLER_43_2004 ();
 sg13g2_decap_8 FILLER_43_2011 ();
 sg13g2_decap_8 FILLER_43_2018 ();
 sg13g2_decap_8 FILLER_43_2025 ();
 sg13g2_decap_8 FILLER_43_2032 ();
 sg13g2_decap_8 FILLER_43_2039 ();
 sg13g2_decap_8 FILLER_43_2046 ();
 sg13g2_decap_8 FILLER_43_2053 ();
 sg13g2_decap_8 FILLER_43_2060 ();
 sg13g2_decap_8 FILLER_43_2067 ();
 sg13g2_decap_8 FILLER_43_2074 ();
 sg13g2_decap_8 FILLER_43_2081 ();
 sg13g2_decap_8 FILLER_43_2096 ();
 sg13g2_decap_8 FILLER_43_2103 ();
 sg13g2_decap_8 FILLER_43_2110 ();
 sg13g2_decap_8 FILLER_43_2117 ();
 sg13g2_decap_8 FILLER_43_2124 ();
 sg13g2_decap_8 FILLER_43_2131 ();
 sg13g2_decap_8 FILLER_43_2138 ();
 sg13g2_decap_8 FILLER_43_2145 ();
 sg13g2_fill_2 FILLER_43_2152 ();
 sg13g2_decap_8 FILLER_43_2159 ();
 sg13g2_decap_8 FILLER_43_2166 ();
 sg13g2_decap_8 FILLER_43_2173 ();
 sg13g2_decap_8 FILLER_43_2180 ();
 sg13g2_decap_8 FILLER_43_2187 ();
 sg13g2_decap_8 FILLER_43_2194 ();
 sg13g2_decap_8 FILLER_43_2201 ();
 sg13g2_decap_8 FILLER_43_2208 ();
 sg13g2_decap_8 FILLER_43_2215 ();
 sg13g2_decap_8 FILLER_43_2222 ();
 sg13g2_decap_8 FILLER_43_2229 ();
 sg13g2_decap_8 FILLER_43_2236 ();
 sg13g2_decap_8 FILLER_43_2243 ();
 sg13g2_decap_8 FILLER_43_2250 ();
 sg13g2_decap_8 FILLER_43_2257 ();
 sg13g2_decap_8 FILLER_43_2264 ();
 sg13g2_decap_8 FILLER_43_2271 ();
 sg13g2_decap_8 FILLER_43_2278 ();
 sg13g2_decap_8 FILLER_43_2285 ();
 sg13g2_decap_8 FILLER_43_2292 ();
 sg13g2_decap_8 FILLER_43_2299 ();
 sg13g2_decap_8 FILLER_43_2306 ();
 sg13g2_decap_8 FILLER_43_2313 ();
 sg13g2_decap_8 FILLER_43_2320 ();
 sg13g2_decap_8 FILLER_43_2327 ();
 sg13g2_decap_8 FILLER_43_2334 ();
 sg13g2_decap_8 FILLER_43_2341 ();
 sg13g2_decap_8 FILLER_43_2348 ();
 sg13g2_decap_8 FILLER_43_2355 ();
 sg13g2_decap_8 FILLER_43_2362 ();
 sg13g2_decap_8 FILLER_43_2369 ();
 sg13g2_decap_8 FILLER_43_2376 ();
 sg13g2_decap_8 FILLER_43_2383 ();
 sg13g2_decap_8 FILLER_43_2390 ();
 sg13g2_decap_8 FILLER_43_2397 ();
 sg13g2_decap_8 FILLER_43_2404 ();
 sg13g2_decap_8 FILLER_43_2411 ();
 sg13g2_decap_8 FILLER_43_2418 ();
 sg13g2_decap_8 FILLER_43_2425 ();
 sg13g2_decap_8 FILLER_43_2432 ();
 sg13g2_decap_8 FILLER_43_2439 ();
 sg13g2_decap_8 FILLER_43_2446 ();
 sg13g2_decap_8 FILLER_43_2453 ();
 sg13g2_decap_8 FILLER_43_2460 ();
 sg13g2_decap_8 FILLER_43_2467 ();
 sg13g2_decap_8 FILLER_43_2474 ();
 sg13g2_decap_8 FILLER_43_2481 ();
 sg13g2_decap_8 FILLER_43_2488 ();
 sg13g2_decap_8 FILLER_43_2495 ();
 sg13g2_decap_8 FILLER_43_2502 ();
 sg13g2_decap_8 FILLER_43_2509 ();
 sg13g2_decap_8 FILLER_43_2516 ();
 sg13g2_decap_8 FILLER_43_2523 ();
 sg13g2_decap_8 FILLER_43_2530 ();
 sg13g2_decap_8 FILLER_43_2537 ();
 sg13g2_decap_8 FILLER_43_2544 ();
 sg13g2_decap_8 FILLER_43_2551 ();
 sg13g2_decap_8 FILLER_43_2558 ();
 sg13g2_decap_8 FILLER_43_2565 ();
 sg13g2_decap_8 FILLER_43_2572 ();
 sg13g2_decap_8 FILLER_43_2579 ();
 sg13g2_decap_8 FILLER_43_2586 ();
 sg13g2_decap_8 FILLER_43_2593 ();
 sg13g2_decap_8 FILLER_43_2600 ();
 sg13g2_decap_8 FILLER_43_2607 ();
 sg13g2_decap_8 FILLER_43_2614 ();
 sg13g2_decap_8 FILLER_43_2621 ();
 sg13g2_decap_8 FILLER_43_2628 ();
 sg13g2_decap_8 FILLER_43_2635 ();
 sg13g2_decap_8 FILLER_43_2642 ();
 sg13g2_decap_8 FILLER_43_2649 ();
 sg13g2_decap_8 FILLER_43_2656 ();
 sg13g2_decap_8 FILLER_43_2663 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_67 ();
 sg13g2_decap_8 FILLER_44_74 ();
 sg13g2_decap_8 FILLER_44_81 ();
 sg13g2_decap_8 FILLER_44_88 ();
 sg13g2_decap_8 FILLER_44_95 ();
 sg13g2_decap_8 FILLER_44_102 ();
 sg13g2_decap_8 FILLER_44_109 ();
 sg13g2_fill_2 FILLER_44_116 ();
 sg13g2_fill_1 FILLER_44_118 ();
 sg13g2_fill_2 FILLER_44_122 ();
 sg13g2_fill_1 FILLER_44_124 ();
 sg13g2_fill_1 FILLER_44_129 ();
 sg13g2_decap_8 FILLER_44_136 ();
 sg13g2_decap_8 FILLER_44_143 ();
 sg13g2_fill_2 FILLER_44_150 ();
 sg13g2_fill_1 FILLER_44_152 ();
 sg13g2_decap_8 FILLER_44_157 ();
 sg13g2_decap_8 FILLER_44_164 ();
 sg13g2_decap_8 FILLER_44_171 ();
 sg13g2_fill_1 FILLER_44_178 ();
 sg13g2_fill_2 FILLER_44_184 ();
 sg13g2_fill_1 FILLER_44_186 ();
 sg13g2_decap_8 FILLER_44_192 ();
 sg13g2_decap_8 FILLER_44_199 ();
 sg13g2_decap_8 FILLER_44_206 ();
 sg13g2_decap_8 FILLER_44_213 ();
 sg13g2_decap_8 FILLER_44_220 ();
 sg13g2_decap_8 FILLER_44_227 ();
 sg13g2_decap_8 FILLER_44_234 ();
 sg13g2_decap_8 FILLER_44_241 ();
 sg13g2_decap_8 FILLER_44_248 ();
 sg13g2_decap_8 FILLER_44_255 ();
 sg13g2_decap_8 FILLER_44_262 ();
 sg13g2_decap_8 FILLER_44_269 ();
 sg13g2_decap_8 FILLER_44_276 ();
 sg13g2_decap_8 FILLER_44_283 ();
 sg13g2_decap_8 FILLER_44_290 ();
 sg13g2_decap_8 FILLER_44_297 ();
 sg13g2_decap_8 FILLER_44_304 ();
 sg13g2_decap_8 FILLER_44_311 ();
 sg13g2_decap_8 FILLER_44_318 ();
 sg13g2_decap_8 FILLER_44_325 ();
 sg13g2_decap_8 FILLER_44_332 ();
 sg13g2_decap_8 FILLER_44_339 ();
 sg13g2_decap_8 FILLER_44_372 ();
 sg13g2_decap_8 FILLER_44_379 ();
 sg13g2_decap_8 FILLER_44_386 ();
 sg13g2_decap_8 FILLER_44_393 ();
 sg13g2_decap_8 FILLER_44_400 ();
 sg13g2_decap_8 FILLER_44_407 ();
 sg13g2_fill_1 FILLER_44_414 ();
 sg13g2_decap_8 FILLER_44_436 ();
 sg13g2_decap_8 FILLER_44_443 ();
 sg13g2_fill_1 FILLER_44_450 ();
 sg13g2_decap_8 FILLER_44_459 ();
 sg13g2_decap_8 FILLER_44_466 ();
 sg13g2_decap_8 FILLER_44_473 ();
 sg13g2_decap_8 FILLER_44_480 ();
 sg13g2_decap_8 FILLER_44_487 ();
 sg13g2_decap_8 FILLER_44_494 ();
 sg13g2_decap_8 FILLER_44_501 ();
 sg13g2_decap_8 FILLER_44_508 ();
 sg13g2_decap_8 FILLER_44_515 ();
 sg13g2_decap_8 FILLER_44_522 ();
 sg13g2_decap_8 FILLER_44_529 ();
 sg13g2_decap_8 FILLER_44_536 ();
 sg13g2_decap_8 FILLER_44_543 ();
 sg13g2_decap_8 FILLER_44_550 ();
 sg13g2_decap_8 FILLER_44_557 ();
 sg13g2_fill_1 FILLER_44_564 ();
 sg13g2_decap_4 FILLER_44_615 ();
 sg13g2_fill_2 FILLER_44_619 ();
 sg13g2_decap_8 FILLER_44_627 ();
 sg13g2_fill_2 FILLER_44_634 ();
 sg13g2_fill_1 FILLER_44_636 ();
 sg13g2_decap_8 FILLER_44_640 ();
 sg13g2_decap_8 FILLER_44_651 ();
 sg13g2_decap_8 FILLER_44_658 ();
 sg13g2_decap_8 FILLER_44_665 ();
 sg13g2_decap_8 FILLER_44_672 ();
 sg13g2_decap_8 FILLER_44_679 ();
 sg13g2_decap_8 FILLER_44_686 ();
 sg13g2_decap_8 FILLER_44_693 ();
 sg13g2_decap_8 FILLER_44_700 ();
 sg13g2_decap_8 FILLER_44_707 ();
 sg13g2_decap_8 FILLER_44_714 ();
 sg13g2_decap_8 FILLER_44_721 ();
 sg13g2_decap_8 FILLER_44_728 ();
 sg13g2_decap_8 FILLER_44_735 ();
 sg13g2_fill_2 FILLER_44_742 ();
 sg13g2_fill_1 FILLER_44_744 ();
 sg13g2_fill_1 FILLER_44_749 ();
 sg13g2_decap_8 FILLER_44_758 ();
 sg13g2_decap_8 FILLER_44_765 ();
 sg13g2_decap_8 FILLER_44_772 ();
 sg13g2_decap_8 FILLER_44_779 ();
 sg13g2_decap_8 FILLER_44_786 ();
 sg13g2_decap_8 FILLER_44_793 ();
 sg13g2_decap_4 FILLER_44_804 ();
 sg13g2_fill_1 FILLER_44_808 ();
 sg13g2_decap_8 FILLER_44_824 ();
 sg13g2_fill_1 FILLER_44_831 ();
 sg13g2_decap_8 FILLER_44_839 ();
 sg13g2_decap_8 FILLER_44_861 ();
 sg13g2_decap_4 FILLER_44_868 ();
 sg13g2_fill_2 FILLER_44_872 ();
 sg13g2_decap_8 FILLER_44_889 ();
 sg13g2_decap_8 FILLER_44_896 ();
 sg13g2_decap_8 FILLER_44_903 ();
 sg13g2_decap_4 FILLER_44_910 ();
 sg13g2_decap_8 FILLER_44_924 ();
 sg13g2_fill_1 FILLER_44_931 ();
 sg13g2_decap_4 FILLER_44_936 ();
 sg13g2_decap_8 FILLER_44_944 ();
 sg13g2_decap_8 FILLER_44_951 ();
 sg13g2_fill_2 FILLER_44_958 ();
 sg13g2_fill_1 FILLER_44_960 ();
 sg13g2_decap_8 FILLER_44_969 ();
 sg13g2_decap_8 FILLER_44_976 ();
 sg13g2_decap_4 FILLER_44_983 ();
 sg13g2_fill_1 FILLER_44_987 ();
 sg13g2_fill_1 FILLER_44_997 ();
 sg13g2_decap_8 FILLER_44_1002 ();
 sg13g2_decap_8 FILLER_44_1009 ();
 sg13g2_decap_8 FILLER_44_1016 ();
 sg13g2_decap_8 FILLER_44_1023 ();
 sg13g2_decap_8 FILLER_44_1030 ();
 sg13g2_decap_8 FILLER_44_1037 ();
 sg13g2_decap_8 FILLER_44_1044 ();
 sg13g2_decap_8 FILLER_44_1051 ();
 sg13g2_decap_8 FILLER_44_1058 ();
 sg13g2_decap_8 FILLER_44_1065 ();
 sg13g2_decap_8 FILLER_44_1072 ();
 sg13g2_decap_8 FILLER_44_1087 ();
 sg13g2_decap_8 FILLER_44_1094 ();
 sg13g2_decap_8 FILLER_44_1101 ();
 sg13g2_decap_8 FILLER_44_1108 ();
 sg13g2_decap_8 FILLER_44_1115 ();
 sg13g2_decap_8 FILLER_44_1122 ();
 sg13g2_decap_8 FILLER_44_1129 ();
 sg13g2_decap_4 FILLER_44_1136 ();
 sg13g2_fill_1 FILLER_44_1140 ();
 sg13g2_decap_8 FILLER_44_1147 ();
 sg13g2_decap_8 FILLER_44_1158 ();
 sg13g2_decap_8 FILLER_44_1165 ();
 sg13g2_decap_8 FILLER_44_1172 ();
 sg13g2_decap_8 FILLER_44_1179 ();
 sg13g2_decap_8 FILLER_44_1186 ();
 sg13g2_decap_4 FILLER_44_1193 ();
 sg13g2_fill_2 FILLER_44_1209 ();
 sg13g2_fill_1 FILLER_44_1211 ();
 sg13g2_decap_8 FILLER_44_1226 ();
 sg13g2_decap_8 FILLER_44_1233 ();
 sg13g2_decap_8 FILLER_44_1240 ();
 sg13g2_decap_8 FILLER_44_1247 ();
 sg13g2_decap_8 FILLER_44_1254 ();
 sg13g2_decap_4 FILLER_44_1261 ();
 sg13g2_fill_1 FILLER_44_1274 ();
 sg13g2_decap_8 FILLER_44_1279 ();
 sg13g2_decap_8 FILLER_44_1286 ();
 sg13g2_decap_8 FILLER_44_1293 ();
 sg13g2_decap_8 FILLER_44_1300 ();
 sg13g2_decap_8 FILLER_44_1307 ();
 sg13g2_decap_8 FILLER_44_1314 ();
 sg13g2_decap_8 FILLER_44_1321 ();
 sg13g2_decap_4 FILLER_44_1328 ();
 sg13g2_fill_1 FILLER_44_1332 ();
 sg13g2_decap_8 FILLER_44_1356 ();
 sg13g2_decap_8 FILLER_44_1363 ();
 sg13g2_decap_8 FILLER_44_1370 ();
 sg13g2_decap_8 FILLER_44_1377 ();
 sg13g2_decap_8 FILLER_44_1384 ();
 sg13g2_decap_8 FILLER_44_1391 ();
 sg13g2_fill_1 FILLER_44_1398 ();
 sg13g2_decap_8 FILLER_44_1405 ();
 sg13g2_decap_8 FILLER_44_1412 ();
 sg13g2_decap_8 FILLER_44_1419 ();
 sg13g2_decap_8 FILLER_44_1426 ();
 sg13g2_decap_8 FILLER_44_1433 ();
 sg13g2_decap_8 FILLER_44_1440 ();
 sg13g2_decap_8 FILLER_44_1447 ();
 sg13g2_decap_4 FILLER_44_1454 ();
 sg13g2_decap_8 FILLER_44_1463 ();
 sg13g2_fill_1 FILLER_44_1470 ();
 sg13g2_decap_8 FILLER_44_1475 ();
 sg13g2_decap_8 FILLER_44_1482 ();
 sg13g2_decap_8 FILLER_44_1489 ();
 sg13g2_decap_8 FILLER_44_1496 ();
 sg13g2_decap_8 FILLER_44_1503 ();
 sg13g2_decap_8 FILLER_44_1510 ();
 sg13g2_decap_8 FILLER_44_1517 ();
 sg13g2_decap_8 FILLER_44_1524 ();
 sg13g2_decap_4 FILLER_44_1531 ();
 sg13g2_decap_8 FILLER_44_1553 ();
 sg13g2_fill_2 FILLER_44_1560 ();
 sg13g2_decap_8 FILLER_44_1566 ();
 sg13g2_decap_8 FILLER_44_1573 ();
 sg13g2_decap_8 FILLER_44_1580 ();
 sg13g2_decap_8 FILLER_44_1587 ();
 sg13g2_decap_8 FILLER_44_1594 ();
 sg13g2_fill_2 FILLER_44_1601 ();
 sg13g2_fill_1 FILLER_44_1603 ();
 sg13g2_decap_8 FILLER_44_1613 ();
 sg13g2_fill_2 FILLER_44_1620 ();
 sg13g2_fill_1 FILLER_44_1622 ();
 sg13g2_decap_8 FILLER_44_1643 ();
 sg13g2_decap_8 FILLER_44_1650 ();
 sg13g2_decap_8 FILLER_44_1657 ();
 sg13g2_fill_2 FILLER_44_1664 ();
 sg13g2_fill_1 FILLER_44_1666 ();
 sg13g2_decap_8 FILLER_44_1675 ();
 sg13g2_fill_2 FILLER_44_1682 ();
 sg13g2_fill_1 FILLER_44_1684 ();
 sg13g2_decap_8 FILLER_44_1688 ();
 sg13g2_fill_1 FILLER_44_1695 ();
 sg13g2_decap_8 FILLER_44_1707 ();
 sg13g2_decap_8 FILLER_44_1714 ();
 sg13g2_fill_1 FILLER_44_1721 ();
 sg13g2_decap_8 FILLER_44_1728 ();
 sg13g2_decap_8 FILLER_44_1735 ();
 sg13g2_decap_8 FILLER_44_1742 ();
 sg13g2_decap_8 FILLER_44_1749 ();
 sg13g2_decap_8 FILLER_44_1756 ();
 sg13g2_decap_8 FILLER_44_1763 ();
 sg13g2_decap_4 FILLER_44_1770 ();
 sg13g2_fill_2 FILLER_44_1774 ();
 sg13g2_decap_8 FILLER_44_1782 ();
 sg13g2_decap_8 FILLER_44_1789 ();
 sg13g2_decap_8 FILLER_44_1796 ();
 sg13g2_decap_4 FILLER_44_1803 ();
 sg13g2_fill_1 FILLER_44_1807 ();
 sg13g2_decap_8 FILLER_44_1821 ();
 sg13g2_decap_8 FILLER_44_1828 ();
 sg13g2_decap_8 FILLER_44_1835 ();
 sg13g2_decap_8 FILLER_44_1842 ();
 sg13g2_decap_8 FILLER_44_1849 ();
 sg13g2_fill_2 FILLER_44_1856 ();
 sg13g2_decap_8 FILLER_44_1871 ();
 sg13g2_decap_8 FILLER_44_1878 ();
 sg13g2_decap_8 FILLER_44_1885 ();
 sg13g2_fill_1 FILLER_44_1892 ();
 sg13g2_decap_8 FILLER_44_1906 ();
 sg13g2_decap_8 FILLER_44_1913 ();
 sg13g2_decap_8 FILLER_44_1920 ();
 sg13g2_decap_8 FILLER_44_1927 ();
 sg13g2_decap_8 FILLER_44_1934 ();
 sg13g2_decap_8 FILLER_44_1941 ();
 sg13g2_decap_8 FILLER_44_1948 ();
 sg13g2_decap_8 FILLER_44_1955 ();
 sg13g2_decap_8 FILLER_44_1962 ();
 sg13g2_decap_8 FILLER_44_1969 ();
 sg13g2_decap_8 FILLER_44_1976 ();
 sg13g2_decap_8 FILLER_44_1983 ();
 sg13g2_decap_8 FILLER_44_1990 ();
 sg13g2_decap_8 FILLER_44_1997 ();
 sg13g2_fill_2 FILLER_44_2004 ();
 sg13g2_decap_8 FILLER_44_2019 ();
 sg13g2_decap_8 FILLER_44_2026 ();
 sg13g2_decap_8 FILLER_44_2033 ();
 sg13g2_decap_8 FILLER_44_2040 ();
 sg13g2_decap_8 FILLER_44_2047 ();
 sg13g2_decap_8 FILLER_44_2054 ();
 sg13g2_decap_8 FILLER_44_2061 ();
 sg13g2_decap_8 FILLER_44_2068 ();
 sg13g2_decap_8 FILLER_44_2075 ();
 sg13g2_decap_8 FILLER_44_2082 ();
 sg13g2_decap_8 FILLER_44_2089 ();
 sg13g2_decap_8 FILLER_44_2096 ();
 sg13g2_decap_8 FILLER_44_2103 ();
 sg13g2_decap_8 FILLER_44_2110 ();
 sg13g2_decap_8 FILLER_44_2117 ();
 sg13g2_decap_8 FILLER_44_2124 ();
 sg13g2_decap_8 FILLER_44_2131 ();
 sg13g2_decap_8 FILLER_44_2138 ();
 sg13g2_decap_8 FILLER_44_2145 ();
 sg13g2_decap_8 FILLER_44_2152 ();
 sg13g2_fill_1 FILLER_44_2159 ();
 sg13g2_decap_8 FILLER_44_2168 ();
 sg13g2_decap_8 FILLER_44_2175 ();
 sg13g2_decap_8 FILLER_44_2182 ();
 sg13g2_decap_8 FILLER_44_2189 ();
 sg13g2_decap_8 FILLER_44_2196 ();
 sg13g2_decap_8 FILLER_44_2203 ();
 sg13g2_decap_8 FILLER_44_2210 ();
 sg13g2_decap_8 FILLER_44_2217 ();
 sg13g2_decap_8 FILLER_44_2224 ();
 sg13g2_decap_8 FILLER_44_2231 ();
 sg13g2_decap_8 FILLER_44_2238 ();
 sg13g2_decap_8 FILLER_44_2245 ();
 sg13g2_decap_8 FILLER_44_2252 ();
 sg13g2_decap_8 FILLER_44_2259 ();
 sg13g2_decap_8 FILLER_44_2266 ();
 sg13g2_decap_8 FILLER_44_2273 ();
 sg13g2_decap_8 FILLER_44_2280 ();
 sg13g2_decap_8 FILLER_44_2287 ();
 sg13g2_decap_8 FILLER_44_2294 ();
 sg13g2_decap_8 FILLER_44_2301 ();
 sg13g2_decap_8 FILLER_44_2308 ();
 sg13g2_decap_8 FILLER_44_2315 ();
 sg13g2_decap_8 FILLER_44_2322 ();
 sg13g2_decap_8 FILLER_44_2329 ();
 sg13g2_decap_8 FILLER_44_2336 ();
 sg13g2_decap_8 FILLER_44_2343 ();
 sg13g2_decap_8 FILLER_44_2350 ();
 sg13g2_decap_8 FILLER_44_2357 ();
 sg13g2_decap_8 FILLER_44_2364 ();
 sg13g2_decap_8 FILLER_44_2371 ();
 sg13g2_decap_8 FILLER_44_2378 ();
 sg13g2_decap_8 FILLER_44_2385 ();
 sg13g2_decap_8 FILLER_44_2392 ();
 sg13g2_decap_8 FILLER_44_2399 ();
 sg13g2_decap_8 FILLER_44_2406 ();
 sg13g2_decap_8 FILLER_44_2413 ();
 sg13g2_decap_8 FILLER_44_2420 ();
 sg13g2_decap_8 FILLER_44_2427 ();
 sg13g2_decap_8 FILLER_44_2434 ();
 sg13g2_decap_8 FILLER_44_2441 ();
 sg13g2_decap_8 FILLER_44_2448 ();
 sg13g2_decap_8 FILLER_44_2455 ();
 sg13g2_decap_8 FILLER_44_2462 ();
 sg13g2_decap_8 FILLER_44_2469 ();
 sg13g2_decap_8 FILLER_44_2476 ();
 sg13g2_decap_8 FILLER_44_2483 ();
 sg13g2_decap_8 FILLER_44_2490 ();
 sg13g2_decap_8 FILLER_44_2497 ();
 sg13g2_decap_8 FILLER_44_2504 ();
 sg13g2_decap_8 FILLER_44_2511 ();
 sg13g2_decap_8 FILLER_44_2518 ();
 sg13g2_decap_8 FILLER_44_2525 ();
 sg13g2_decap_8 FILLER_44_2532 ();
 sg13g2_decap_8 FILLER_44_2539 ();
 sg13g2_decap_8 FILLER_44_2546 ();
 sg13g2_decap_8 FILLER_44_2553 ();
 sg13g2_decap_8 FILLER_44_2560 ();
 sg13g2_decap_8 FILLER_44_2567 ();
 sg13g2_decap_8 FILLER_44_2574 ();
 sg13g2_decap_8 FILLER_44_2581 ();
 sg13g2_decap_8 FILLER_44_2588 ();
 sg13g2_decap_8 FILLER_44_2595 ();
 sg13g2_decap_8 FILLER_44_2602 ();
 sg13g2_decap_8 FILLER_44_2609 ();
 sg13g2_decap_8 FILLER_44_2616 ();
 sg13g2_decap_8 FILLER_44_2623 ();
 sg13g2_decap_8 FILLER_44_2630 ();
 sg13g2_decap_8 FILLER_44_2637 ();
 sg13g2_decap_8 FILLER_44_2644 ();
 sg13g2_decap_8 FILLER_44_2651 ();
 sg13g2_decap_8 FILLER_44_2658 ();
 sg13g2_decap_4 FILLER_44_2665 ();
 sg13g2_fill_1 FILLER_44_2669 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_4 FILLER_45_70 ();
 sg13g2_fill_1 FILLER_45_74 ();
 sg13g2_decap_8 FILLER_45_86 ();
 sg13g2_decap_8 FILLER_45_93 ();
 sg13g2_decap_8 FILLER_45_100 ();
 sg13g2_decap_8 FILLER_45_107 ();
 sg13g2_decap_8 FILLER_45_114 ();
 sg13g2_decap_8 FILLER_45_121 ();
 sg13g2_decap_8 FILLER_45_128 ();
 sg13g2_decap_8 FILLER_45_135 ();
 sg13g2_decap_8 FILLER_45_142 ();
 sg13g2_decap_8 FILLER_45_149 ();
 sg13g2_decap_8 FILLER_45_156 ();
 sg13g2_decap_8 FILLER_45_163 ();
 sg13g2_decap_8 FILLER_45_170 ();
 sg13g2_decap_8 FILLER_45_177 ();
 sg13g2_decap_8 FILLER_45_184 ();
 sg13g2_decap_8 FILLER_45_191 ();
 sg13g2_decap_8 FILLER_45_198 ();
 sg13g2_decap_8 FILLER_45_205 ();
 sg13g2_decap_8 FILLER_45_212 ();
 sg13g2_decap_8 FILLER_45_219 ();
 sg13g2_decap_8 FILLER_45_226 ();
 sg13g2_decap_8 FILLER_45_233 ();
 sg13g2_fill_2 FILLER_45_240 ();
 sg13g2_fill_1 FILLER_45_242 ();
 sg13g2_decap_8 FILLER_45_247 ();
 sg13g2_decap_8 FILLER_45_254 ();
 sg13g2_decap_8 FILLER_45_261 ();
 sg13g2_decap_8 FILLER_45_268 ();
 sg13g2_decap_8 FILLER_45_275 ();
 sg13g2_decap_8 FILLER_45_282 ();
 sg13g2_decap_8 FILLER_45_289 ();
 sg13g2_decap_8 FILLER_45_296 ();
 sg13g2_decap_8 FILLER_45_303 ();
 sg13g2_decap_8 FILLER_45_310 ();
 sg13g2_decap_8 FILLER_45_317 ();
 sg13g2_decap_8 FILLER_45_324 ();
 sg13g2_decap_8 FILLER_45_331 ();
 sg13g2_decap_8 FILLER_45_338 ();
 sg13g2_decap_4 FILLER_45_345 ();
 sg13g2_fill_2 FILLER_45_349 ();
 sg13g2_decap_8 FILLER_45_355 ();
 sg13g2_decap_8 FILLER_45_362 ();
 sg13g2_decap_8 FILLER_45_369 ();
 sg13g2_decap_8 FILLER_45_376 ();
 sg13g2_decap_8 FILLER_45_383 ();
 sg13g2_decap_8 FILLER_45_390 ();
 sg13g2_decap_8 FILLER_45_397 ();
 sg13g2_decap_8 FILLER_45_404 ();
 sg13g2_decap_8 FILLER_45_411 ();
 sg13g2_decap_4 FILLER_45_418 ();
 sg13g2_fill_2 FILLER_45_422 ();
 sg13g2_fill_2 FILLER_45_428 ();
 sg13g2_decap_8 FILLER_45_438 ();
 sg13g2_decap_8 FILLER_45_445 ();
 sg13g2_decap_8 FILLER_45_452 ();
 sg13g2_decap_8 FILLER_45_459 ();
 sg13g2_decap_8 FILLER_45_471 ();
 sg13g2_decap_8 FILLER_45_478 ();
 sg13g2_decap_8 FILLER_45_485 ();
 sg13g2_decap_8 FILLER_45_492 ();
 sg13g2_decap_8 FILLER_45_499 ();
 sg13g2_decap_8 FILLER_45_506 ();
 sg13g2_decap_4 FILLER_45_513 ();
 sg13g2_fill_2 FILLER_45_517 ();
 sg13g2_decap_8 FILLER_45_524 ();
 sg13g2_fill_2 FILLER_45_531 ();
 sg13g2_fill_1 FILLER_45_533 ();
 sg13g2_decap_8 FILLER_45_539 ();
 sg13g2_decap_8 FILLER_45_546 ();
 sg13g2_decap_8 FILLER_45_553 ();
 sg13g2_decap_8 FILLER_45_560 ();
 sg13g2_decap_8 FILLER_45_567 ();
 sg13g2_decap_8 FILLER_45_585 ();
 sg13g2_decap_8 FILLER_45_592 ();
 sg13g2_decap_8 FILLER_45_599 ();
 sg13g2_decap_4 FILLER_45_606 ();
 sg13g2_fill_2 FILLER_45_610 ();
 sg13g2_fill_2 FILLER_45_635 ();
 sg13g2_fill_1 FILLER_45_646 ();
 sg13g2_decap_8 FILLER_45_653 ();
 sg13g2_fill_1 FILLER_45_660 ();
 sg13g2_decap_8 FILLER_45_665 ();
 sg13g2_decap_8 FILLER_45_672 ();
 sg13g2_decap_8 FILLER_45_679 ();
 sg13g2_decap_8 FILLER_45_686 ();
 sg13g2_decap_8 FILLER_45_693 ();
 sg13g2_decap_8 FILLER_45_700 ();
 sg13g2_fill_2 FILLER_45_707 ();
 sg13g2_fill_1 FILLER_45_709 ();
 sg13g2_fill_1 FILLER_45_726 ();
 sg13g2_decap_8 FILLER_45_735 ();
 sg13g2_decap_8 FILLER_45_742 ();
 sg13g2_decap_8 FILLER_45_749 ();
 sg13g2_fill_2 FILLER_45_756 ();
 sg13g2_decap_8 FILLER_45_762 ();
 sg13g2_decap_8 FILLER_45_769 ();
 sg13g2_decap_8 FILLER_45_776 ();
 sg13g2_decap_8 FILLER_45_783 ();
 sg13g2_decap_8 FILLER_45_790 ();
 sg13g2_decap_8 FILLER_45_797 ();
 sg13g2_decap_8 FILLER_45_804 ();
 sg13g2_fill_1 FILLER_45_811 ();
 sg13g2_decap_8 FILLER_45_818 ();
 sg13g2_decap_8 FILLER_45_825 ();
 sg13g2_decap_8 FILLER_45_832 ();
 sg13g2_decap_4 FILLER_45_839 ();
 sg13g2_fill_1 FILLER_45_854 ();
 sg13g2_fill_2 FILLER_45_874 ();
 sg13g2_fill_1 FILLER_45_876 ();
 sg13g2_decap_8 FILLER_45_882 ();
 sg13g2_decap_8 FILLER_45_889 ();
 sg13g2_decap_8 FILLER_45_896 ();
 sg13g2_decap_8 FILLER_45_903 ();
 sg13g2_decap_8 FILLER_45_910 ();
 sg13g2_decap_8 FILLER_45_917 ();
 sg13g2_decap_8 FILLER_45_924 ();
 sg13g2_decap_8 FILLER_45_937 ();
 sg13g2_decap_8 FILLER_45_944 ();
 sg13g2_decap_8 FILLER_45_951 ();
 sg13g2_decap_8 FILLER_45_958 ();
 sg13g2_decap_8 FILLER_45_965 ();
 sg13g2_decap_8 FILLER_45_972 ();
 sg13g2_decap_8 FILLER_45_979 ();
 sg13g2_decap_4 FILLER_45_986 ();
 sg13g2_fill_2 FILLER_45_990 ();
 sg13g2_decap_8 FILLER_45_995 ();
 sg13g2_decap_8 FILLER_45_1002 ();
 sg13g2_decap_8 FILLER_45_1009 ();
 sg13g2_decap_8 FILLER_45_1016 ();
 sg13g2_decap_8 FILLER_45_1023 ();
 sg13g2_decap_8 FILLER_45_1030 ();
 sg13g2_decap_4 FILLER_45_1037 ();
 sg13g2_fill_1 FILLER_45_1041 ();
 sg13g2_decap_8 FILLER_45_1047 ();
 sg13g2_decap_8 FILLER_45_1054 ();
 sg13g2_decap_8 FILLER_45_1061 ();
 sg13g2_decap_8 FILLER_45_1068 ();
 sg13g2_decap_4 FILLER_45_1075 ();
 sg13g2_decap_8 FILLER_45_1084 ();
 sg13g2_decap_8 FILLER_45_1091 ();
 sg13g2_decap_8 FILLER_45_1098 ();
 sg13g2_decap_8 FILLER_45_1105 ();
 sg13g2_decap_8 FILLER_45_1112 ();
 sg13g2_fill_2 FILLER_45_1119 ();
 sg13g2_fill_1 FILLER_45_1121 ();
 sg13g2_decap_8 FILLER_45_1137 ();
 sg13g2_decap_8 FILLER_45_1144 ();
 sg13g2_decap_8 FILLER_45_1151 ();
 sg13g2_decap_8 FILLER_45_1158 ();
 sg13g2_decap_8 FILLER_45_1165 ();
 sg13g2_decap_8 FILLER_45_1182 ();
 sg13g2_decap_8 FILLER_45_1189 ();
 sg13g2_decap_8 FILLER_45_1196 ();
 sg13g2_decap_8 FILLER_45_1203 ();
 sg13g2_decap_8 FILLER_45_1210 ();
 sg13g2_decap_8 FILLER_45_1217 ();
 sg13g2_decap_8 FILLER_45_1224 ();
 sg13g2_decap_8 FILLER_45_1231 ();
 sg13g2_decap_8 FILLER_45_1238 ();
 sg13g2_decap_8 FILLER_45_1245 ();
 sg13g2_decap_8 FILLER_45_1256 ();
 sg13g2_decap_8 FILLER_45_1263 ();
 sg13g2_decap_8 FILLER_45_1270 ();
 sg13g2_decap_8 FILLER_45_1277 ();
 sg13g2_decap_8 FILLER_45_1284 ();
 sg13g2_decap_8 FILLER_45_1291 ();
 sg13g2_decap_8 FILLER_45_1298 ();
 sg13g2_decap_8 FILLER_45_1305 ();
 sg13g2_decap_8 FILLER_45_1312 ();
 sg13g2_decap_8 FILLER_45_1319 ();
 sg13g2_decap_8 FILLER_45_1326 ();
 sg13g2_decap_8 FILLER_45_1333 ();
 sg13g2_fill_2 FILLER_45_1348 ();
 sg13g2_decap_8 FILLER_45_1355 ();
 sg13g2_decap_8 FILLER_45_1362 ();
 sg13g2_decap_8 FILLER_45_1369 ();
 sg13g2_decap_8 FILLER_45_1376 ();
 sg13g2_decap_8 FILLER_45_1383 ();
 sg13g2_decap_4 FILLER_45_1395 ();
 sg13g2_decap_8 FILLER_45_1403 ();
 sg13g2_decap_8 FILLER_45_1410 ();
 sg13g2_decap_8 FILLER_45_1417 ();
 sg13g2_decap_8 FILLER_45_1424 ();
 sg13g2_decap_8 FILLER_45_1431 ();
 sg13g2_decap_8 FILLER_45_1438 ();
 sg13g2_decap_8 FILLER_45_1445 ();
 sg13g2_fill_2 FILLER_45_1452 ();
 sg13g2_decap_8 FILLER_45_1459 ();
 sg13g2_decap_8 FILLER_45_1466 ();
 sg13g2_decap_8 FILLER_45_1473 ();
 sg13g2_decap_8 FILLER_45_1480 ();
 sg13g2_decap_8 FILLER_45_1487 ();
 sg13g2_decap_8 FILLER_45_1494 ();
 sg13g2_decap_8 FILLER_45_1501 ();
 sg13g2_decap_8 FILLER_45_1508 ();
 sg13g2_decap_8 FILLER_45_1515 ();
 sg13g2_decap_8 FILLER_45_1522 ();
 sg13g2_decap_4 FILLER_45_1529 ();
 sg13g2_fill_2 FILLER_45_1533 ();
 sg13g2_decap_8 FILLER_45_1551 ();
 sg13g2_decap_8 FILLER_45_1558 ();
 sg13g2_decap_8 FILLER_45_1565 ();
 sg13g2_decap_8 FILLER_45_1572 ();
 sg13g2_decap_8 FILLER_45_1579 ();
 sg13g2_decap_8 FILLER_45_1586 ();
 sg13g2_decap_8 FILLER_45_1593 ();
 sg13g2_decap_8 FILLER_45_1600 ();
 sg13g2_decap_8 FILLER_45_1607 ();
 sg13g2_decap_8 FILLER_45_1614 ();
 sg13g2_decap_8 FILLER_45_1621 ();
 sg13g2_fill_1 FILLER_45_1628 ();
 sg13g2_fill_1 FILLER_45_1638 ();
 sg13g2_decap_8 FILLER_45_1643 ();
 sg13g2_decap_8 FILLER_45_1650 ();
 sg13g2_decap_8 FILLER_45_1657 ();
 sg13g2_decap_8 FILLER_45_1664 ();
 sg13g2_decap_8 FILLER_45_1671 ();
 sg13g2_decap_8 FILLER_45_1678 ();
 sg13g2_decap_8 FILLER_45_1685 ();
 sg13g2_decap_8 FILLER_45_1692 ();
 sg13g2_decap_8 FILLER_45_1699 ();
 sg13g2_decap_8 FILLER_45_1706 ();
 sg13g2_decap_8 FILLER_45_1747 ();
 sg13g2_decap_8 FILLER_45_1754 ();
 sg13g2_decap_8 FILLER_45_1761 ();
 sg13g2_decap_8 FILLER_45_1768 ();
 sg13g2_decap_8 FILLER_45_1775 ();
 sg13g2_decap_8 FILLER_45_1782 ();
 sg13g2_decap_8 FILLER_45_1789 ();
 sg13g2_decap_8 FILLER_45_1796 ();
 sg13g2_decap_8 FILLER_45_1803 ();
 sg13g2_decap_8 FILLER_45_1810 ();
 sg13g2_decap_8 FILLER_45_1817 ();
 sg13g2_decap_8 FILLER_45_1824 ();
 sg13g2_decap_8 FILLER_45_1831 ();
 sg13g2_decap_8 FILLER_45_1838 ();
 sg13g2_decap_8 FILLER_45_1845 ();
 sg13g2_decap_8 FILLER_45_1852 ();
 sg13g2_decap_8 FILLER_45_1859 ();
 sg13g2_decap_8 FILLER_45_1866 ();
 sg13g2_decap_8 FILLER_45_1873 ();
 sg13g2_decap_8 FILLER_45_1880 ();
 sg13g2_decap_8 FILLER_45_1887 ();
 sg13g2_decap_8 FILLER_45_1894 ();
 sg13g2_decap_8 FILLER_45_1901 ();
 sg13g2_decap_8 FILLER_45_1908 ();
 sg13g2_decap_8 FILLER_45_1915 ();
 sg13g2_decap_8 FILLER_45_1922 ();
 sg13g2_decap_8 FILLER_45_1929 ();
 sg13g2_decap_8 FILLER_45_1936 ();
 sg13g2_decap_8 FILLER_45_1943 ();
 sg13g2_decap_8 FILLER_45_1950 ();
 sg13g2_decap_8 FILLER_45_1957 ();
 sg13g2_decap_8 FILLER_45_1964 ();
 sg13g2_fill_1 FILLER_45_1971 ();
 sg13g2_decap_8 FILLER_45_1981 ();
 sg13g2_decap_8 FILLER_45_1988 ();
 sg13g2_decap_8 FILLER_45_1995 ();
 sg13g2_decap_8 FILLER_45_2007 ();
 sg13g2_decap_8 FILLER_45_2014 ();
 sg13g2_decap_8 FILLER_45_2021 ();
 sg13g2_decap_8 FILLER_45_2028 ();
 sg13g2_decap_8 FILLER_45_2035 ();
 sg13g2_decap_8 FILLER_45_2042 ();
 sg13g2_decap_8 FILLER_45_2049 ();
 sg13g2_decap_8 FILLER_45_2056 ();
 sg13g2_decap_8 FILLER_45_2063 ();
 sg13g2_decap_8 FILLER_45_2070 ();
 sg13g2_decap_8 FILLER_45_2077 ();
 sg13g2_decap_8 FILLER_45_2084 ();
 sg13g2_decap_8 FILLER_45_2091 ();
 sg13g2_decap_8 FILLER_45_2098 ();
 sg13g2_decap_8 FILLER_45_2105 ();
 sg13g2_decap_8 FILLER_45_2112 ();
 sg13g2_decap_8 FILLER_45_2119 ();
 sg13g2_decap_8 FILLER_45_2126 ();
 sg13g2_decap_8 FILLER_45_2133 ();
 sg13g2_decap_8 FILLER_45_2140 ();
 sg13g2_decap_8 FILLER_45_2147 ();
 sg13g2_decap_8 FILLER_45_2154 ();
 sg13g2_decap_8 FILLER_45_2161 ();
 sg13g2_decap_8 FILLER_45_2168 ();
 sg13g2_decap_8 FILLER_45_2175 ();
 sg13g2_decap_8 FILLER_45_2182 ();
 sg13g2_decap_8 FILLER_45_2189 ();
 sg13g2_decap_8 FILLER_45_2196 ();
 sg13g2_decap_8 FILLER_45_2203 ();
 sg13g2_decap_8 FILLER_45_2210 ();
 sg13g2_decap_8 FILLER_45_2217 ();
 sg13g2_decap_8 FILLER_45_2224 ();
 sg13g2_decap_8 FILLER_45_2231 ();
 sg13g2_decap_8 FILLER_45_2238 ();
 sg13g2_decap_8 FILLER_45_2245 ();
 sg13g2_decap_8 FILLER_45_2252 ();
 sg13g2_decap_8 FILLER_45_2259 ();
 sg13g2_decap_8 FILLER_45_2266 ();
 sg13g2_decap_8 FILLER_45_2273 ();
 sg13g2_decap_8 FILLER_45_2280 ();
 sg13g2_decap_8 FILLER_45_2287 ();
 sg13g2_decap_8 FILLER_45_2294 ();
 sg13g2_decap_8 FILLER_45_2301 ();
 sg13g2_decap_8 FILLER_45_2308 ();
 sg13g2_decap_8 FILLER_45_2315 ();
 sg13g2_decap_8 FILLER_45_2322 ();
 sg13g2_decap_8 FILLER_45_2329 ();
 sg13g2_decap_8 FILLER_45_2336 ();
 sg13g2_decap_8 FILLER_45_2343 ();
 sg13g2_decap_8 FILLER_45_2350 ();
 sg13g2_decap_8 FILLER_45_2357 ();
 sg13g2_decap_8 FILLER_45_2364 ();
 sg13g2_decap_8 FILLER_45_2371 ();
 sg13g2_decap_8 FILLER_45_2378 ();
 sg13g2_decap_8 FILLER_45_2385 ();
 sg13g2_decap_8 FILLER_45_2392 ();
 sg13g2_decap_8 FILLER_45_2399 ();
 sg13g2_decap_8 FILLER_45_2406 ();
 sg13g2_decap_8 FILLER_45_2413 ();
 sg13g2_decap_8 FILLER_45_2420 ();
 sg13g2_decap_8 FILLER_45_2427 ();
 sg13g2_decap_8 FILLER_45_2434 ();
 sg13g2_decap_8 FILLER_45_2441 ();
 sg13g2_decap_8 FILLER_45_2448 ();
 sg13g2_decap_8 FILLER_45_2455 ();
 sg13g2_decap_8 FILLER_45_2462 ();
 sg13g2_decap_8 FILLER_45_2469 ();
 sg13g2_decap_8 FILLER_45_2476 ();
 sg13g2_decap_8 FILLER_45_2483 ();
 sg13g2_decap_8 FILLER_45_2490 ();
 sg13g2_decap_8 FILLER_45_2497 ();
 sg13g2_decap_8 FILLER_45_2504 ();
 sg13g2_decap_8 FILLER_45_2511 ();
 sg13g2_decap_8 FILLER_45_2518 ();
 sg13g2_decap_8 FILLER_45_2525 ();
 sg13g2_decap_8 FILLER_45_2532 ();
 sg13g2_decap_8 FILLER_45_2539 ();
 sg13g2_decap_8 FILLER_45_2546 ();
 sg13g2_decap_8 FILLER_45_2553 ();
 sg13g2_decap_8 FILLER_45_2560 ();
 sg13g2_decap_8 FILLER_45_2567 ();
 sg13g2_decap_8 FILLER_45_2574 ();
 sg13g2_decap_8 FILLER_45_2581 ();
 sg13g2_decap_8 FILLER_45_2588 ();
 sg13g2_decap_8 FILLER_45_2595 ();
 sg13g2_decap_8 FILLER_45_2602 ();
 sg13g2_decap_8 FILLER_45_2609 ();
 sg13g2_decap_8 FILLER_45_2616 ();
 sg13g2_decap_8 FILLER_45_2623 ();
 sg13g2_decap_8 FILLER_45_2630 ();
 sg13g2_decap_8 FILLER_45_2637 ();
 sg13g2_decap_8 FILLER_45_2644 ();
 sg13g2_decap_8 FILLER_45_2651 ();
 sg13g2_decap_8 FILLER_45_2658 ();
 sg13g2_decap_4 FILLER_45_2665 ();
 sg13g2_fill_1 FILLER_45_2669 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_4 FILLER_46_56 ();
 sg13g2_fill_2 FILLER_46_60 ();
 sg13g2_decap_8 FILLER_46_65 ();
 sg13g2_decap_8 FILLER_46_72 ();
 sg13g2_decap_8 FILLER_46_79 ();
 sg13g2_decap_8 FILLER_46_86 ();
 sg13g2_decap_8 FILLER_46_93 ();
 sg13g2_decap_8 FILLER_46_100 ();
 sg13g2_fill_1 FILLER_46_107 ();
 sg13g2_fill_2 FILLER_46_112 ();
 sg13g2_fill_1 FILLER_46_114 ();
 sg13g2_fill_1 FILLER_46_125 ();
 sg13g2_fill_2 FILLER_46_131 ();
 sg13g2_fill_1 FILLER_46_137 ();
 sg13g2_decap_8 FILLER_46_141 ();
 sg13g2_decap_8 FILLER_46_148 ();
 sg13g2_decap_8 FILLER_46_155 ();
 sg13g2_decap_8 FILLER_46_162 ();
 sg13g2_decap_8 FILLER_46_169 ();
 sg13g2_decap_8 FILLER_46_176 ();
 sg13g2_fill_2 FILLER_46_183 ();
 sg13g2_fill_1 FILLER_46_185 ();
 sg13g2_decap_8 FILLER_46_190 ();
 sg13g2_decap_8 FILLER_46_197 ();
 sg13g2_decap_8 FILLER_46_204 ();
 sg13g2_decap_8 FILLER_46_211 ();
 sg13g2_decap_8 FILLER_46_218 ();
 sg13g2_decap_8 FILLER_46_225 ();
 sg13g2_decap_4 FILLER_46_232 ();
 sg13g2_decap_8 FILLER_46_262 ();
 sg13g2_decap_8 FILLER_46_269 ();
 sg13g2_decap_8 FILLER_46_276 ();
 sg13g2_decap_8 FILLER_46_283 ();
 sg13g2_decap_8 FILLER_46_290 ();
 sg13g2_decap_8 FILLER_46_297 ();
 sg13g2_decap_8 FILLER_46_304 ();
 sg13g2_decap_8 FILLER_46_311 ();
 sg13g2_decap_8 FILLER_46_318 ();
 sg13g2_decap_8 FILLER_46_325 ();
 sg13g2_decap_8 FILLER_46_332 ();
 sg13g2_decap_8 FILLER_46_339 ();
 sg13g2_decap_8 FILLER_46_346 ();
 sg13g2_decap_8 FILLER_46_353 ();
 sg13g2_decap_8 FILLER_46_360 ();
 sg13g2_decap_8 FILLER_46_367 ();
 sg13g2_decap_8 FILLER_46_374 ();
 sg13g2_decap_8 FILLER_46_381 ();
 sg13g2_decap_8 FILLER_46_388 ();
 sg13g2_decap_8 FILLER_46_395 ();
 sg13g2_decap_8 FILLER_46_402 ();
 sg13g2_decap_8 FILLER_46_409 ();
 sg13g2_decap_8 FILLER_46_416 ();
 sg13g2_decap_8 FILLER_46_423 ();
 sg13g2_decap_8 FILLER_46_430 ();
 sg13g2_decap_8 FILLER_46_437 ();
 sg13g2_fill_2 FILLER_46_444 ();
 sg13g2_decap_8 FILLER_46_461 ();
 sg13g2_decap_8 FILLER_46_468 ();
 sg13g2_decap_8 FILLER_46_475 ();
 sg13g2_decap_4 FILLER_46_482 ();
 sg13g2_fill_1 FILLER_46_486 ();
 sg13g2_decap_8 FILLER_46_491 ();
 sg13g2_decap_8 FILLER_46_498 ();
 sg13g2_decap_8 FILLER_46_505 ();
 sg13g2_decap_8 FILLER_46_512 ();
 sg13g2_decap_4 FILLER_46_519 ();
 sg13g2_decap_8 FILLER_46_527 ();
 sg13g2_decap_8 FILLER_46_534 ();
 sg13g2_decap_8 FILLER_46_541 ();
 sg13g2_fill_2 FILLER_46_548 ();
 sg13g2_decap_8 FILLER_46_562 ();
 sg13g2_decap_8 FILLER_46_569 ();
 sg13g2_fill_1 FILLER_46_576 ();
 sg13g2_decap_8 FILLER_46_586 ();
 sg13g2_decap_8 FILLER_46_593 ();
 sg13g2_decap_8 FILLER_46_600 ();
 sg13g2_decap_8 FILLER_46_607 ();
 sg13g2_decap_8 FILLER_46_614 ();
 sg13g2_decap_8 FILLER_46_621 ();
 sg13g2_decap_8 FILLER_46_628 ();
 sg13g2_decap_8 FILLER_46_635 ();
 sg13g2_fill_1 FILLER_46_642 ();
 sg13g2_decap_8 FILLER_46_651 ();
 sg13g2_decap_8 FILLER_46_658 ();
 sg13g2_decap_8 FILLER_46_665 ();
 sg13g2_decap_8 FILLER_46_672 ();
 sg13g2_decap_8 FILLER_46_679 ();
 sg13g2_decap_8 FILLER_46_686 ();
 sg13g2_decap_8 FILLER_46_693 ();
 sg13g2_decap_8 FILLER_46_700 ();
 sg13g2_decap_8 FILLER_46_707 ();
 sg13g2_decap_8 FILLER_46_714 ();
 sg13g2_decap_4 FILLER_46_721 ();
 sg13g2_fill_2 FILLER_46_725 ();
 sg13g2_decap_8 FILLER_46_734 ();
 sg13g2_decap_8 FILLER_46_741 ();
 sg13g2_decap_8 FILLER_46_748 ();
 sg13g2_decap_8 FILLER_46_755 ();
 sg13g2_fill_2 FILLER_46_762 ();
 sg13g2_decap_8 FILLER_46_772 ();
 sg13g2_decap_8 FILLER_46_779 ();
 sg13g2_decap_8 FILLER_46_786 ();
 sg13g2_decap_8 FILLER_46_793 ();
 sg13g2_decap_8 FILLER_46_800 ();
 sg13g2_decap_8 FILLER_46_807 ();
 sg13g2_decap_8 FILLER_46_814 ();
 sg13g2_decap_8 FILLER_46_821 ();
 sg13g2_decap_8 FILLER_46_828 ();
 sg13g2_decap_8 FILLER_46_835 ();
 sg13g2_decap_4 FILLER_46_842 ();
 sg13g2_fill_2 FILLER_46_850 ();
 sg13g2_decap_4 FILLER_46_872 ();
 sg13g2_fill_1 FILLER_46_876 ();
 sg13g2_decap_8 FILLER_46_880 ();
 sg13g2_decap_4 FILLER_46_887 ();
 sg13g2_fill_2 FILLER_46_891 ();
 sg13g2_decap_4 FILLER_46_896 ();
 sg13g2_fill_1 FILLER_46_900 ();
 sg13g2_decap_8 FILLER_46_905 ();
 sg13g2_decap_8 FILLER_46_912 ();
 sg13g2_decap_8 FILLER_46_919 ();
 sg13g2_decap_8 FILLER_46_926 ();
 sg13g2_fill_2 FILLER_46_933 ();
 sg13g2_decap_8 FILLER_46_940 ();
 sg13g2_decap_8 FILLER_46_947 ();
 sg13g2_decap_8 FILLER_46_954 ();
 sg13g2_decap_8 FILLER_46_961 ();
 sg13g2_decap_8 FILLER_46_968 ();
 sg13g2_decap_8 FILLER_46_975 ();
 sg13g2_decap_8 FILLER_46_982 ();
 sg13g2_decap_8 FILLER_46_989 ();
 sg13g2_fill_2 FILLER_46_996 ();
 sg13g2_fill_1 FILLER_46_998 ();
 sg13g2_decap_8 FILLER_46_1003 ();
 sg13g2_decap_4 FILLER_46_1010 ();
 sg13g2_decap_8 FILLER_46_1018 ();
 sg13g2_decap_8 FILLER_46_1025 ();
 sg13g2_decap_8 FILLER_46_1032 ();
 sg13g2_decap_4 FILLER_46_1039 ();
 sg13g2_fill_2 FILLER_46_1043 ();
 sg13g2_decap_8 FILLER_46_1065 ();
 sg13g2_decap_8 FILLER_46_1072 ();
 sg13g2_fill_1 FILLER_46_1079 ();
 sg13g2_decap_8 FILLER_46_1084 ();
 sg13g2_decap_8 FILLER_46_1091 ();
 sg13g2_decap_8 FILLER_46_1098 ();
 sg13g2_decap_8 FILLER_46_1105 ();
 sg13g2_decap_8 FILLER_46_1112 ();
 sg13g2_decap_4 FILLER_46_1119 ();
 sg13g2_fill_2 FILLER_46_1123 ();
 sg13g2_decap_8 FILLER_46_1130 ();
 sg13g2_decap_8 FILLER_46_1137 ();
 sg13g2_decap_8 FILLER_46_1144 ();
 sg13g2_decap_8 FILLER_46_1151 ();
 sg13g2_decap_8 FILLER_46_1158 ();
 sg13g2_decap_8 FILLER_46_1165 ();
 sg13g2_decap_8 FILLER_46_1172 ();
 sg13g2_decap_8 FILLER_46_1179 ();
 sg13g2_decap_8 FILLER_46_1186 ();
 sg13g2_decap_8 FILLER_46_1193 ();
 sg13g2_decap_8 FILLER_46_1200 ();
 sg13g2_decap_8 FILLER_46_1207 ();
 sg13g2_decap_8 FILLER_46_1214 ();
 sg13g2_decap_8 FILLER_46_1221 ();
 sg13g2_decap_8 FILLER_46_1228 ();
 sg13g2_decap_8 FILLER_46_1235 ();
 sg13g2_decap_8 FILLER_46_1242 ();
 sg13g2_decap_8 FILLER_46_1254 ();
 sg13g2_decap_8 FILLER_46_1261 ();
 sg13g2_decap_8 FILLER_46_1268 ();
 sg13g2_decap_8 FILLER_46_1275 ();
 sg13g2_fill_2 FILLER_46_1282 ();
 sg13g2_fill_1 FILLER_46_1284 ();
 sg13g2_decap_8 FILLER_46_1289 ();
 sg13g2_decap_8 FILLER_46_1296 ();
 sg13g2_decap_4 FILLER_46_1303 ();
 sg13g2_fill_2 FILLER_46_1307 ();
 sg13g2_decap_8 FILLER_46_1313 ();
 sg13g2_decap_8 FILLER_46_1320 ();
 sg13g2_decap_8 FILLER_46_1327 ();
 sg13g2_decap_4 FILLER_46_1334 ();
 sg13g2_fill_2 FILLER_46_1338 ();
 sg13g2_decap_8 FILLER_46_1345 ();
 sg13g2_decap_8 FILLER_46_1352 ();
 sg13g2_decap_8 FILLER_46_1359 ();
 sg13g2_decap_8 FILLER_46_1372 ();
 sg13g2_decap_8 FILLER_46_1379 ();
 sg13g2_decap_8 FILLER_46_1386 ();
 sg13g2_decap_8 FILLER_46_1393 ();
 sg13g2_decap_8 FILLER_46_1400 ();
 sg13g2_fill_2 FILLER_46_1407 ();
 sg13g2_fill_1 FILLER_46_1409 ();
 sg13g2_decap_8 FILLER_46_1416 ();
 sg13g2_decap_8 FILLER_46_1423 ();
 sg13g2_decap_8 FILLER_46_1430 ();
 sg13g2_fill_2 FILLER_46_1437 ();
 sg13g2_decap_8 FILLER_46_1442 ();
 sg13g2_decap_4 FILLER_46_1449 ();
 sg13g2_decap_8 FILLER_46_1457 ();
 sg13g2_decap_8 FILLER_46_1464 ();
 sg13g2_decap_8 FILLER_46_1471 ();
 sg13g2_decap_4 FILLER_46_1482 ();
 sg13g2_decap_8 FILLER_46_1490 ();
 sg13g2_decap_8 FILLER_46_1497 ();
 sg13g2_decap_8 FILLER_46_1504 ();
 sg13g2_decap_4 FILLER_46_1511 ();
 sg13g2_decap_8 FILLER_46_1525 ();
 sg13g2_decap_8 FILLER_46_1532 ();
 sg13g2_fill_1 FILLER_46_1539 ();
 sg13g2_decap_4 FILLER_46_1543 ();
 sg13g2_fill_2 FILLER_46_1547 ();
 sg13g2_decap_8 FILLER_46_1553 ();
 sg13g2_decap_4 FILLER_46_1560 ();
 sg13g2_fill_1 FILLER_46_1564 ();
 sg13g2_decap_8 FILLER_46_1571 ();
 sg13g2_fill_2 FILLER_46_1578 ();
 sg13g2_decap_8 FILLER_46_1588 ();
 sg13g2_decap_8 FILLER_46_1595 ();
 sg13g2_decap_8 FILLER_46_1602 ();
 sg13g2_decap_8 FILLER_46_1609 ();
 sg13g2_decap_8 FILLER_46_1616 ();
 sg13g2_decap_8 FILLER_46_1623 ();
 sg13g2_decap_8 FILLER_46_1630 ();
 sg13g2_decap_8 FILLER_46_1637 ();
 sg13g2_decap_8 FILLER_46_1644 ();
 sg13g2_decap_8 FILLER_46_1651 ();
 sg13g2_decap_8 FILLER_46_1658 ();
 sg13g2_decap_4 FILLER_46_1665 ();
 sg13g2_fill_2 FILLER_46_1669 ();
 sg13g2_fill_1 FILLER_46_1675 ();
 sg13g2_fill_2 FILLER_46_1685 ();
 sg13g2_decap_8 FILLER_46_1693 ();
 sg13g2_decap_8 FILLER_46_1704 ();
 sg13g2_decap_8 FILLER_46_1711 ();
 sg13g2_decap_4 FILLER_46_1718 ();
 sg13g2_fill_1 FILLER_46_1722 ();
 sg13g2_decap_8 FILLER_46_1736 ();
 sg13g2_decap_8 FILLER_46_1743 ();
 sg13g2_decap_8 FILLER_46_1758 ();
 sg13g2_decap_8 FILLER_46_1765 ();
 sg13g2_decap_8 FILLER_46_1772 ();
 sg13g2_decap_8 FILLER_46_1779 ();
 sg13g2_decap_8 FILLER_46_1786 ();
 sg13g2_decap_8 FILLER_46_1793 ();
 sg13g2_decap_8 FILLER_46_1800 ();
 sg13g2_decap_8 FILLER_46_1807 ();
 sg13g2_decap_8 FILLER_46_1814 ();
 sg13g2_decap_8 FILLER_46_1821 ();
 sg13g2_decap_8 FILLER_46_1828 ();
 sg13g2_decap_8 FILLER_46_1835 ();
 sg13g2_decap_8 FILLER_46_1842 ();
 sg13g2_decap_8 FILLER_46_1849 ();
 sg13g2_decap_8 FILLER_46_1856 ();
 sg13g2_decap_8 FILLER_46_1863 ();
 sg13g2_decap_8 FILLER_46_1870 ();
 sg13g2_decap_8 FILLER_46_1877 ();
 sg13g2_decap_8 FILLER_46_1884 ();
 sg13g2_decap_8 FILLER_46_1891 ();
 sg13g2_decap_8 FILLER_46_1898 ();
 sg13g2_decap_8 FILLER_46_1905 ();
 sg13g2_decap_8 FILLER_46_1912 ();
 sg13g2_decap_8 FILLER_46_1919 ();
 sg13g2_decap_8 FILLER_46_1926 ();
 sg13g2_decap_8 FILLER_46_1933 ();
 sg13g2_decap_8 FILLER_46_1940 ();
 sg13g2_decap_8 FILLER_46_1947 ();
 sg13g2_decap_8 FILLER_46_1954 ();
 sg13g2_decap_8 FILLER_46_1961 ();
 sg13g2_fill_2 FILLER_46_1968 ();
 sg13g2_fill_1 FILLER_46_1970 ();
 sg13g2_decap_8 FILLER_46_1976 ();
 sg13g2_decap_8 FILLER_46_1983 ();
 sg13g2_decap_8 FILLER_46_1990 ();
 sg13g2_fill_2 FILLER_46_1997 ();
 sg13g2_decap_8 FILLER_46_2016 ();
 sg13g2_decap_8 FILLER_46_2023 ();
 sg13g2_decap_8 FILLER_46_2030 ();
 sg13g2_decap_8 FILLER_46_2037 ();
 sg13g2_decap_8 FILLER_46_2044 ();
 sg13g2_decap_8 FILLER_46_2051 ();
 sg13g2_decap_8 FILLER_46_2058 ();
 sg13g2_decap_8 FILLER_46_2065 ();
 sg13g2_decap_8 FILLER_46_2072 ();
 sg13g2_decap_8 FILLER_46_2079 ();
 sg13g2_decap_8 FILLER_46_2086 ();
 sg13g2_decap_8 FILLER_46_2093 ();
 sg13g2_decap_8 FILLER_46_2100 ();
 sg13g2_decap_8 FILLER_46_2107 ();
 sg13g2_decap_8 FILLER_46_2114 ();
 sg13g2_decap_4 FILLER_46_2121 ();
 sg13g2_fill_2 FILLER_46_2125 ();
 sg13g2_decap_8 FILLER_46_2131 ();
 sg13g2_decap_8 FILLER_46_2138 ();
 sg13g2_decap_8 FILLER_46_2145 ();
 sg13g2_decap_8 FILLER_46_2152 ();
 sg13g2_decap_8 FILLER_46_2159 ();
 sg13g2_decap_8 FILLER_46_2166 ();
 sg13g2_decap_8 FILLER_46_2173 ();
 sg13g2_decap_8 FILLER_46_2180 ();
 sg13g2_decap_8 FILLER_46_2187 ();
 sg13g2_decap_4 FILLER_46_2194 ();
 sg13g2_fill_1 FILLER_46_2198 ();
 sg13g2_decap_8 FILLER_46_2203 ();
 sg13g2_decap_8 FILLER_46_2210 ();
 sg13g2_decap_8 FILLER_46_2217 ();
 sg13g2_decap_8 FILLER_46_2224 ();
 sg13g2_decap_8 FILLER_46_2231 ();
 sg13g2_decap_8 FILLER_46_2238 ();
 sg13g2_decap_8 FILLER_46_2245 ();
 sg13g2_decap_8 FILLER_46_2252 ();
 sg13g2_decap_8 FILLER_46_2259 ();
 sg13g2_decap_8 FILLER_46_2266 ();
 sg13g2_decap_8 FILLER_46_2273 ();
 sg13g2_decap_8 FILLER_46_2280 ();
 sg13g2_decap_8 FILLER_46_2287 ();
 sg13g2_decap_8 FILLER_46_2294 ();
 sg13g2_decap_8 FILLER_46_2301 ();
 sg13g2_decap_8 FILLER_46_2308 ();
 sg13g2_decap_8 FILLER_46_2315 ();
 sg13g2_decap_8 FILLER_46_2322 ();
 sg13g2_decap_8 FILLER_46_2329 ();
 sg13g2_decap_8 FILLER_46_2336 ();
 sg13g2_decap_8 FILLER_46_2343 ();
 sg13g2_decap_8 FILLER_46_2350 ();
 sg13g2_decap_8 FILLER_46_2357 ();
 sg13g2_decap_8 FILLER_46_2364 ();
 sg13g2_decap_8 FILLER_46_2371 ();
 sg13g2_decap_8 FILLER_46_2378 ();
 sg13g2_decap_8 FILLER_46_2385 ();
 sg13g2_decap_8 FILLER_46_2392 ();
 sg13g2_decap_8 FILLER_46_2399 ();
 sg13g2_decap_8 FILLER_46_2406 ();
 sg13g2_decap_8 FILLER_46_2413 ();
 sg13g2_decap_8 FILLER_46_2420 ();
 sg13g2_decap_8 FILLER_46_2427 ();
 sg13g2_decap_8 FILLER_46_2434 ();
 sg13g2_decap_8 FILLER_46_2441 ();
 sg13g2_decap_8 FILLER_46_2448 ();
 sg13g2_decap_8 FILLER_46_2455 ();
 sg13g2_decap_8 FILLER_46_2462 ();
 sg13g2_decap_8 FILLER_46_2469 ();
 sg13g2_decap_8 FILLER_46_2476 ();
 sg13g2_decap_8 FILLER_46_2483 ();
 sg13g2_decap_8 FILLER_46_2490 ();
 sg13g2_decap_8 FILLER_46_2497 ();
 sg13g2_decap_8 FILLER_46_2504 ();
 sg13g2_decap_8 FILLER_46_2511 ();
 sg13g2_decap_8 FILLER_46_2518 ();
 sg13g2_decap_8 FILLER_46_2525 ();
 sg13g2_decap_8 FILLER_46_2532 ();
 sg13g2_decap_8 FILLER_46_2539 ();
 sg13g2_decap_8 FILLER_46_2546 ();
 sg13g2_decap_8 FILLER_46_2553 ();
 sg13g2_decap_8 FILLER_46_2560 ();
 sg13g2_decap_8 FILLER_46_2567 ();
 sg13g2_decap_8 FILLER_46_2574 ();
 sg13g2_decap_8 FILLER_46_2581 ();
 sg13g2_decap_8 FILLER_46_2588 ();
 sg13g2_decap_8 FILLER_46_2595 ();
 sg13g2_decap_8 FILLER_46_2602 ();
 sg13g2_decap_8 FILLER_46_2609 ();
 sg13g2_decap_8 FILLER_46_2616 ();
 sg13g2_decap_8 FILLER_46_2623 ();
 sg13g2_decap_8 FILLER_46_2630 ();
 sg13g2_decap_8 FILLER_46_2637 ();
 sg13g2_decap_8 FILLER_46_2644 ();
 sg13g2_decap_8 FILLER_46_2651 ();
 sg13g2_decap_8 FILLER_46_2658 ();
 sg13g2_decap_4 FILLER_46_2665 ();
 sg13g2_fill_1 FILLER_46_2669 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_4 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_120 ();
 sg13g2_decap_8 FILLER_47_127 ();
 sg13g2_decap_8 FILLER_47_134 ();
 sg13g2_fill_1 FILLER_47_141 ();
 sg13g2_decap_8 FILLER_47_147 ();
 sg13g2_decap_8 FILLER_47_154 ();
 sg13g2_decap_8 FILLER_47_161 ();
 sg13g2_decap_8 FILLER_47_168 ();
 sg13g2_decap_4 FILLER_47_175 ();
 sg13g2_fill_1 FILLER_47_179 ();
 sg13g2_decap_8 FILLER_47_189 ();
 sg13g2_decap_8 FILLER_47_196 ();
 sg13g2_decap_8 FILLER_47_203 ();
 sg13g2_decap_8 FILLER_47_210 ();
 sg13g2_decap_8 FILLER_47_217 ();
 sg13g2_decap_8 FILLER_47_224 ();
 sg13g2_decap_8 FILLER_47_231 ();
 sg13g2_decap_8 FILLER_47_238 ();
 sg13g2_decap_8 FILLER_47_245 ();
 sg13g2_decap_8 FILLER_47_252 ();
 sg13g2_decap_8 FILLER_47_259 ();
 sg13g2_decap_8 FILLER_47_266 ();
 sg13g2_decap_8 FILLER_47_273 ();
 sg13g2_decap_8 FILLER_47_280 ();
 sg13g2_decap_8 FILLER_47_287 ();
 sg13g2_decap_8 FILLER_47_294 ();
 sg13g2_decap_8 FILLER_47_301 ();
 sg13g2_decap_8 FILLER_47_308 ();
 sg13g2_decap_8 FILLER_47_315 ();
 sg13g2_decap_8 FILLER_47_322 ();
 sg13g2_decap_8 FILLER_47_329 ();
 sg13g2_decap_8 FILLER_47_336 ();
 sg13g2_decap_8 FILLER_47_343 ();
 sg13g2_decap_8 FILLER_47_350 ();
 sg13g2_decap_8 FILLER_47_357 ();
 sg13g2_decap_8 FILLER_47_364 ();
 sg13g2_decap_8 FILLER_47_371 ();
 sg13g2_decap_8 FILLER_47_378 ();
 sg13g2_decap_8 FILLER_47_398 ();
 sg13g2_decap_8 FILLER_47_405 ();
 sg13g2_decap_8 FILLER_47_412 ();
 sg13g2_decap_8 FILLER_47_424 ();
 sg13g2_decap_8 FILLER_47_431 ();
 sg13g2_decap_4 FILLER_47_438 ();
 sg13g2_fill_1 FILLER_47_442 ();
 sg13g2_fill_2 FILLER_47_447 ();
 sg13g2_decap_8 FILLER_47_454 ();
 sg13g2_fill_2 FILLER_47_461 ();
 sg13g2_fill_1 FILLER_47_463 ();
 sg13g2_decap_8 FILLER_47_468 ();
 sg13g2_decap_4 FILLER_47_475 ();
 sg13g2_fill_2 FILLER_47_479 ();
 sg13g2_decap_4 FILLER_47_485 ();
 sg13g2_fill_1 FILLER_47_489 ();
 sg13g2_decap_8 FILLER_47_499 ();
 sg13g2_decap_8 FILLER_47_506 ();
 sg13g2_decap_8 FILLER_47_513 ();
 sg13g2_decap_8 FILLER_47_520 ();
 sg13g2_decap_8 FILLER_47_527 ();
 sg13g2_decap_8 FILLER_47_534 ();
 sg13g2_decap_8 FILLER_47_541 ();
 sg13g2_fill_2 FILLER_47_548 ();
 sg13g2_decap_4 FILLER_47_554 ();
 sg13g2_decap_8 FILLER_47_563 ();
 sg13g2_decap_4 FILLER_47_570 ();
 sg13g2_fill_1 FILLER_47_574 ();
 sg13g2_fill_2 FILLER_47_578 ();
 sg13g2_decap_8 FILLER_47_587 ();
 sg13g2_fill_2 FILLER_47_594 ();
 sg13g2_fill_1 FILLER_47_596 ();
 sg13g2_decap_8 FILLER_47_602 ();
 sg13g2_decap_8 FILLER_47_609 ();
 sg13g2_decap_8 FILLER_47_616 ();
 sg13g2_fill_1 FILLER_47_623 ();
 sg13g2_decap_8 FILLER_47_629 ();
 sg13g2_decap_8 FILLER_47_636 ();
 sg13g2_decap_8 FILLER_47_643 ();
 sg13g2_decap_8 FILLER_47_650 ();
 sg13g2_decap_4 FILLER_47_657 ();
 sg13g2_fill_1 FILLER_47_661 ();
 sg13g2_decap_8 FILLER_47_678 ();
 sg13g2_decap_4 FILLER_47_685 ();
 sg13g2_fill_2 FILLER_47_689 ();
 sg13g2_decap_8 FILLER_47_697 ();
 sg13g2_decap_8 FILLER_47_704 ();
 sg13g2_decap_8 FILLER_47_711 ();
 sg13g2_decap_8 FILLER_47_718 ();
 sg13g2_decap_8 FILLER_47_725 ();
 sg13g2_decap_8 FILLER_47_732 ();
 sg13g2_decap_8 FILLER_47_739 ();
 sg13g2_decap_8 FILLER_47_746 ();
 sg13g2_decap_8 FILLER_47_753 ();
 sg13g2_decap_8 FILLER_47_760 ();
 sg13g2_decap_8 FILLER_47_767 ();
 sg13g2_decap_8 FILLER_47_774 ();
 sg13g2_decap_4 FILLER_47_781 ();
 sg13g2_fill_1 FILLER_47_785 ();
 sg13g2_decap_8 FILLER_47_801 ();
 sg13g2_decap_8 FILLER_47_808 ();
 sg13g2_decap_8 FILLER_47_815 ();
 sg13g2_decap_8 FILLER_47_822 ();
 sg13g2_decap_8 FILLER_47_833 ();
 sg13g2_decap_8 FILLER_47_840 ();
 sg13g2_decap_8 FILLER_47_847 ();
 sg13g2_decap_8 FILLER_47_854 ();
 sg13g2_decap_8 FILLER_47_861 ();
 sg13g2_decap_8 FILLER_47_868 ();
 sg13g2_decap_8 FILLER_47_875 ();
 sg13g2_decap_8 FILLER_47_882 ();
 sg13g2_decap_8 FILLER_47_889 ();
 sg13g2_decap_8 FILLER_47_896 ();
 sg13g2_decap_8 FILLER_47_903 ();
 sg13g2_decap_8 FILLER_47_910 ();
 sg13g2_decap_8 FILLER_47_917 ();
 sg13g2_decap_8 FILLER_47_924 ();
 sg13g2_decap_8 FILLER_47_931 ();
 sg13g2_decap_8 FILLER_47_938 ();
 sg13g2_decap_8 FILLER_47_945 ();
 sg13g2_decap_8 FILLER_47_952 ();
 sg13g2_decap_8 FILLER_47_959 ();
 sg13g2_decap_8 FILLER_47_966 ();
 sg13g2_decap_8 FILLER_47_973 ();
 sg13g2_decap_8 FILLER_47_980 ();
 sg13g2_decap_8 FILLER_47_987 ();
 sg13g2_decap_4 FILLER_47_994 ();
 sg13g2_fill_1 FILLER_47_998 ();
 sg13g2_decap_8 FILLER_47_1003 ();
 sg13g2_decap_8 FILLER_47_1010 ();
 sg13g2_decap_8 FILLER_47_1017 ();
 sg13g2_decap_8 FILLER_47_1024 ();
 sg13g2_decap_8 FILLER_47_1031 ();
 sg13g2_decap_8 FILLER_47_1038 ();
 sg13g2_decap_8 FILLER_47_1045 ();
 sg13g2_fill_2 FILLER_47_1052 ();
 sg13g2_decap_8 FILLER_47_1066 ();
 sg13g2_decap_4 FILLER_47_1073 ();
 sg13g2_fill_1 FILLER_47_1077 ();
 sg13g2_decap_8 FILLER_47_1082 ();
 sg13g2_decap_8 FILLER_47_1089 ();
 sg13g2_decap_8 FILLER_47_1096 ();
 sg13g2_decap_8 FILLER_47_1103 ();
 sg13g2_decap_8 FILLER_47_1110 ();
 sg13g2_decap_8 FILLER_47_1117 ();
 sg13g2_decap_4 FILLER_47_1124 ();
 sg13g2_fill_1 FILLER_47_1128 ();
 sg13g2_decap_8 FILLER_47_1140 ();
 sg13g2_decap_4 FILLER_47_1147 ();
 sg13g2_fill_1 FILLER_47_1151 ();
 sg13g2_decap_8 FILLER_47_1158 ();
 sg13g2_decap_8 FILLER_47_1165 ();
 sg13g2_decap_8 FILLER_47_1172 ();
 sg13g2_decap_8 FILLER_47_1179 ();
 sg13g2_decap_8 FILLER_47_1186 ();
 sg13g2_decap_8 FILLER_47_1193 ();
 sg13g2_decap_8 FILLER_47_1200 ();
 sg13g2_decap_8 FILLER_47_1207 ();
 sg13g2_decap_8 FILLER_47_1214 ();
 sg13g2_decap_8 FILLER_47_1221 ();
 sg13g2_decap_8 FILLER_47_1228 ();
 sg13g2_decap_8 FILLER_47_1235 ();
 sg13g2_decap_8 FILLER_47_1242 ();
 sg13g2_decap_8 FILLER_47_1253 ();
 sg13g2_decap_8 FILLER_47_1260 ();
 sg13g2_decap_4 FILLER_47_1267 ();
 sg13g2_fill_2 FILLER_47_1271 ();
 sg13g2_decap_8 FILLER_47_1277 ();
 sg13g2_decap_8 FILLER_47_1284 ();
 sg13g2_decap_8 FILLER_47_1291 ();
 sg13g2_decap_8 FILLER_47_1298 ();
 sg13g2_decap_8 FILLER_47_1305 ();
 sg13g2_decap_8 FILLER_47_1312 ();
 sg13g2_decap_8 FILLER_47_1319 ();
 sg13g2_decap_8 FILLER_47_1326 ();
 sg13g2_decap_8 FILLER_47_1333 ();
 sg13g2_decap_8 FILLER_47_1344 ();
 sg13g2_decap_8 FILLER_47_1351 ();
 sg13g2_decap_8 FILLER_47_1358 ();
 sg13g2_decap_8 FILLER_47_1365 ();
 sg13g2_decap_8 FILLER_47_1372 ();
 sg13g2_decap_8 FILLER_47_1379 ();
 sg13g2_decap_8 FILLER_47_1386 ();
 sg13g2_decap_8 FILLER_47_1393 ();
 sg13g2_decap_8 FILLER_47_1400 ();
 sg13g2_decap_8 FILLER_47_1407 ();
 sg13g2_decap_8 FILLER_47_1414 ();
 sg13g2_decap_4 FILLER_47_1421 ();
 sg13g2_fill_2 FILLER_47_1425 ();
 sg13g2_decap_8 FILLER_47_1431 ();
 sg13g2_decap_8 FILLER_47_1438 ();
 sg13g2_decap_8 FILLER_47_1445 ();
 sg13g2_decap_8 FILLER_47_1452 ();
 sg13g2_fill_1 FILLER_47_1459 ();
 sg13g2_decap_8 FILLER_47_1463 ();
 sg13g2_decap_8 FILLER_47_1470 ();
 sg13g2_decap_8 FILLER_47_1477 ();
 sg13g2_decap_8 FILLER_47_1484 ();
 sg13g2_decap_8 FILLER_47_1491 ();
 sg13g2_decap_8 FILLER_47_1498 ();
 sg13g2_decap_8 FILLER_47_1505 ();
 sg13g2_decap_8 FILLER_47_1512 ();
 sg13g2_decap_8 FILLER_47_1519 ();
 sg13g2_decap_8 FILLER_47_1526 ();
 sg13g2_decap_8 FILLER_47_1533 ();
 sg13g2_decap_8 FILLER_47_1540 ();
 sg13g2_decap_4 FILLER_47_1547 ();
 sg13g2_fill_1 FILLER_47_1551 ();
 sg13g2_decap_8 FILLER_47_1556 ();
 sg13g2_decap_4 FILLER_47_1563 ();
 sg13g2_fill_1 FILLER_47_1567 ();
 sg13g2_decap_8 FILLER_47_1583 ();
 sg13g2_decap_8 FILLER_47_1590 ();
 sg13g2_decap_8 FILLER_47_1597 ();
 sg13g2_decap_8 FILLER_47_1604 ();
 sg13g2_decap_8 FILLER_47_1611 ();
 sg13g2_decap_8 FILLER_47_1618 ();
 sg13g2_decap_8 FILLER_47_1625 ();
 sg13g2_decap_8 FILLER_47_1632 ();
 sg13g2_decap_8 FILLER_47_1639 ();
 sg13g2_fill_2 FILLER_47_1646 ();
 sg13g2_decap_4 FILLER_47_1657 ();
 sg13g2_decap_4 FILLER_47_1673 ();
 sg13g2_fill_2 FILLER_47_1677 ();
 sg13g2_decap_8 FILLER_47_1691 ();
 sg13g2_decap_8 FILLER_47_1698 ();
 sg13g2_decap_8 FILLER_47_1705 ();
 sg13g2_decap_8 FILLER_47_1712 ();
 sg13g2_fill_1 FILLER_47_1719 ();
 sg13g2_decap_8 FILLER_47_1724 ();
 sg13g2_decap_8 FILLER_47_1731 ();
 sg13g2_fill_2 FILLER_47_1738 ();
 sg13g2_fill_1 FILLER_47_1740 ();
 sg13g2_fill_2 FILLER_47_1753 ();
 sg13g2_decap_8 FILLER_47_1761 ();
 sg13g2_decap_8 FILLER_47_1768 ();
 sg13g2_decap_8 FILLER_47_1775 ();
 sg13g2_decap_8 FILLER_47_1782 ();
 sg13g2_fill_2 FILLER_47_1789 ();
 sg13g2_decap_8 FILLER_47_1799 ();
 sg13g2_decap_8 FILLER_47_1806 ();
 sg13g2_decap_8 FILLER_47_1813 ();
 sg13g2_decap_8 FILLER_47_1820 ();
 sg13g2_decap_4 FILLER_47_1827 ();
 sg13g2_decap_8 FILLER_47_1844 ();
 sg13g2_decap_8 FILLER_47_1851 ();
 sg13g2_decap_8 FILLER_47_1858 ();
 sg13g2_decap_8 FILLER_47_1865 ();
 sg13g2_decap_8 FILLER_47_1872 ();
 sg13g2_decap_8 FILLER_47_1879 ();
 sg13g2_decap_8 FILLER_47_1886 ();
 sg13g2_decap_8 FILLER_47_1893 ();
 sg13g2_decap_8 FILLER_47_1900 ();
 sg13g2_decap_8 FILLER_47_1907 ();
 sg13g2_decap_8 FILLER_47_1914 ();
 sg13g2_decap_8 FILLER_47_1921 ();
 sg13g2_decap_8 FILLER_47_1928 ();
 sg13g2_decap_8 FILLER_47_1935 ();
 sg13g2_decap_8 FILLER_47_1942 ();
 sg13g2_decap_8 FILLER_47_1949 ();
 sg13g2_decap_8 FILLER_47_1956 ();
 sg13g2_decap_8 FILLER_47_1963 ();
 sg13g2_decap_8 FILLER_47_1970 ();
 sg13g2_fill_1 FILLER_47_1977 ();
 sg13g2_decap_8 FILLER_47_1982 ();
 sg13g2_decap_8 FILLER_47_1989 ();
 sg13g2_decap_4 FILLER_47_1996 ();
 sg13g2_fill_2 FILLER_47_2000 ();
 sg13g2_decap_8 FILLER_47_2007 ();
 sg13g2_decap_8 FILLER_47_2014 ();
 sg13g2_decap_8 FILLER_47_2021 ();
 sg13g2_decap_8 FILLER_47_2028 ();
 sg13g2_decap_8 FILLER_47_2035 ();
 sg13g2_decap_8 FILLER_47_2042 ();
 sg13g2_decap_8 FILLER_47_2049 ();
 sg13g2_decap_8 FILLER_47_2056 ();
 sg13g2_decap_4 FILLER_47_2063 ();
 sg13g2_fill_1 FILLER_47_2067 ();
 sg13g2_decap_8 FILLER_47_2072 ();
 sg13g2_decap_8 FILLER_47_2079 ();
 sg13g2_fill_2 FILLER_47_2086 ();
 sg13g2_fill_1 FILLER_47_2088 ();
 sg13g2_decap_4 FILLER_47_2094 ();
 sg13g2_fill_2 FILLER_47_2098 ();
 sg13g2_decap_8 FILLER_47_2104 ();
 sg13g2_decap_8 FILLER_47_2111 ();
 sg13g2_decap_4 FILLER_47_2118 ();
 sg13g2_fill_2 FILLER_47_2122 ();
 sg13g2_fill_2 FILLER_47_2129 ();
 sg13g2_fill_1 FILLER_47_2131 ();
 sg13g2_decap_8 FILLER_47_2158 ();
 sg13g2_decap_8 FILLER_47_2165 ();
 sg13g2_decap_8 FILLER_47_2172 ();
 sg13g2_decap_4 FILLER_47_2179 ();
 sg13g2_fill_1 FILLER_47_2183 ();
 sg13g2_fill_1 FILLER_47_2193 ();
 sg13g2_decap_8 FILLER_47_2220 ();
 sg13g2_decap_8 FILLER_47_2227 ();
 sg13g2_decap_8 FILLER_47_2234 ();
 sg13g2_decap_8 FILLER_47_2241 ();
 sg13g2_decap_8 FILLER_47_2248 ();
 sg13g2_decap_8 FILLER_47_2255 ();
 sg13g2_decap_8 FILLER_47_2262 ();
 sg13g2_decap_8 FILLER_47_2269 ();
 sg13g2_decap_8 FILLER_47_2276 ();
 sg13g2_decap_8 FILLER_47_2283 ();
 sg13g2_decap_8 FILLER_47_2290 ();
 sg13g2_decap_8 FILLER_47_2297 ();
 sg13g2_decap_8 FILLER_47_2304 ();
 sg13g2_decap_8 FILLER_47_2311 ();
 sg13g2_decap_8 FILLER_47_2318 ();
 sg13g2_decap_8 FILLER_47_2325 ();
 sg13g2_decap_8 FILLER_47_2332 ();
 sg13g2_decap_8 FILLER_47_2339 ();
 sg13g2_decap_8 FILLER_47_2346 ();
 sg13g2_decap_8 FILLER_47_2353 ();
 sg13g2_decap_8 FILLER_47_2360 ();
 sg13g2_decap_8 FILLER_47_2367 ();
 sg13g2_decap_8 FILLER_47_2374 ();
 sg13g2_decap_8 FILLER_47_2381 ();
 sg13g2_decap_8 FILLER_47_2388 ();
 sg13g2_decap_8 FILLER_47_2395 ();
 sg13g2_decap_8 FILLER_47_2402 ();
 sg13g2_decap_8 FILLER_47_2409 ();
 sg13g2_decap_8 FILLER_47_2416 ();
 sg13g2_decap_8 FILLER_47_2423 ();
 sg13g2_decap_8 FILLER_47_2430 ();
 sg13g2_decap_8 FILLER_47_2437 ();
 sg13g2_decap_8 FILLER_47_2444 ();
 sg13g2_decap_8 FILLER_47_2451 ();
 sg13g2_decap_8 FILLER_47_2458 ();
 sg13g2_decap_8 FILLER_47_2465 ();
 sg13g2_decap_8 FILLER_47_2472 ();
 sg13g2_decap_8 FILLER_47_2479 ();
 sg13g2_decap_8 FILLER_47_2486 ();
 sg13g2_decap_8 FILLER_47_2493 ();
 sg13g2_decap_8 FILLER_47_2500 ();
 sg13g2_decap_8 FILLER_47_2507 ();
 sg13g2_decap_8 FILLER_47_2514 ();
 sg13g2_decap_8 FILLER_47_2521 ();
 sg13g2_decap_8 FILLER_47_2528 ();
 sg13g2_decap_8 FILLER_47_2535 ();
 sg13g2_decap_8 FILLER_47_2542 ();
 sg13g2_decap_8 FILLER_47_2549 ();
 sg13g2_decap_8 FILLER_47_2556 ();
 sg13g2_decap_8 FILLER_47_2563 ();
 sg13g2_decap_8 FILLER_47_2570 ();
 sg13g2_decap_8 FILLER_47_2577 ();
 sg13g2_decap_8 FILLER_47_2584 ();
 sg13g2_decap_8 FILLER_47_2591 ();
 sg13g2_decap_8 FILLER_47_2598 ();
 sg13g2_decap_8 FILLER_47_2605 ();
 sg13g2_decap_8 FILLER_47_2612 ();
 sg13g2_decap_8 FILLER_47_2619 ();
 sg13g2_decap_8 FILLER_47_2626 ();
 sg13g2_decap_8 FILLER_47_2633 ();
 sg13g2_decap_8 FILLER_47_2640 ();
 sg13g2_decap_8 FILLER_47_2647 ();
 sg13g2_decap_8 FILLER_47_2654 ();
 sg13g2_decap_8 FILLER_47_2661 ();
 sg13g2_fill_2 FILLER_47_2668 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_4 FILLER_48_56 ();
 sg13g2_fill_1 FILLER_48_60 ();
 sg13g2_decap_8 FILLER_48_67 ();
 sg13g2_decap_4 FILLER_48_74 ();
 sg13g2_fill_2 FILLER_48_78 ();
 sg13g2_decap_4 FILLER_48_83 ();
 sg13g2_fill_1 FILLER_48_87 ();
 sg13g2_decap_8 FILLER_48_93 ();
 sg13g2_decap_4 FILLER_48_100 ();
 sg13g2_fill_2 FILLER_48_104 ();
 sg13g2_decap_8 FILLER_48_111 ();
 sg13g2_decap_8 FILLER_48_118 ();
 sg13g2_decap_8 FILLER_48_125 ();
 sg13g2_decap_4 FILLER_48_132 ();
 sg13g2_decap_8 FILLER_48_139 ();
 sg13g2_decap_8 FILLER_48_146 ();
 sg13g2_decap_8 FILLER_48_153 ();
 sg13g2_decap_8 FILLER_48_160 ();
 sg13g2_decap_8 FILLER_48_167 ();
 sg13g2_decap_8 FILLER_48_174 ();
 sg13g2_fill_1 FILLER_48_181 ();
 sg13g2_fill_2 FILLER_48_187 ();
 sg13g2_decap_8 FILLER_48_194 ();
 sg13g2_decap_8 FILLER_48_201 ();
 sg13g2_decap_8 FILLER_48_208 ();
 sg13g2_decap_8 FILLER_48_215 ();
 sg13g2_decap_8 FILLER_48_222 ();
 sg13g2_decap_8 FILLER_48_229 ();
 sg13g2_decap_8 FILLER_48_236 ();
 sg13g2_decap_8 FILLER_48_243 ();
 sg13g2_decap_8 FILLER_48_250 ();
 sg13g2_decap_8 FILLER_48_257 ();
 sg13g2_decap_8 FILLER_48_264 ();
 sg13g2_decap_8 FILLER_48_271 ();
 sg13g2_fill_1 FILLER_48_278 ();
 sg13g2_decap_8 FILLER_48_305 ();
 sg13g2_decap_8 FILLER_48_312 ();
 sg13g2_decap_8 FILLER_48_319 ();
 sg13g2_decap_8 FILLER_48_326 ();
 sg13g2_decap_8 FILLER_48_333 ();
 sg13g2_decap_8 FILLER_48_340 ();
 sg13g2_decap_8 FILLER_48_347 ();
 sg13g2_decap_8 FILLER_48_354 ();
 sg13g2_decap_8 FILLER_48_361 ();
 sg13g2_decap_8 FILLER_48_368 ();
 sg13g2_decap_8 FILLER_48_375 ();
 sg13g2_decap_8 FILLER_48_382 ();
 sg13g2_decap_8 FILLER_48_389 ();
 sg13g2_decap_8 FILLER_48_396 ();
 sg13g2_decap_8 FILLER_48_403 ();
 sg13g2_decap_8 FILLER_48_410 ();
 sg13g2_decap_8 FILLER_48_417 ();
 sg13g2_decap_8 FILLER_48_424 ();
 sg13g2_decap_8 FILLER_48_431 ();
 sg13g2_fill_2 FILLER_48_438 ();
 sg13g2_fill_1 FILLER_48_440 ();
 sg13g2_fill_2 FILLER_48_446 ();
 sg13g2_fill_1 FILLER_48_448 ();
 sg13g2_decap_8 FILLER_48_455 ();
 sg13g2_decap_8 FILLER_48_462 ();
 sg13g2_decap_8 FILLER_48_469 ();
 sg13g2_decap_8 FILLER_48_476 ();
 sg13g2_decap_8 FILLER_48_483 ();
 sg13g2_decap_8 FILLER_48_490 ();
 sg13g2_decap_8 FILLER_48_497 ();
 sg13g2_decap_8 FILLER_48_504 ();
 sg13g2_decap_8 FILLER_48_511 ();
 sg13g2_decap_8 FILLER_48_518 ();
 sg13g2_decap_8 FILLER_48_525 ();
 sg13g2_decap_8 FILLER_48_532 ();
 sg13g2_decap_8 FILLER_48_539 ();
 sg13g2_decap_8 FILLER_48_546 ();
 sg13g2_decap_8 FILLER_48_553 ();
 sg13g2_decap_4 FILLER_48_560 ();
 sg13g2_fill_2 FILLER_48_564 ();
 sg13g2_decap_4 FILLER_48_583 ();
 sg13g2_fill_2 FILLER_48_587 ();
 sg13g2_decap_8 FILLER_48_604 ();
 sg13g2_decap_8 FILLER_48_611 ();
 sg13g2_decap_8 FILLER_48_618 ();
 sg13g2_decap_8 FILLER_48_625 ();
 sg13g2_decap_8 FILLER_48_632 ();
 sg13g2_decap_8 FILLER_48_639 ();
 sg13g2_decap_8 FILLER_48_646 ();
 sg13g2_decap_8 FILLER_48_653 ();
 sg13g2_decap_4 FILLER_48_660 ();
 sg13g2_fill_1 FILLER_48_664 ();
 sg13g2_decap_8 FILLER_48_680 ();
 sg13g2_decap_4 FILLER_48_687 ();
 sg13g2_fill_1 FILLER_48_691 ();
 sg13g2_decap_8 FILLER_48_695 ();
 sg13g2_decap_8 FILLER_48_702 ();
 sg13g2_decap_4 FILLER_48_709 ();
 sg13g2_fill_2 FILLER_48_713 ();
 sg13g2_decap_8 FILLER_48_718 ();
 sg13g2_decap_8 FILLER_48_725 ();
 sg13g2_decap_8 FILLER_48_732 ();
 sg13g2_decap_8 FILLER_48_739 ();
 sg13g2_decap_8 FILLER_48_746 ();
 sg13g2_decap_8 FILLER_48_753 ();
 sg13g2_decap_8 FILLER_48_760 ();
 sg13g2_decap_8 FILLER_48_767 ();
 sg13g2_decap_8 FILLER_48_774 ();
 sg13g2_decap_8 FILLER_48_781 ();
 sg13g2_fill_1 FILLER_48_788 ();
 sg13g2_decap_8 FILLER_48_794 ();
 sg13g2_decap_8 FILLER_48_801 ();
 sg13g2_decap_8 FILLER_48_808 ();
 sg13g2_decap_8 FILLER_48_815 ();
 sg13g2_decap_8 FILLER_48_822 ();
 sg13g2_decap_8 FILLER_48_829 ();
 sg13g2_decap_8 FILLER_48_836 ();
 sg13g2_decap_8 FILLER_48_843 ();
 sg13g2_decap_8 FILLER_48_850 ();
 sg13g2_decap_4 FILLER_48_857 ();
 sg13g2_fill_2 FILLER_48_861 ();
 sg13g2_fill_1 FILLER_48_866 ();
 sg13g2_fill_2 FILLER_48_870 ();
 sg13g2_decap_8 FILLER_48_881 ();
 sg13g2_decap_8 FILLER_48_888 ();
 sg13g2_decap_8 FILLER_48_895 ();
 sg13g2_decap_8 FILLER_48_902 ();
 sg13g2_decap_8 FILLER_48_909 ();
 sg13g2_decap_4 FILLER_48_916 ();
 sg13g2_fill_2 FILLER_48_920 ();
 sg13g2_decap_4 FILLER_48_925 ();
 sg13g2_fill_1 FILLER_48_929 ();
 sg13g2_decap_8 FILLER_48_942 ();
 sg13g2_decap_8 FILLER_48_949 ();
 sg13g2_fill_2 FILLER_48_956 ();
 sg13g2_decap_8 FILLER_48_961 ();
 sg13g2_decap_8 FILLER_48_968 ();
 sg13g2_decap_8 FILLER_48_975 ();
 sg13g2_decap_8 FILLER_48_982 ();
 sg13g2_decap_8 FILLER_48_989 ();
 sg13g2_decap_4 FILLER_48_996 ();
 sg13g2_fill_2 FILLER_48_1011 ();
 sg13g2_decap_8 FILLER_48_1017 ();
 sg13g2_decap_8 FILLER_48_1024 ();
 sg13g2_decap_8 FILLER_48_1031 ();
 sg13g2_decap_4 FILLER_48_1038 ();
 sg13g2_fill_2 FILLER_48_1057 ();
 sg13g2_decap_8 FILLER_48_1064 ();
 sg13g2_decap_8 FILLER_48_1071 ();
 sg13g2_decap_8 FILLER_48_1078 ();
 sg13g2_decap_8 FILLER_48_1085 ();
 sg13g2_decap_8 FILLER_48_1092 ();
 sg13g2_decap_8 FILLER_48_1099 ();
 sg13g2_decap_8 FILLER_48_1106 ();
 sg13g2_decap_8 FILLER_48_1113 ();
 sg13g2_fill_2 FILLER_48_1120 ();
 sg13g2_decap_8 FILLER_48_1128 ();
 sg13g2_decap_8 FILLER_48_1135 ();
 sg13g2_decap_8 FILLER_48_1142 ();
 sg13g2_decap_8 FILLER_48_1149 ();
 sg13g2_decap_8 FILLER_48_1156 ();
 sg13g2_decap_8 FILLER_48_1163 ();
 sg13g2_fill_2 FILLER_48_1170 ();
 sg13g2_fill_1 FILLER_48_1172 ();
 sg13g2_decap_8 FILLER_48_1176 ();
 sg13g2_decap_8 FILLER_48_1183 ();
 sg13g2_decap_8 FILLER_48_1190 ();
 sg13g2_decap_8 FILLER_48_1197 ();
 sg13g2_decap_8 FILLER_48_1204 ();
 sg13g2_decap_8 FILLER_48_1211 ();
 sg13g2_decap_8 FILLER_48_1218 ();
 sg13g2_decap_8 FILLER_48_1225 ();
 sg13g2_decap_8 FILLER_48_1232 ();
 sg13g2_decap_8 FILLER_48_1239 ();
 sg13g2_decap_8 FILLER_48_1246 ();
 sg13g2_decap_8 FILLER_48_1253 ();
 sg13g2_decap_8 FILLER_48_1260 ();
 sg13g2_decap_8 FILLER_48_1267 ();
 sg13g2_decap_8 FILLER_48_1274 ();
 sg13g2_decap_8 FILLER_48_1281 ();
 sg13g2_decap_8 FILLER_48_1288 ();
 sg13g2_decap_8 FILLER_48_1295 ();
 sg13g2_decap_8 FILLER_48_1302 ();
 sg13g2_decap_8 FILLER_48_1309 ();
 sg13g2_decap_8 FILLER_48_1316 ();
 sg13g2_decap_8 FILLER_48_1323 ();
 sg13g2_decap_8 FILLER_48_1330 ();
 sg13g2_decap_8 FILLER_48_1337 ();
 sg13g2_decap_8 FILLER_48_1344 ();
 sg13g2_decap_8 FILLER_48_1351 ();
 sg13g2_decap_8 FILLER_48_1358 ();
 sg13g2_decap_8 FILLER_48_1365 ();
 sg13g2_decap_8 FILLER_48_1372 ();
 sg13g2_fill_1 FILLER_48_1379 ();
 sg13g2_decap_8 FILLER_48_1392 ();
 sg13g2_decap_8 FILLER_48_1399 ();
 sg13g2_decap_8 FILLER_48_1406 ();
 sg13g2_fill_1 FILLER_48_1413 ();
 sg13g2_decap_8 FILLER_48_1419 ();
 sg13g2_decap_4 FILLER_48_1426 ();
 sg13g2_fill_2 FILLER_48_1430 ();
 sg13g2_decap_8 FILLER_48_1436 ();
 sg13g2_decap_8 FILLER_48_1443 ();
 sg13g2_decap_8 FILLER_48_1450 ();
 sg13g2_fill_2 FILLER_48_1457 ();
 sg13g2_fill_1 FILLER_48_1459 ();
 sg13g2_decap_8 FILLER_48_1475 ();
 sg13g2_decap_8 FILLER_48_1482 ();
 sg13g2_decap_8 FILLER_48_1489 ();
 sg13g2_decap_8 FILLER_48_1496 ();
 sg13g2_decap_8 FILLER_48_1503 ();
 sg13g2_decap_8 FILLER_48_1510 ();
 sg13g2_decap_8 FILLER_48_1517 ();
 sg13g2_fill_2 FILLER_48_1524 ();
 sg13g2_fill_1 FILLER_48_1526 ();
 sg13g2_fill_2 FILLER_48_1542 ();
 sg13g2_decap_8 FILLER_48_1550 ();
 sg13g2_decap_8 FILLER_48_1557 ();
 sg13g2_decap_4 FILLER_48_1564 ();
 sg13g2_fill_2 FILLER_48_1574 ();
 sg13g2_decap_8 FILLER_48_1584 ();
 sg13g2_decap_8 FILLER_48_1591 ();
 sg13g2_decap_8 FILLER_48_1598 ();
 sg13g2_decap_8 FILLER_48_1605 ();
 sg13g2_decap_8 FILLER_48_1612 ();
 sg13g2_fill_2 FILLER_48_1619 ();
 sg13g2_fill_1 FILLER_48_1621 ();
 sg13g2_decap_8 FILLER_48_1625 ();
 sg13g2_decap_8 FILLER_48_1632 ();
 sg13g2_decap_8 FILLER_48_1639 ();
 sg13g2_fill_2 FILLER_48_1646 ();
 sg13g2_decap_4 FILLER_48_1653 ();
 sg13g2_fill_1 FILLER_48_1657 ();
 sg13g2_decap_8 FILLER_48_1667 ();
 sg13g2_decap_8 FILLER_48_1674 ();
 sg13g2_decap_8 FILLER_48_1681 ();
 sg13g2_decap_8 FILLER_48_1688 ();
 sg13g2_decap_8 FILLER_48_1695 ();
 sg13g2_decap_8 FILLER_48_1702 ();
 sg13g2_decap_8 FILLER_48_1709 ();
 sg13g2_decap_8 FILLER_48_1716 ();
 sg13g2_decap_8 FILLER_48_1723 ();
 sg13g2_decap_8 FILLER_48_1730 ();
 sg13g2_fill_1 FILLER_48_1737 ();
 sg13g2_decap_8 FILLER_48_1748 ();
 sg13g2_decap_8 FILLER_48_1755 ();
 sg13g2_decap_8 FILLER_48_1762 ();
 sg13g2_decap_8 FILLER_48_1769 ();
 sg13g2_decap_8 FILLER_48_1776 ();
 sg13g2_decap_8 FILLER_48_1783 ();
 sg13g2_decap_8 FILLER_48_1790 ();
 sg13g2_decap_8 FILLER_48_1797 ();
 sg13g2_decap_8 FILLER_48_1804 ();
 sg13g2_decap_8 FILLER_48_1811 ();
 sg13g2_decap_8 FILLER_48_1818 ();
 sg13g2_decap_8 FILLER_48_1825 ();
 sg13g2_decap_8 FILLER_48_1832 ();
 sg13g2_decap_8 FILLER_48_1839 ();
 sg13g2_decap_8 FILLER_48_1846 ();
 sg13g2_decap_8 FILLER_48_1853 ();
 sg13g2_fill_2 FILLER_48_1860 ();
 sg13g2_decap_8 FILLER_48_1875 ();
 sg13g2_decap_8 FILLER_48_1882 ();
 sg13g2_decap_8 FILLER_48_1889 ();
 sg13g2_decap_8 FILLER_48_1896 ();
 sg13g2_decap_8 FILLER_48_1903 ();
 sg13g2_decap_8 FILLER_48_1910 ();
 sg13g2_decap_8 FILLER_48_1917 ();
 sg13g2_fill_2 FILLER_48_1924 ();
 sg13g2_decap_8 FILLER_48_1939 ();
 sg13g2_decap_8 FILLER_48_1946 ();
 sg13g2_decap_8 FILLER_48_1953 ();
 sg13g2_decap_8 FILLER_48_1960 ();
 sg13g2_fill_2 FILLER_48_1967 ();
 sg13g2_fill_1 FILLER_48_1969 ();
 sg13g2_decap_8 FILLER_48_1996 ();
 sg13g2_decap_8 FILLER_48_2003 ();
 sg13g2_decap_8 FILLER_48_2010 ();
 sg13g2_decap_8 FILLER_48_2017 ();
 sg13g2_decap_8 FILLER_48_2024 ();
 sg13g2_decap_8 FILLER_48_2031 ();
 sg13g2_decap_8 FILLER_48_2038 ();
 sg13g2_decap_8 FILLER_48_2045 ();
 sg13g2_decap_8 FILLER_48_2052 ();
 sg13g2_fill_2 FILLER_48_2059 ();
 sg13g2_decap_8 FILLER_48_2092 ();
 sg13g2_decap_8 FILLER_48_2099 ();
 sg13g2_decap_8 FILLER_48_2106 ();
 sg13g2_decap_8 FILLER_48_2113 ();
 sg13g2_fill_2 FILLER_48_2120 ();
 sg13g2_decap_8 FILLER_48_2126 ();
 sg13g2_decap_8 FILLER_48_2133 ();
 sg13g2_decap_8 FILLER_48_2140 ();
 sg13g2_decap_8 FILLER_48_2147 ();
 sg13g2_decap_8 FILLER_48_2154 ();
 sg13g2_decap_8 FILLER_48_2161 ();
 sg13g2_decap_8 FILLER_48_2168 ();
 sg13g2_decap_4 FILLER_48_2175 ();
 sg13g2_fill_2 FILLER_48_2179 ();
 sg13g2_fill_1 FILLER_48_2185 ();
 sg13g2_decap_8 FILLER_48_2190 ();
 sg13g2_decap_8 FILLER_48_2197 ();
 sg13g2_decap_8 FILLER_48_2204 ();
 sg13g2_decap_8 FILLER_48_2211 ();
 sg13g2_decap_8 FILLER_48_2218 ();
 sg13g2_decap_8 FILLER_48_2225 ();
 sg13g2_decap_8 FILLER_48_2232 ();
 sg13g2_decap_8 FILLER_48_2239 ();
 sg13g2_decap_8 FILLER_48_2246 ();
 sg13g2_decap_8 FILLER_48_2253 ();
 sg13g2_decap_8 FILLER_48_2260 ();
 sg13g2_decap_8 FILLER_48_2267 ();
 sg13g2_decap_8 FILLER_48_2274 ();
 sg13g2_decap_8 FILLER_48_2281 ();
 sg13g2_decap_8 FILLER_48_2288 ();
 sg13g2_decap_8 FILLER_48_2295 ();
 sg13g2_decap_8 FILLER_48_2302 ();
 sg13g2_decap_8 FILLER_48_2309 ();
 sg13g2_decap_8 FILLER_48_2316 ();
 sg13g2_decap_8 FILLER_48_2323 ();
 sg13g2_decap_8 FILLER_48_2330 ();
 sg13g2_decap_8 FILLER_48_2337 ();
 sg13g2_decap_8 FILLER_48_2344 ();
 sg13g2_decap_8 FILLER_48_2351 ();
 sg13g2_decap_8 FILLER_48_2358 ();
 sg13g2_decap_8 FILLER_48_2365 ();
 sg13g2_decap_8 FILLER_48_2372 ();
 sg13g2_decap_8 FILLER_48_2379 ();
 sg13g2_decap_8 FILLER_48_2386 ();
 sg13g2_decap_8 FILLER_48_2393 ();
 sg13g2_decap_8 FILLER_48_2400 ();
 sg13g2_decap_8 FILLER_48_2407 ();
 sg13g2_decap_8 FILLER_48_2414 ();
 sg13g2_decap_8 FILLER_48_2421 ();
 sg13g2_decap_8 FILLER_48_2428 ();
 sg13g2_decap_8 FILLER_48_2435 ();
 sg13g2_decap_8 FILLER_48_2442 ();
 sg13g2_decap_8 FILLER_48_2449 ();
 sg13g2_decap_8 FILLER_48_2456 ();
 sg13g2_decap_8 FILLER_48_2463 ();
 sg13g2_decap_8 FILLER_48_2470 ();
 sg13g2_decap_8 FILLER_48_2477 ();
 sg13g2_decap_8 FILLER_48_2484 ();
 sg13g2_decap_8 FILLER_48_2491 ();
 sg13g2_decap_8 FILLER_48_2498 ();
 sg13g2_decap_8 FILLER_48_2505 ();
 sg13g2_decap_8 FILLER_48_2512 ();
 sg13g2_decap_8 FILLER_48_2519 ();
 sg13g2_decap_8 FILLER_48_2526 ();
 sg13g2_decap_8 FILLER_48_2533 ();
 sg13g2_decap_8 FILLER_48_2540 ();
 sg13g2_decap_8 FILLER_48_2547 ();
 sg13g2_decap_8 FILLER_48_2554 ();
 sg13g2_decap_8 FILLER_48_2561 ();
 sg13g2_decap_8 FILLER_48_2568 ();
 sg13g2_decap_8 FILLER_48_2575 ();
 sg13g2_decap_8 FILLER_48_2582 ();
 sg13g2_decap_8 FILLER_48_2589 ();
 sg13g2_decap_8 FILLER_48_2596 ();
 sg13g2_decap_8 FILLER_48_2603 ();
 sg13g2_decap_8 FILLER_48_2610 ();
 sg13g2_decap_8 FILLER_48_2617 ();
 sg13g2_decap_8 FILLER_48_2624 ();
 sg13g2_decap_8 FILLER_48_2631 ();
 sg13g2_decap_8 FILLER_48_2638 ();
 sg13g2_decap_8 FILLER_48_2645 ();
 sg13g2_decap_8 FILLER_48_2652 ();
 sg13g2_decap_8 FILLER_48_2659 ();
 sg13g2_decap_4 FILLER_48_2666 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_fill_1 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_65 ();
 sg13g2_decap_8 FILLER_49_72 ();
 sg13g2_decap_8 FILLER_49_79 ();
 sg13g2_decap_8 FILLER_49_86 ();
 sg13g2_decap_8 FILLER_49_93 ();
 sg13g2_decap_8 FILLER_49_100 ();
 sg13g2_fill_2 FILLER_49_107 ();
 sg13g2_decap_8 FILLER_49_113 ();
 sg13g2_decap_8 FILLER_49_120 ();
 sg13g2_decap_8 FILLER_49_127 ();
 sg13g2_fill_2 FILLER_49_134 ();
 sg13g2_fill_1 FILLER_49_136 ();
 sg13g2_decap_8 FILLER_49_141 ();
 sg13g2_decap_8 FILLER_49_148 ();
 sg13g2_decap_8 FILLER_49_155 ();
 sg13g2_decap_8 FILLER_49_162 ();
 sg13g2_decap_8 FILLER_49_169 ();
 sg13g2_decap_8 FILLER_49_176 ();
 sg13g2_decap_8 FILLER_49_191 ();
 sg13g2_decap_8 FILLER_49_198 ();
 sg13g2_decap_8 FILLER_49_205 ();
 sg13g2_decap_8 FILLER_49_212 ();
 sg13g2_decap_8 FILLER_49_219 ();
 sg13g2_decap_8 FILLER_49_226 ();
 sg13g2_decap_8 FILLER_49_233 ();
 sg13g2_decap_8 FILLER_49_240 ();
 sg13g2_decap_8 FILLER_49_247 ();
 sg13g2_decap_8 FILLER_49_254 ();
 sg13g2_decap_8 FILLER_49_261 ();
 sg13g2_decap_8 FILLER_49_268 ();
 sg13g2_decap_8 FILLER_49_275 ();
 sg13g2_fill_2 FILLER_49_282 ();
 sg13g2_fill_1 FILLER_49_284 ();
 sg13g2_decap_8 FILLER_49_289 ();
 sg13g2_decap_8 FILLER_49_296 ();
 sg13g2_decap_8 FILLER_49_303 ();
 sg13g2_decap_8 FILLER_49_310 ();
 sg13g2_decap_8 FILLER_49_317 ();
 sg13g2_decap_8 FILLER_49_324 ();
 sg13g2_decap_8 FILLER_49_331 ();
 sg13g2_decap_8 FILLER_49_338 ();
 sg13g2_decap_8 FILLER_49_345 ();
 sg13g2_decap_8 FILLER_49_352 ();
 sg13g2_fill_2 FILLER_49_359 ();
 sg13g2_fill_1 FILLER_49_361 ();
 sg13g2_decap_8 FILLER_49_388 ();
 sg13g2_decap_8 FILLER_49_395 ();
 sg13g2_decap_8 FILLER_49_402 ();
 sg13g2_decap_8 FILLER_49_409 ();
 sg13g2_decap_8 FILLER_49_416 ();
 sg13g2_decap_8 FILLER_49_423 ();
 sg13g2_decap_8 FILLER_49_430 ();
 sg13g2_decap_4 FILLER_49_437 ();
 sg13g2_decap_8 FILLER_49_447 ();
 sg13g2_decap_8 FILLER_49_454 ();
 sg13g2_fill_2 FILLER_49_461 ();
 sg13g2_fill_1 FILLER_49_463 ();
 sg13g2_decap_8 FILLER_49_476 ();
 sg13g2_decap_4 FILLER_49_483 ();
 sg13g2_fill_2 FILLER_49_487 ();
 sg13g2_decap_8 FILLER_49_493 ();
 sg13g2_decap_8 FILLER_49_500 ();
 sg13g2_decap_8 FILLER_49_507 ();
 sg13g2_decap_8 FILLER_49_514 ();
 sg13g2_decap_4 FILLER_49_521 ();
 sg13g2_fill_1 FILLER_49_525 ();
 sg13g2_decap_8 FILLER_49_529 ();
 sg13g2_decap_8 FILLER_49_536 ();
 sg13g2_decap_8 FILLER_49_543 ();
 sg13g2_fill_1 FILLER_49_550 ();
 sg13g2_decap_8 FILLER_49_555 ();
 sg13g2_decap_8 FILLER_49_562 ();
 sg13g2_decap_8 FILLER_49_569 ();
 sg13g2_fill_1 FILLER_49_576 ();
 sg13g2_decap_8 FILLER_49_600 ();
 sg13g2_decap_8 FILLER_49_607 ();
 sg13g2_decap_8 FILLER_49_614 ();
 sg13g2_fill_2 FILLER_49_621 ();
 sg13g2_fill_1 FILLER_49_623 ();
 sg13g2_decap_8 FILLER_49_636 ();
 sg13g2_decap_8 FILLER_49_643 ();
 sg13g2_decap_8 FILLER_49_650 ();
 sg13g2_decap_8 FILLER_49_657 ();
 sg13g2_decap_4 FILLER_49_664 ();
 sg13g2_decap_8 FILLER_49_674 ();
 sg13g2_decap_8 FILLER_49_681 ();
 sg13g2_fill_1 FILLER_49_688 ();
 sg13g2_decap_8 FILLER_49_698 ();
 sg13g2_decap_8 FILLER_49_705 ();
 sg13g2_decap_8 FILLER_49_712 ();
 sg13g2_decap_8 FILLER_49_719 ();
 sg13g2_decap_8 FILLER_49_726 ();
 sg13g2_decap_8 FILLER_49_733 ();
 sg13g2_decap_8 FILLER_49_740 ();
 sg13g2_decap_8 FILLER_49_747 ();
 sg13g2_fill_2 FILLER_49_754 ();
 sg13g2_decap_8 FILLER_49_771 ();
 sg13g2_decap_8 FILLER_49_778 ();
 sg13g2_decap_8 FILLER_49_785 ();
 sg13g2_decap_8 FILLER_49_792 ();
 sg13g2_decap_8 FILLER_49_799 ();
 sg13g2_decap_8 FILLER_49_806 ();
 sg13g2_decap_8 FILLER_49_813 ();
 sg13g2_decap_8 FILLER_49_820 ();
 sg13g2_fill_1 FILLER_49_827 ();
 sg13g2_decap_4 FILLER_49_831 ();
 sg13g2_decap_4 FILLER_49_854 ();
 sg13g2_fill_2 FILLER_49_858 ();
 sg13g2_decap_8 FILLER_49_890 ();
 sg13g2_decap_8 FILLER_49_897 ();
 sg13g2_decap_8 FILLER_49_904 ();
 sg13g2_decap_8 FILLER_49_911 ();
 sg13g2_decap_8 FILLER_49_918 ();
 sg13g2_decap_4 FILLER_49_925 ();
 sg13g2_fill_1 FILLER_49_929 ();
 sg13g2_decap_8 FILLER_49_934 ();
 sg13g2_decap_8 FILLER_49_970 ();
 sg13g2_decap_4 FILLER_49_977 ();
 sg13g2_fill_2 FILLER_49_981 ();
 sg13g2_decap_8 FILLER_49_987 ();
 sg13g2_decap_8 FILLER_49_994 ();
 sg13g2_decap_8 FILLER_49_1001 ();
 sg13g2_decap_8 FILLER_49_1008 ();
 sg13g2_decap_8 FILLER_49_1015 ();
 sg13g2_decap_8 FILLER_49_1022 ();
 sg13g2_decap_8 FILLER_49_1029 ();
 sg13g2_decap_8 FILLER_49_1036 ();
 sg13g2_decap_8 FILLER_49_1043 ();
 sg13g2_decap_4 FILLER_49_1050 ();
 sg13g2_fill_1 FILLER_49_1058 ();
 sg13g2_decap_8 FILLER_49_1063 ();
 sg13g2_decap_8 FILLER_49_1070 ();
 sg13g2_decap_8 FILLER_49_1077 ();
 sg13g2_decap_8 FILLER_49_1093 ();
 sg13g2_decap_8 FILLER_49_1100 ();
 sg13g2_decap_8 FILLER_49_1107 ();
 sg13g2_decap_4 FILLER_49_1114 ();
 sg13g2_fill_1 FILLER_49_1118 ();
 sg13g2_decap_8 FILLER_49_1124 ();
 sg13g2_decap_8 FILLER_49_1131 ();
 sg13g2_decap_8 FILLER_49_1138 ();
 sg13g2_decap_8 FILLER_49_1145 ();
 sg13g2_decap_8 FILLER_49_1152 ();
 sg13g2_decap_8 FILLER_49_1159 ();
 sg13g2_decap_4 FILLER_49_1166 ();
 sg13g2_fill_1 FILLER_49_1185 ();
 sg13g2_fill_2 FILLER_49_1190 ();
 sg13g2_fill_1 FILLER_49_1192 ();
 sg13g2_decap_8 FILLER_49_1208 ();
 sg13g2_decap_8 FILLER_49_1215 ();
 sg13g2_decap_8 FILLER_49_1222 ();
 sg13g2_decap_8 FILLER_49_1229 ();
 sg13g2_decap_8 FILLER_49_1236 ();
 sg13g2_decap_8 FILLER_49_1243 ();
 sg13g2_decap_8 FILLER_49_1250 ();
 sg13g2_decap_8 FILLER_49_1257 ();
 sg13g2_decap_8 FILLER_49_1264 ();
 sg13g2_decap_4 FILLER_49_1271 ();
 sg13g2_fill_2 FILLER_49_1275 ();
 sg13g2_decap_8 FILLER_49_1292 ();
 sg13g2_decap_8 FILLER_49_1299 ();
 sg13g2_fill_2 FILLER_49_1306 ();
 sg13g2_fill_1 FILLER_49_1308 ();
 sg13g2_decap_4 FILLER_49_1315 ();
 sg13g2_fill_2 FILLER_49_1319 ();
 sg13g2_decap_8 FILLER_49_1327 ();
 sg13g2_decap_8 FILLER_49_1334 ();
 sg13g2_fill_2 FILLER_49_1341 ();
 sg13g2_decap_8 FILLER_49_1347 ();
 sg13g2_decap_8 FILLER_49_1354 ();
 sg13g2_decap_8 FILLER_49_1361 ();
 sg13g2_fill_2 FILLER_49_1368 ();
 sg13g2_fill_1 FILLER_49_1370 ();
 sg13g2_decap_8 FILLER_49_1391 ();
 sg13g2_decap_8 FILLER_49_1398 ();
 sg13g2_decap_8 FILLER_49_1405 ();
 sg13g2_decap_8 FILLER_49_1412 ();
 sg13g2_decap_8 FILLER_49_1419 ();
 sg13g2_decap_8 FILLER_49_1426 ();
 sg13g2_decap_8 FILLER_49_1433 ();
 sg13g2_decap_8 FILLER_49_1440 ();
 sg13g2_decap_8 FILLER_49_1447 ();
 sg13g2_decap_8 FILLER_49_1480 ();
 sg13g2_decap_8 FILLER_49_1487 ();
 sg13g2_decap_8 FILLER_49_1494 ();
 sg13g2_decap_8 FILLER_49_1501 ();
 sg13g2_decap_8 FILLER_49_1508 ();
 sg13g2_decap_8 FILLER_49_1515 ();
 sg13g2_decap_4 FILLER_49_1522 ();
 sg13g2_fill_1 FILLER_49_1526 ();
 sg13g2_decap_8 FILLER_49_1532 ();
 sg13g2_decap_8 FILLER_49_1539 ();
 sg13g2_decap_8 FILLER_49_1546 ();
 sg13g2_decap_8 FILLER_49_1553 ();
 sg13g2_decap_4 FILLER_49_1560 ();
 sg13g2_fill_2 FILLER_49_1564 ();
 sg13g2_decap_8 FILLER_49_1575 ();
 sg13g2_decap_8 FILLER_49_1582 ();
 sg13g2_decap_8 FILLER_49_1589 ();
 sg13g2_decap_8 FILLER_49_1596 ();
 sg13g2_decap_8 FILLER_49_1603 ();
 sg13g2_decap_4 FILLER_49_1610 ();
 sg13g2_fill_2 FILLER_49_1614 ();
 sg13g2_fill_1 FILLER_49_1629 ();
 sg13g2_decap_4 FILLER_49_1642 ();
 sg13g2_fill_1 FILLER_49_1646 ();
 sg13g2_decap_4 FILLER_49_1655 ();
 sg13g2_fill_2 FILLER_49_1659 ();
 sg13g2_fill_1 FILLER_49_1664 ();
 sg13g2_decap_8 FILLER_49_1668 ();
 sg13g2_decap_8 FILLER_49_1675 ();
 sg13g2_decap_8 FILLER_49_1682 ();
 sg13g2_decap_8 FILLER_49_1689 ();
 sg13g2_decap_8 FILLER_49_1696 ();
 sg13g2_decap_8 FILLER_49_1703 ();
 sg13g2_decap_8 FILLER_49_1710 ();
 sg13g2_decap_8 FILLER_49_1717 ();
 sg13g2_decap_8 FILLER_49_1730 ();
 sg13g2_decap_8 FILLER_49_1737 ();
 sg13g2_decap_8 FILLER_49_1750 ();
 sg13g2_decap_8 FILLER_49_1757 ();
 sg13g2_decap_8 FILLER_49_1764 ();
 sg13g2_decap_8 FILLER_49_1771 ();
 sg13g2_decap_8 FILLER_49_1778 ();
 sg13g2_decap_8 FILLER_49_1785 ();
 sg13g2_decap_8 FILLER_49_1792 ();
 sg13g2_decap_4 FILLER_49_1799 ();
 sg13g2_decap_8 FILLER_49_1808 ();
 sg13g2_decap_8 FILLER_49_1815 ();
 sg13g2_decap_8 FILLER_49_1826 ();
 sg13g2_decap_8 FILLER_49_1833 ();
 sg13g2_decap_8 FILLER_49_1840 ();
 sg13g2_decap_8 FILLER_49_1847 ();
 sg13g2_decap_8 FILLER_49_1854 ();
 sg13g2_decap_8 FILLER_49_1861 ();
 sg13g2_decap_8 FILLER_49_1868 ();
 sg13g2_decap_8 FILLER_49_1875 ();
 sg13g2_decap_8 FILLER_49_1882 ();
 sg13g2_decap_8 FILLER_49_1889 ();
 sg13g2_decap_8 FILLER_49_1896 ();
 sg13g2_decap_8 FILLER_49_1903 ();
 sg13g2_decap_8 FILLER_49_1910 ();
 sg13g2_decap_8 FILLER_49_1917 ();
 sg13g2_decap_8 FILLER_49_1924 ();
 sg13g2_decap_8 FILLER_49_1931 ();
 sg13g2_decap_8 FILLER_49_1938 ();
 sg13g2_decap_8 FILLER_49_1945 ();
 sg13g2_decap_8 FILLER_49_1952 ();
 sg13g2_decap_8 FILLER_49_1959 ();
 sg13g2_decap_8 FILLER_49_1966 ();
 sg13g2_decap_8 FILLER_49_1973 ();
 sg13g2_decap_8 FILLER_49_1980 ();
 sg13g2_decap_8 FILLER_49_1987 ();
 sg13g2_decap_8 FILLER_49_1994 ();
 sg13g2_decap_8 FILLER_49_2001 ();
 sg13g2_decap_8 FILLER_49_2008 ();
 sg13g2_decap_8 FILLER_49_2015 ();
 sg13g2_decap_8 FILLER_49_2022 ();
 sg13g2_decap_8 FILLER_49_2029 ();
 sg13g2_decap_8 FILLER_49_2036 ();
 sg13g2_decap_8 FILLER_49_2043 ();
 sg13g2_decap_8 FILLER_49_2050 ();
 sg13g2_decap_8 FILLER_49_2057 ();
 sg13g2_decap_8 FILLER_49_2064 ();
 sg13g2_decap_8 FILLER_49_2071 ();
 sg13g2_decap_8 FILLER_49_2078 ();
 sg13g2_decap_8 FILLER_49_2085 ();
 sg13g2_decap_8 FILLER_49_2092 ();
 sg13g2_decap_8 FILLER_49_2099 ();
 sg13g2_decap_8 FILLER_49_2106 ();
 sg13g2_decap_8 FILLER_49_2113 ();
 sg13g2_decap_8 FILLER_49_2120 ();
 sg13g2_decap_8 FILLER_49_2127 ();
 sg13g2_decap_8 FILLER_49_2134 ();
 sg13g2_decap_8 FILLER_49_2141 ();
 sg13g2_decap_8 FILLER_49_2148 ();
 sg13g2_decap_8 FILLER_49_2155 ();
 sg13g2_decap_8 FILLER_49_2162 ();
 sg13g2_decap_8 FILLER_49_2169 ();
 sg13g2_decap_4 FILLER_49_2176 ();
 sg13g2_fill_1 FILLER_49_2180 ();
 sg13g2_decap_8 FILLER_49_2187 ();
 sg13g2_decap_8 FILLER_49_2194 ();
 sg13g2_decap_8 FILLER_49_2201 ();
 sg13g2_decap_8 FILLER_49_2208 ();
 sg13g2_decap_8 FILLER_49_2215 ();
 sg13g2_decap_8 FILLER_49_2222 ();
 sg13g2_decap_8 FILLER_49_2229 ();
 sg13g2_decap_8 FILLER_49_2236 ();
 sg13g2_decap_8 FILLER_49_2243 ();
 sg13g2_decap_8 FILLER_49_2250 ();
 sg13g2_decap_8 FILLER_49_2257 ();
 sg13g2_decap_8 FILLER_49_2264 ();
 sg13g2_decap_8 FILLER_49_2271 ();
 sg13g2_decap_8 FILLER_49_2278 ();
 sg13g2_decap_8 FILLER_49_2285 ();
 sg13g2_decap_8 FILLER_49_2292 ();
 sg13g2_decap_8 FILLER_49_2299 ();
 sg13g2_decap_8 FILLER_49_2306 ();
 sg13g2_decap_8 FILLER_49_2313 ();
 sg13g2_decap_8 FILLER_49_2320 ();
 sg13g2_decap_8 FILLER_49_2327 ();
 sg13g2_decap_8 FILLER_49_2334 ();
 sg13g2_decap_8 FILLER_49_2341 ();
 sg13g2_decap_8 FILLER_49_2348 ();
 sg13g2_decap_8 FILLER_49_2355 ();
 sg13g2_decap_8 FILLER_49_2362 ();
 sg13g2_decap_8 FILLER_49_2369 ();
 sg13g2_decap_8 FILLER_49_2376 ();
 sg13g2_decap_8 FILLER_49_2383 ();
 sg13g2_decap_8 FILLER_49_2390 ();
 sg13g2_decap_8 FILLER_49_2397 ();
 sg13g2_decap_8 FILLER_49_2404 ();
 sg13g2_decap_8 FILLER_49_2411 ();
 sg13g2_decap_8 FILLER_49_2418 ();
 sg13g2_decap_8 FILLER_49_2425 ();
 sg13g2_decap_8 FILLER_49_2432 ();
 sg13g2_decap_8 FILLER_49_2439 ();
 sg13g2_decap_8 FILLER_49_2446 ();
 sg13g2_decap_8 FILLER_49_2453 ();
 sg13g2_decap_8 FILLER_49_2460 ();
 sg13g2_decap_8 FILLER_49_2467 ();
 sg13g2_decap_8 FILLER_49_2474 ();
 sg13g2_decap_8 FILLER_49_2481 ();
 sg13g2_decap_8 FILLER_49_2488 ();
 sg13g2_decap_8 FILLER_49_2495 ();
 sg13g2_decap_8 FILLER_49_2502 ();
 sg13g2_decap_8 FILLER_49_2509 ();
 sg13g2_decap_8 FILLER_49_2516 ();
 sg13g2_decap_8 FILLER_49_2523 ();
 sg13g2_decap_8 FILLER_49_2530 ();
 sg13g2_decap_8 FILLER_49_2537 ();
 sg13g2_decap_8 FILLER_49_2544 ();
 sg13g2_decap_8 FILLER_49_2551 ();
 sg13g2_decap_8 FILLER_49_2558 ();
 sg13g2_decap_8 FILLER_49_2565 ();
 sg13g2_decap_8 FILLER_49_2572 ();
 sg13g2_decap_8 FILLER_49_2579 ();
 sg13g2_decap_8 FILLER_49_2586 ();
 sg13g2_decap_8 FILLER_49_2593 ();
 sg13g2_decap_8 FILLER_49_2600 ();
 sg13g2_decap_8 FILLER_49_2607 ();
 sg13g2_decap_8 FILLER_49_2614 ();
 sg13g2_decap_8 FILLER_49_2621 ();
 sg13g2_decap_8 FILLER_49_2628 ();
 sg13g2_decap_8 FILLER_49_2635 ();
 sg13g2_decap_8 FILLER_49_2642 ();
 sg13g2_decap_8 FILLER_49_2649 ();
 sg13g2_decap_8 FILLER_49_2656 ();
 sg13g2_decap_8 FILLER_49_2663 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_4 FILLER_50_42 ();
 sg13g2_fill_2 FILLER_50_46 ();
 sg13g2_decap_8 FILLER_50_52 ();
 sg13g2_decap_4 FILLER_50_59 ();
 sg13g2_decap_8 FILLER_50_67 ();
 sg13g2_decap_8 FILLER_50_74 ();
 sg13g2_decap_8 FILLER_50_81 ();
 sg13g2_decap_8 FILLER_50_88 ();
 sg13g2_decap_4 FILLER_50_95 ();
 sg13g2_fill_2 FILLER_50_99 ();
 sg13g2_decap_8 FILLER_50_111 ();
 sg13g2_decap_8 FILLER_50_118 ();
 sg13g2_decap_8 FILLER_50_125 ();
 sg13g2_decap_8 FILLER_50_132 ();
 sg13g2_decap_8 FILLER_50_139 ();
 sg13g2_fill_1 FILLER_50_146 ();
 sg13g2_decap_8 FILLER_50_152 ();
 sg13g2_decap_8 FILLER_50_159 ();
 sg13g2_decap_8 FILLER_50_166 ();
 sg13g2_decap_8 FILLER_50_173 ();
 sg13g2_decap_8 FILLER_50_180 ();
 sg13g2_decap_8 FILLER_50_187 ();
 sg13g2_decap_8 FILLER_50_194 ();
 sg13g2_decap_8 FILLER_50_201 ();
 sg13g2_decap_8 FILLER_50_208 ();
 sg13g2_decap_8 FILLER_50_215 ();
 sg13g2_decap_8 FILLER_50_222 ();
 sg13g2_decap_8 FILLER_50_229 ();
 sg13g2_decap_8 FILLER_50_236 ();
 sg13g2_decap_8 FILLER_50_243 ();
 sg13g2_decap_8 FILLER_50_250 ();
 sg13g2_decap_8 FILLER_50_257 ();
 sg13g2_decap_8 FILLER_50_264 ();
 sg13g2_decap_8 FILLER_50_271 ();
 sg13g2_decap_8 FILLER_50_278 ();
 sg13g2_decap_4 FILLER_50_285 ();
 sg13g2_fill_2 FILLER_50_289 ();
 sg13g2_decap_8 FILLER_50_302 ();
 sg13g2_decap_8 FILLER_50_309 ();
 sg13g2_decap_8 FILLER_50_316 ();
 sg13g2_decap_8 FILLER_50_323 ();
 sg13g2_decap_8 FILLER_50_330 ();
 sg13g2_decap_8 FILLER_50_337 ();
 sg13g2_decap_8 FILLER_50_344 ();
 sg13g2_decap_8 FILLER_50_351 ();
 sg13g2_decap_8 FILLER_50_358 ();
 sg13g2_decap_8 FILLER_50_365 ();
 sg13g2_decap_8 FILLER_50_372 ();
 sg13g2_decap_8 FILLER_50_379 ();
 sg13g2_decap_8 FILLER_50_386 ();
 sg13g2_decap_8 FILLER_50_393 ();
 sg13g2_decap_8 FILLER_50_400 ();
 sg13g2_decap_8 FILLER_50_407 ();
 sg13g2_decap_8 FILLER_50_414 ();
 sg13g2_decap_8 FILLER_50_421 ();
 sg13g2_decap_8 FILLER_50_428 ();
 sg13g2_decap_4 FILLER_50_435 ();
 sg13g2_fill_2 FILLER_50_439 ();
 sg13g2_decap_8 FILLER_50_446 ();
 sg13g2_fill_2 FILLER_50_453 ();
 sg13g2_decap_8 FILLER_50_472 ();
 sg13g2_decap_4 FILLER_50_479 ();
 sg13g2_fill_2 FILLER_50_483 ();
 sg13g2_decap_8 FILLER_50_490 ();
 sg13g2_decap_8 FILLER_50_497 ();
 sg13g2_decap_8 FILLER_50_504 ();
 sg13g2_decap_8 FILLER_50_511 ();
 sg13g2_decap_8 FILLER_50_518 ();
 sg13g2_fill_1 FILLER_50_525 ();
 sg13g2_decap_8 FILLER_50_530 ();
 sg13g2_decap_8 FILLER_50_537 ();
 sg13g2_decap_8 FILLER_50_544 ();
 sg13g2_decap_8 FILLER_50_551 ();
 sg13g2_decap_8 FILLER_50_558 ();
 sg13g2_decap_8 FILLER_50_565 ();
 sg13g2_decap_8 FILLER_50_572 ();
 sg13g2_decap_8 FILLER_50_579 ();
 sg13g2_decap_8 FILLER_50_586 ();
 sg13g2_decap_8 FILLER_50_593 ();
 sg13g2_decap_8 FILLER_50_600 ();
 sg13g2_decap_8 FILLER_50_607 ();
 sg13g2_fill_1 FILLER_50_614 ();
 sg13g2_fill_1 FILLER_50_628 ();
 sg13g2_decap_8 FILLER_50_644 ();
 sg13g2_decap_8 FILLER_50_651 ();
 sg13g2_decap_4 FILLER_50_658 ();
 sg13g2_fill_1 FILLER_50_662 ();
 sg13g2_decap_4 FILLER_50_687 ();
 sg13g2_decap_8 FILLER_50_706 ();
 sg13g2_decap_8 FILLER_50_713 ();
 sg13g2_decap_8 FILLER_50_720 ();
 sg13g2_decap_8 FILLER_50_727 ();
 sg13g2_decap_8 FILLER_50_734 ();
 sg13g2_decap_8 FILLER_50_741 ();
 sg13g2_fill_2 FILLER_50_748 ();
 sg13g2_decap_8 FILLER_50_766 ();
 sg13g2_decap_4 FILLER_50_773 ();
 sg13g2_decap_4 FILLER_50_781 ();
 sg13g2_fill_1 FILLER_50_785 ();
 sg13g2_decap_8 FILLER_50_792 ();
 sg13g2_decap_8 FILLER_50_799 ();
 sg13g2_decap_8 FILLER_50_806 ();
 sg13g2_decap_8 FILLER_50_813 ();
 sg13g2_decap_8 FILLER_50_820 ();
 sg13g2_fill_1 FILLER_50_827 ();
 sg13g2_decap_4 FILLER_50_833 ();
 sg13g2_fill_2 FILLER_50_837 ();
 sg13g2_fill_1 FILLER_50_843 ();
 sg13g2_decap_8 FILLER_50_849 ();
 sg13g2_decap_8 FILLER_50_856 ();
 sg13g2_fill_2 FILLER_50_863 ();
 sg13g2_fill_1 FILLER_50_865 ();
 sg13g2_fill_2 FILLER_50_873 ();
 sg13g2_fill_1 FILLER_50_875 ();
 sg13g2_decap_8 FILLER_50_881 ();
 sg13g2_decap_8 FILLER_50_888 ();
 sg13g2_fill_2 FILLER_50_895 ();
 sg13g2_decap_8 FILLER_50_900 ();
 sg13g2_decap_8 FILLER_50_907 ();
 sg13g2_decap_8 FILLER_50_914 ();
 sg13g2_decap_8 FILLER_50_921 ();
 sg13g2_decap_8 FILLER_50_928 ();
 sg13g2_decap_8 FILLER_50_935 ();
 sg13g2_decap_8 FILLER_50_942 ();
 sg13g2_decap_8 FILLER_50_963 ();
 sg13g2_decap_8 FILLER_50_970 ();
 sg13g2_decap_4 FILLER_50_977 ();
 sg13g2_decap_8 FILLER_50_996 ();
 sg13g2_decap_8 FILLER_50_1003 ();
 sg13g2_decap_8 FILLER_50_1010 ();
 sg13g2_decap_8 FILLER_50_1017 ();
 sg13g2_decap_8 FILLER_50_1024 ();
 sg13g2_decap_8 FILLER_50_1031 ();
 sg13g2_decap_8 FILLER_50_1038 ();
 sg13g2_decap_8 FILLER_50_1045 ();
 sg13g2_fill_2 FILLER_50_1052 ();
 sg13g2_decap_8 FILLER_50_1061 ();
 sg13g2_decap_8 FILLER_50_1068 ();
 sg13g2_decap_8 FILLER_50_1075 ();
 sg13g2_fill_2 FILLER_50_1082 ();
 sg13g2_decap_8 FILLER_50_1089 ();
 sg13g2_decap_8 FILLER_50_1096 ();
 sg13g2_decap_8 FILLER_50_1103 ();
 sg13g2_decap_8 FILLER_50_1110 ();
 sg13g2_decap_8 FILLER_50_1117 ();
 sg13g2_decap_8 FILLER_50_1124 ();
 sg13g2_decap_8 FILLER_50_1131 ();
 sg13g2_decap_8 FILLER_50_1138 ();
 sg13g2_decap_8 FILLER_50_1145 ();
 sg13g2_decap_8 FILLER_50_1152 ();
 sg13g2_decap_8 FILLER_50_1159 ();
 sg13g2_decap_8 FILLER_50_1166 ();
 sg13g2_decap_8 FILLER_50_1177 ();
 sg13g2_fill_2 FILLER_50_1184 ();
 sg13g2_fill_2 FILLER_50_1194 ();
 sg13g2_decap_8 FILLER_50_1205 ();
 sg13g2_fill_2 FILLER_50_1212 ();
 sg13g2_fill_1 FILLER_50_1214 ();
 sg13g2_decap_8 FILLER_50_1219 ();
 sg13g2_decap_4 FILLER_50_1226 ();
 sg13g2_fill_1 FILLER_50_1230 ();
 sg13g2_decap_8 FILLER_50_1236 ();
 sg13g2_decap_8 FILLER_50_1243 ();
 sg13g2_decap_8 FILLER_50_1250 ();
 sg13g2_decap_8 FILLER_50_1257 ();
 sg13g2_decap_8 FILLER_50_1264 ();
 sg13g2_decap_4 FILLER_50_1275 ();
 sg13g2_fill_1 FILLER_50_1279 ();
 sg13g2_decap_8 FILLER_50_1288 ();
 sg13g2_decap_4 FILLER_50_1295 ();
 sg13g2_decap_8 FILLER_50_1304 ();
 sg13g2_decap_8 FILLER_50_1311 ();
 sg13g2_decap_8 FILLER_50_1318 ();
 sg13g2_decap_8 FILLER_50_1325 ();
 sg13g2_fill_2 FILLER_50_1332 ();
 sg13g2_fill_1 FILLER_50_1334 ();
 sg13g2_decap_4 FILLER_50_1339 ();
 sg13g2_fill_2 FILLER_50_1343 ();
 sg13g2_decap_8 FILLER_50_1360 ();
 sg13g2_decap_4 FILLER_50_1367 ();
 sg13g2_decap_4 FILLER_50_1379 ();
 sg13g2_fill_1 FILLER_50_1383 ();
 sg13g2_decap_8 FILLER_50_1389 ();
 sg13g2_decap_8 FILLER_50_1396 ();
 sg13g2_decap_8 FILLER_50_1403 ();
 sg13g2_decap_8 FILLER_50_1410 ();
 sg13g2_decap_8 FILLER_50_1417 ();
 sg13g2_decap_8 FILLER_50_1424 ();
 sg13g2_decap_8 FILLER_50_1431 ();
 sg13g2_decap_8 FILLER_50_1438 ();
 sg13g2_decap_8 FILLER_50_1445 ();
 sg13g2_decap_8 FILLER_50_1452 ();
 sg13g2_fill_1 FILLER_50_1459 ();
 sg13g2_decap_8 FILLER_50_1475 ();
 sg13g2_decap_8 FILLER_50_1482 ();
 sg13g2_decap_8 FILLER_50_1489 ();
 sg13g2_decap_8 FILLER_50_1496 ();
 sg13g2_decap_4 FILLER_50_1503 ();
 sg13g2_fill_2 FILLER_50_1516 ();
 sg13g2_fill_1 FILLER_50_1526 ();
 sg13g2_decap_8 FILLER_50_1534 ();
 sg13g2_decap_8 FILLER_50_1541 ();
 sg13g2_decap_8 FILLER_50_1548 ();
 sg13g2_decap_8 FILLER_50_1555 ();
 sg13g2_decap_8 FILLER_50_1570 ();
 sg13g2_decap_8 FILLER_50_1577 ();
 sg13g2_decap_8 FILLER_50_1584 ();
 sg13g2_decap_8 FILLER_50_1591 ();
 sg13g2_decap_4 FILLER_50_1598 ();
 sg13g2_fill_1 FILLER_50_1602 ();
 sg13g2_decap_8 FILLER_50_1607 ();
 sg13g2_decap_8 FILLER_50_1626 ();
 sg13g2_decap_8 FILLER_50_1633 ();
 sg13g2_decap_8 FILLER_50_1640 ();
 sg13g2_decap_8 FILLER_50_1647 ();
 sg13g2_decap_8 FILLER_50_1654 ();
 sg13g2_decap_8 FILLER_50_1669 ();
 sg13g2_decap_8 FILLER_50_1676 ();
 sg13g2_decap_8 FILLER_50_1683 ();
 sg13g2_decap_8 FILLER_50_1690 ();
 sg13g2_decap_8 FILLER_50_1697 ();
 sg13g2_decap_8 FILLER_50_1704 ();
 sg13g2_decap_8 FILLER_50_1711 ();
 sg13g2_decap_8 FILLER_50_1718 ();
 sg13g2_decap_8 FILLER_50_1725 ();
 sg13g2_decap_8 FILLER_50_1732 ();
 sg13g2_decap_8 FILLER_50_1739 ();
 sg13g2_decap_8 FILLER_50_1746 ();
 sg13g2_decap_8 FILLER_50_1753 ();
 sg13g2_decap_8 FILLER_50_1760 ();
 sg13g2_decap_8 FILLER_50_1767 ();
 sg13g2_decap_8 FILLER_50_1774 ();
 sg13g2_decap_8 FILLER_50_1781 ();
 sg13g2_decap_8 FILLER_50_1788 ();
 sg13g2_decap_8 FILLER_50_1795 ();
 sg13g2_decap_8 FILLER_50_1802 ();
 sg13g2_decap_8 FILLER_50_1809 ();
 sg13g2_decap_8 FILLER_50_1816 ();
 sg13g2_decap_8 FILLER_50_1823 ();
 sg13g2_decap_8 FILLER_50_1830 ();
 sg13g2_decap_8 FILLER_50_1837 ();
 sg13g2_decap_4 FILLER_50_1844 ();
 sg13g2_fill_1 FILLER_50_1848 ();
 sg13g2_decap_8 FILLER_50_1862 ();
 sg13g2_decap_8 FILLER_50_1869 ();
 sg13g2_decap_8 FILLER_50_1876 ();
 sg13g2_decap_8 FILLER_50_1883 ();
 sg13g2_decap_8 FILLER_50_1890 ();
 sg13g2_decap_8 FILLER_50_1897 ();
 sg13g2_decap_8 FILLER_50_1904 ();
 sg13g2_decap_8 FILLER_50_1911 ();
 sg13g2_decap_8 FILLER_50_1918 ();
 sg13g2_decap_8 FILLER_50_1925 ();
 sg13g2_decap_8 FILLER_50_1932 ();
 sg13g2_decap_8 FILLER_50_1939 ();
 sg13g2_decap_8 FILLER_50_1946 ();
 sg13g2_decap_8 FILLER_50_1953 ();
 sg13g2_decap_8 FILLER_50_1960 ();
 sg13g2_decap_8 FILLER_50_1967 ();
 sg13g2_decap_8 FILLER_50_1974 ();
 sg13g2_decap_8 FILLER_50_1981 ();
 sg13g2_decap_8 FILLER_50_1988 ();
 sg13g2_decap_8 FILLER_50_1995 ();
 sg13g2_decap_4 FILLER_50_2002 ();
 sg13g2_decap_8 FILLER_50_2010 ();
 sg13g2_decap_8 FILLER_50_2017 ();
 sg13g2_decap_8 FILLER_50_2024 ();
 sg13g2_decap_8 FILLER_50_2031 ();
 sg13g2_decap_8 FILLER_50_2038 ();
 sg13g2_decap_8 FILLER_50_2045 ();
 sg13g2_decap_8 FILLER_50_2052 ();
 sg13g2_decap_8 FILLER_50_2059 ();
 sg13g2_decap_8 FILLER_50_2066 ();
 sg13g2_decap_8 FILLER_50_2073 ();
 sg13g2_decap_8 FILLER_50_2080 ();
 sg13g2_fill_2 FILLER_50_2087 ();
 sg13g2_fill_1 FILLER_50_2089 ();
 sg13g2_decap_8 FILLER_50_2093 ();
 sg13g2_decap_8 FILLER_50_2100 ();
 sg13g2_decap_8 FILLER_50_2107 ();
 sg13g2_decap_8 FILLER_50_2114 ();
 sg13g2_decap_8 FILLER_50_2121 ();
 sg13g2_decap_8 FILLER_50_2128 ();
 sg13g2_decap_8 FILLER_50_2135 ();
 sg13g2_decap_8 FILLER_50_2142 ();
 sg13g2_decap_8 FILLER_50_2149 ();
 sg13g2_decap_8 FILLER_50_2156 ();
 sg13g2_decap_8 FILLER_50_2163 ();
 sg13g2_decap_8 FILLER_50_2170 ();
 sg13g2_decap_8 FILLER_50_2177 ();
 sg13g2_decap_8 FILLER_50_2184 ();
 sg13g2_decap_8 FILLER_50_2191 ();
 sg13g2_decap_8 FILLER_50_2198 ();
 sg13g2_decap_8 FILLER_50_2205 ();
 sg13g2_decap_8 FILLER_50_2212 ();
 sg13g2_decap_8 FILLER_50_2219 ();
 sg13g2_decap_8 FILLER_50_2226 ();
 sg13g2_decap_8 FILLER_50_2233 ();
 sg13g2_decap_8 FILLER_50_2240 ();
 sg13g2_decap_8 FILLER_50_2247 ();
 sg13g2_decap_8 FILLER_50_2254 ();
 sg13g2_decap_8 FILLER_50_2261 ();
 sg13g2_decap_8 FILLER_50_2268 ();
 sg13g2_decap_8 FILLER_50_2275 ();
 sg13g2_decap_8 FILLER_50_2282 ();
 sg13g2_decap_8 FILLER_50_2289 ();
 sg13g2_decap_8 FILLER_50_2296 ();
 sg13g2_decap_8 FILLER_50_2303 ();
 sg13g2_decap_8 FILLER_50_2310 ();
 sg13g2_decap_8 FILLER_50_2317 ();
 sg13g2_decap_8 FILLER_50_2324 ();
 sg13g2_decap_8 FILLER_50_2331 ();
 sg13g2_decap_8 FILLER_50_2338 ();
 sg13g2_decap_8 FILLER_50_2345 ();
 sg13g2_decap_8 FILLER_50_2352 ();
 sg13g2_decap_8 FILLER_50_2359 ();
 sg13g2_decap_8 FILLER_50_2366 ();
 sg13g2_decap_8 FILLER_50_2373 ();
 sg13g2_decap_8 FILLER_50_2380 ();
 sg13g2_decap_8 FILLER_50_2387 ();
 sg13g2_decap_8 FILLER_50_2394 ();
 sg13g2_decap_8 FILLER_50_2401 ();
 sg13g2_decap_8 FILLER_50_2408 ();
 sg13g2_decap_8 FILLER_50_2415 ();
 sg13g2_decap_8 FILLER_50_2422 ();
 sg13g2_decap_8 FILLER_50_2429 ();
 sg13g2_decap_8 FILLER_50_2436 ();
 sg13g2_decap_8 FILLER_50_2443 ();
 sg13g2_decap_8 FILLER_50_2450 ();
 sg13g2_decap_8 FILLER_50_2457 ();
 sg13g2_decap_8 FILLER_50_2464 ();
 sg13g2_decap_8 FILLER_50_2471 ();
 sg13g2_decap_8 FILLER_50_2478 ();
 sg13g2_decap_8 FILLER_50_2485 ();
 sg13g2_decap_8 FILLER_50_2492 ();
 sg13g2_decap_8 FILLER_50_2499 ();
 sg13g2_decap_8 FILLER_50_2506 ();
 sg13g2_decap_8 FILLER_50_2513 ();
 sg13g2_decap_8 FILLER_50_2520 ();
 sg13g2_decap_8 FILLER_50_2527 ();
 sg13g2_decap_8 FILLER_50_2534 ();
 sg13g2_decap_8 FILLER_50_2541 ();
 sg13g2_decap_8 FILLER_50_2548 ();
 sg13g2_decap_8 FILLER_50_2555 ();
 sg13g2_decap_8 FILLER_50_2562 ();
 sg13g2_decap_8 FILLER_50_2569 ();
 sg13g2_decap_8 FILLER_50_2576 ();
 sg13g2_decap_8 FILLER_50_2583 ();
 sg13g2_decap_8 FILLER_50_2590 ();
 sg13g2_decap_8 FILLER_50_2597 ();
 sg13g2_decap_8 FILLER_50_2604 ();
 sg13g2_decap_8 FILLER_50_2611 ();
 sg13g2_decap_8 FILLER_50_2618 ();
 sg13g2_decap_8 FILLER_50_2625 ();
 sg13g2_decap_8 FILLER_50_2632 ();
 sg13g2_decap_8 FILLER_50_2639 ();
 sg13g2_decap_8 FILLER_50_2646 ();
 sg13g2_decap_8 FILLER_50_2653 ();
 sg13g2_decap_8 FILLER_50_2660 ();
 sg13g2_fill_2 FILLER_50_2667 ();
 sg13g2_fill_1 FILLER_50_2669 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_4 FILLER_51_56 ();
 sg13g2_fill_1 FILLER_51_60 ();
 sg13g2_fill_2 FILLER_51_65 ();
 sg13g2_decap_8 FILLER_51_71 ();
 sg13g2_decap_8 FILLER_51_78 ();
 sg13g2_decap_8 FILLER_51_85 ();
 sg13g2_decap_8 FILLER_51_92 ();
 sg13g2_fill_1 FILLER_51_99 ();
 sg13g2_decap_8 FILLER_51_104 ();
 sg13g2_decap_8 FILLER_51_111 ();
 sg13g2_decap_8 FILLER_51_118 ();
 sg13g2_decap_8 FILLER_51_125 ();
 sg13g2_decap_8 FILLER_51_132 ();
 sg13g2_decap_8 FILLER_51_139 ();
 sg13g2_decap_8 FILLER_51_146 ();
 sg13g2_fill_2 FILLER_51_153 ();
 sg13g2_decap_8 FILLER_51_159 ();
 sg13g2_decap_8 FILLER_51_166 ();
 sg13g2_decap_8 FILLER_51_173 ();
 sg13g2_decap_8 FILLER_51_180 ();
 sg13g2_decap_8 FILLER_51_187 ();
 sg13g2_decap_8 FILLER_51_194 ();
 sg13g2_decap_8 FILLER_51_201 ();
 sg13g2_decap_8 FILLER_51_208 ();
 sg13g2_decap_8 FILLER_51_215 ();
 sg13g2_decap_8 FILLER_51_222 ();
 sg13g2_decap_8 FILLER_51_229 ();
 sg13g2_decap_8 FILLER_51_236 ();
 sg13g2_decap_8 FILLER_51_243 ();
 sg13g2_decap_8 FILLER_51_254 ();
 sg13g2_decap_8 FILLER_51_261 ();
 sg13g2_decap_8 FILLER_51_268 ();
 sg13g2_decap_8 FILLER_51_275 ();
 sg13g2_decap_8 FILLER_51_282 ();
 sg13g2_decap_8 FILLER_51_289 ();
 sg13g2_decap_8 FILLER_51_296 ();
 sg13g2_decap_8 FILLER_51_303 ();
 sg13g2_decap_8 FILLER_51_310 ();
 sg13g2_decap_8 FILLER_51_317 ();
 sg13g2_decap_8 FILLER_51_324 ();
 sg13g2_decap_8 FILLER_51_331 ();
 sg13g2_decap_8 FILLER_51_338 ();
 sg13g2_decap_8 FILLER_51_345 ();
 sg13g2_decap_8 FILLER_51_352 ();
 sg13g2_decap_8 FILLER_51_359 ();
 sg13g2_fill_2 FILLER_51_366 ();
 sg13g2_decap_8 FILLER_51_372 ();
 sg13g2_decap_8 FILLER_51_379 ();
 sg13g2_decap_8 FILLER_51_386 ();
 sg13g2_decap_8 FILLER_51_393 ();
 sg13g2_decap_8 FILLER_51_400 ();
 sg13g2_decap_8 FILLER_51_407 ();
 sg13g2_decap_8 FILLER_51_414 ();
 sg13g2_decap_8 FILLER_51_421 ();
 sg13g2_decap_8 FILLER_51_428 ();
 sg13g2_decap_8 FILLER_51_435 ();
 sg13g2_decap_8 FILLER_51_442 ();
 sg13g2_decap_8 FILLER_51_449 ();
 sg13g2_decap_8 FILLER_51_456 ();
 sg13g2_decap_8 FILLER_51_463 ();
 sg13g2_decap_8 FILLER_51_470 ();
 sg13g2_decap_8 FILLER_51_477 ();
 sg13g2_decap_8 FILLER_51_489 ();
 sg13g2_decap_8 FILLER_51_496 ();
 sg13g2_decap_8 FILLER_51_503 ();
 sg13g2_decap_4 FILLER_51_510 ();
 sg13g2_fill_2 FILLER_51_514 ();
 sg13g2_decap_8 FILLER_51_521 ();
 sg13g2_decap_8 FILLER_51_528 ();
 sg13g2_decap_8 FILLER_51_550 ();
 sg13g2_decap_8 FILLER_51_557 ();
 sg13g2_decap_8 FILLER_51_564 ();
 sg13g2_decap_8 FILLER_51_571 ();
 sg13g2_decap_4 FILLER_51_578 ();
 sg13g2_fill_1 FILLER_51_582 ();
 sg13g2_decap_8 FILLER_51_598 ();
 sg13g2_decap_8 FILLER_51_605 ();
 sg13g2_decap_4 FILLER_51_612 ();
 sg13g2_decap_8 FILLER_51_646 ();
 sg13g2_decap_8 FILLER_51_653 ();
 sg13g2_decap_8 FILLER_51_660 ();
 sg13g2_fill_2 FILLER_51_673 ();
 sg13g2_decap_8 FILLER_51_679 ();
 sg13g2_decap_8 FILLER_51_686 ();
 sg13g2_fill_1 FILLER_51_693 ();
 sg13g2_decap_8 FILLER_51_700 ();
 sg13g2_fill_2 FILLER_51_707 ();
 sg13g2_fill_1 FILLER_51_709 ();
 sg13g2_fill_1 FILLER_51_719 ();
 sg13g2_decap_8 FILLER_51_758 ();
 sg13g2_decap_4 FILLER_51_765 ();
 sg13g2_decap_8 FILLER_51_772 ();
 sg13g2_decap_8 FILLER_51_779 ();
 sg13g2_decap_8 FILLER_51_786 ();
 sg13g2_decap_8 FILLER_51_793 ();
 sg13g2_decap_8 FILLER_51_800 ();
 sg13g2_decap_8 FILLER_51_807 ();
 sg13g2_decap_8 FILLER_51_814 ();
 sg13g2_decap_8 FILLER_51_821 ();
 sg13g2_decap_4 FILLER_51_831 ();
 sg13g2_fill_1 FILLER_51_835 ();
 sg13g2_decap_8 FILLER_51_840 ();
 sg13g2_decap_8 FILLER_51_847 ();
 sg13g2_decap_8 FILLER_51_854 ();
 sg13g2_decap_8 FILLER_51_861 ();
 sg13g2_fill_1 FILLER_51_868 ();
 sg13g2_decap_8 FILLER_51_875 ();
 sg13g2_decap_8 FILLER_51_882 ();
 sg13g2_decap_4 FILLER_51_889 ();
 sg13g2_fill_1 FILLER_51_893 ();
 sg13g2_decap_8 FILLER_51_904 ();
 sg13g2_decap_8 FILLER_51_911 ();
 sg13g2_decap_8 FILLER_51_918 ();
 sg13g2_decap_8 FILLER_51_925 ();
 sg13g2_fill_1 FILLER_51_932 ();
 sg13g2_decap_4 FILLER_51_948 ();
 sg13g2_fill_2 FILLER_51_952 ();
 sg13g2_decap_8 FILLER_51_958 ();
 sg13g2_decap_8 FILLER_51_965 ();
 sg13g2_decap_8 FILLER_51_991 ();
 sg13g2_decap_8 FILLER_51_998 ();
 sg13g2_decap_8 FILLER_51_1005 ();
 sg13g2_decap_8 FILLER_51_1012 ();
 sg13g2_decap_8 FILLER_51_1019 ();
 sg13g2_decap_8 FILLER_51_1026 ();
 sg13g2_decap_8 FILLER_51_1033 ();
 sg13g2_decap_8 FILLER_51_1040 ();
 sg13g2_decap_8 FILLER_51_1047 ();
 sg13g2_decap_8 FILLER_51_1054 ();
 sg13g2_decap_8 FILLER_51_1061 ();
 sg13g2_decap_8 FILLER_51_1068 ();
 sg13g2_decap_8 FILLER_51_1075 ();
 sg13g2_decap_8 FILLER_51_1082 ();
 sg13g2_decap_8 FILLER_51_1089 ();
 sg13g2_fill_1 FILLER_51_1100 ();
 sg13g2_decap_8 FILLER_51_1113 ();
 sg13g2_decap_8 FILLER_51_1120 ();
 sg13g2_decap_8 FILLER_51_1127 ();
 sg13g2_decap_8 FILLER_51_1134 ();
 sg13g2_decap_4 FILLER_51_1141 ();
 sg13g2_decap_8 FILLER_51_1154 ();
 sg13g2_decap_8 FILLER_51_1161 ();
 sg13g2_fill_1 FILLER_51_1168 ();
 sg13g2_decap_8 FILLER_51_1179 ();
 sg13g2_decap_8 FILLER_51_1186 ();
 sg13g2_decap_8 FILLER_51_1193 ();
 sg13g2_decap_8 FILLER_51_1200 ();
 sg13g2_decap_8 FILLER_51_1207 ();
 sg13g2_decap_8 FILLER_51_1214 ();
 sg13g2_decap_8 FILLER_51_1233 ();
 sg13g2_decap_8 FILLER_51_1240 ();
 sg13g2_decap_8 FILLER_51_1247 ();
 sg13g2_decap_8 FILLER_51_1254 ();
 sg13g2_decap_8 FILLER_51_1261 ();
 sg13g2_decap_8 FILLER_51_1268 ();
 sg13g2_decap_8 FILLER_51_1275 ();
 sg13g2_decap_8 FILLER_51_1282 ();
 sg13g2_decap_8 FILLER_51_1289 ();
 sg13g2_decap_8 FILLER_51_1296 ();
 sg13g2_decap_8 FILLER_51_1303 ();
 sg13g2_decap_8 FILLER_51_1310 ();
 sg13g2_decap_8 FILLER_51_1317 ();
 sg13g2_decap_8 FILLER_51_1324 ();
 sg13g2_decap_8 FILLER_51_1331 ();
 sg13g2_decap_4 FILLER_51_1338 ();
 sg13g2_decap_8 FILLER_51_1350 ();
 sg13g2_decap_8 FILLER_51_1357 ();
 sg13g2_decap_8 FILLER_51_1364 ();
 sg13g2_decap_8 FILLER_51_1371 ();
 sg13g2_decap_8 FILLER_51_1378 ();
 sg13g2_decap_8 FILLER_51_1385 ();
 sg13g2_decap_8 FILLER_51_1392 ();
 sg13g2_decap_8 FILLER_51_1399 ();
 sg13g2_decap_8 FILLER_51_1406 ();
 sg13g2_decap_8 FILLER_51_1413 ();
 sg13g2_decap_8 FILLER_51_1420 ();
 sg13g2_decap_4 FILLER_51_1427 ();
 sg13g2_fill_1 FILLER_51_1431 ();
 sg13g2_fill_1 FILLER_51_1441 ();
 sg13g2_decap_8 FILLER_51_1463 ();
 sg13g2_decap_8 FILLER_51_1470 ();
 sg13g2_decap_8 FILLER_51_1477 ();
 sg13g2_decap_8 FILLER_51_1484 ();
 sg13g2_decap_8 FILLER_51_1491 ();
 sg13g2_decap_8 FILLER_51_1498 ();
 sg13g2_fill_2 FILLER_51_1505 ();
 sg13g2_fill_1 FILLER_51_1511 ();
 sg13g2_decap_8 FILLER_51_1516 ();
 sg13g2_decap_8 FILLER_51_1523 ();
 sg13g2_decap_8 FILLER_51_1530 ();
 sg13g2_decap_8 FILLER_51_1537 ();
 sg13g2_decap_8 FILLER_51_1544 ();
 sg13g2_decap_8 FILLER_51_1551 ();
 sg13g2_decap_8 FILLER_51_1558 ();
 sg13g2_decap_8 FILLER_51_1565 ();
 sg13g2_decap_8 FILLER_51_1572 ();
 sg13g2_decap_8 FILLER_51_1579 ();
 sg13g2_decap_8 FILLER_51_1586 ();
 sg13g2_decap_8 FILLER_51_1593 ();
 sg13g2_decap_4 FILLER_51_1600 ();
 sg13g2_fill_1 FILLER_51_1604 ();
 sg13g2_decap_8 FILLER_51_1609 ();
 sg13g2_decap_8 FILLER_51_1616 ();
 sg13g2_fill_2 FILLER_51_1623 ();
 sg13g2_fill_1 FILLER_51_1625 ();
 sg13g2_decap_8 FILLER_51_1641 ();
 sg13g2_decap_8 FILLER_51_1648 ();
 sg13g2_decap_8 FILLER_51_1655 ();
 sg13g2_decap_8 FILLER_51_1662 ();
 sg13g2_decap_8 FILLER_51_1669 ();
 sg13g2_decap_8 FILLER_51_1676 ();
 sg13g2_decap_8 FILLER_51_1683 ();
 sg13g2_fill_2 FILLER_51_1690 ();
 sg13g2_fill_1 FILLER_51_1692 ();
 sg13g2_decap_8 FILLER_51_1708 ();
 sg13g2_decap_8 FILLER_51_1715 ();
 sg13g2_decap_8 FILLER_51_1722 ();
 sg13g2_decap_8 FILLER_51_1729 ();
 sg13g2_decap_8 FILLER_51_1736 ();
 sg13g2_fill_1 FILLER_51_1743 ();
 sg13g2_decap_8 FILLER_51_1748 ();
 sg13g2_decap_8 FILLER_51_1755 ();
 sg13g2_decap_8 FILLER_51_1762 ();
 sg13g2_fill_2 FILLER_51_1769 ();
 sg13g2_decap_8 FILLER_51_1776 ();
 sg13g2_decap_8 FILLER_51_1792 ();
 sg13g2_decap_8 FILLER_51_1799 ();
 sg13g2_decap_8 FILLER_51_1806 ();
 sg13g2_decap_8 FILLER_51_1813 ();
 sg13g2_decap_8 FILLER_51_1820 ();
 sg13g2_decap_8 FILLER_51_1827 ();
 sg13g2_decap_8 FILLER_51_1834 ();
 sg13g2_decap_8 FILLER_51_1841 ();
 sg13g2_decap_8 FILLER_51_1848 ();
 sg13g2_decap_8 FILLER_51_1855 ();
 sg13g2_decap_8 FILLER_51_1862 ();
 sg13g2_decap_8 FILLER_51_1869 ();
 sg13g2_decap_8 FILLER_51_1876 ();
 sg13g2_decap_8 FILLER_51_1883 ();
 sg13g2_decap_8 FILLER_51_1890 ();
 sg13g2_decap_8 FILLER_51_1897 ();
 sg13g2_decap_8 FILLER_51_1904 ();
 sg13g2_decap_8 FILLER_51_1911 ();
 sg13g2_decap_8 FILLER_51_1918 ();
 sg13g2_decap_8 FILLER_51_1925 ();
 sg13g2_decap_8 FILLER_51_1932 ();
 sg13g2_decap_8 FILLER_51_1939 ();
 sg13g2_decap_8 FILLER_51_1946 ();
 sg13g2_decap_8 FILLER_51_1953 ();
 sg13g2_decap_8 FILLER_51_1960 ();
 sg13g2_decap_8 FILLER_51_1967 ();
 sg13g2_decap_8 FILLER_51_1974 ();
 sg13g2_decap_8 FILLER_51_1981 ();
 sg13g2_decap_8 FILLER_51_1988 ();
 sg13g2_decap_4 FILLER_51_1995 ();
 sg13g2_decap_8 FILLER_51_2025 ();
 sg13g2_decap_8 FILLER_51_2032 ();
 sg13g2_decap_8 FILLER_51_2039 ();
 sg13g2_decap_8 FILLER_51_2046 ();
 sg13g2_decap_8 FILLER_51_2053 ();
 sg13g2_decap_8 FILLER_51_2060 ();
 sg13g2_decap_8 FILLER_51_2067 ();
 sg13g2_decap_8 FILLER_51_2074 ();
 sg13g2_decap_8 FILLER_51_2081 ();
 sg13g2_decap_8 FILLER_51_2088 ();
 sg13g2_decap_8 FILLER_51_2095 ();
 sg13g2_decap_8 FILLER_51_2106 ();
 sg13g2_decap_8 FILLER_51_2113 ();
 sg13g2_fill_2 FILLER_51_2120 ();
 sg13g2_decap_8 FILLER_51_2130 ();
 sg13g2_decap_8 FILLER_51_2137 ();
 sg13g2_decap_8 FILLER_51_2144 ();
 sg13g2_decap_8 FILLER_51_2151 ();
 sg13g2_decap_8 FILLER_51_2158 ();
 sg13g2_fill_2 FILLER_51_2165 ();
 sg13g2_decap_8 FILLER_51_2170 ();
 sg13g2_decap_8 FILLER_51_2177 ();
 sg13g2_decap_4 FILLER_51_2184 ();
 sg13g2_fill_1 FILLER_51_2188 ();
 sg13g2_decap_8 FILLER_51_2193 ();
 sg13g2_decap_8 FILLER_51_2200 ();
 sg13g2_decap_8 FILLER_51_2207 ();
 sg13g2_decap_8 FILLER_51_2214 ();
 sg13g2_decap_8 FILLER_51_2221 ();
 sg13g2_decap_8 FILLER_51_2228 ();
 sg13g2_decap_8 FILLER_51_2235 ();
 sg13g2_decap_8 FILLER_51_2242 ();
 sg13g2_decap_8 FILLER_51_2249 ();
 sg13g2_decap_8 FILLER_51_2256 ();
 sg13g2_decap_8 FILLER_51_2263 ();
 sg13g2_decap_8 FILLER_51_2270 ();
 sg13g2_decap_8 FILLER_51_2277 ();
 sg13g2_decap_8 FILLER_51_2284 ();
 sg13g2_decap_8 FILLER_51_2291 ();
 sg13g2_decap_8 FILLER_51_2298 ();
 sg13g2_decap_8 FILLER_51_2305 ();
 sg13g2_decap_8 FILLER_51_2312 ();
 sg13g2_decap_8 FILLER_51_2319 ();
 sg13g2_decap_8 FILLER_51_2326 ();
 sg13g2_decap_8 FILLER_51_2333 ();
 sg13g2_decap_8 FILLER_51_2340 ();
 sg13g2_decap_8 FILLER_51_2347 ();
 sg13g2_decap_8 FILLER_51_2354 ();
 sg13g2_decap_8 FILLER_51_2361 ();
 sg13g2_decap_8 FILLER_51_2368 ();
 sg13g2_decap_8 FILLER_51_2375 ();
 sg13g2_decap_8 FILLER_51_2382 ();
 sg13g2_decap_8 FILLER_51_2389 ();
 sg13g2_decap_8 FILLER_51_2396 ();
 sg13g2_decap_8 FILLER_51_2403 ();
 sg13g2_decap_8 FILLER_51_2410 ();
 sg13g2_decap_8 FILLER_51_2417 ();
 sg13g2_decap_8 FILLER_51_2424 ();
 sg13g2_decap_8 FILLER_51_2431 ();
 sg13g2_decap_8 FILLER_51_2438 ();
 sg13g2_decap_8 FILLER_51_2445 ();
 sg13g2_decap_8 FILLER_51_2452 ();
 sg13g2_decap_8 FILLER_51_2459 ();
 sg13g2_decap_8 FILLER_51_2466 ();
 sg13g2_decap_8 FILLER_51_2473 ();
 sg13g2_decap_8 FILLER_51_2480 ();
 sg13g2_decap_8 FILLER_51_2487 ();
 sg13g2_decap_8 FILLER_51_2494 ();
 sg13g2_decap_8 FILLER_51_2501 ();
 sg13g2_decap_8 FILLER_51_2508 ();
 sg13g2_decap_8 FILLER_51_2515 ();
 sg13g2_decap_8 FILLER_51_2522 ();
 sg13g2_decap_8 FILLER_51_2529 ();
 sg13g2_decap_8 FILLER_51_2536 ();
 sg13g2_decap_8 FILLER_51_2543 ();
 sg13g2_decap_8 FILLER_51_2550 ();
 sg13g2_decap_8 FILLER_51_2557 ();
 sg13g2_decap_8 FILLER_51_2564 ();
 sg13g2_decap_8 FILLER_51_2571 ();
 sg13g2_decap_8 FILLER_51_2578 ();
 sg13g2_decap_8 FILLER_51_2585 ();
 sg13g2_decap_8 FILLER_51_2592 ();
 sg13g2_decap_8 FILLER_51_2599 ();
 sg13g2_decap_8 FILLER_51_2606 ();
 sg13g2_decap_8 FILLER_51_2613 ();
 sg13g2_decap_8 FILLER_51_2620 ();
 sg13g2_decap_8 FILLER_51_2627 ();
 sg13g2_decap_8 FILLER_51_2634 ();
 sg13g2_decap_8 FILLER_51_2641 ();
 sg13g2_decap_8 FILLER_51_2648 ();
 sg13g2_decap_8 FILLER_51_2655 ();
 sg13g2_decap_8 FILLER_51_2662 ();
 sg13g2_fill_1 FILLER_51_2669 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_8 FILLER_52_91 ();
 sg13g2_fill_2 FILLER_52_98 ();
 sg13g2_decap_8 FILLER_52_103 ();
 sg13g2_decap_8 FILLER_52_110 ();
 sg13g2_decap_8 FILLER_52_117 ();
 sg13g2_decap_8 FILLER_52_124 ();
 sg13g2_decap_8 FILLER_52_131 ();
 sg13g2_decap_8 FILLER_52_138 ();
 sg13g2_decap_8 FILLER_52_145 ();
 sg13g2_decap_8 FILLER_52_152 ();
 sg13g2_decap_8 FILLER_52_162 ();
 sg13g2_decap_4 FILLER_52_169 ();
 sg13g2_decap_8 FILLER_52_178 ();
 sg13g2_decap_8 FILLER_52_185 ();
 sg13g2_decap_8 FILLER_52_192 ();
 sg13g2_decap_8 FILLER_52_199 ();
 sg13g2_decap_8 FILLER_52_206 ();
 sg13g2_decap_8 FILLER_52_213 ();
 sg13g2_decap_8 FILLER_52_220 ();
 sg13g2_decap_8 FILLER_52_227 ();
 sg13g2_decap_8 FILLER_52_234 ();
 sg13g2_fill_2 FILLER_52_241 ();
 sg13g2_decap_8 FILLER_52_269 ();
 sg13g2_decap_8 FILLER_52_276 ();
 sg13g2_decap_8 FILLER_52_283 ();
 sg13g2_decap_8 FILLER_52_290 ();
 sg13g2_decap_8 FILLER_52_297 ();
 sg13g2_decap_8 FILLER_52_304 ();
 sg13g2_decap_8 FILLER_52_311 ();
 sg13g2_decap_8 FILLER_52_318 ();
 sg13g2_decap_8 FILLER_52_325 ();
 sg13g2_decap_8 FILLER_52_332 ();
 sg13g2_decap_8 FILLER_52_339 ();
 sg13g2_decap_8 FILLER_52_346 ();
 sg13g2_decap_8 FILLER_52_353 ();
 sg13g2_decap_8 FILLER_52_360 ();
 sg13g2_decap_8 FILLER_52_367 ();
 sg13g2_decap_8 FILLER_52_374 ();
 sg13g2_decap_8 FILLER_52_381 ();
 sg13g2_decap_8 FILLER_52_388 ();
 sg13g2_decap_8 FILLER_52_395 ();
 sg13g2_fill_1 FILLER_52_402 ();
 sg13g2_decap_8 FILLER_52_408 ();
 sg13g2_decap_4 FILLER_52_415 ();
 sg13g2_fill_1 FILLER_52_419 ();
 sg13g2_decap_8 FILLER_52_424 ();
 sg13g2_decap_4 FILLER_52_431 ();
 sg13g2_fill_2 FILLER_52_435 ();
 sg13g2_decap_8 FILLER_52_441 ();
 sg13g2_decap_8 FILLER_52_448 ();
 sg13g2_decap_8 FILLER_52_455 ();
 sg13g2_decap_8 FILLER_52_462 ();
 sg13g2_decap_8 FILLER_52_469 ();
 sg13g2_decap_8 FILLER_52_476 ();
 sg13g2_decap_8 FILLER_52_483 ();
 sg13g2_decap_8 FILLER_52_490 ();
 sg13g2_decap_8 FILLER_52_497 ();
 sg13g2_decap_8 FILLER_52_504 ();
 sg13g2_decap_8 FILLER_52_511 ();
 sg13g2_decap_8 FILLER_52_518 ();
 sg13g2_fill_1 FILLER_52_525 ();
 sg13g2_decap_4 FILLER_52_545 ();
 sg13g2_fill_1 FILLER_52_549 ();
 sg13g2_decap_8 FILLER_52_559 ();
 sg13g2_decap_8 FILLER_52_566 ();
 sg13g2_decap_8 FILLER_52_573 ();
 sg13g2_fill_1 FILLER_52_580 ();
 sg13g2_decap_8 FILLER_52_590 ();
 sg13g2_decap_8 FILLER_52_597 ();
 sg13g2_fill_1 FILLER_52_633 ();
 sg13g2_decap_8 FILLER_52_640 ();
 sg13g2_decap_8 FILLER_52_647 ();
 sg13g2_decap_8 FILLER_52_654 ();
 sg13g2_decap_8 FILLER_52_661 ();
 sg13g2_decap_8 FILLER_52_668 ();
 sg13g2_decap_8 FILLER_52_675 ();
 sg13g2_decap_8 FILLER_52_682 ();
 sg13g2_decap_8 FILLER_52_689 ();
 sg13g2_decap_4 FILLER_52_696 ();
 sg13g2_fill_1 FILLER_52_700 ();
 sg13g2_decap_8 FILLER_52_720 ();
 sg13g2_decap_4 FILLER_52_727 ();
 sg13g2_fill_1 FILLER_52_731 ();
 sg13g2_decap_4 FILLER_52_740 ();
 sg13g2_fill_2 FILLER_52_744 ();
 sg13g2_fill_1 FILLER_52_751 ();
 sg13g2_fill_2 FILLER_52_767 ();
 sg13g2_decap_8 FILLER_52_779 ();
 sg13g2_decap_8 FILLER_52_786 ();
 sg13g2_decap_8 FILLER_52_793 ();
 sg13g2_fill_2 FILLER_52_800 ();
 sg13g2_fill_1 FILLER_52_806 ();
 sg13g2_decap_8 FILLER_52_812 ();
 sg13g2_decap_8 FILLER_52_819 ();
 sg13g2_decap_8 FILLER_52_826 ();
 sg13g2_decap_8 FILLER_52_833 ();
 sg13g2_decap_8 FILLER_52_840 ();
 sg13g2_decap_8 FILLER_52_847 ();
 sg13g2_decap_4 FILLER_52_854 ();
 sg13g2_fill_1 FILLER_52_858 ();
 sg13g2_decap_8 FILLER_52_863 ();
 sg13g2_decap_8 FILLER_52_870 ();
 sg13g2_decap_8 FILLER_52_877 ();
 sg13g2_decap_8 FILLER_52_884 ();
 sg13g2_decap_4 FILLER_52_891 ();
 sg13g2_fill_2 FILLER_52_895 ();
 sg13g2_decap_8 FILLER_52_904 ();
 sg13g2_decap_8 FILLER_52_911 ();
 sg13g2_decap_8 FILLER_52_918 ();
 sg13g2_decap_8 FILLER_52_925 ();
 sg13g2_decap_4 FILLER_52_932 ();
 sg13g2_decap_8 FILLER_52_940 ();
 sg13g2_decap_8 FILLER_52_947 ();
 sg13g2_decap_8 FILLER_52_954 ();
 sg13g2_decap_8 FILLER_52_961 ();
 sg13g2_decap_8 FILLER_52_968 ();
 sg13g2_decap_8 FILLER_52_975 ();
 sg13g2_decap_8 FILLER_52_982 ();
 sg13g2_decap_8 FILLER_52_989 ();
 sg13g2_decap_8 FILLER_52_996 ();
 sg13g2_decap_8 FILLER_52_1003 ();
 sg13g2_decap_8 FILLER_52_1014 ();
 sg13g2_decap_8 FILLER_52_1021 ();
 sg13g2_fill_2 FILLER_52_1028 ();
 sg13g2_decap_8 FILLER_52_1035 ();
 sg13g2_decap_8 FILLER_52_1042 ();
 sg13g2_decap_8 FILLER_52_1049 ();
 sg13g2_fill_2 FILLER_52_1056 ();
 sg13g2_fill_1 FILLER_52_1058 ();
 sg13g2_decap_8 FILLER_52_1063 ();
 sg13g2_decap_8 FILLER_52_1070 ();
 sg13g2_decap_8 FILLER_52_1077 ();
 sg13g2_decap_8 FILLER_52_1084 ();
 sg13g2_fill_2 FILLER_52_1091 ();
 sg13g2_decap_8 FILLER_52_1106 ();
 sg13g2_decap_8 FILLER_52_1113 ();
 sg13g2_decap_8 FILLER_52_1120 ();
 sg13g2_decap_8 FILLER_52_1127 ();
 sg13g2_fill_1 FILLER_52_1134 ();
 sg13g2_decap_8 FILLER_52_1139 ();
 sg13g2_fill_2 FILLER_52_1146 ();
 sg13g2_decap_8 FILLER_52_1156 ();
 sg13g2_decap_4 FILLER_52_1163 ();
 sg13g2_fill_2 FILLER_52_1167 ();
 sg13g2_decap_8 FILLER_52_1184 ();
 sg13g2_decap_8 FILLER_52_1191 ();
 sg13g2_decap_8 FILLER_52_1198 ();
 sg13g2_decap_8 FILLER_52_1205 ();
 sg13g2_decap_8 FILLER_52_1228 ();
 sg13g2_decap_8 FILLER_52_1235 ();
 sg13g2_decap_8 FILLER_52_1242 ();
 sg13g2_decap_8 FILLER_52_1249 ();
 sg13g2_decap_8 FILLER_52_1256 ();
 sg13g2_decap_8 FILLER_52_1263 ();
 sg13g2_decap_8 FILLER_52_1270 ();
 sg13g2_decap_8 FILLER_52_1277 ();
 sg13g2_decap_4 FILLER_52_1284 ();
 sg13g2_decap_8 FILLER_52_1292 ();
 sg13g2_decap_8 FILLER_52_1299 ();
 sg13g2_decap_8 FILLER_52_1306 ();
 sg13g2_decap_8 FILLER_52_1313 ();
 sg13g2_decap_8 FILLER_52_1320 ();
 sg13g2_decap_8 FILLER_52_1327 ();
 sg13g2_decap_8 FILLER_52_1334 ();
 sg13g2_decap_8 FILLER_52_1341 ();
 sg13g2_decap_8 FILLER_52_1348 ();
 sg13g2_decap_8 FILLER_52_1355 ();
 sg13g2_decap_8 FILLER_52_1362 ();
 sg13g2_decap_8 FILLER_52_1369 ();
 sg13g2_fill_1 FILLER_52_1376 ();
 sg13g2_decap_8 FILLER_52_1386 ();
 sg13g2_decap_8 FILLER_52_1399 ();
 sg13g2_fill_1 FILLER_52_1406 ();
 sg13g2_decap_8 FILLER_52_1410 ();
 sg13g2_decap_8 FILLER_52_1417 ();
 sg13g2_decap_8 FILLER_52_1424 ();
 sg13g2_fill_1 FILLER_52_1431 ();
 sg13g2_decap_8 FILLER_52_1447 ();
 sg13g2_decap_8 FILLER_52_1454 ();
 sg13g2_decap_8 FILLER_52_1461 ();
 sg13g2_decap_8 FILLER_52_1468 ();
 sg13g2_decap_4 FILLER_52_1475 ();
 sg13g2_decap_8 FILLER_52_1485 ();
 sg13g2_decap_8 FILLER_52_1492 ();
 sg13g2_decap_8 FILLER_52_1499 ();
 sg13g2_decap_4 FILLER_52_1506 ();
 sg13g2_fill_2 FILLER_52_1510 ();
 sg13g2_decap_8 FILLER_52_1515 ();
 sg13g2_decap_8 FILLER_52_1522 ();
 sg13g2_fill_1 FILLER_52_1529 ();
 sg13g2_decap_8 FILLER_52_1545 ();
 sg13g2_decap_8 FILLER_52_1552 ();
 sg13g2_decap_8 FILLER_52_1559 ();
 sg13g2_decap_8 FILLER_52_1566 ();
 sg13g2_decap_8 FILLER_52_1573 ();
 sg13g2_decap_8 FILLER_52_1580 ();
 sg13g2_decap_8 FILLER_52_1587 ();
 sg13g2_decap_8 FILLER_52_1594 ();
 sg13g2_decap_8 FILLER_52_1601 ();
 sg13g2_decap_8 FILLER_52_1608 ();
 sg13g2_decap_8 FILLER_52_1615 ();
 sg13g2_decap_4 FILLER_52_1622 ();
 sg13g2_decap_4 FILLER_52_1631 ();
 sg13g2_fill_1 FILLER_52_1635 ();
 sg13g2_decap_8 FILLER_52_1644 ();
 sg13g2_decap_8 FILLER_52_1651 ();
 sg13g2_decap_8 FILLER_52_1658 ();
 sg13g2_decap_8 FILLER_52_1665 ();
 sg13g2_decap_8 FILLER_52_1672 ();
 sg13g2_decap_8 FILLER_52_1679 ();
 sg13g2_decap_8 FILLER_52_1686 ();
 sg13g2_fill_1 FILLER_52_1701 ();
 sg13g2_fill_2 FILLER_52_1722 ();
 sg13g2_fill_2 FILLER_52_1728 ();
 sg13g2_fill_1 FILLER_52_1730 ();
 sg13g2_decap_8 FILLER_52_1739 ();
 sg13g2_decap_8 FILLER_52_1746 ();
 sg13g2_decap_8 FILLER_52_1753 ();
 sg13g2_decap_8 FILLER_52_1760 ();
 sg13g2_decap_4 FILLER_52_1767 ();
 sg13g2_fill_2 FILLER_52_1771 ();
 sg13g2_decap_8 FILLER_52_1789 ();
 sg13g2_decap_8 FILLER_52_1796 ();
 sg13g2_decap_8 FILLER_52_1803 ();
 sg13g2_decap_8 FILLER_52_1810 ();
 sg13g2_decap_8 FILLER_52_1817 ();
 sg13g2_decap_8 FILLER_52_1824 ();
 sg13g2_decap_8 FILLER_52_1831 ();
 sg13g2_decap_8 FILLER_52_1838 ();
 sg13g2_decap_8 FILLER_52_1845 ();
 sg13g2_decap_8 FILLER_52_1852 ();
 sg13g2_decap_8 FILLER_52_1859 ();
 sg13g2_decap_8 FILLER_52_1866 ();
 sg13g2_decap_8 FILLER_52_1873 ();
 sg13g2_decap_8 FILLER_52_1880 ();
 sg13g2_decap_8 FILLER_52_1887 ();
 sg13g2_decap_8 FILLER_52_1894 ();
 sg13g2_decap_8 FILLER_52_1901 ();
 sg13g2_decap_8 FILLER_52_1908 ();
 sg13g2_decap_8 FILLER_52_1915 ();
 sg13g2_decap_8 FILLER_52_1922 ();
 sg13g2_decap_8 FILLER_52_1929 ();
 sg13g2_decap_8 FILLER_52_1936 ();
 sg13g2_decap_8 FILLER_52_1943 ();
 sg13g2_decap_8 FILLER_52_1950 ();
 sg13g2_decap_8 FILLER_52_1957 ();
 sg13g2_decap_8 FILLER_52_1964 ();
 sg13g2_decap_8 FILLER_52_1971 ();
 sg13g2_decap_8 FILLER_52_1978 ();
 sg13g2_decap_8 FILLER_52_1985 ();
 sg13g2_decap_8 FILLER_52_1992 ();
 sg13g2_decap_8 FILLER_52_1999 ();
 sg13g2_decap_8 FILLER_52_2006 ();
 sg13g2_decap_8 FILLER_52_2013 ();
 sg13g2_decap_8 FILLER_52_2020 ();
 sg13g2_decap_8 FILLER_52_2027 ();
 sg13g2_decap_8 FILLER_52_2034 ();
 sg13g2_decap_8 FILLER_52_2041 ();
 sg13g2_decap_8 FILLER_52_2048 ();
 sg13g2_decap_8 FILLER_52_2055 ();
 sg13g2_decap_8 FILLER_52_2062 ();
 sg13g2_decap_8 FILLER_52_2069 ();
 sg13g2_decap_8 FILLER_52_2076 ();
 sg13g2_decap_8 FILLER_52_2083 ();
 sg13g2_decap_8 FILLER_52_2090 ();
 sg13g2_decap_8 FILLER_52_2097 ();
 sg13g2_decap_8 FILLER_52_2104 ();
 sg13g2_decap_8 FILLER_52_2111 ();
 sg13g2_decap_8 FILLER_52_2130 ();
 sg13g2_decap_8 FILLER_52_2137 ();
 sg13g2_decap_8 FILLER_52_2144 ();
 sg13g2_decap_8 FILLER_52_2151 ();
 sg13g2_fill_2 FILLER_52_2158 ();
 sg13g2_decap_8 FILLER_52_2166 ();
 sg13g2_decap_8 FILLER_52_2173 ();
 sg13g2_decap_8 FILLER_52_2180 ();
 sg13g2_fill_1 FILLER_52_2187 ();
 sg13g2_decap_8 FILLER_52_2223 ();
 sg13g2_decap_8 FILLER_52_2230 ();
 sg13g2_decap_8 FILLER_52_2237 ();
 sg13g2_decap_8 FILLER_52_2244 ();
 sg13g2_decap_8 FILLER_52_2251 ();
 sg13g2_decap_8 FILLER_52_2258 ();
 sg13g2_decap_8 FILLER_52_2265 ();
 sg13g2_decap_8 FILLER_52_2272 ();
 sg13g2_decap_8 FILLER_52_2279 ();
 sg13g2_decap_8 FILLER_52_2286 ();
 sg13g2_decap_8 FILLER_52_2293 ();
 sg13g2_decap_8 FILLER_52_2300 ();
 sg13g2_decap_8 FILLER_52_2307 ();
 sg13g2_decap_8 FILLER_52_2314 ();
 sg13g2_decap_8 FILLER_52_2321 ();
 sg13g2_decap_8 FILLER_52_2328 ();
 sg13g2_decap_8 FILLER_52_2335 ();
 sg13g2_decap_8 FILLER_52_2342 ();
 sg13g2_decap_8 FILLER_52_2349 ();
 sg13g2_decap_8 FILLER_52_2356 ();
 sg13g2_decap_8 FILLER_52_2363 ();
 sg13g2_decap_8 FILLER_52_2370 ();
 sg13g2_decap_8 FILLER_52_2377 ();
 sg13g2_decap_8 FILLER_52_2384 ();
 sg13g2_decap_8 FILLER_52_2391 ();
 sg13g2_decap_8 FILLER_52_2398 ();
 sg13g2_decap_8 FILLER_52_2405 ();
 sg13g2_decap_8 FILLER_52_2412 ();
 sg13g2_decap_8 FILLER_52_2419 ();
 sg13g2_decap_8 FILLER_52_2426 ();
 sg13g2_decap_8 FILLER_52_2433 ();
 sg13g2_decap_8 FILLER_52_2440 ();
 sg13g2_decap_8 FILLER_52_2447 ();
 sg13g2_decap_8 FILLER_52_2454 ();
 sg13g2_decap_8 FILLER_52_2461 ();
 sg13g2_decap_8 FILLER_52_2468 ();
 sg13g2_decap_8 FILLER_52_2475 ();
 sg13g2_decap_8 FILLER_52_2482 ();
 sg13g2_decap_8 FILLER_52_2489 ();
 sg13g2_decap_8 FILLER_52_2496 ();
 sg13g2_decap_8 FILLER_52_2503 ();
 sg13g2_decap_8 FILLER_52_2510 ();
 sg13g2_decap_8 FILLER_52_2517 ();
 sg13g2_decap_8 FILLER_52_2524 ();
 sg13g2_decap_8 FILLER_52_2531 ();
 sg13g2_decap_8 FILLER_52_2538 ();
 sg13g2_decap_8 FILLER_52_2545 ();
 sg13g2_decap_8 FILLER_52_2552 ();
 sg13g2_decap_8 FILLER_52_2559 ();
 sg13g2_decap_8 FILLER_52_2566 ();
 sg13g2_decap_8 FILLER_52_2573 ();
 sg13g2_decap_8 FILLER_52_2580 ();
 sg13g2_decap_8 FILLER_52_2587 ();
 sg13g2_decap_8 FILLER_52_2594 ();
 sg13g2_decap_8 FILLER_52_2601 ();
 sg13g2_decap_8 FILLER_52_2608 ();
 sg13g2_decap_8 FILLER_52_2615 ();
 sg13g2_decap_8 FILLER_52_2622 ();
 sg13g2_decap_8 FILLER_52_2629 ();
 sg13g2_decap_8 FILLER_52_2636 ();
 sg13g2_decap_8 FILLER_52_2643 ();
 sg13g2_decap_8 FILLER_52_2650 ();
 sg13g2_decap_8 FILLER_52_2657 ();
 sg13g2_decap_4 FILLER_52_2664 ();
 sg13g2_fill_2 FILLER_52_2668 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_4 FILLER_53_28 ();
 sg13g2_fill_2 FILLER_53_32 ();
 sg13g2_decap_8 FILLER_53_50 ();
 sg13g2_decap_8 FILLER_53_57 ();
 sg13g2_fill_1 FILLER_53_64 ();
 sg13g2_decap_8 FILLER_53_74 ();
 sg13g2_decap_8 FILLER_53_81 ();
 sg13g2_decap_8 FILLER_53_88 ();
 sg13g2_decap_8 FILLER_53_95 ();
 sg13g2_fill_2 FILLER_53_102 ();
 sg13g2_fill_1 FILLER_53_104 ();
 sg13g2_decap_8 FILLER_53_109 ();
 sg13g2_decap_8 FILLER_53_116 ();
 sg13g2_decap_4 FILLER_53_123 ();
 sg13g2_fill_1 FILLER_53_127 ();
 sg13g2_fill_2 FILLER_53_132 ();
 sg13g2_decap_4 FILLER_53_139 ();
 sg13g2_fill_2 FILLER_53_143 ();
 sg13g2_fill_2 FILLER_53_148 ();
 sg13g2_fill_1 FILLER_53_150 ();
 sg13g2_decap_8 FILLER_53_155 ();
 sg13g2_decap_8 FILLER_53_162 ();
 sg13g2_decap_8 FILLER_53_169 ();
 sg13g2_decap_8 FILLER_53_176 ();
 sg13g2_decap_4 FILLER_53_183 ();
 sg13g2_decap_8 FILLER_53_191 ();
 sg13g2_decap_8 FILLER_53_198 ();
 sg13g2_decap_8 FILLER_53_205 ();
 sg13g2_decap_8 FILLER_53_212 ();
 sg13g2_decap_8 FILLER_53_219 ();
 sg13g2_decap_8 FILLER_53_226 ();
 sg13g2_decap_8 FILLER_53_233 ();
 sg13g2_decap_8 FILLER_53_240 ();
 sg13g2_decap_8 FILLER_53_247 ();
 sg13g2_decap_8 FILLER_53_254 ();
 sg13g2_decap_8 FILLER_53_261 ();
 sg13g2_decap_8 FILLER_53_268 ();
 sg13g2_decap_8 FILLER_53_275 ();
 sg13g2_decap_8 FILLER_53_282 ();
 sg13g2_decap_8 FILLER_53_289 ();
 sg13g2_decap_8 FILLER_53_296 ();
 sg13g2_decap_8 FILLER_53_303 ();
 sg13g2_decap_8 FILLER_53_310 ();
 sg13g2_decap_8 FILLER_53_317 ();
 sg13g2_decap_8 FILLER_53_324 ();
 sg13g2_decap_8 FILLER_53_331 ();
 sg13g2_decap_8 FILLER_53_338 ();
 sg13g2_decap_8 FILLER_53_345 ();
 sg13g2_decap_8 FILLER_53_352 ();
 sg13g2_decap_8 FILLER_53_359 ();
 sg13g2_decap_8 FILLER_53_366 ();
 sg13g2_decap_8 FILLER_53_373 ();
 sg13g2_decap_8 FILLER_53_380 ();
 sg13g2_decap_8 FILLER_53_387 ();
 sg13g2_decap_4 FILLER_53_394 ();
 sg13g2_fill_2 FILLER_53_398 ();
 sg13g2_decap_8 FILLER_53_409 ();
 sg13g2_decap_8 FILLER_53_416 ();
 sg13g2_decap_8 FILLER_53_423 ();
 sg13g2_decap_8 FILLER_53_430 ();
 sg13g2_decap_8 FILLER_53_437 ();
 sg13g2_decap_8 FILLER_53_444 ();
 sg13g2_decap_8 FILLER_53_451 ();
 sg13g2_decap_4 FILLER_53_458 ();
 sg13g2_decap_8 FILLER_53_466 ();
 sg13g2_fill_1 FILLER_53_473 ();
 sg13g2_decap_8 FILLER_53_483 ();
 sg13g2_decap_8 FILLER_53_490 ();
 sg13g2_decap_8 FILLER_53_497 ();
 sg13g2_decap_8 FILLER_53_504 ();
 sg13g2_decap_8 FILLER_53_511 ();
 sg13g2_decap_8 FILLER_53_518 ();
 sg13g2_fill_1 FILLER_53_525 ();
 sg13g2_decap_8 FILLER_53_535 ();
 sg13g2_decap_4 FILLER_53_542 ();
 sg13g2_fill_1 FILLER_53_546 ();
 sg13g2_fill_2 FILLER_53_550 ();
 sg13g2_fill_1 FILLER_53_552 ();
 sg13g2_decap_8 FILLER_53_558 ();
 sg13g2_decap_8 FILLER_53_565 ();
 sg13g2_decap_8 FILLER_53_572 ();
 sg13g2_fill_2 FILLER_53_579 ();
 sg13g2_fill_2 FILLER_53_584 ();
 sg13g2_fill_1 FILLER_53_586 ();
 sg13g2_decap_8 FILLER_53_591 ();
 sg13g2_decap_8 FILLER_53_598 ();
 sg13g2_decap_8 FILLER_53_605 ();
 sg13g2_decap_4 FILLER_53_612 ();
 sg13g2_decap_4 FILLER_53_620 ();
 sg13g2_decap_8 FILLER_53_627 ();
 sg13g2_decap_8 FILLER_53_634 ();
 sg13g2_decap_8 FILLER_53_641 ();
 sg13g2_decap_8 FILLER_53_648 ();
 sg13g2_decap_8 FILLER_53_655 ();
 sg13g2_decap_8 FILLER_53_662 ();
 sg13g2_decap_8 FILLER_53_669 ();
 sg13g2_decap_8 FILLER_53_676 ();
 sg13g2_decap_8 FILLER_53_683 ();
 sg13g2_decap_8 FILLER_53_690 ();
 sg13g2_decap_8 FILLER_53_697 ();
 sg13g2_decap_8 FILLER_53_708 ();
 sg13g2_decap_8 FILLER_53_715 ();
 sg13g2_decap_8 FILLER_53_722 ();
 sg13g2_decap_8 FILLER_53_729 ();
 sg13g2_decap_4 FILLER_53_736 ();
 sg13g2_decap_8 FILLER_53_773 ();
 sg13g2_decap_8 FILLER_53_780 ();
 sg13g2_decap_8 FILLER_53_787 ();
 sg13g2_decap_8 FILLER_53_794 ();
 sg13g2_decap_4 FILLER_53_801 ();
 sg13g2_fill_2 FILLER_53_805 ();
 sg13g2_decap_8 FILLER_53_825 ();
 sg13g2_decap_8 FILLER_53_832 ();
 sg13g2_decap_8 FILLER_53_839 ();
 sg13g2_decap_8 FILLER_53_846 ();
 sg13g2_decap_8 FILLER_53_853 ();
 sg13g2_decap_8 FILLER_53_860 ();
 sg13g2_decap_8 FILLER_53_867 ();
 sg13g2_decap_8 FILLER_53_874 ();
 sg13g2_decap_4 FILLER_53_881 ();
 sg13g2_fill_1 FILLER_53_885 ();
 sg13g2_fill_2 FILLER_53_894 ();
 sg13g2_decap_8 FILLER_53_901 ();
 sg13g2_decap_4 FILLER_53_908 ();
 sg13g2_fill_2 FILLER_53_912 ();
 sg13g2_decap_8 FILLER_53_920 ();
 sg13g2_decap_8 FILLER_53_927 ();
 sg13g2_decap_8 FILLER_53_934 ();
 sg13g2_decap_8 FILLER_53_941 ();
 sg13g2_decap_8 FILLER_53_948 ();
 sg13g2_decap_8 FILLER_53_955 ();
 sg13g2_decap_8 FILLER_53_962 ();
 sg13g2_decap_8 FILLER_53_969 ();
 sg13g2_decap_8 FILLER_53_976 ();
 sg13g2_decap_8 FILLER_53_983 ();
 sg13g2_decap_8 FILLER_53_990 ();
 sg13g2_decap_8 FILLER_53_997 ();
 sg13g2_decap_8 FILLER_53_1004 ();
 sg13g2_decap_8 FILLER_53_1011 ();
 sg13g2_decap_8 FILLER_53_1018 ();
 sg13g2_decap_8 FILLER_53_1025 ();
 sg13g2_decap_8 FILLER_53_1032 ();
 sg13g2_decap_8 FILLER_53_1039 ();
 sg13g2_decap_8 FILLER_53_1046 ();
 sg13g2_fill_1 FILLER_53_1053 ();
 sg13g2_decap_8 FILLER_53_1081 ();
 sg13g2_decap_8 FILLER_53_1088 ();
 sg13g2_decap_8 FILLER_53_1095 ();
 sg13g2_decap_8 FILLER_53_1102 ();
 sg13g2_decap_8 FILLER_53_1109 ();
 sg13g2_decap_8 FILLER_53_1116 ();
 sg13g2_decap_8 FILLER_53_1123 ();
 sg13g2_decap_8 FILLER_53_1130 ();
 sg13g2_decap_8 FILLER_53_1137 ();
 sg13g2_decap_8 FILLER_53_1144 ();
 sg13g2_decap_8 FILLER_53_1154 ();
 sg13g2_decap_8 FILLER_53_1161 ();
 sg13g2_fill_2 FILLER_53_1168 ();
 sg13g2_decap_8 FILLER_53_1175 ();
 sg13g2_decap_8 FILLER_53_1194 ();
 sg13g2_fill_2 FILLER_53_1201 ();
 sg13g2_decap_4 FILLER_53_1209 ();
 sg13g2_fill_2 FILLER_53_1213 ();
 sg13g2_decap_4 FILLER_53_1224 ();
 sg13g2_decap_8 FILLER_53_1231 ();
 sg13g2_decap_8 FILLER_53_1238 ();
 sg13g2_decap_8 FILLER_53_1245 ();
 sg13g2_decap_8 FILLER_53_1252 ();
 sg13g2_decap_8 FILLER_53_1259 ();
 sg13g2_decap_8 FILLER_53_1266 ();
 sg13g2_decap_4 FILLER_53_1273 ();
 sg13g2_fill_1 FILLER_53_1277 ();
 sg13g2_decap_8 FILLER_53_1282 ();
 sg13g2_decap_8 FILLER_53_1289 ();
 sg13g2_fill_2 FILLER_53_1296 ();
 sg13g2_fill_1 FILLER_53_1298 ();
 sg13g2_decap_8 FILLER_53_1318 ();
 sg13g2_decap_8 FILLER_53_1325 ();
 sg13g2_decap_8 FILLER_53_1332 ();
 sg13g2_fill_1 FILLER_53_1339 ();
 sg13g2_decap_8 FILLER_53_1355 ();
 sg13g2_decap_8 FILLER_53_1362 ();
 sg13g2_fill_2 FILLER_53_1369 ();
 sg13g2_fill_1 FILLER_53_1371 ();
 sg13g2_decap_8 FILLER_53_1381 ();
 sg13g2_decap_4 FILLER_53_1388 ();
 sg13g2_fill_1 FILLER_53_1392 ();
 sg13g2_decap_8 FILLER_53_1397 ();
 sg13g2_decap_8 FILLER_53_1404 ();
 sg13g2_decap_8 FILLER_53_1411 ();
 sg13g2_decap_8 FILLER_53_1418 ();
 sg13g2_decap_8 FILLER_53_1425 ();
 sg13g2_decap_8 FILLER_53_1432 ();
 sg13g2_decap_8 FILLER_53_1439 ();
 sg13g2_decap_8 FILLER_53_1446 ();
 sg13g2_fill_1 FILLER_53_1453 ();
 sg13g2_decap_4 FILLER_53_1464 ();
 sg13g2_fill_1 FILLER_53_1468 ();
 sg13g2_decap_4 FILLER_53_1474 ();
 sg13g2_fill_1 FILLER_53_1478 ();
 sg13g2_decap_4 FILLER_53_1483 ();
 sg13g2_fill_1 FILLER_53_1487 ();
 sg13g2_decap_8 FILLER_53_1494 ();
 sg13g2_decap_4 FILLER_53_1501 ();
 sg13g2_fill_1 FILLER_53_1505 ();
 sg13g2_decap_8 FILLER_53_1514 ();
 sg13g2_decap_8 FILLER_53_1521 ();
 sg13g2_fill_2 FILLER_53_1528 ();
 sg13g2_decap_8 FILLER_53_1535 ();
 sg13g2_decap_8 FILLER_53_1542 ();
 sg13g2_decap_8 FILLER_53_1549 ();
 sg13g2_decap_4 FILLER_53_1556 ();
 sg13g2_fill_2 FILLER_53_1560 ();
 sg13g2_decap_8 FILLER_53_1566 ();
 sg13g2_decap_8 FILLER_53_1573 ();
 sg13g2_decap_8 FILLER_53_1580 ();
 sg13g2_decap_8 FILLER_53_1587 ();
 sg13g2_decap_8 FILLER_53_1594 ();
 sg13g2_fill_2 FILLER_53_1606 ();
 sg13g2_decap_8 FILLER_53_1612 ();
 sg13g2_decap_8 FILLER_53_1619 ();
 sg13g2_decap_8 FILLER_53_1626 ();
 sg13g2_decap_8 FILLER_53_1633 ();
 sg13g2_decap_4 FILLER_53_1640 ();
 sg13g2_fill_1 FILLER_53_1644 ();
 sg13g2_decap_4 FILLER_53_1660 ();
 sg13g2_decap_8 FILLER_53_1668 ();
 sg13g2_decap_8 FILLER_53_1675 ();
 sg13g2_decap_8 FILLER_53_1682 ();
 sg13g2_decap_4 FILLER_53_1689 ();
 sg13g2_decap_8 FILLER_53_1696 ();
 sg13g2_decap_4 FILLER_53_1703 ();
 sg13g2_decap_8 FILLER_53_1714 ();
 sg13g2_decap_4 FILLER_53_1721 ();
 sg13g2_fill_1 FILLER_53_1725 ();
 sg13g2_decap_8 FILLER_53_1730 ();
 sg13g2_decap_8 FILLER_53_1737 ();
 sg13g2_decap_8 FILLER_53_1744 ();
 sg13g2_decap_8 FILLER_53_1751 ();
 sg13g2_decap_8 FILLER_53_1758 ();
 sg13g2_decap_8 FILLER_53_1765 ();
 sg13g2_decap_4 FILLER_53_1772 ();
 sg13g2_fill_1 FILLER_53_1776 ();
 sg13g2_fill_1 FILLER_53_1786 ();
 sg13g2_decap_8 FILLER_53_1795 ();
 sg13g2_decap_8 FILLER_53_1802 ();
 sg13g2_decap_8 FILLER_53_1809 ();
 sg13g2_decap_4 FILLER_53_1816 ();
 sg13g2_fill_2 FILLER_53_1820 ();
 sg13g2_decap_8 FILLER_53_1835 ();
 sg13g2_fill_2 FILLER_53_1842 ();
 sg13g2_decap_8 FILLER_53_1856 ();
 sg13g2_decap_8 FILLER_53_1863 ();
 sg13g2_decap_8 FILLER_53_1870 ();
 sg13g2_decap_8 FILLER_53_1877 ();
 sg13g2_decap_8 FILLER_53_1884 ();
 sg13g2_decap_8 FILLER_53_1891 ();
 sg13g2_decap_8 FILLER_53_1898 ();
 sg13g2_decap_8 FILLER_53_1905 ();
 sg13g2_decap_8 FILLER_53_1912 ();
 sg13g2_decap_8 FILLER_53_1919 ();
 sg13g2_decap_8 FILLER_53_1926 ();
 sg13g2_decap_8 FILLER_53_1933 ();
 sg13g2_decap_8 FILLER_53_1940 ();
 sg13g2_decap_8 FILLER_53_1947 ();
 sg13g2_decap_8 FILLER_53_1954 ();
 sg13g2_decap_8 FILLER_53_1961 ();
 sg13g2_decap_8 FILLER_53_1968 ();
 sg13g2_decap_8 FILLER_53_1975 ();
 sg13g2_decap_8 FILLER_53_1982 ();
 sg13g2_decap_8 FILLER_53_1989 ();
 sg13g2_decap_8 FILLER_53_1996 ();
 sg13g2_decap_8 FILLER_53_2003 ();
 sg13g2_decap_8 FILLER_53_2010 ();
 sg13g2_decap_8 FILLER_53_2017 ();
 sg13g2_decap_8 FILLER_53_2024 ();
 sg13g2_decap_8 FILLER_53_2031 ();
 sg13g2_decap_8 FILLER_53_2038 ();
 sg13g2_decap_8 FILLER_53_2045 ();
 sg13g2_decap_8 FILLER_53_2056 ();
 sg13g2_decap_8 FILLER_53_2063 ();
 sg13g2_decap_8 FILLER_53_2070 ();
 sg13g2_decap_8 FILLER_53_2077 ();
 sg13g2_decap_8 FILLER_53_2084 ();
 sg13g2_decap_8 FILLER_53_2091 ();
 sg13g2_decap_8 FILLER_53_2098 ();
 sg13g2_decap_8 FILLER_53_2105 ();
 sg13g2_decap_8 FILLER_53_2112 ();
 sg13g2_decap_8 FILLER_53_2119 ();
 sg13g2_decap_8 FILLER_53_2126 ();
 sg13g2_decap_8 FILLER_53_2133 ();
 sg13g2_decap_8 FILLER_53_2140 ();
 sg13g2_decap_8 FILLER_53_2147 ();
 sg13g2_decap_8 FILLER_53_2154 ();
 sg13g2_decap_8 FILLER_53_2161 ();
 sg13g2_decap_8 FILLER_53_2168 ();
 sg13g2_decap_8 FILLER_53_2175 ();
 sg13g2_decap_8 FILLER_53_2182 ();
 sg13g2_decap_8 FILLER_53_2189 ();
 sg13g2_decap_8 FILLER_53_2196 ();
 sg13g2_decap_8 FILLER_53_2203 ();
 sg13g2_decap_8 FILLER_53_2210 ();
 sg13g2_decap_8 FILLER_53_2217 ();
 sg13g2_decap_8 FILLER_53_2224 ();
 sg13g2_decap_8 FILLER_53_2231 ();
 sg13g2_decap_8 FILLER_53_2238 ();
 sg13g2_decap_8 FILLER_53_2245 ();
 sg13g2_decap_8 FILLER_53_2252 ();
 sg13g2_decap_8 FILLER_53_2259 ();
 sg13g2_decap_8 FILLER_53_2266 ();
 sg13g2_decap_8 FILLER_53_2273 ();
 sg13g2_decap_8 FILLER_53_2280 ();
 sg13g2_decap_8 FILLER_53_2287 ();
 sg13g2_decap_8 FILLER_53_2294 ();
 sg13g2_decap_8 FILLER_53_2301 ();
 sg13g2_decap_8 FILLER_53_2308 ();
 sg13g2_decap_8 FILLER_53_2315 ();
 sg13g2_decap_8 FILLER_53_2322 ();
 sg13g2_decap_8 FILLER_53_2329 ();
 sg13g2_decap_8 FILLER_53_2336 ();
 sg13g2_decap_8 FILLER_53_2343 ();
 sg13g2_decap_8 FILLER_53_2350 ();
 sg13g2_decap_8 FILLER_53_2357 ();
 sg13g2_decap_8 FILLER_53_2364 ();
 sg13g2_decap_8 FILLER_53_2371 ();
 sg13g2_decap_8 FILLER_53_2378 ();
 sg13g2_decap_8 FILLER_53_2385 ();
 sg13g2_decap_8 FILLER_53_2392 ();
 sg13g2_decap_8 FILLER_53_2399 ();
 sg13g2_decap_8 FILLER_53_2406 ();
 sg13g2_decap_8 FILLER_53_2413 ();
 sg13g2_decap_8 FILLER_53_2420 ();
 sg13g2_decap_8 FILLER_53_2427 ();
 sg13g2_decap_8 FILLER_53_2434 ();
 sg13g2_decap_8 FILLER_53_2441 ();
 sg13g2_decap_8 FILLER_53_2448 ();
 sg13g2_decap_8 FILLER_53_2455 ();
 sg13g2_decap_8 FILLER_53_2462 ();
 sg13g2_decap_8 FILLER_53_2469 ();
 sg13g2_decap_8 FILLER_53_2476 ();
 sg13g2_decap_8 FILLER_53_2483 ();
 sg13g2_decap_8 FILLER_53_2490 ();
 sg13g2_decap_8 FILLER_53_2497 ();
 sg13g2_decap_8 FILLER_53_2504 ();
 sg13g2_decap_8 FILLER_53_2511 ();
 sg13g2_decap_8 FILLER_53_2518 ();
 sg13g2_decap_8 FILLER_53_2525 ();
 sg13g2_decap_8 FILLER_53_2532 ();
 sg13g2_decap_8 FILLER_53_2539 ();
 sg13g2_decap_8 FILLER_53_2546 ();
 sg13g2_decap_8 FILLER_53_2553 ();
 sg13g2_decap_8 FILLER_53_2560 ();
 sg13g2_decap_8 FILLER_53_2567 ();
 sg13g2_decap_8 FILLER_53_2574 ();
 sg13g2_decap_8 FILLER_53_2581 ();
 sg13g2_decap_8 FILLER_53_2588 ();
 sg13g2_decap_8 FILLER_53_2595 ();
 sg13g2_decap_8 FILLER_53_2602 ();
 sg13g2_decap_8 FILLER_53_2609 ();
 sg13g2_decap_8 FILLER_53_2616 ();
 sg13g2_decap_8 FILLER_53_2623 ();
 sg13g2_decap_8 FILLER_53_2630 ();
 sg13g2_decap_8 FILLER_53_2637 ();
 sg13g2_decap_8 FILLER_53_2644 ();
 sg13g2_decap_8 FILLER_53_2651 ();
 sg13g2_decap_8 FILLER_53_2658 ();
 sg13g2_decap_4 FILLER_53_2665 ();
 sg13g2_fill_1 FILLER_53_2669 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_4 FILLER_54_91 ();
 sg13g2_fill_2 FILLER_54_95 ();
 sg13g2_decap_8 FILLER_54_101 ();
 sg13g2_decap_8 FILLER_54_118 ();
 sg13g2_decap_4 FILLER_54_125 ();
 sg13g2_fill_1 FILLER_54_129 ();
 sg13g2_decap_8 FILLER_54_134 ();
 sg13g2_decap_8 FILLER_54_141 ();
 sg13g2_decap_8 FILLER_54_148 ();
 sg13g2_decap_8 FILLER_54_155 ();
 sg13g2_decap_8 FILLER_54_162 ();
 sg13g2_fill_2 FILLER_54_169 ();
 sg13g2_fill_1 FILLER_54_171 ();
 sg13g2_decap_8 FILLER_54_187 ();
 sg13g2_decap_8 FILLER_54_194 ();
 sg13g2_decap_8 FILLER_54_201 ();
 sg13g2_decap_8 FILLER_54_208 ();
 sg13g2_decap_8 FILLER_54_215 ();
 sg13g2_decap_8 FILLER_54_222 ();
 sg13g2_decap_8 FILLER_54_229 ();
 sg13g2_decap_8 FILLER_54_236 ();
 sg13g2_decap_8 FILLER_54_243 ();
 sg13g2_decap_8 FILLER_54_250 ();
 sg13g2_decap_8 FILLER_54_257 ();
 sg13g2_decap_8 FILLER_54_264 ();
 sg13g2_decap_8 FILLER_54_271 ();
 sg13g2_decap_8 FILLER_54_278 ();
 sg13g2_decap_8 FILLER_54_285 ();
 sg13g2_decap_8 FILLER_54_292 ();
 sg13g2_decap_8 FILLER_54_299 ();
 sg13g2_decap_8 FILLER_54_306 ();
 sg13g2_decap_8 FILLER_54_317 ();
 sg13g2_decap_8 FILLER_54_324 ();
 sg13g2_decap_8 FILLER_54_331 ();
 sg13g2_fill_1 FILLER_54_338 ();
 sg13g2_decap_8 FILLER_54_343 ();
 sg13g2_decap_8 FILLER_54_350 ();
 sg13g2_decap_8 FILLER_54_357 ();
 sg13g2_decap_8 FILLER_54_364 ();
 sg13g2_decap_8 FILLER_54_371 ();
 sg13g2_decap_8 FILLER_54_378 ();
 sg13g2_decap_8 FILLER_54_385 ();
 sg13g2_decap_8 FILLER_54_392 ();
 sg13g2_decap_8 FILLER_54_399 ();
 sg13g2_decap_8 FILLER_54_406 ();
 sg13g2_decap_4 FILLER_54_413 ();
 sg13g2_fill_1 FILLER_54_417 ();
 sg13g2_decap_8 FILLER_54_422 ();
 sg13g2_decap_8 FILLER_54_429 ();
 sg13g2_decap_8 FILLER_54_436 ();
 sg13g2_decap_8 FILLER_54_443 ();
 sg13g2_decap_8 FILLER_54_450 ();
 sg13g2_decap_8 FILLER_54_457 ();
 sg13g2_decap_8 FILLER_54_464 ();
 sg13g2_decap_8 FILLER_54_471 ();
 sg13g2_decap_8 FILLER_54_478 ();
 sg13g2_decap_8 FILLER_54_485 ();
 sg13g2_decap_8 FILLER_54_492 ();
 sg13g2_fill_1 FILLER_54_499 ();
 sg13g2_decap_8 FILLER_54_506 ();
 sg13g2_fill_2 FILLER_54_513 ();
 sg13g2_fill_1 FILLER_54_515 ();
 sg13g2_decap_4 FILLER_54_522 ();
 sg13g2_decap_8 FILLER_54_530 ();
 sg13g2_decap_8 FILLER_54_537 ();
 sg13g2_fill_2 FILLER_54_544 ();
 sg13g2_fill_1 FILLER_54_546 ();
 sg13g2_decap_8 FILLER_54_552 ();
 sg13g2_decap_8 FILLER_54_559 ();
 sg13g2_decap_8 FILLER_54_566 ();
 sg13g2_decap_8 FILLER_54_573 ();
 sg13g2_fill_1 FILLER_54_580 ();
 sg13g2_decap_8 FILLER_54_584 ();
 sg13g2_decap_8 FILLER_54_591 ();
 sg13g2_decap_8 FILLER_54_598 ();
 sg13g2_decap_8 FILLER_54_605 ();
 sg13g2_decap_8 FILLER_54_612 ();
 sg13g2_decap_8 FILLER_54_619 ();
 sg13g2_decap_8 FILLER_54_626 ();
 sg13g2_decap_8 FILLER_54_633 ();
 sg13g2_decap_8 FILLER_54_640 ();
 sg13g2_decap_8 FILLER_54_647 ();
 sg13g2_decap_8 FILLER_54_654 ();
 sg13g2_decap_8 FILLER_54_661 ();
 sg13g2_decap_8 FILLER_54_668 ();
 sg13g2_decap_8 FILLER_54_675 ();
 sg13g2_decap_8 FILLER_54_682 ();
 sg13g2_decap_8 FILLER_54_689 ();
 sg13g2_decap_8 FILLER_54_696 ();
 sg13g2_fill_1 FILLER_54_703 ();
 sg13g2_decap_8 FILLER_54_707 ();
 sg13g2_fill_1 FILLER_54_714 ();
 sg13g2_fill_1 FILLER_54_718 ();
 sg13g2_decap_8 FILLER_54_723 ();
 sg13g2_decap_8 FILLER_54_730 ();
 sg13g2_decap_8 FILLER_54_737 ();
 sg13g2_fill_1 FILLER_54_767 ();
 sg13g2_decap_8 FILLER_54_773 ();
 sg13g2_decap_4 FILLER_54_780 ();
 sg13g2_decap_8 FILLER_54_788 ();
 sg13g2_decap_8 FILLER_54_795 ();
 sg13g2_decap_4 FILLER_54_802 ();
 sg13g2_fill_2 FILLER_54_806 ();
 sg13g2_decap_4 FILLER_54_817 ();
 sg13g2_fill_1 FILLER_54_821 ();
 sg13g2_decap_8 FILLER_54_831 ();
 sg13g2_decap_8 FILLER_54_838 ();
 sg13g2_decap_8 FILLER_54_845 ();
 sg13g2_decap_8 FILLER_54_852 ();
 sg13g2_decap_8 FILLER_54_859 ();
 sg13g2_decap_8 FILLER_54_866 ();
 sg13g2_decap_8 FILLER_54_873 ();
 sg13g2_decap_8 FILLER_54_880 ();
 sg13g2_decap_8 FILLER_54_887 ();
 sg13g2_decap_8 FILLER_54_894 ();
 sg13g2_decap_8 FILLER_54_901 ();
 sg13g2_decap_8 FILLER_54_908 ();
 sg13g2_decap_8 FILLER_54_915 ();
 sg13g2_decap_8 FILLER_54_922 ();
 sg13g2_decap_4 FILLER_54_929 ();
 sg13g2_fill_1 FILLER_54_933 ();
 sg13g2_decap_4 FILLER_54_942 ();
 sg13g2_decap_8 FILLER_54_955 ();
 sg13g2_decap_8 FILLER_54_962 ();
 sg13g2_decap_8 FILLER_54_969 ();
 sg13g2_decap_8 FILLER_54_976 ();
 sg13g2_fill_2 FILLER_54_983 ();
 sg13g2_decap_8 FILLER_54_994 ();
 sg13g2_decap_8 FILLER_54_1001 ();
 sg13g2_decap_8 FILLER_54_1008 ();
 sg13g2_decap_8 FILLER_54_1015 ();
 sg13g2_decap_4 FILLER_54_1022 ();
 sg13g2_fill_1 FILLER_54_1026 ();
 sg13g2_decap_8 FILLER_54_1031 ();
 sg13g2_fill_2 FILLER_54_1038 ();
 sg13g2_decap_8 FILLER_54_1045 ();
 sg13g2_fill_2 FILLER_54_1052 ();
 sg13g2_decap_8 FILLER_54_1076 ();
 sg13g2_decap_8 FILLER_54_1083 ();
 sg13g2_decap_4 FILLER_54_1090 ();
 sg13g2_fill_1 FILLER_54_1094 ();
 sg13g2_decap_8 FILLER_54_1100 ();
 sg13g2_decap_8 FILLER_54_1107 ();
 sg13g2_decap_8 FILLER_54_1114 ();
 sg13g2_decap_8 FILLER_54_1121 ();
 sg13g2_decap_8 FILLER_54_1128 ();
 sg13g2_decap_8 FILLER_54_1135 ();
 sg13g2_decap_8 FILLER_54_1148 ();
 sg13g2_decap_8 FILLER_54_1155 ();
 sg13g2_decap_4 FILLER_54_1162 ();
 sg13g2_fill_1 FILLER_54_1166 ();
 sg13g2_decap_8 FILLER_54_1189 ();
 sg13g2_decap_8 FILLER_54_1196 ();
 sg13g2_decap_8 FILLER_54_1203 ();
 sg13g2_decap_8 FILLER_54_1210 ();
 sg13g2_fill_1 FILLER_54_1217 ();
 sg13g2_decap_4 FILLER_54_1224 ();
 sg13g2_decap_8 FILLER_54_1233 ();
 sg13g2_fill_2 FILLER_54_1240 ();
 sg13g2_fill_1 FILLER_54_1247 ();
 sg13g2_decap_8 FILLER_54_1252 ();
 sg13g2_decap_8 FILLER_54_1259 ();
 sg13g2_decap_8 FILLER_54_1266 ();
 sg13g2_decap_4 FILLER_54_1273 ();
 sg13g2_decap_8 FILLER_54_1281 ();
 sg13g2_fill_2 FILLER_54_1288 ();
 sg13g2_fill_1 FILLER_54_1290 ();
 sg13g2_decap_8 FILLER_54_1299 ();
 sg13g2_fill_2 FILLER_54_1306 ();
 sg13g2_decap_8 FILLER_54_1313 ();
 sg13g2_fill_2 FILLER_54_1320 ();
 sg13g2_fill_1 FILLER_54_1322 ();
 sg13g2_fill_2 FILLER_54_1338 ();
 sg13g2_decap_8 FILLER_54_1348 ();
 sg13g2_fill_1 FILLER_54_1355 ();
 sg13g2_fill_1 FILLER_54_1362 ();
 sg13g2_decap_8 FILLER_54_1368 ();
 sg13g2_decap_4 FILLER_54_1375 ();
 sg13g2_fill_1 FILLER_54_1379 ();
 sg13g2_decap_8 FILLER_54_1383 ();
 sg13g2_decap_8 FILLER_54_1390 ();
 sg13g2_decap_8 FILLER_54_1397 ();
 sg13g2_decap_8 FILLER_54_1404 ();
 sg13g2_decap_8 FILLER_54_1411 ();
 sg13g2_fill_1 FILLER_54_1418 ();
 sg13g2_decap_8 FILLER_54_1423 ();
 sg13g2_decap_8 FILLER_54_1430 ();
 sg13g2_decap_8 FILLER_54_1437 ();
 sg13g2_decap_8 FILLER_54_1444 ();
 sg13g2_decap_8 FILLER_54_1451 ();
 sg13g2_decap_8 FILLER_54_1458 ();
 sg13g2_decap_8 FILLER_54_1465 ();
 sg13g2_decap_8 FILLER_54_1472 ();
 sg13g2_decap_8 FILLER_54_1479 ();
 sg13g2_decap_8 FILLER_54_1486 ();
 sg13g2_decap_8 FILLER_54_1493 ();
 sg13g2_decap_8 FILLER_54_1500 ();
 sg13g2_decap_8 FILLER_54_1507 ();
 sg13g2_decap_8 FILLER_54_1514 ();
 sg13g2_decap_8 FILLER_54_1521 ();
 sg13g2_fill_2 FILLER_54_1528 ();
 sg13g2_decap_8 FILLER_54_1535 ();
 sg13g2_decap_8 FILLER_54_1542 ();
 sg13g2_fill_2 FILLER_54_1549 ();
 sg13g2_decap_8 FILLER_54_1556 ();
 sg13g2_decap_8 FILLER_54_1563 ();
 sg13g2_decap_8 FILLER_54_1570 ();
 sg13g2_decap_4 FILLER_54_1577 ();
 sg13g2_fill_2 FILLER_54_1581 ();
 sg13g2_decap_8 FILLER_54_1588 ();
 sg13g2_fill_2 FILLER_54_1595 ();
 sg13g2_fill_2 FILLER_54_1601 ();
 sg13g2_fill_1 FILLER_54_1603 ();
 sg13g2_decap_8 FILLER_54_1608 ();
 sg13g2_decap_8 FILLER_54_1615 ();
 sg13g2_decap_4 FILLER_54_1622 ();
 sg13g2_fill_2 FILLER_54_1626 ();
 sg13g2_decap_4 FILLER_54_1640 ();
 sg13g2_fill_1 FILLER_54_1644 ();
 sg13g2_decap_8 FILLER_54_1649 ();
 sg13g2_decap_8 FILLER_54_1656 ();
 sg13g2_fill_1 FILLER_54_1663 ();
 sg13g2_decap_8 FILLER_54_1668 ();
 sg13g2_decap_8 FILLER_54_1679 ();
 sg13g2_decap_8 FILLER_54_1686 ();
 sg13g2_fill_2 FILLER_54_1693 ();
 sg13g2_decap_8 FILLER_54_1708 ();
 sg13g2_decap_8 FILLER_54_1715 ();
 sg13g2_decap_4 FILLER_54_1722 ();
 sg13g2_decap_8 FILLER_54_1730 ();
 sg13g2_decap_8 FILLER_54_1737 ();
 sg13g2_decap_8 FILLER_54_1744 ();
 sg13g2_decap_8 FILLER_54_1751 ();
 sg13g2_decap_8 FILLER_54_1758 ();
 sg13g2_decap_4 FILLER_54_1765 ();
 sg13g2_fill_2 FILLER_54_1769 ();
 sg13g2_fill_1 FILLER_54_1785 ();
 sg13g2_decap_8 FILLER_54_1808 ();
 sg13g2_decap_8 FILLER_54_1815 ();
 sg13g2_decap_8 FILLER_54_1822 ();
 sg13g2_decap_8 FILLER_54_1829 ();
 sg13g2_decap_8 FILLER_54_1836 ();
 sg13g2_decap_8 FILLER_54_1843 ();
 sg13g2_decap_8 FILLER_54_1850 ();
 sg13g2_decap_8 FILLER_54_1857 ();
 sg13g2_fill_1 FILLER_54_1864 ();
 sg13g2_decap_8 FILLER_54_1878 ();
 sg13g2_decap_8 FILLER_54_1885 ();
 sg13g2_decap_8 FILLER_54_1892 ();
 sg13g2_decap_8 FILLER_54_1899 ();
 sg13g2_decap_8 FILLER_54_1906 ();
 sg13g2_decap_8 FILLER_54_1913 ();
 sg13g2_decap_8 FILLER_54_1920 ();
 sg13g2_decap_8 FILLER_54_1927 ();
 sg13g2_decap_8 FILLER_54_1934 ();
 sg13g2_fill_2 FILLER_54_1941 ();
 sg13g2_fill_1 FILLER_54_1943 ();
 sg13g2_decap_8 FILLER_54_1957 ();
 sg13g2_decap_8 FILLER_54_1964 ();
 sg13g2_decap_8 FILLER_54_1971 ();
 sg13g2_decap_8 FILLER_54_1978 ();
 sg13g2_decap_8 FILLER_54_1985 ();
 sg13g2_decap_8 FILLER_54_1992 ();
 sg13g2_decap_8 FILLER_54_1999 ();
 sg13g2_decap_8 FILLER_54_2006 ();
 sg13g2_decap_8 FILLER_54_2013 ();
 sg13g2_fill_2 FILLER_54_2020 ();
 sg13g2_decap_8 FILLER_54_2035 ();
 sg13g2_decap_4 FILLER_54_2042 ();
 sg13g2_decap_8 FILLER_54_2072 ();
 sg13g2_decap_8 FILLER_54_2079 ();
 sg13g2_decap_8 FILLER_54_2086 ();
 sg13g2_decap_8 FILLER_54_2093 ();
 sg13g2_decap_8 FILLER_54_2100 ();
 sg13g2_decap_8 FILLER_54_2107 ();
 sg13g2_decap_8 FILLER_54_2114 ();
 sg13g2_decap_8 FILLER_54_2121 ();
 sg13g2_decap_8 FILLER_54_2128 ();
 sg13g2_decap_8 FILLER_54_2135 ();
 sg13g2_decap_4 FILLER_54_2142 ();
 sg13g2_decap_8 FILLER_54_2149 ();
 sg13g2_decap_4 FILLER_54_2156 ();
 sg13g2_fill_1 FILLER_54_2164 ();
 sg13g2_decap_8 FILLER_54_2168 ();
 sg13g2_decap_8 FILLER_54_2175 ();
 sg13g2_decap_8 FILLER_54_2182 ();
 sg13g2_decap_8 FILLER_54_2189 ();
 sg13g2_decap_8 FILLER_54_2196 ();
 sg13g2_decap_8 FILLER_54_2203 ();
 sg13g2_decap_8 FILLER_54_2210 ();
 sg13g2_decap_8 FILLER_54_2217 ();
 sg13g2_decap_8 FILLER_54_2224 ();
 sg13g2_decap_8 FILLER_54_2231 ();
 sg13g2_decap_8 FILLER_54_2238 ();
 sg13g2_decap_8 FILLER_54_2245 ();
 sg13g2_decap_8 FILLER_54_2252 ();
 sg13g2_decap_8 FILLER_54_2259 ();
 sg13g2_decap_8 FILLER_54_2266 ();
 sg13g2_decap_8 FILLER_54_2273 ();
 sg13g2_decap_8 FILLER_54_2280 ();
 sg13g2_decap_8 FILLER_54_2287 ();
 sg13g2_decap_8 FILLER_54_2294 ();
 sg13g2_decap_8 FILLER_54_2301 ();
 sg13g2_decap_8 FILLER_54_2308 ();
 sg13g2_decap_8 FILLER_54_2315 ();
 sg13g2_decap_8 FILLER_54_2322 ();
 sg13g2_decap_8 FILLER_54_2329 ();
 sg13g2_decap_8 FILLER_54_2336 ();
 sg13g2_decap_8 FILLER_54_2343 ();
 sg13g2_decap_8 FILLER_54_2350 ();
 sg13g2_decap_8 FILLER_54_2357 ();
 sg13g2_decap_8 FILLER_54_2364 ();
 sg13g2_decap_8 FILLER_54_2371 ();
 sg13g2_decap_8 FILLER_54_2378 ();
 sg13g2_decap_8 FILLER_54_2385 ();
 sg13g2_decap_8 FILLER_54_2392 ();
 sg13g2_decap_8 FILLER_54_2399 ();
 sg13g2_decap_8 FILLER_54_2406 ();
 sg13g2_decap_8 FILLER_54_2413 ();
 sg13g2_decap_8 FILLER_54_2420 ();
 sg13g2_decap_8 FILLER_54_2427 ();
 sg13g2_decap_8 FILLER_54_2434 ();
 sg13g2_decap_8 FILLER_54_2441 ();
 sg13g2_decap_8 FILLER_54_2448 ();
 sg13g2_decap_8 FILLER_54_2455 ();
 sg13g2_decap_8 FILLER_54_2462 ();
 sg13g2_decap_8 FILLER_54_2469 ();
 sg13g2_decap_8 FILLER_54_2476 ();
 sg13g2_decap_8 FILLER_54_2483 ();
 sg13g2_decap_8 FILLER_54_2490 ();
 sg13g2_decap_8 FILLER_54_2497 ();
 sg13g2_decap_8 FILLER_54_2504 ();
 sg13g2_decap_8 FILLER_54_2511 ();
 sg13g2_decap_8 FILLER_54_2518 ();
 sg13g2_decap_8 FILLER_54_2525 ();
 sg13g2_decap_8 FILLER_54_2532 ();
 sg13g2_decap_8 FILLER_54_2539 ();
 sg13g2_decap_8 FILLER_54_2546 ();
 sg13g2_decap_8 FILLER_54_2553 ();
 sg13g2_decap_8 FILLER_54_2560 ();
 sg13g2_decap_8 FILLER_54_2567 ();
 sg13g2_decap_8 FILLER_54_2574 ();
 sg13g2_decap_8 FILLER_54_2581 ();
 sg13g2_decap_8 FILLER_54_2588 ();
 sg13g2_decap_8 FILLER_54_2595 ();
 sg13g2_decap_8 FILLER_54_2602 ();
 sg13g2_decap_8 FILLER_54_2609 ();
 sg13g2_decap_8 FILLER_54_2616 ();
 sg13g2_decap_8 FILLER_54_2623 ();
 sg13g2_decap_8 FILLER_54_2630 ();
 sg13g2_decap_8 FILLER_54_2637 ();
 sg13g2_decap_8 FILLER_54_2644 ();
 sg13g2_decap_8 FILLER_54_2651 ();
 sg13g2_decap_8 FILLER_54_2658 ();
 sg13g2_decap_4 FILLER_54_2665 ();
 sg13g2_fill_1 FILLER_54_2669 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_fill_1 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_46 ();
 sg13g2_decap_8 FILLER_55_53 ();
 sg13g2_decap_8 FILLER_55_60 ();
 sg13g2_decap_8 FILLER_55_67 ();
 sg13g2_decap_4 FILLER_55_74 ();
 sg13g2_fill_1 FILLER_55_78 ();
 sg13g2_decap_8 FILLER_55_89 ();
 sg13g2_decap_8 FILLER_55_96 ();
 sg13g2_decap_8 FILLER_55_103 ();
 sg13g2_decap_8 FILLER_55_110 ();
 sg13g2_decap_8 FILLER_55_117 ();
 sg13g2_decap_8 FILLER_55_124 ();
 sg13g2_decap_8 FILLER_55_131 ();
 sg13g2_decap_8 FILLER_55_138 ();
 sg13g2_decap_8 FILLER_55_145 ();
 sg13g2_decap_8 FILLER_55_152 ();
 sg13g2_decap_8 FILLER_55_159 ();
 sg13g2_decap_4 FILLER_55_166 ();
 sg13g2_fill_2 FILLER_55_170 ();
 sg13g2_decap_8 FILLER_55_183 ();
 sg13g2_decap_8 FILLER_55_190 ();
 sg13g2_decap_8 FILLER_55_197 ();
 sg13g2_decap_8 FILLER_55_204 ();
 sg13g2_decap_8 FILLER_55_211 ();
 sg13g2_decap_8 FILLER_55_218 ();
 sg13g2_decap_8 FILLER_55_225 ();
 sg13g2_decap_8 FILLER_55_232 ();
 sg13g2_decap_8 FILLER_55_239 ();
 sg13g2_decap_8 FILLER_55_246 ();
 sg13g2_decap_8 FILLER_55_253 ();
 sg13g2_decap_8 FILLER_55_260 ();
 sg13g2_decap_8 FILLER_55_267 ();
 sg13g2_decap_8 FILLER_55_274 ();
 sg13g2_decap_8 FILLER_55_281 ();
 sg13g2_decap_8 FILLER_55_288 ();
 sg13g2_decap_8 FILLER_55_295 ();
 sg13g2_decap_8 FILLER_55_302 ();
 sg13g2_decap_4 FILLER_55_309 ();
 sg13g2_fill_2 FILLER_55_313 ();
 sg13g2_decap_8 FILLER_55_341 ();
 sg13g2_decap_8 FILLER_55_348 ();
 sg13g2_decap_8 FILLER_55_355 ();
 sg13g2_decap_8 FILLER_55_362 ();
 sg13g2_decap_8 FILLER_55_369 ();
 sg13g2_decap_8 FILLER_55_376 ();
 sg13g2_decap_8 FILLER_55_383 ();
 sg13g2_decap_8 FILLER_55_390 ();
 sg13g2_decap_8 FILLER_55_397 ();
 sg13g2_decap_4 FILLER_55_404 ();
 sg13g2_decap_8 FILLER_55_412 ();
 sg13g2_decap_8 FILLER_55_419 ();
 sg13g2_decap_8 FILLER_55_426 ();
 sg13g2_decap_4 FILLER_55_433 ();
 sg13g2_fill_1 FILLER_55_437 ();
 sg13g2_decap_8 FILLER_55_442 ();
 sg13g2_decap_8 FILLER_55_449 ();
 sg13g2_decap_8 FILLER_55_456 ();
 sg13g2_decap_8 FILLER_55_463 ();
 sg13g2_decap_8 FILLER_55_470 ();
 sg13g2_decap_8 FILLER_55_477 ();
 sg13g2_decap_4 FILLER_55_484 ();
 sg13g2_decap_8 FILLER_55_492 ();
 sg13g2_decap_8 FILLER_55_499 ();
 sg13g2_decap_8 FILLER_55_506 ();
 sg13g2_decap_8 FILLER_55_513 ();
 sg13g2_decap_8 FILLER_55_520 ();
 sg13g2_decap_4 FILLER_55_527 ();
 sg13g2_fill_2 FILLER_55_531 ();
 sg13g2_decap_8 FILLER_55_552 ();
 sg13g2_decap_8 FILLER_55_559 ();
 sg13g2_decap_8 FILLER_55_566 ();
 sg13g2_fill_2 FILLER_55_573 ();
 sg13g2_fill_1 FILLER_55_575 ();
 sg13g2_decap_8 FILLER_55_591 ();
 sg13g2_decap_8 FILLER_55_598 ();
 sg13g2_fill_2 FILLER_55_605 ();
 sg13g2_decap_4 FILLER_55_619 ();
 sg13g2_fill_2 FILLER_55_623 ();
 sg13g2_decap_8 FILLER_55_635 ();
 sg13g2_decap_8 FILLER_55_642 ();
 sg13g2_decap_8 FILLER_55_649 ();
 sg13g2_decap_8 FILLER_55_656 ();
 sg13g2_fill_2 FILLER_55_663 ();
 sg13g2_fill_1 FILLER_55_665 ();
 sg13g2_fill_2 FILLER_55_681 ();
 sg13g2_fill_1 FILLER_55_688 ();
 sg13g2_decap_8 FILLER_55_699 ();
 sg13g2_decap_8 FILLER_55_706 ();
 sg13g2_decap_8 FILLER_55_713 ();
 sg13g2_decap_8 FILLER_55_720 ();
 sg13g2_decap_8 FILLER_55_727 ();
 sg13g2_decap_8 FILLER_55_734 ();
 sg13g2_decap_8 FILLER_55_746 ();
 sg13g2_decap_4 FILLER_55_753 ();
 sg13g2_fill_1 FILLER_55_757 ();
 sg13g2_decap_4 FILLER_55_762 ();
 sg13g2_fill_2 FILLER_55_766 ();
 sg13g2_decap_8 FILLER_55_774 ();
 sg13g2_decap_8 FILLER_55_781 ();
 sg13g2_decap_8 FILLER_55_788 ();
 sg13g2_decap_8 FILLER_55_795 ();
 sg13g2_decap_8 FILLER_55_802 ();
 sg13g2_decap_8 FILLER_55_809 ();
 sg13g2_fill_1 FILLER_55_819 ();
 sg13g2_decap_8 FILLER_55_829 ();
 sg13g2_decap_8 FILLER_55_836 ();
 sg13g2_decap_8 FILLER_55_843 ();
 sg13g2_decap_8 FILLER_55_850 ();
 sg13g2_decap_8 FILLER_55_857 ();
 sg13g2_decap_4 FILLER_55_864 ();
 sg13g2_fill_2 FILLER_55_868 ();
 sg13g2_decap_8 FILLER_55_879 ();
 sg13g2_fill_2 FILLER_55_886 ();
 sg13g2_fill_2 FILLER_55_891 ();
 sg13g2_fill_1 FILLER_55_893 ();
 sg13g2_decap_8 FILLER_55_899 ();
 sg13g2_decap_8 FILLER_55_906 ();
 sg13g2_decap_8 FILLER_55_913 ();
 sg13g2_decap_8 FILLER_55_920 ();
 sg13g2_decap_8 FILLER_55_927 ();
 sg13g2_decap_8 FILLER_55_934 ();
 sg13g2_decap_8 FILLER_55_941 ();
 sg13g2_fill_2 FILLER_55_948 ();
 sg13g2_decap_8 FILLER_55_956 ();
 sg13g2_decap_8 FILLER_55_963 ();
 sg13g2_decap_8 FILLER_55_970 ();
 sg13g2_decap_8 FILLER_55_977 ();
 sg13g2_decap_8 FILLER_55_984 ();
 sg13g2_decap_8 FILLER_55_991 ();
 sg13g2_fill_1 FILLER_55_998 ();
 sg13g2_decap_8 FILLER_55_1003 ();
 sg13g2_decap_8 FILLER_55_1010 ();
 sg13g2_decap_8 FILLER_55_1017 ();
 sg13g2_decap_8 FILLER_55_1024 ();
 sg13g2_decap_8 FILLER_55_1031 ();
 sg13g2_decap_8 FILLER_55_1038 ();
 sg13g2_decap_8 FILLER_55_1045 ();
 sg13g2_decap_8 FILLER_55_1052 ();
 sg13g2_decap_8 FILLER_55_1059 ();
 sg13g2_decap_8 FILLER_55_1069 ();
 sg13g2_decap_8 FILLER_55_1076 ();
 sg13g2_decap_8 FILLER_55_1083 ();
 sg13g2_decap_8 FILLER_55_1090 ();
 sg13g2_decap_8 FILLER_55_1097 ();
 sg13g2_decap_8 FILLER_55_1104 ();
 sg13g2_decap_8 FILLER_55_1111 ();
 sg13g2_decap_8 FILLER_55_1118 ();
 sg13g2_decap_8 FILLER_55_1125 ();
 sg13g2_decap_4 FILLER_55_1132 ();
 sg13g2_decap_8 FILLER_55_1151 ();
 sg13g2_decap_8 FILLER_55_1158 ();
 sg13g2_decap_8 FILLER_55_1165 ();
 sg13g2_fill_1 FILLER_55_1172 ();
 sg13g2_fill_2 FILLER_55_1180 ();
 sg13g2_decap_8 FILLER_55_1191 ();
 sg13g2_decap_8 FILLER_55_1198 ();
 sg13g2_decap_8 FILLER_55_1205 ();
 sg13g2_decap_8 FILLER_55_1212 ();
 sg13g2_decap_8 FILLER_55_1219 ();
 sg13g2_decap_8 FILLER_55_1226 ();
 sg13g2_decap_8 FILLER_55_1233 ();
 sg13g2_decap_8 FILLER_55_1240 ();
 sg13g2_decap_8 FILLER_55_1247 ();
 sg13g2_decap_8 FILLER_55_1260 ();
 sg13g2_decap_8 FILLER_55_1267 ();
 sg13g2_decap_8 FILLER_55_1274 ();
 sg13g2_decap_8 FILLER_55_1281 ();
 sg13g2_decap_8 FILLER_55_1288 ();
 sg13g2_decap_8 FILLER_55_1295 ();
 sg13g2_fill_2 FILLER_55_1302 ();
 sg13g2_fill_1 FILLER_55_1304 ();
 sg13g2_decap_4 FILLER_55_1320 ();
 sg13g2_fill_1 FILLER_55_1324 ();
 sg13g2_decap_8 FILLER_55_1328 ();
 sg13g2_decap_8 FILLER_55_1339 ();
 sg13g2_decap_8 FILLER_55_1346 ();
 sg13g2_fill_2 FILLER_55_1353 ();
 sg13g2_fill_1 FILLER_55_1355 ();
 sg13g2_decap_8 FILLER_55_1360 ();
 sg13g2_decap_8 FILLER_55_1367 ();
 sg13g2_decap_4 FILLER_55_1374 ();
 sg13g2_fill_2 FILLER_55_1378 ();
 sg13g2_decap_4 FILLER_55_1385 ();
 sg13g2_fill_1 FILLER_55_1389 ();
 sg13g2_fill_2 FILLER_55_1394 ();
 sg13g2_fill_1 FILLER_55_1396 ();
 sg13g2_decap_8 FILLER_55_1403 ();
 sg13g2_decap_8 FILLER_55_1410 ();
 sg13g2_decap_4 FILLER_55_1417 ();
 sg13g2_decap_8 FILLER_55_1425 ();
 sg13g2_decap_8 FILLER_55_1432 ();
 sg13g2_decap_8 FILLER_55_1439 ();
 sg13g2_decap_8 FILLER_55_1446 ();
 sg13g2_decap_8 FILLER_55_1453 ();
 sg13g2_decap_8 FILLER_55_1460 ();
 sg13g2_decap_8 FILLER_55_1467 ();
 sg13g2_decap_8 FILLER_55_1474 ();
 sg13g2_decap_8 FILLER_55_1481 ();
 sg13g2_decap_8 FILLER_55_1488 ();
 sg13g2_decap_8 FILLER_55_1495 ();
 sg13g2_decap_8 FILLER_55_1502 ();
 sg13g2_decap_8 FILLER_55_1509 ();
 sg13g2_decap_8 FILLER_55_1516 ();
 sg13g2_decap_8 FILLER_55_1523 ();
 sg13g2_fill_2 FILLER_55_1530 ();
 sg13g2_decap_8 FILLER_55_1544 ();
 sg13g2_fill_2 FILLER_55_1551 ();
 sg13g2_fill_1 FILLER_55_1553 ();
 sg13g2_decap_8 FILLER_55_1560 ();
 sg13g2_decap_8 FILLER_55_1567 ();
 sg13g2_decap_8 FILLER_55_1574 ();
 sg13g2_decap_8 FILLER_55_1581 ();
 sg13g2_decap_8 FILLER_55_1588 ();
 sg13g2_decap_8 FILLER_55_1595 ();
 sg13g2_decap_8 FILLER_55_1602 ();
 sg13g2_decap_8 FILLER_55_1609 ();
 sg13g2_decap_8 FILLER_55_1616 ();
 sg13g2_decap_8 FILLER_55_1623 ();
 sg13g2_decap_8 FILLER_55_1630 ();
 sg13g2_decap_8 FILLER_55_1637 ();
 sg13g2_fill_1 FILLER_55_1644 ();
 sg13g2_decap_8 FILLER_55_1651 ();
 sg13g2_decap_8 FILLER_55_1658 ();
 sg13g2_decap_8 FILLER_55_1665 ();
 sg13g2_decap_8 FILLER_55_1672 ();
 sg13g2_decap_8 FILLER_55_1679 ();
 sg13g2_fill_2 FILLER_55_1686 ();
 sg13g2_fill_1 FILLER_55_1688 ();
 sg13g2_fill_2 FILLER_55_1703 ();
 sg13g2_decap_8 FILLER_55_1713 ();
 sg13g2_decap_8 FILLER_55_1720 ();
 sg13g2_decap_8 FILLER_55_1727 ();
 sg13g2_decap_8 FILLER_55_1734 ();
 sg13g2_decap_8 FILLER_55_1741 ();
 sg13g2_decap_8 FILLER_55_1748 ();
 sg13g2_decap_8 FILLER_55_1755 ();
 sg13g2_decap_8 FILLER_55_1762 ();
 sg13g2_decap_8 FILLER_55_1769 ();
 sg13g2_decap_8 FILLER_55_1776 ();
 sg13g2_decap_8 FILLER_55_1783 ();
 sg13g2_decap_8 FILLER_55_1790 ();
 sg13g2_decap_8 FILLER_55_1797 ();
 sg13g2_decap_8 FILLER_55_1804 ();
 sg13g2_decap_8 FILLER_55_1811 ();
 sg13g2_decap_8 FILLER_55_1818 ();
 sg13g2_decap_8 FILLER_55_1825 ();
 sg13g2_decap_8 FILLER_55_1832 ();
 sg13g2_decap_8 FILLER_55_1839 ();
 sg13g2_decap_8 FILLER_55_1846 ();
 sg13g2_decap_4 FILLER_55_1853 ();
 sg13g2_fill_2 FILLER_55_1857 ();
 sg13g2_decap_8 FILLER_55_1867 ();
 sg13g2_decap_8 FILLER_55_1874 ();
 sg13g2_decap_8 FILLER_55_1881 ();
 sg13g2_decap_8 FILLER_55_1888 ();
 sg13g2_decap_8 FILLER_55_1895 ();
 sg13g2_decap_8 FILLER_55_1902 ();
 sg13g2_decap_8 FILLER_55_1909 ();
 sg13g2_decap_8 FILLER_55_1916 ();
 sg13g2_decap_8 FILLER_55_1923 ();
 sg13g2_decap_8 FILLER_55_1930 ();
 sg13g2_decap_8 FILLER_55_1937 ();
 sg13g2_decap_8 FILLER_55_1944 ();
 sg13g2_decap_8 FILLER_55_1951 ();
 sg13g2_decap_8 FILLER_55_1958 ();
 sg13g2_decap_8 FILLER_55_1965 ();
 sg13g2_decap_8 FILLER_55_1972 ();
 sg13g2_decap_8 FILLER_55_1979 ();
 sg13g2_decap_8 FILLER_55_1986 ();
 sg13g2_decap_8 FILLER_55_1993 ();
 sg13g2_fill_2 FILLER_55_2000 ();
 sg13g2_fill_1 FILLER_55_2002 ();
 sg13g2_decap_8 FILLER_55_2007 ();
 sg13g2_decap_8 FILLER_55_2014 ();
 sg13g2_decap_8 FILLER_55_2021 ();
 sg13g2_decap_8 FILLER_55_2028 ();
 sg13g2_decap_8 FILLER_55_2035 ();
 sg13g2_decap_8 FILLER_55_2042 ();
 sg13g2_fill_1 FILLER_55_2049 ();
 sg13g2_decap_8 FILLER_55_2054 ();
 sg13g2_decap_4 FILLER_55_2061 ();
 sg13g2_fill_1 FILLER_55_2065 ();
 sg13g2_decap_8 FILLER_55_2074 ();
 sg13g2_decap_4 FILLER_55_2081 ();
 sg13g2_decap_8 FILLER_55_2091 ();
 sg13g2_decap_8 FILLER_55_2098 ();
 sg13g2_decap_8 FILLER_55_2105 ();
 sg13g2_decap_8 FILLER_55_2112 ();
 sg13g2_decap_8 FILLER_55_2119 ();
 sg13g2_decap_8 FILLER_55_2126 ();
 sg13g2_decap_8 FILLER_55_2133 ();
 sg13g2_decap_8 FILLER_55_2140 ();
 sg13g2_decap_8 FILLER_55_2147 ();
 sg13g2_decap_8 FILLER_55_2154 ();
 sg13g2_decap_4 FILLER_55_2161 ();
 sg13g2_fill_2 FILLER_55_2165 ();
 sg13g2_decap_8 FILLER_55_2177 ();
 sg13g2_decap_8 FILLER_55_2184 ();
 sg13g2_decap_4 FILLER_55_2191 ();
 sg13g2_fill_1 FILLER_55_2195 ();
 sg13g2_fill_2 FILLER_55_2204 ();
 sg13g2_decap_8 FILLER_55_2210 ();
 sg13g2_decap_8 FILLER_55_2217 ();
 sg13g2_fill_2 FILLER_55_2224 ();
 sg13g2_decap_8 FILLER_55_2256 ();
 sg13g2_decap_8 FILLER_55_2263 ();
 sg13g2_decap_8 FILLER_55_2270 ();
 sg13g2_decap_8 FILLER_55_2277 ();
 sg13g2_decap_8 FILLER_55_2284 ();
 sg13g2_decap_8 FILLER_55_2291 ();
 sg13g2_decap_8 FILLER_55_2298 ();
 sg13g2_decap_8 FILLER_55_2305 ();
 sg13g2_decap_8 FILLER_55_2312 ();
 sg13g2_decap_8 FILLER_55_2319 ();
 sg13g2_decap_8 FILLER_55_2326 ();
 sg13g2_decap_8 FILLER_55_2333 ();
 sg13g2_decap_8 FILLER_55_2340 ();
 sg13g2_decap_8 FILLER_55_2347 ();
 sg13g2_decap_8 FILLER_55_2354 ();
 sg13g2_decap_8 FILLER_55_2361 ();
 sg13g2_decap_8 FILLER_55_2368 ();
 sg13g2_decap_8 FILLER_55_2375 ();
 sg13g2_decap_8 FILLER_55_2382 ();
 sg13g2_decap_8 FILLER_55_2389 ();
 sg13g2_decap_8 FILLER_55_2396 ();
 sg13g2_decap_8 FILLER_55_2403 ();
 sg13g2_decap_8 FILLER_55_2410 ();
 sg13g2_decap_8 FILLER_55_2417 ();
 sg13g2_decap_8 FILLER_55_2424 ();
 sg13g2_decap_8 FILLER_55_2431 ();
 sg13g2_decap_8 FILLER_55_2438 ();
 sg13g2_decap_8 FILLER_55_2445 ();
 sg13g2_decap_8 FILLER_55_2452 ();
 sg13g2_decap_8 FILLER_55_2459 ();
 sg13g2_decap_8 FILLER_55_2466 ();
 sg13g2_decap_8 FILLER_55_2473 ();
 sg13g2_decap_8 FILLER_55_2480 ();
 sg13g2_decap_8 FILLER_55_2487 ();
 sg13g2_decap_8 FILLER_55_2494 ();
 sg13g2_decap_8 FILLER_55_2501 ();
 sg13g2_decap_8 FILLER_55_2508 ();
 sg13g2_decap_8 FILLER_55_2515 ();
 sg13g2_decap_8 FILLER_55_2522 ();
 sg13g2_decap_8 FILLER_55_2529 ();
 sg13g2_decap_8 FILLER_55_2536 ();
 sg13g2_decap_8 FILLER_55_2543 ();
 sg13g2_decap_8 FILLER_55_2550 ();
 sg13g2_decap_8 FILLER_55_2557 ();
 sg13g2_decap_8 FILLER_55_2564 ();
 sg13g2_decap_8 FILLER_55_2571 ();
 sg13g2_decap_8 FILLER_55_2578 ();
 sg13g2_decap_8 FILLER_55_2585 ();
 sg13g2_decap_8 FILLER_55_2592 ();
 sg13g2_decap_8 FILLER_55_2599 ();
 sg13g2_decap_8 FILLER_55_2606 ();
 sg13g2_decap_8 FILLER_55_2613 ();
 sg13g2_decap_8 FILLER_55_2620 ();
 sg13g2_decap_8 FILLER_55_2627 ();
 sg13g2_decap_8 FILLER_55_2634 ();
 sg13g2_decap_8 FILLER_55_2641 ();
 sg13g2_decap_8 FILLER_55_2648 ();
 sg13g2_decap_8 FILLER_55_2655 ();
 sg13g2_decap_8 FILLER_55_2662 ();
 sg13g2_fill_1 FILLER_55_2669 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_4 FILLER_56_35 ();
 sg13g2_fill_2 FILLER_56_39 ();
 sg13g2_decap_8 FILLER_56_46 ();
 sg13g2_fill_1 FILLER_56_53 ();
 sg13g2_decap_8 FILLER_56_58 ();
 sg13g2_decap_8 FILLER_56_65 ();
 sg13g2_decap_8 FILLER_56_72 ();
 sg13g2_fill_2 FILLER_56_79 ();
 sg13g2_decap_8 FILLER_56_86 ();
 sg13g2_decap_8 FILLER_56_93 ();
 sg13g2_decap_8 FILLER_56_100 ();
 sg13g2_decap_8 FILLER_56_107 ();
 sg13g2_decap_8 FILLER_56_114 ();
 sg13g2_decap_8 FILLER_56_121 ();
 sg13g2_fill_1 FILLER_56_128 ();
 sg13g2_decap_8 FILLER_56_133 ();
 sg13g2_decap_8 FILLER_56_140 ();
 sg13g2_decap_8 FILLER_56_147 ();
 sg13g2_decap_8 FILLER_56_154 ();
 sg13g2_decap_8 FILLER_56_161 ();
 sg13g2_decap_8 FILLER_56_168 ();
 sg13g2_decap_8 FILLER_56_175 ();
 sg13g2_decap_4 FILLER_56_182 ();
 sg13g2_fill_2 FILLER_56_186 ();
 sg13g2_decap_8 FILLER_56_197 ();
 sg13g2_decap_8 FILLER_56_204 ();
 sg13g2_decap_8 FILLER_56_211 ();
 sg13g2_decap_8 FILLER_56_218 ();
 sg13g2_decap_8 FILLER_56_225 ();
 sg13g2_decap_8 FILLER_56_232 ();
 sg13g2_decap_8 FILLER_56_239 ();
 sg13g2_decap_8 FILLER_56_246 ();
 sg13g2_decap_8 FILLER_56_253 ();
 sg13g2_decap_8 FILLER_56_260 ();
 sg13g2_decap_8 FILLER_56_267 ();
 sg13g2_decap_8 FILLER_56_274 ();
 sg13g2_decap_8 FILLER_56_281 ();
 sg13g2_decap_8 FILLER_56_288 ();
 sg13g2_decap_8 FILLER_56_295 ();
 sg13g2_decap_8 FILLER_56_302 ();
 sg13g2_decap_8 FILLER_56_309 ();
 sg13g2_decap_8 FILLER_56_316 ();
 sg13g2_decap_8 FILLER_56_323 ();
 sg13g2_decap_8 FILLER_56_330 ();
 sg13g2_decap_8 FILLER_56_337 ();
 sg13g2_decap_8 FILLER_56_344 ();
 sg13g2_decap_8 FILLER_56_351 ();
 sg13g2_decap_8 FILLER_56_358 ();
 sg13g2_decap_8 FILLER_56_365 ();
 sg13g2_decap_8 FILLER_56_372 ();
 sg13g2_decap_8 FILLER_56_379 ();
 sg13g2_decap_8 FILLER_56_386 ();
 sg13g2_decap_8 FILLER_56_393 ();
 sg13g2_decap_4 FILLER_56_400 ();
 sg13g2_fill_2 FILLER_56_407 ();
 sg13g2_decap_8 FILLER_56_420 ();
 sg13g2_decap_8 FILLER_56_427 ();
 sg13g2_decap_8 FILLER_56_434 ();
 sg13g2_decap_8 FILLER_56_441 ();
 sg13g2_decap_8 FILLER_56_448 ();
 sg13g2_decap_8 FILLER_56_455 ();
 sg13g2_decap_8 FILLER_56_462 ();
 sg13g2_decap_8 FILLER_56_469 ();
 sg13g2_decap_8 FILLER_56_476 ();
 sg13g2_decap_8 FILLER_56_483 ();
 sg13g2_decap_8 FILLER_56_490 ();
 sg13g2_decap_8 FILLER_56_497 ();
 sg13g2_decap_8 FILLER_56_504 ();
 sg13g2_decap_4 FILLER_56_511 ();
 sg13g2_fill_1 FILLER_56_515 ();
 sg13g2_decap_8 FILLER_56_531 ();
 sg13g2_decap_8 FILLER_56_538 ();
 sg13g2_decap_8 FILLER_56_545 ();
 sg13g2_decap_8 FILLER_56_557 ();
 sg13g2_decap_8 FILLER_56_564 ();
 sg13g2_decap_8 FILLER_56_571 ();
 sg13g2_fill_1 FILLER_56_578 ();
 sg13g2_decap_8 FILLER_56_584 ();
 sg13g2_decap_8 FILLER_56_591 ();
 sg13g2_fill_2 FILLER_56_598 ();
 sg13g2_fill_1 FILLER_56_600 ();
 sg13g2_decap_8 FILLER_56_611 ();
 sg13g2_decap_8 FILLER_56_618 ();
 sg13g2_decap_8 FILLER_56_625 ();
 sg13g2_decap_8 FILLER_56_632 ();
 sg13g2_decap_8 FILLER_56_639 ();
 sg13g2_decap_8 FILLER_56_646 ();
 sg13g2_decap_8 FILLER_56_653 ();
 sg13g2_decap_8 FILLER_56_660 ();
 sg13g2_decap_8 FILLER_56_667 ();
 sg13g2_fill_1 FILLER_56_674 ();
 sg13g2_fill_2 FILLER_56_680 ();
 sg13g2_decap_4 FILLER_56_694 ();
 sg13g2_decap_8 FILLER_56_713 ();
 sg13g2_decap_8 FILLER_56_720 ();
 sg13g2_decap_8 FILLER_56_727 ();
 sg13g2_fill_2 FILLER_56_734 ();
 sg13g2_decap_8 FILLER_56_741 ();
 sg13g2_decap_4 FILLER_56_748 ();
 sg13g2_decap_8 FILLER_56_756 ();
 sg13g2_decap_4 FILLER_56_763 ();
 sg13g2_fill_1 FILLER_56_767 ();
 sg13g2_decap_8 FILLER_56_771 ();
 sg13g2_decap_8 FILLER_56_778 ();
 sg13g2_decap_8 FILLER_56_785 ();
 sg13g2_decap_8 FILLER_56_792 ();
 sg13g2_decap_8 FILLER_56_799 ();
 sg13g2_decap_4 FILLER_56_806 ();
 sg13g2_fill_1 FILLER_56_810 ();
 sg13g2_fill_2 FILLER_56_814 ();
 sg13g2_fill_1 FILLER_56_816 ();
 sg13g2_decap_8 FILLER_56_832 ();
 sg13g2_decap_8 FILLER_56_839 ();
 sg13g2_decap_8 FILLER_56_846 ();
 sg13g2_decap_8 FILLER_56_853 ();
 sg13g2_decap_8 FILLER_56_860 ();
 sg13g2_fill_2 FILLER_56_867 ();
 sg13g2_fill_1 FILLER_56_869 ();
 sg13g2_decap_8 FILLER_56_874 ();
 sg13g2_decap_8 FILLER_56_881 ();
 sg13g2_decap_8 FILLER_56_888 ();
 sg13g2_decap_8 FILLER_56_895 ();
 sg13g2_decap_4 FILLER_56_902 ();
 sg13g2_decap_8 FILLER_56_921 ();
 sg13g2_decap_8 FILLER_56_928 ();
 sg13g2_decap_8 FILLER_56_935 ();
 sg13g2_decap_8 FILLER_56_942 ();
 sg13g2_decap_8 FILLER_56_949 ();
 sg13g2_decap_8 FILLER_56_956 ();
 sg13g2_decap_8 FILLER_56_963 ();
 sg13g2_decap_8 FILLER_56_970 ();
 sg13g2_decap_8 FILLER_56_977 ();
 sg13g2_decap_8 FILLER_56_984 ();
 sg13g2_decap_4 FILLER_56_991 ();
 sg13g2_fill_2 FILLER_56_995 ();
 sg13g2_decap_8 FILLER_56_1009 ();
 sg13g2_decap_8 FILLER_56_1016 ();
 sg13g2_decap_8 FILLER_56_1023 ();
 sg13g2_decap_8 FILLER_56_1030 ();
 sg13g2_decap_8 FILLER_56_1037 ();
 sg13g2_decap_8 FILLER_56_1044 ();
 sg13g2_fill_2 FILLER_56_1051 ();
 sg13g2_decap_8 FILLER_56_1063 ();
 sg13g2_decap_8 FILLER_56_1070 ();
 sg13g2_decap_8 FILLER_56_1081 ();
 sg13g2_decap_8 FILLER_56_1088 ();
 sg13g2_decap_8 FILLER_56_1095 ();
 sg13g2_fill_2 FILLER_56_1102 ();
 sg13g2_fill_1 FILLER_56_1104 ();
 sg13g2_fill_2 FILLER_56_1110 ();
 sg13g2_decap_8 FILLER_56_1127 ();
 sg13g2_decap_4 FILLER_56_1134 ();
 sg13g2_fill_1 FILLER_56_1138 ();
 sg13g2_decap_8 FILLER_56_1144 ();
 sg13g2_decap_8 FILLER_56_1151 ();
 sg13g2_decap_8 FILLER_56_1158 ();
 sg13g2_decap_4 FILLER_56_1165 ();
 sg13g2_fill_2 FILLER_56_1174 ();
 sg13g2_decap_8 FILLER_56_1179 ();
 sg13g2_decap_8 FILLER_56_1186 ();
 sg13g2_decap_4 FILLER_56_1193 ();
 sg13g2_fill_2 FILLER_56_1197 ();
 sg13g2_decap_4 FILLER_56_1214 ();
 sg13g2_fill_1 FILLER_56_1218 ();
 sg13g2_fill_2 FILLER_56_1222 ();
 sg13g2_fill_1 FILLER_56_1224 ();
 sg13g2_decap_8 FILLER_56_1240 ();
 sg13g2_decap_8 FILLER_56_1247 ();
 sg13g2_decap_8 FILLER_56_1254 ();
 sg13g2_decap_8 FILLER_56_1261 ();
 sg13g2_decap_8 FILLER_56_1268 ();
 sg13g2_decap_8 FILLER_56_1275 ();
 sg13g2_decap_8 FILLER_56_1282 ();
 sg13g2_decap_8 FILLER_56_1289 ();
 sg13g2_decap_8 FILLER_56_1296 ();
 sg13g2_fill_2 FILLER_56_1303 ();
 sg13g2_decap_8 FILLER_56_1312 ();
 sg13g2_decap_8 FILLER_56_1319 ();
 sg13g2_decap_8 FILLER_56_1326 ();
 sg13g2_decap_4 FILLER_56_1333 ();
 sg13g2_decap_8 FILLER_56_1341 ();
 sg13g2_decap_8 FILLER_56_1348 ();
 sg13g2_decap_8 FILLER_56_1355 ();
 sg13g2_decap_8 FILLER_56_1362 ();
 sg13g2_decap_8 FILLER_56_1369 ();
 sg13g2_decap_8 FILLER_56_1376 ();
 sg13g2_decap_8 FILLER_56_1383 ();
 sg13g2_decap_8 FILLER_56_1390 ();
 sg13g2_decap_8 FILLER_56_1397 ();
 sg13g2_decap_8 FILLER_56_1404 ();
 sg13g2_decap_8 FILLER_56_1411 ();
 sg13g2_decap_8 FILLER_56_1418 ();
 sg13g2_decap_8 FILLER_56_1425 ();
 sg13g2_decap_4 FILLER_56_1432 ();
 sg13g2_decap_8 FILLER_56_1440 ();
 sg13g2_decap_8 FILLER_56_1447 ();
 sg13g2_fill_2 FILLER_56_1454 ();
 sg13g2_decap_4 FILLER_56_1471 ();
 sg13g2_fill_2 FILLER_56_1475 ();
 sg13g2_fill_1 FILLER_56_1488 ();
 sg13g2_decap_8 FILLER_56_1493 ();
 sg13g2_decap_8 FILLER_56_1500 ();
 sg13g2_decap_8 FILLER_56_1507 ();
 sg13g2_decap_8 FILLER_56_1514 ();
 sg13g2_decap_8 FILLER_56_1521 ();
 sg13g2_fill_1 FILLER_56_1528 ();
 sg13g2_decap_8 FILLER_56_1544 ();
 sg13g2_decap_8 FILLER_56_1551 ();
 sg13g2_decap_8 FILLER_56_1558 ();
 sg13g2_decap_8 FILLER_56_1565 ();
 sg13g2_decap_8 FILLER_56_1572 ();
 sg13g2_decap_8 FILLER_56_1579 ();
 sg13g2_decap_8 FILLER_56_1586 ();
 sg13g2_decap_8 FILLER_56_1593 ();
 sg13g2_decap_8 FILLER_56_1600 ();
 sg13g2_decap_8 FILLER_56_1607 ();
 sg13g2_decap_8 FILLER_56_1614 ();
 sg13g2_decap_8 FILLER_56_1621 ();
 sg13g2_decap_4 FILLER_56_1628 ();
 sg13g2_decap_8 FILLER_56_1647 ();
 sg13g2_decap_8 FILLER_56_1654 ();
 sg13g2_decap_8 FILLER_56_1661 ();
 sg13g2_decap_8 FILLER_56_1668 ();
 sg13g2_decap_8 FILLER_56_1675 ();
 sg13g2_decap_8 FILLER_56_1682 ();
 sg13g2_decap_8 FILLER_56_1689 ();
 sg13g2_decap_8 FILLER_56_1696 ();
 sg13g2_decap_8 FILLER_56_1703 ();
 sg13g2_decap_8 FILLER_56_1710 ();
 sg13g2_decap_8 FILLER_56_1717 ();
 sg13g2_decap_8 FILLER_56_1724 ();
 sg13g2_decap_8 FILLER_56_1731 ();
 sg13g2_decap_8 FILLER_56_1738 ();
 sg13g2_fill_2 FILLER_56_1745 ();
 sg13g2_fill_1 FILLER_56_1747 ();
 sg13g2_decap_8 FILLER_56_1751 ();
 sg13g2_decap_8 FILLER_56_1758 ();
 sg13g2_decap_8 FILLER_56_1765 ();
 sg13g2_decap_8 FILLER_56_1772 ();
 sg13g2_decap_8 FILLER_56_1779 ();
 sg13g2_decap_8 FILLER_56_1786 ();
 sg13g2_decap_8 FILLER_56_1793 ();
 sg13g2_decap_8 FILLER_56_1800 ();
 sg13g2_decap_8 FILLER_56_1807 ();
 sg13g2_decap_8 FILLER_56_1814 ();
 sg13g2_decap_8 FILLER_56_1821 ();
 sg13g2_decap_8 FILLER_56_1828 ();
 sg13g2_decap_8 FILLER_56_1835 ();
 sg13g2_decap_8 FILLER_56_1842 ();
 sg13g2_decap_4 FILLER_56_1849 ();
 sg13g2_decap_8 FILLER_56_1856 ();
 sg13g2_decap_8 FILLER_56_1863 ();
 sg13g2_decap_8 FILLER_56_1870 ();
 sg13g2_decap_8 FILLER_56_1877 ();
 sg13g2_decap_8 FILLER_56_1884 ();
 sg13g2_decap_8 FILLER_56_1891 ();
 sg13g2_decap_8 FILLER_56_1898 ();
 sg13g2_decap_8 FILLER_56_1905 ();
 sg13g2_decap_8 FILLER_56_1912 ();
 sg13g2_decap_8 FILLER_56_1919 ();
 sg13g2_decap_8 FILLER_56_1926 ();
 sg13g2_decap_8 FILLER_56_1933 ();
 sg13g2_decap_8 FILLER_56_1940 ();
 sg13g2_decap_8 FILLER_56_1947 ();
 sg13g2_decap_8 FILLER_56_1954 ();
 sg13g2_decap_8 FILLER_56_1961 ();
 sg13g2_decap_8 FILLER_56_1968 ();
 sg13g2_decap_8 FILLER_56_1975 ();
 sg13g2_decap_8 FILLER_56_1982 ();
 sg13g2_decap_8 FILLER_56_1989 ();
 sg13g2_fill_2 FILLER_56_2022 ();
 sg13g2_fill_1 FILLER_56_2024 ();
 sg13g2_decap_8 FILLER_56_2029 ();
 sg13g2_decap_8 FILLER_56_2036 ();
 sg13g2_decap_8 FILLER_56_2043 ();
 sg13g2_decap_8 FILLER_56_2050 ();
 sg13g2_decap_8 FILLER_56_2057 ();
 sg13g2_decap_8 FILLER_56_2064 ();
 sg13g2_decap_8 FILLER_56_2071 ();
 sg13g2_decap_8 FILLER_56_2078 ();
 sg13g2_decap_8 FILLER_56_2085 ();
 sg13g2_decap_8 FILLER_56_2092 ();
 sg13g2_decap_8 FILLER_56_2099 ();
 sg13g2_decap_8 FILLER_56_2106 ();
 sg13g2_decap_8 FILLER_56_2113 ();
 sg13g2_decap_8 FILLER_56_2120 ();
 sg13g2_decap_8 FILLER_56_2127 ();
 sg13g2_decap_8 FILLER_56_2134 ();
 sg13g2_decap_8 FILLER_56_2141 ();
 sg13g2_decap_8 FILLER_56_2148 ();
 sg13g2_decap_8 FILLER_56_2155 ();
 sg13g2_fill_2 FILLER_56_2162 ();
 sg13g2_fill_1 FILLER_56_2164 ();
 sg13g2_fill_1 FILLER_56_2170 ();
 sg13g2_decap_8 FILLER_56_2174 ();
 sg13g2_decap_4 FILLER_56_2181 ();
 sg13g2_fill_2 FILLER_56_2185 ();
 sg13g2_decap_4 FILLER_56_2192 ();
 sg13g2_fill_1 FILLER_56_2196 ();
 sg13g2_decap_8 FILLER_56_2200 ();
 sg13g2_decap_8 FILLER_56_2207 ();
 sg13g2_decap_8 FILLER_56_2214 ();
 sg13g2_decap_8 FILLER_56_2221 ();
 sg13g2_decap_8 FILLER_56_2228 ();
 sg13g2_decap_8 FILLER_56_2235 ();
 sg13g2_decap_8 FILLER_56_2242 ();
 sg13g2_decap_8 FILLER_56_2249 ();
 sg13g2_decap_8 FILLER_56_2256 ();
 sg13g2_decap_8 FILLER_56_2263 ();
 sg13g2_decap_8 FILLER_56_2270 ();
 sg13g2_decap_8 FILLER_56_2277 ();
 sg13g2_decap_8 FILLER_56_2284 ();
 sg13g2_decap_8 FILLER_56_2291 ();
 sg13g2_decap_8 FILLER_56_2298 ();
 sg13g2_decap_8 FILLER_56_2305 ();
 sg13g2_decap_8 FILLER_56_2312 ();
 sg13g2_decap_8 FILLER_56_2319 ();
 sg13g2_decap_8 FILLER_56_2326 ();
 sg13g2_decap_8 FILLER_56_2333 ();
 sg13g2_decap_8 FILLER_56_2340 ();
 sg13g2_decap_8 FILLER_56_2347 ();
 sg13g2_decap_8 FILLER_56_2354 ();
 sg13g2_decap_8 FILLER_56_2361 ();
 sg13g2_decap_8 FILLER_56_2368 ();
 sg13g2_decap_8 FILLER_56_2375 ();
 sg13g2_decap_8 FILLER_56_2382 ();
 sg13g2_decap_8 FILLER_56_2389 ();
 sg13g2_decap_8 FILLER_56_2396 ();
 sg13g2_decap_8 FILLER_56_2403 ();
 sg13g2_decap_8 FILLER_56_2410 ();
 sg13g2_decap_8 FILLER_56_2417 ();
 sg13g2_decap_8 FILLER_56_2424 ();
 sg13g2_decap_8 FILLER_56_2431 ();
 sg13g2_decap_8 FILLER_56_2438 ();
 sg13g2_decap_8 FILLER_56_2445 ();
 sg13g2_decap_8 FILLER_56_2452 ();
 sg13g2_decap_8 FILLER_56_2459 ();
 sg13g2_decap_8 FILLER_56_2466 ();
 sg13g2_decap_8 FILLER_56_2473 ();
 sg13g2_decap_8 FILLER_56_2480 ();
 sg13g2_decap_8 FILLER_56_2487 ();
 sg13g2_decap_8 FILLER_56_2494 ();
 sg13g2_decap_8 FILLER_56_2501 ();
 sg13g2_decap_8 FILLER_56_2508 ();
 sg13g2_decap_8 FILLER_56_2515 ();
 sg13g2_decap_8 FILLER_56_2522 ();
 sg13g2_decap_8 FILLER_56_2529 ();
 sg13g2_decap_8 FILLER_56_2536 ();
 sg13g2_decap_8 FILLER_56_2543 ();
 sg13g2_decap_8 FILLER_56_2550 ();
 sg13g2_decap_8 FILLER_56_2557 ();
 sg13g2_decap_8 FILLER_56_2564 ();
 sg13g2_decap_8 FILLER_56_2571 ();
 sg13g2_decap_8 FILLER_56_2578 ();
 sg13g2_decap_8 FILLER_56_2585 ();
 sg13g2_decap_8 FILLER_56_2592 ();
 sg13g2_decap_8 FILLER_56_2599 ();
 sg13g2_decap_8 FILLER_56_2606 ();
 sg13g2_decap_8 FILLER_56_2613 ();
 sg13g2_decap_8 FILLER_56_2620 ();
 sg13g2_decap_8 FILLER_56_2627 ();
 sg13g2_decap_8 FILLER_56_2634 ();
 sg13g2_decap_8 FILLER_56_2641 ();
 sg13g2_decap_8 FILLER_56_2648 ();
 sg13g2_decap_8 FILLER_56_2655 ();
 sg13g2_decap_8 FILLER_56_2662 ();
 sg13g2_fill_1 FILLER_56_2669 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_fill_2 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_65 ();
 sg13g2_decap_8 FILLER_57_72 ();
 sg13g2_fill_2 FILLER_57_79 ();
 sg13g2_decap_8 FILLER_57_87 ();
 sg13g2_decap_8 FILLER_57_94 ();
 sg13g2_decap_8 FILLER_57_101 ();
 sg13g2_decap_8 FILLER_57_108 ();
 sg13g2_decap_8 FILLER_57_115 ();
 sg13g2_decap_8 FILLER_57_122 ();
 sg13g2_decap_8 FILLER_57_129 ();
 sg13g2_decap_4 FILLER_57_140 ();
 sg13g2_fill_1 FILLER_57_144 ();
 sg13g2_decap_8 FILLER_57_150 ();
 sg13g2_decap_8 FILLER_57_157 ();
 sg13g2_fill_1 FILLER_57_164 ();
 sg13g2_decap_8 FILLER_57_170 ();
 sg13g2_decap_8 FILLER_57_177 ();
 sg13g2_decap_8 FILLER_57_184 ();
 sg13g2_decap_8 FILLER_57_191 ();
 sg13g2_decap_8 FILLER_57_198 ();
 sg13g2_decap_8 FILLER_57_205 ();
 sg13g2_decap_8 FILLER_57_212 ();
 sg13g2_decap_8 FILLER_57_219 ();
 sg13g2_decap_8 FILLER_57_226 ();
 sg13g2_decap_8 FILLER_57_233 ();
 sg13g2_fill_1 FILLER_57_240 ();
 sg13g2_decap_8 FILLER_57_267 ();
 sg13g2_decap_8 FILLER_57_274 ();
 sg13g2_decap_8 FILLER_57_281 ();
 sg13g2_decap_8 FILLER_57_288 ();
 sg13g2_decap_8 FILLER_57_295 ();
 sg13g2_decap_8 FILLER_57_302 ();
 sg13g2_decap_8 FILLER_57_309 ();
 sg13g2_decap_8 FILLER_57_316 ();
 sg13g2_decap_8 FILLER_57_323 ();
 sg13g2_decap_8 FILLER_57_330 ();
 sg13g2_fill_2 FILLER_57_337 ();
 sg13g2_decap_8 FILLER_57_344 ();
 sg13g2_decap_8 FILLER_57_351 ();
 sg13g2_decap_8 FILLER_57_358 ();
 sg13g2_decap_8 FILLER_57_365 ();
 sg13g2_decap_8 FILLER_57_372 ();
 sg13g2_fill_2 FILLER_57_379 ();
 sg13g2_fill_2 FILLER_57_388 ();
 sg13g2_fill_2 FILLER_57_407 ();
 sg13g2_decap_8 FILLER_57_416 ();
 sg13g2_decap_8 FILLER_57_423 ();
 sg13g2_decap_8 FILLER_57_430 ();
 sg13g2_decap_8 FILLER_57_437 ();
 sg13g2_fill_2 FILLER_57_444 ();
 sg13g2_fill_1 FILLER_57_446 ();
 sg13g2_decap_8 FILLER_57_457 ();
 sg13g2_decap_8 FILLER_57_464 ();
 sg13g2_decap_8 FILLER_57_471 ();
 sg13g2_decap_8 FILLER_57_478 ();
 sg13g2_decap_8 FILLER_57_485 ();
 sg13g2_decap_8 FILLER_57_492 ();
 sg13g2_decap_8 FILLER_57_499 ();
 sg13g2_decap_8 FILLER_57_506 ();
 sg13g2_decap_4 FILLER_57_513 ();
 sg13g2_fill_2 FILLER_57_517 ();
 sg13g2_decap_8 FILLER_57_525 ();
 sg13g2_decap_8 FILLER_57_532 ();
 sg13g2_decap_8 FILLER_57_539 ();
 sg13g2_decap_8 FILLER_57_546 ();
 sg13g2_decap_8 FILLER_57_553 ();
 sg13g2_decap_8 FILLER_57_560 ();
 sg13g2_decap_8 FILLER_57_567 ();
 sg13g2_decap_4 FILLER_57_574 ();
 sg13g2_fill_1 FILLER_57_578 ();
 sg13g2_decap_8 FILLER_57_586 ();
 sg13g2_decap_8 FILLER_57_593 ();
 sg13g2_decap_8 FILLER_57_600 ();
 sg13g2_decap_8 FILLER_57_607 ();
 sg13g2_decap_8 FILLER_57_614 ();
 sg13g2_decap_8 FILLER_57_621 ();
 sg13g2_decap_8 FILLER_57_628 ();
 sg13g2_decap_8 FILLER_57_635 ();
 sg13g2_decap_8 FILLER_57_642 ();
 sg13g2_fill_2 FILLER_57_649 ();
 sg13g2_fill_1 FILLER_57_651 ();
 sg13g2_decap_8 FILLER_57_657 ();
 sg13g2_fill_2 FILLER_57_664 ();
 sg13g2_fill_1 FILLER_57_681 ();
 sg13g2_decap_8 FILLER_57_685 ();
 sg13g2_decap_4 FILLER_57_692 ();
 sg13g2_fill_2 FILLER_57_696 ();
 sg13g2_decap_8 FILLER_57_713 ();
 sg13g2_decap_8 FILLER_57_720 ();
 sg13g2_decap_8 FILLER_57_727 ();
 sg13g2_decap_8 FILLER_57_734 ();
 sg13g2_decap_8 FILLER_57_741 ();
 sg13g2_decap_8 FILLER_57_748 ();
 sg13g2_decap_8 FILLER_57_755 ();
 sg13g2_decap_8 FILLER_57_762 ();
 sg13g2_decap_8 FILLER_57_769 ();
 sg13g2_decap_8 FILLER_57_776 ();
 sg13g2_decap_4 FILLER_57_783 ();
 sg13g2_fill_2 FILLER_57_790 ();
 sg13g2_fill_1 FILLER_57_792 ();
 sg13g2_decap_8 FILLER_57_834 ();
 sg13g2_decap_8 FILLER_57_841 ();
 sg13g2_decap_8 FILLER_57_848 ();
 sg13g2_decap_8 FILLER_57_855 ();
 sg13g2_decap_8 FILLER_57_862 ();
 sg13g2_fill_1 FILLER_57_869 ();
 sg13g2_decap_8 FILLER_57_873 ();
 sg13g2_decap_4 FILLER_57_880 ();
 sg13g2_decap_8 FILLER_57_887 ();
 sg13g2_decap_8 FILLER_57_894 ();
 sg13g2_decap_8 FILLER_57_901 ();
 sg13g2_fill_1 FILLER_57_908 ();
 sg13g2_decap_8 FILLER_57_915 ();
 sg13g2_decap_8 FILLER_57_922 ();
 sg13g2_decap_8 FILLER_57_929 ();
 sg13g2_decap_8 FILLER_57_936 ();
 sg13g2_decap_8 FILLER_57_943 ();
 sg13g2_decap_8 FILLER_57_950 ();
 sg13g2_decap_8 FILLER_57_957 ();
 sg13g2_decap_8 FILLER_57_964 ();
 sg13g2_decap_8 FILLER_57_971 ();
 sg13g2_decap_8 FILLER_57_978 ();
 sg13g2_decap_8 FILLER_57_985 ();
 sg13g2_fill_2 FILLER_57_992 ();
 sg13g2_decap_8 FILLER_57_1007 ();
 sg13g2_decap_8 FILLER_57_1014 ();
 sg13g2_decap_8 FILLER_57_1021 ();
 sg13g2_decap_8 FILLER_57_1058 ();
 sg13g2_decap_8 FILLER_57_1065 ();
 sg13g2_decap_8 FILLER_57_1072 ();
 sg13g2_decap_8 FILLER_57_1079 ();
 sg13g2_decap_8 FILLER_57_1086 ();
 sg13g2_decap_8 FILLER_57_1093 ();
 sg13g2_decap_8 FILLER_57_1100 ();
 sg13g2_decap_8 FILLER_57_1107 ();
 sg13g2_fill_1 FILLER_57_1114 ();
 sg13g2_decap_8 FILLER_57_1123 ();
 sg13g2_decap_8 FILLER_57_1130 ();
 sg13g2_decap_8 FILLER_57_1137 ();
 sg13g2_decap_8 FILLER_57_1144 ();
 sg13g2_decap_8 FILLER_57_1151 ();
 sg13g2_decap_8 FILLER_57_1158 ();
 sg13g2_decap_8 FILLER_57_1165 ();
 sg13g2_fill_1 FILLER_57_1172 ();
 sg13g2_decap_8 FILLER_57_1181 ();
 sg13g2_decap_8 FILLER_57_1188 ();
 sg13g2_fill_1 FILLER_57_1195 ();
 sg13g2_fill_2 FILLER_57_1210 ();
 sg13g2_fill_1 FILLER_57_1212 ();
 sg13g2_decap_8 FILLER_57_1236 ();
 sg13g2_decap_8 FILLER_57_1243 ();
 sg13g2_decap_8 FILLER_57_1250 ();
 sg13g2_decap_8 FILLER_57_1257 ();
 sg13g2_fill_1 FILLER_57_1264 ();
 sg13g2_decap_8 FILLER_57_1280 ();
 sg13g2_decap_8 FILLER_57_1287 ();
 sg13g2_decap_8 FILLER_57_1294 ();
 sg13g2_fill_2 FILLER_57_1301 ();
 sg13g2_fill_2 FILLER_57_1311 ();
 sg13g2_fill_1 FILLER_57_1318 ();
 sg13g2_decap_8 FILLER_57_1324 ();
 sg13g2_decap_8 FILLER_57_1331 ();
 sg13g2_decap_8 FILLER_57_1338 ();
 sg13g2_decap_8 FILLER_57_1345 ();
 sg13g2_decap_8 FILLER_57_1352 ();
 sg13g2_decap_8 FILLER_57_1359 ();
 sg13g2_decap_8 FILLER_57_1366 ();
 sg13g2_decap_4 FILLER_57_1373 ();
 sg13g2_fill_2 FILLER_57_1377 ();
 sg13g2_decap_8 FILLER_57_1383 ();
 sg13g2_decap_8 FILLER_57_1390 ();
 sg13g2_decap_8 FILLER_57_1397 ();
 sg13g2_decap_8 FILLER_57_1404 ();
 sg13g2_decap_8 FILLER_57_1411 ();
 sg13g2_decap_8 FILLER_57_1418 ();
 sg13g2_decap_8 FILLER_57_1425 ();
 sg13g2_decap_8 FILLER_57_1432 ();
 sg13g2_decap_8 FILLER_57_1439 ();
 sg13g2_decap_8 FILLER_57_1446 ();
 sg13g2_fill_2 FILLER_57_1453 ();
 sg13g2_fill_1 FILLER_57_1455 ();
 sg13g2_decap_8 FILLER_57_1460 ();
 sg13g2_decap_8 FILLER_57_1467 ();
 sg13g2_fill_2 FILLER_57_1474 ();
 sg13g2_fill_1 FILLER_57_1476 ();
 sg13g2_decap_8 FILLER_57_1481 ();
 sg13g2_decap_8 FILLER_57_1488 ();
 sg13g2_decap_8 FILLER_57_1495 ();
 sg13g2_decap_8 FILLER_57_1502 ();
 sg13g2_decap_8 FILLER_57_1509 ();
 sg13g2_decap_8 FILLER_57_1516 ();
 sg13g2_decap_8 FILLER_57_1523 ();
 sg13g2_decap_8 FILLER_57_1530 ();
 sg13g2_decap_8 FILLER_57_1537 ();
 sg13g2_decap_8 FILLER_57_1544 ();
 sg13g2_decap_8 FILLER_57_1551 ();
 sg13g2_decap_8 FILLER_57_1558 ();
 sg13g2_decap_4 FILLER_57_1565 ();
 sg13g2_decap_8 FILLER_57_1574 ();
 sg13g2_decap_8 FILLER_57_1581 ();
 sg13g2_decap_8 FILLER_57_1588 ();
 sg13g2_decap_8 FILLER_57_1595 ();
 sg13g2_decap_8 FILLER_57_1602 ();
 sg13g2_decap_4 FILLER_57_1609 ();
 sg13g2_fill_1 FILLER_57_1613 ();
 sg13g2_fill_2 FILLER_57_1629 ();
 sg13g2_fill_1 FILLER_57_1631 ();
 sg13g2_decap_8 FILLER_57_1637 ();
 sg13g2_decap_8 FILLER_57_1644 ();
 sg13g2_decap_8 FILLER_57_1651 ();
 sg13g2_decap_8 FILLER_57_1658 ();
 sg13g2_decap_4 FILLER_57_1665 ();
 sg13g2_fill_1 FILLER_57_1669 ();
 sg13g2_decap_8 FILLER_57_1685 ();
 sg13g2_decap_8 FILLER_57_1692 ();
 sg13g2_decap_8 FILLER_57_1699 ();
 sg13g2_decap_8 FILLER_57_1706 ();
 sg13g2_decap_8 FILLER_57_1713 ();
 sg13g2_decap_8 FILLER_57_1720 ();
 sg13g2_decap_8 FILLER_57_1727 ();
 sg13g2_fill_2 FILLER_57_1734 ();
 sg13g2_decap_4 FILLER_57_1744 ();
 sg13g2_decap_8 FILLER_57_1753 ();
 sg13g2_decap_8 FILLER_57_1760 ();
 sg13g2_decap_8 FILLER_57_1767 ();
 sg13g2_decap_8 FILLER_57_1774 ();
 sg13g2_decap_8 FILLER_57_1781 ();
 sg13g2_decap_8 FILLER_57_1788 ();
 sg13g2_decap_8 FILLER_57_1795 ();
 sg13g2_decap_8 FILLER_57_1802 ();
 sg13g2_decap_8 FILLER_57_1809 ();
 sg13g2_fill_2 FILLER_57_1816 ();
 sg13g2_fill_1 FILLER_57_1818 ();
 sg13g2_decap_8 FILLER_57_1824 ();
 sg13g2_decap_8 FILLER_57_1831 ();
 sg13g2_fill_1 FILLER_57_1838 ();
 sg13g2_decap_4 FILLER_57_1849 ();
 sg13g2_decap_8 FILLER_57_1857 ();
 sg13g2_decap_8 FILLER_57_1864 ();
 sg13g2_decap_8 FILLER_57_1871 ();
 sg13g2_decap_8 FILLER_57_1878 ();
 sg13g2_decap_8 FILLER_57_1885 ();
 sg13g2_decap_8 FILLER_57_1892 ();
 sg13g2_decap_8 FILLER_57_1899 ();
 sg13g2_decap_8 FILLER_57_1906 ();
 sg13g2_decap_8 FILLER_57_1913 ();
 sg13g2_decap_8 FILLER_57_1920 ();
 sg13g2_decap_8 FILLER_57_1927 ();
 sg13g2_decap_8 FILLER_57_1934 ();
 sg13g2_decap_8 FILLER_57_1941 ();
 sg13g2_decap_8 FILLER_57_1948 ();
 sg13g2_decap_8 FILLER_57_1955 ();
 sg13g2_fill_2 FILLER_57_1962 ();
 sg13g2_decap_8 FILLER_57_1968 ();
 sg13g2_decap_8 FILLER_57_1975 ();
 sg13g2_decap_8 FILLER_57_1982 ();
 sg13g2_decap_8 FILLER_57_1989 ();
 sg13g2_decap_4 FILLER_57_1996 ();
 sg13g2_decap_8 FILLER_57_2004 ();
 sg13g2_decap_8 FILLER_57_2011 ();
 sg13g2_decap_8 FILLER_57_2018 ();
 sg13g2_decap_4 FILLER_57_2025 ();
 sg13g2_decap_8 FILLER_57_2032 ();
 sg13g2_decap_8 FILLER_57_2039 ();
 sg13g2_decap_8 FILLER_57_2046 ();
 sg13g2_decap_8 FILLER_57_2053 ();
 sg13g2_decap_8 FILLER_57_2060 ();
 sg13g2_decap_8 FILLER_57_2067 ();
 sg13g2_decap_8 FILLER_57_2074 ();
 sg13g2_decap_8 FILLER_57_2081 ();
 sg13g2_decap_8 FILLER_57_2088 ();
 sg13g2_decap_8 FILLER_57_2095 ();
 sg13g2_decap_8 FILLER_57_2102 ();
 sg13g2_decap_8 FILLER_57_2109 ();
 sg13g2_decap_8 FILLER_57_2116 ();
 sg13g2_decap_8 FILLER_57_2123 ();
 sg13g2_decap_8 FILLER_57_2130 ();
 sg13g2_decap_8 FILLER_57_2137 ();
 sg13g2_decap_8 FILLER_57_2144 ();
 sg13g2_decap_8 FILLER_57_2151 ();
 sg13g2_decap_8 FILLER_57_2158 ();
 sg13g2_decap_8 FILLER_57_2169 ();
 sg13g2_decap_8 FILLER_57_2176 ();
 sg13g2_decap_8 FILLER_57_2183 ();
 sg13g2_decap_8 FILLER_57_2190 ();
 sg13g2_decap_8 FILLER_57_2202 ();
 sg13g2_decap_8 FILLER_57_2209 ();
 sg13g2_decap_8 FILLER_57_2216 ();
 sg13g2_decap_8 FILLER_57_2223 ();
 sg13g2_decap_8 FILLER_57_2230 ();
 sg13g2_decap_8 FILLER_57_2237 ();
 sg13g2_decap_8 FILLER_57_2244 ();
 sg13g2_decap_8 FILLER_57_2251 ();
 sg13g2_decap_8 FILLER_57_2258 ();
 sg13g2_decap_8 FILLER_57_2265 ();
 sg13g2_decap_8 FILLER_57_2272 ();
 sg13g2_decap_8 FILLER_57_2279 ();
 sg13g2_decap_8 FILLER_57_2286 ();
 sg13g2_decap_8 FILLER_57_2293 ();
 sg13g2_decap_8 FILLER_57_2300 ();
 sg13g2_decap_8 FILLER_57_2307 ();
 sg13g2_decap_8 FILLER_57_2314 ();
 sg13g2_decap_8 FILLER_57_2321 ();
 sg13g2_decap_8 FILLER_57_2328 ();
 sg13g2_decap_8 FILLER_57_2335 ();
 sg13g2_decap_8 FILLER_57_2342 ();
 sg13g2_decap_8 FILLER_57_2349 ();
 sg13g2_decap_8 FILLER_57_2356 ();
 sg13g2_decap_8 FILLER_57_2363 ();
 sg13g2_decap_8 FILLER_57_2370 ();
 sg13g2_decap_8 FILLER_57_2377 ();
 sg13g2_decap_8 FILLER_57_2384 ();
 sg13g2_decap_8 FILLER_57_2391 ();
 sg13g2_decap_8 FILLER_57_2398 ();
 sg13g2_decap_8 FILLER_57_2405 ();
 sg13g2_decap_8 FILLER_57_2412 ();
 sg13g2_decap_8 FILLER_57_2419 ();
 sg13g2_decap_8 FILLER_57_2426 ();
 sg13g2_decap_8 FILLER_57_2433 ();
 sg13g2_decap_8 FILLER_57_2440 ();
 sg13g2_decap_8 FILLER_57_2447 ();
 sg13g2_decap_8 FILLER_57_2454 ();
 sg13g2_decap_8 FILLER_57_2461 ();
 sg13g2_decap_8 FILLER_57_2468 ();
 sg13g2_decap_8 FILLER_57_2475 ();
 sg13g2_decap_8 FILLER_57_2482 ();
 sg13g2_decap_8 FILLER_57_2489 ();
 sg13g2_decap_8 FILLER_57_2496 ();
 sg13g2_decap_8 FILLER_57_2503 ();
 sg13g2_decap_8 FILLER_57_2510 ();
 sg13g2_decap_8 FILLER_57_2517 ();
 sg13g2_decap_8 FILLER_57_2524 ();
 sg13g2_decap_8 FILLER_57_2531 ();
 sg13g2_decap_8 FILLER_57_2538 ();
 sg13g2_decap_8 FILLER_57_2545 ();
 sg13g2_decap_8 FILLER_57_2552 ();
 sg13g2_decap_8 FILLER_57_2559 ();
 sg13g2_decap_8 FILLER_57_2566 ();
 sg13g2_decap_8 FILLER_57_2573 ();
 sg13g2_decap_8 FILLER_57_2580 ();
 sg13g2_decap_8 FILLER_57_2587 ();
 sg13g2_decap_8 FILLER_57_2594 ();
 sg13g2_decap_8 FILLER_57_2601 ();
 sg13g2_decap_8 FILLER_57_2608 ();
 sg13g2_decap_8 FILLER_57_2615 ();
 sg13g2_decap_8 FILLER_57_2622 ();
 sg13g2_decap_8 FILLER_57_2629 ();
 sg13g2_decap_8 FILLER_57_2636 ();
 sg13g2_decap_8 FILLER_57_2643 ();
 sg13g2_decap_8 FILLER_57_2650 ();
 sg13g2_decap_8 FILLER_57_2657 ();
 sg13g2_decap_4 FILLER_57_2664 ();
 sg13g2_fill_2 FILLER_57_2668 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_4 FILLER_58_42 ();
 sg13g2_fill_1 FILLER_58_46 ();
 sg13g2_decap_8 FILLER_58_52 ();
 sg13g2_decap_8 FILLER_58_59 ();
 sg13g2_decap_8 FILLER_58_66 ();
 sg13g2_decap_8 FILLER_58_73 ();
 sg13g2_decap_8 FILLER_58_80 ();
 sg13g2_decap_4 FILLER_58_87 ();
 sg13g2_fill_1 FILLER_58_91 ();
 sg13g2_decap_8 FILLER_58_96 ();
 sg13g2_fill_1 FILLER_58_103 ();
 sg13g2_decap_8 FILLER_58_117 ();
 sg13g2_decap_8 FILLER_58_124 ();
 sg13g2_decap_8 FILLER_58_131 ();
 sg13g2_decap_8 FILLER_58_138 ();
 sg13g2_decap_8 FILLER_58_145 ();
 sg13g2_decap_8 FILLER_58_152 ();
 sg13g2_decap_8 FILLER_58_159 ();
 sg13g2_decap_8 FILLER_58_166 ();
 sg13g2_decap_8 FILLER_58_173 ();
 sg13g2_decap_8 FILLER_58_180 ();
 sg13g2_decap_8 FILLER_58_187 ();
 sg13g2_decap_8 FILLER_58_194 ();
 sg13g2_decap_8 FILLER_58_201 ();
 sg13g2_decap_8 FILLER_58_208 ();
 sg13g2_decap_4 FILLER_58_215 ();
 sg13g2_fill_2 FILLER_58_219 ();
 sg13g2_decap_8 FILLER_58_229 ();
 sg13g2_decap_8 FILLER_58_236 ();
 sg13g2_decap_4 FILLER_58_243 ();
 sg13g2_fill_2 FILLER_58_247 ();
 sg13g2_decap_8 FILLER_58_253 ();
 sg13g2_decap_8 FILLER_58_260 ();
 sg13g2_decap_8 FILLER_58_267 ();
 sg13g2_decap_8 FILLER_58_274 ();
 sg13g2_decap_8 FILLER_58_281 ();
 sg13g2_decap_8 FILLER_58_288 ();
 sg13g2_decap_8 FILLER_58_295 ();
 sg13g2_decap_8 FILLER_58_302 ();
 sg13g2_decap_8 FILLER_58_309 ();
 sg13g2_decap_8 FILLER_58_316 ();
 sg13g2_decap_8 FILLER_58_323 ();
 sg13g2_decap_8 FILLER_58_330 ();
 sg13g2_decap_8 FILLER_58_337 ();
 sg13g2_decap_8 FILLER_58_344 ();
 sg13g2_decap_8 FILLER_58_351 ();
 sg13g2_decap_8 FILLER_58_358 ();
 sg13g2_decap_8 FILLER_58_365 ();
 sg13g2_decap_8 FILLER_58_372 ();
 sg13g2_fill_2 FILLER_58_379 ();
 sg13g2_decap_8 FILLER_58_385 ();
 sg13g2_decap_8 FILLER_58_412 ();
 sg13g2_decap_8 FILLER_58_419 ();
 sg13g2_decap_8 FILLER_58_426 ();
 sg13g2_fill_2 FILLER_58_433 ();
 sg13g2_fill_1 FILLER_58_435 ();
 sg13g2_decap_8 FILLER_58_459 ();
 sg13g2_decap_8 FILLER_58_466 ();
 sg13g2_decap_8 FILLER_58_473 ();
 sg13g2_decap_4 FILLER_58_480 ();
 sg13g2_fill_1 FILLER_58_484 ();
 sg13g2_decap_8 FILLER_58_495 ();
 sg13g2_decap_8 FILLER_58_502 ();
 sg13g2_decap_8 FILLER_58_509 ();
 sg13g2_fill_2 FILLER_58_519 ();
 sg13g2_decap_8 FILLER_58_524 ();
 sg13g2_decap_8 FILLER_58_531 ();
 sg13g2_decap_8 FILLER_58_538 ();
 sg13g2_decap_8 FILLER_58_545 ();
 sg13g2_decap_8 FILLER_58_552 ();
 sg13g2_fill_1 FILLER_58_559 ();
 sg13g2_fill_2 FILLER_58_575 ();
 sg13g2_fill_1 FILLER_58_577 ();
 sg13g2_decap_8 FILLER_58_593 ();
 sg13g2_decap_8 FILLER_58_600 ();
 sg13g2_decap_8 FILLER_58_607 ();
 sg13g2_decap_8 FILLER_58_614 ();
 sg13g2_decap_8 FILLER_58_621 ();
 sg13g2_decap_8 FILLER_58_628 ();
 sg13g2_decap_8 FILLER_58_635 ();
 sg13g2_decap_8 FILLER_58_642 ();
 sg13g2_decap_8 FILLER_58_649 ();
 sg13g2_decap_4 FILLER_58_656 ();
 sg13g2_fill_2 FILLER_58_660 ();
 sg13g2_fill_1 FILLER_58_667 ();
 sg13g2_decap_8 FILLER_58_684 ();
 sg13g2_decap_8 FILLER_58_691 ();
 sg13g2_fill_2 FILLER_58_698 ();
 sg13g2_fill_1 FILLER_58_700 ();
 sg13g2_decap_8 FILLER_58_706 ();
 sg13g2_decap_8 FILLER_58_713 ();
 sg13g2_decap_8 FILLER_58_720 ();
 sg13g2_decap_8 FILLER_58_727 ();
 sg13g2_decap_8 FILLER_58_734 ();
 sg13g2_fill_1 FILLER_58_741 ();
 sg13g2_fill_1 FILLER_58_748 ();
 sg13g2_fill_1 FILLER_58_752 ();
 sg13g2_fill_2 FILLER_58_765 ();
 sg13g2_fill_1 FILLER_58_767 ();
 sg13g2_decap_4 FILLER_58_791 ();
 sg13g2_fill_1 FILLER_58_795 ();
 sg13g2_fill_2 FILLER_58_808 ();
 sg13g2_fill_1 FILLER_58_817 ();
 sg13g2_decap_8 FILLER_58_828 ();
 sg13g2_decap_8 FILLER_58_835 ();
 sg13g2_decap_8 FILLER_58_842 ();
 sg13g2_decap_8 FILLER_58_849 ();
 sg13g2_decap_8 FILLER_58_856 ();
 sg13g2_decap_8 FILLER_58_863 ();
 sg13g2_decap_8 FILLER_58_870 ();
 sg13g2_decap_4 FILLER_58_877 ();
 sg13g2_decap_8 FILLER_58_888 ();
 sg13g2_fill_1 FILLER_58_895 ();
 sg13g2_fill_1 FILLER_58_908 ();
 sg13g2_decap_8 FILLER_58_915 ();
 sg13g2_decap_8 FILLER_58_922 ();
 sg13g2_fill_1 FILLER_58_929 ();
 sg13g2_decap_8 FILLER_58_948 ();
 sg13g2_decap_8 FILLER_58_955 ();
 sg13g2_decap_4 FILLER_58_962 ();
 sg13g2_fill_2 FILLER_58_966 ();
 sg13g2_decap_8 FILLER_58_1007 ();
 sg13g2_decap_8 FILLER_58_1014 ();
 sg13g2_decap_8 FILLER_58_1021 ();
 sg13g2_decap_4 FILLER_58_1028 ();
 sg13g2_fill_2 FILLER_58_1032 ();
 sg13g2_fill_1 FILLER_58_1039 ();
 sg13g2_decap_8 FILLER_58_1051 ();
 sg13g2_decap_8 FILLER_58_1058 ();
 sg13g2_decap_8 FILLER_58_1065 ();
 sg13g2_decap_8 FILLER_58_1072 ();
 sg13g2_decap_8 FILLER_58_1079 ();
 sg13g2_decap_8 FILLER_58_1086 ();
 sg13g2_decap_8 FILLER_58_1093 ();
 sg13g2_decap_8 FILLER_58_1100 ();
 sg13g2_decap_8 FILLER_58_1107 ();
 sg13g2_decap_8 FILLER_58_1114 ();
 sg13g2_decap_8 FILLER_58_1121 ();
 sg13g2_decap_8 FILLER_58_1128 ();
 sg13g2_fill_2 FILLER_58_1135 ();
 sg13g2_fill_1 FILLER_58_1137 ();
 sg13g2_decap_8 FILLER_58_1142 ();
 sg13g2_fill_2 FILLER_58_1149 ();
 sg13g2_decap_8 FILLER_58_1156 ();
 sg13g2_decap_8 FILLER_58_1163 ();
 sg13g2_decap_4 FILLER_58_1170 ();
 sg13g2_fill_1 FILLER_58_1174 ();
 sg13g2_decap_8 FILLER_58_1180 ();
 sg13g2_decap_8 FILLER_58_1187 ();
 sg13g2_decap_8 FILLER_58_1194 ();
 sg13g2_decap_8 FILLER_58_1201 ();
 sg13g2_decap_8 FILLER_58_1208 ();
 sg13g2_decap_8 FILLER_58_1215 ();
 sg13g2_decap_8 FILLER_58_1222 ();
 sg13g2_decap_8 FILLER_58_1229 ();
 sg13g2_decap_8 FILLER_58_1236 ();
 sg13g2_decap_8 FILLER_58_1243 ();
 sg13g2_decap_8 FILLER_58_1250 ();
 sg13g2_decap_8 FILLER_58_1257 ();
 sg13g2_fill_1 FILLER_58_1264 ();
 sg13g2_fill_2 FILLER_58_1284 ();
 sg13g2_fill_2 FILLER_58_1289 ();
 sg13g2_decap_8 FILLER_58_1297 ();
 sg13g2_decap_8 FILLER_58_1304 ();
 sg13g2_decap_8 FILLER_58_1311 ();
 sg13g2_decap_8 FILLER_58_1318 ();
 sg13g2_decap_8 FILLER_58_1325 ();
 sg13g2_decap_8 FILLER_58_1332 ();
 sg13g2_decap_4 FILLER_58_1339 ();
 sg13g2_fill_1 FILLER_58_1343 ();
 sg13g2_decap_8 FILLER_58_1356 ();
 sg13g2_decap_4 FILLER_58_1363 ();
 sg13g2_fill_2 FILLER_58_1367 ();
 sg13g2_fill_2 FILLER_58_1376 ();
 sg13g2_fill_2 FILLER_58_1381 ();
 sg13g2_decap_8 FILLER_58_1398 ();
 sg13g2_decap_8 FILLER_58_1405 ();
 sg13g2_decap_8 FILLER_58_1412 ();
 sg13g2_decap_8 FILLER_58_1419 ();
 sg13g2_decap_4 FILLER_58_1426 ();
 sg13g2_fill_2 FILLER_58_1445 ();
 sg13g2_decap_8 FILLER_58_1457 ();
 sg13g2_decap_4 FILLER_58_1464 ();
 sg13g2_decap_8 FILLER_58_1474 ();
 sg13g2_decap_8 FILLER_58_1481 ();
 sg13g2_decap_8 FILLER_58_1488 ();
 sg13g2_decap_8 FILLER_58_1495 ();
 sg13g2_decap_8 FILLER_58_1502 ();
 sg13g2_decap_8 FILLER_58_1509 ();
 sg13g2_decap_8 FILLER_58_1516 ();
 sg13g2_decap_8 FILLER_58_1523 ();
 sg13g2_decap_8 FILLER_58_1530 ();
 sg13g2_decap_8 FILLER_58_1537 ();
 sg13g2_decap_8 FILLER_58_1544 ();
 sg13g2_decap_8 FILLER_58_1551 ();
 sg13g2_fill_2 FILLER_58_1558 ();
 sg13g2_decap_8 FILLER_58_1567 ();
 sg13g2_decap_8 FILLER_58_1574 ();
 sg13g2_decap_8 FILLER_58_1581 ();
 sg13g2_decap_8 FILLER_58_1588 ();
 sg13g2_decap_8 FILLER_58_1595 ();
 sg13g2_decap_8 FILLER_58_1602 ();
 sg13g2_fill_2 FILLER_58_1609 ();
 sg13g2_decap_4 FILLER_58_1618 ();
 sg13g2_fill_2 FILLER_58_1622 ();
 sg13g2_fill_2 FILLER_58_1635 ();
 sg13g2_decap_8 FILLER_58_1652 ();
 sg13g2_decap_8 FILLER_58_1659 ();
 sg13g2_decap_4 FILLER_58_1666 ();
 sg13g2_decap_8 FILLER_58_1674 ();
 sg13g2_decap_8 FILLER_58_1681 ();
 sg13g2_decap_8 FILLER_58_1688 ();
 sg13g2_decap_8 FILLER_58_1695 ();
 sg13g2_decap_8 FILLER_58_1702 ();
 sg13g2_decap_8 FILLER_58_1709 ();
 sg13g2_decap_8 FILLER_58_1716 ();
 sg13g2_fill_2 FILLER_58_1723 ();
 sg13g2_fill_2 FILLER_58_1730 ();
 sg13g2_decap_8 FILLER_58_1738 ();
 sg13g2_decap_8 FILLER_58_1745 ();
 sg13g2_decap_8 FILLER_58_1752 ();
 sg13g2_decap_8 FILLER_58_1759 ();
 sg13g2_decap_4 FILLER_58_1766 ();
 sg13g2_fill_1 FILLER_58_1770 ();
 sg13g2_decap_8 FILLER_58_1775 ();
 sg13g2_decap_8 FILLER_58_1782 ();
 sg13g2_decap_8 FILLER_58_1789 ();
 sg13g2_decap_8 FILLER_58_1796 ();
 sg13g2_decap_8 FILLER_58_1803 ();
 sg13g2_decap_8 FILLER_58_1810 ();
 sg13g2_decap_8 FILLER_58_1817 ();
 sg13g2_decap_8 FILLER_58_1824 ();
 sg13g2_decap_8 FILLER_58_1831 ();
 sg13g2_decap_8 FILLER_58_1838 ();
 sg13g2_decap_8 FILLER_58_1845 ();
 sg13g2_decap_8 FILLER_58_1852 ();
 sg13g2_decap_8 FILLER_58_1859 ();
 sg13g2_decap_8 FILLER_58_1866 ();
 sg13g2_decap_8 FILLER_58_1873 ();
 sg13g2_decap_8 FILLER_58_1880 ();
 sg13g2_decap_8 FILLER_58_1887 ();
 sg13g2_decap_8 FILLER_58_1894 ();
 sg13g2_decap_8 FILLER_58_1901 ();
 sg13g2_decap_8 FILLER_58_1908 ();
 sg13g2_decap_8 FILLER_58_1915 ();
 sg13g2_decap_8 FILLER_58_1922 ();
 sg13g2_decap_8 FILLER_58_1929 ();
 sg13g2_decap_8 FILLER_58_1936 ();
 sg13g2_decap_8 FILLER_58_1943 ();
 sg13g2_decap_8 FILLER_58_1950 ();
 sg13g2_decap_8 FILLER_58_1957 ();
 sg13g2_decap_8 FILLER_58_1964 ();
 sg13g2_decap_8 FILLER_58_1971 ();
 sg13g2_decap_8 FILLER_58_1978 ();
 sg13g2_decap_8 FILLER_58_1985 ();
 sg13g2_decap_8 FILLER_58_1992 ();
 sg13g2_decap_4 FILLER_58_1999 ();
 sg13g2_fill_1 FILLER_58_2003 ();
 sg13g2_decap_8 FILLER_58_2009 ();
 sg13g2_decap_8 FILLER_58_2016 ();
 sg13g2_decap_8 FILLER_58_2023 ();
 sg13g2_decap_8 FILLER_58_2038 ();
 sg13g2_decap_8 FILLER_58_2045 ();
 sg13g2_decap_8 FILLER_58_2052 ();
 sg13g2_decap_8 FILLER_58_2064 ();
 sg13g2_decap_8 FILLER_58_2071 ();
 sg13g2_decap_8 FILLER_58_2078 ();
 sg13g2_decap_8 FILLER_58_2085 ();
 sg13g2_decap_8 FILLER_58_2092 ();
 sg13g2_decap_8 FILLER_58_2099 ();
 sg13g2_decap_8 FILLER_58_2106 ();
 sg13g2_decap_8 FILLER_58_2113 ();
 sg13g2_decap_8 FILLER_58_2120 ();
 sg13g2_decap_8 FILLER_58_2127 ();
 sg13g2_decap_8 FILLER_58_2134 ();
 sg13g2_decap_8 FILLER_58_2141 ();
 sg13g2_decap_8 FILLER_58_2148 ();
 sg13g2_decap_8 FILLER_58_2155 ();
 sg13g2_decap_8 FILLER_58_2162 ();
 sg13g2_decap_8 FILLER_58_2169 ();
 sg13g2_decap_8 FILLER_58_2176 ();
 sg13g2_decap_8 FILLER_58_2183 ();
 sg13g2_decap_8 FILLER_58_2190 ();
 sg13g2_decap_8 FILLER_58_2197 ();
 sg13g2_decap_8 FILLER_58_2204 ();
 sg13g2_decap_8 FILLER_58_2211 ();
 sg13g2_decap_8 FILLER_58_2218 ();
 sg13g2_decap_8 FILLER_58_2225 ();
 sg13g2_decap_8 FILLER_58_2232 ();
 sg13g2_decap_8 FILLER_58_2239 ();
 sg13g2_decap_8 FILLER_58_2246 ();
 sg13g2_decap_8 FILLER_58_2253 ();
 sg13g2_decap_8 FILLER_58_2260 ();
 sg13g2_decap_8 FILLER_58_2267 ();
 sg13g2_decap_8 FILLER_58_2274 ();
 sg13g2_decap_8 FILLER_58_2281 ();
 sg13g2_decap_8 FILLER_58_2288 ();
 sg13g2_decap_8 FILLER_58_2295 ();
 sg13g2_decap_8 FILLER_58_2302 ();
 sg13g2_decap_8 FILLER_58_2309 ();
 sg13g2_decap_8 FILLER_58_2316 ();
 sg13g2_decap_8 FILLER_58_2323 ();
 sg13g2_decap_8 FILLER_58_2330 ();
 sg13g2_decap_8 FILLER_58_2337 ();
 sg13g2_decap_8 FILLER_58_2344 ();
 sg13g2_decap_8 FILLER_58_2351 ();
 sg13g2_decap_8 FILLER_58_2358 ();
 sg13g2_decap_8 FILLER_58_2365 ();
 sg13g2_decap_8 FILLER_58_2372 ();
 sg13g2_decap_8 FILLER_58_2379 ();
 sg13g2_decap_8 FILLER_58_2386 ();
 sg13g2_decap_8 FILLER_58_2393 ();
 sg13g2_decap_8 FILLER_58_2400 ();
 sg13g2_decap_8 FILLER_58_2407 ();
 sg13g2_decap_8 FILLER_58_2414 ();
 sg13g2_decap_8 FILLER_58_2421 ();
 sg13g2_decap_8 FILLER_58_2428 ();
 sg13g2_decap_8 FILLER_58_2435 ();
 sg13g2_decap_8 FILLER_58_2442 ();
 sg13g2_decap_8 FILLER_58_2449 ();
 sg13g2_decap_8 FILLER_58_2456 ();
 sg13g2_decap_8 FILLER_58_2463 ();
 sg13g2_decap_8 FILLER_58_2470 ();
 sg13g2_decap_8 FILLER_58_2477 ();
 sg13g2_decap_8 FILLER_58_2484 ();
 sg13g2_decap_8 FILLER_58_2491 ();
 sg13g2_decap_8 FILLER_58_2498 ();
 sg13g2_decap_8 FILLER_58_2505 ();
 sg13g2_decap_8 FILLER_58_2512 ();
 sg13g2_decap_8 FILLER_58_2519 ();
 sg13g2_decap_8 FILLER_58_2526 ();
 sg13g2_decap_8 FILLER_58_2533 ();
 sg13g2_decap_8 FILLER_58_2540 ();
 sg13g2_decap_8 FILLER_58_2547 ();
 sg13g2_decap_8 FILLER_58_2554 ();
 sg13g2_decap_8 FILLER_58_2561 ();
 sg13g2_decap_8 FILLER_58_2568 ();
 sg13g2_decap_8 FILLER_58_2575 ();
 sg13g2_decap_8 FILLER_58_2582 ();
 sg13g2_decap_8 FILLER_58_2589 ();
 sg13g2_decap_8 FILLER_58_2596 ();
 sg13g2_decap_8 FILLER_58_2603 ();
 sg13g2_decap_8 FILLER_58_2610 ();
 sg13g2_decap_8 FILLER_58_2617 ();
 sg13g2_decap_8 FILLER_58_2624 ();
 sg13g2_decap_8 FILLER_58_2631 ();
 sg13g2_decap_8 FILLER_58_2638 ();
 sg13g2_decap_8 FILLER_58_2645 ();
 sg13g2_decap_8 FILLER_58_2652 ();
 sg13g2_decap_8 FILLER_58_2659 ();
 sg13g2_decap_4 FILLER_58_2666 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_4 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_57 ();
 sg13g2_decap_8 FILLER_59_64 ();
 sg13g2_decap_8 FILLER_59_71 ();
 sg13g2_decap_8 FILLER_59_78 ();
 sg13g2_fill_2 FILLER_59_85 ();
 sg13g2_decap_8 FILLER_59_91 ();
 sg13g2_decap_8 FILLER_59_98 ();
 sg13g2_decap_8 FILLER_59_105 ();
 sg13g2_decap_8 FILLER_59_112 ();
 sg13g2_decap_8 FILLER_59_119 ();
 sg13g2_decap_8 FILLER_59_126 ();
 sg13g2_decap_8 FILLER_59_133 ();
 sg13g2_fill_2 FILLER_59_140 ();
 sg13g2_fill_1 FILLER_59_142 ();
 sg13g2_decap_8 FILLER_59_147 ();
 sg13g2_decap_8 FILLER_59_154 ();
 sg13g2_decap_8 FILLER_59_161 ();
 sg13g2_fill_2 FILLER_59_168 ();
 sg13g2_fill_1 FILLER_59_170 ();
 sg13g2_decap_8 FILLER_59_174 ();
 sg13g2_decap_8 FILLER_59_181 ();
 sg13g2_fill_1 FILLER_59_188 ();
 sg13g2_decap_8 FILLER_59_192 ();
 sg13g2_decap_8 FILLER_59_199 ();
 sg13g2_decap_8 FILLER_59_206 ();
 sg13g2_decap_8 FILLER_59_213 ();
 sg13g2_decap_8 FILLER_59_220 ();
 sg13g2_decap_8 FILLER_59_227 ();
 sg13g2_decap_8 FILLER_59_234 ();
 sg13g2_decap_8 FILLER_59_241 ();
 sg13g2_decap_8 FILLER_59_248 ();
 sg13g2_decap_8 FILLER_59_255 ();
 sg13g2_decap_8 FILLER_59_262 ();
 sg13g2_decap_8 FILLER_59_269 ();
 sg13g2_decap_8 FILLER_59_276 ();
 sg13g2_decap_8 FILLER_59_283 ();
 sg13g2_decap_8 FILLER_59_290 ();
 sg13g2_decap_8 FILLER_59_297 ();
 sg13g2_decap_8 FILLER_59_304 ();
 sg13g2_decap_8 FILLER_59_311 ();
 sg13g2_decap_8 FILLER_59_318 ();
 sg13g2_decap_8 FILLER_59_325 ();
 sg13g2_fill_2 FILLER_59_332 ();
 sg13g2_decap_8 FILLER_59_346 ();
 sg13g2_decap_8 FILLER_59_353 ();
 sg13g2_decap_8 FILLER_59_360 ();
 sg13g2_decap_8 FILLER_59_367 ();
 sg13g2_decap_8 FILLER_59_374 ();
 sg13g2_decap_8 FILLER_59_381 ();
 sg13g2_decap_8 FILLER_59_388 ();
 sg13g2_decap_8 FILLER_59_395 ();
 sg13g2_fill_2 FILLER_59_402 ();
 sg13g2_decap_8 FILLER_59_407 ();
 sg13g2_decap_8 FILLER_59_414 ();
 sg13g2_decap_8 FILLER_59_421 ();
 sg13g2_decap_8 FILLER_59_428 ();
 sg13g2_fill_2 FILLER_59_435 ();
 sg13g2_decap_8 FILLER_59_446 ();
 sg13g2_decap_8 FILLER_59_453 ();
 sg13g2_decap_8 FILLER_59_460 ();
 sg13g2_decap_8 FILLER_59_467 ();
 sg13g2_decap_8 FILLER_59_474 ();
 sg13g2_decap_8 FILLER_59_481 ();
 sg13g2_decap_8 FILLER_59_488 ();
 sg13g2_decap_8 FILLER_59_495 ();
 sg13g2_decap_8 FILLER_59_502 ();
 sg13g2_decap_4 FILLER_59_509 ();
 sg13g2_decap_8 FILLER_59_532 ();
 sg13g2_decap_4 FILLER_59_539 ();
 sg13g2_decap_4 FILLER_59_547 ();
 sg13g2_decap_8 FILLER_59_556 ();
 sg13g2_decap_8 FILLER_59_568 ();
 sg13g2_decap_4 FILLER_59_575 ();
 sg13g2_fill_2 FILLER_59_579 ();
 sg13g2_decap_8 FILLER_59_586 ();
 sg13g2_decap_8 FILLER_59_593 ();
 sg13g2_decap_8 FILLER_59_600 ();
 sg13g2_decap_8 FILLER_59_607 ();
 sg13g2_decap_8 FILLER_59_614 ();
 sg13g2_decap_4 FILLER_59_621 ();
 sg13g2_fill_2 FILLER_59_625 ();
 sg13g2_decap_8 FILLER_59_634 ();
 sg13g2_decap_8 FILLER_59_641 ();
 sg13g2_decap_4 FILLER_59_648 ();
 sg13g2_fill_2 FILLER_59_657 ();
 sg13g2_decap_8 FILLER_59_682 ();
 sg13g2_decap_8 FILLER_59_689 ();
 sg13g2_fill_2 FILLER_59_696 ();
 sg13g2_decap_4 FILLER_59_716 ();
 sg13g2_decap_4 FILLER_59_725 ();
 sg13g2_fill_2 FILLER_59_729 ();
 sg13g2_fill_2 FILLER_59_745 ();
 sg13g2_decap_8 FILLER_59_760 ();
 sg13g2_decap_8 FILLER_59_767 ();
 sg13g2_decap_8 FILLER_59_774 ();
 sg13g2_decap_4 FILLER_59_781 ();
 sg13g2_fill_2 FILLER_59_785 ();
 sg13g2_decap_8 FILLER_59_790 ();
 sg13g2_decap_4 FILLER_59_797 ();
 sg13g2_fill_1 FILLER_59_801 ();
 sg13g2_decap_8 FILLER_59_828 ();
 sg13g2_decap_8 FILLER_59_835 ();
 sg13g2_decap_8 FILLER_59_842 ();
 sg13g2_decap_8 FILLER_59_849 ();
 sg13g2_fill_2 FILLER_59_856 ();
 sg13g2_fill_1 FILLER_59_858 ();
 sg13g2_fill_1 FILLER_59_874 ();
 sg13g2_decap_8 FILLER_59_893 ();
 sg13g2_decap_4 FILLER_59_900 ();
 sg13g2_fill_1 FILLER_59_904 ();
 sg13g2_decap_8 FILLER_59_911 ();
 sg13g2_decap_8 FILLER_59_918 ();
 sg13g2_fill_2 FILLER_59_925 ();
 sg13g2_decap_8 FILLER_59_944 ();
 sg13g2_decap_8 FILLER_59_951 ();
 sg13g2_decap_4 FILLER_59_958 ();
 sg13g2_fill_2 FILLER_59_962 ();
 sg13g2_fill_2 FILLER_59_969 ();
 sg13g2_decap_8 FILLER_59_987 ();
 sg13g2_fill_2 FILLER_59_994 ();
 sg13g2_decap_8 FILLER_59_1011 ();
 sg13g2_decap_8 FILLER_59_1018 ();
 sg13g2_decap_8 FILLER_59_1025 ();
 sg13g2_decap_8 FILLER_59_1032 ();
 sg13g2_decap_8 FILLER_59_1039 ();
 sg13g2_decap_8 FILLER_59_1046 ();
 sg13g2_decap_8 FILLER_59_1053 ();
 sg13g2_fill_2 FILLER_59_1060 ();
 sg13g2_fill_1 FILLER_59_1062 ();
 sg13g2_decap_8 FILLER_59_1080 ();
 sg13g2_decap_8 FILLER_59_1087 ();
 sg13g2_decap_8 FILLER_59_1094 ();
 sg13g2_decap_8 FILLER_59_1101 ();
 sg13g2_fill_2 FILLER_59_1108 ();
 sg13g2_fill_1 FILLER_59_1110 ();
 sg13g2_fill_2 FILLER_59_1123 ();
 sg13g2_fill_1 FILLER_59_1125 ();
 sg13g2_decap_8 FILLER_59_1131 ();
 sg13g2_decap_8 FILLER_59_1138 ();
 sg13g2_decap_8 FILLER_59_1145 ();
 sg13g2_decap_8 FILLER_59_1152 ();
 sg13g2_decap_8 FILLER_59_1159 ();
 sg13g2_decap_8 FILLER_59_1166 ();
 sg13g2_decap_8 FILLER_59_1173 ();
 sg13g2_decap_8 FILLER_59_1180 ();
 sg13g2_decap_8 FILLER_59_1187 ();
 sg13g2_decap_8 FILLER_59_1194 ();
 sg13g2_decap_4 FILLER_59_1201 ();
 sg13g2_fill_2 FILLER_59_1205 ();
 sg13g2_fill_2 FILLER_59_1216 ();
 sg13g2_fill_1 FILLER_59_1218 ();
 sg13g2_decap_8 FILLER_59_1225 ();
 sg13g2_decap_8 FILLER_59_1232 ();
 sg13g2_decap_8 FILLER_59_1239 ();
 sg13g2_decap_8 FILLER_59_1246 ();
 sg13g2_decap_8 FILLER_59_1253 ();
 sg13g2_fill_2 FILLER_59_1260 ();
 sg13g2_fill_1 FILLER_59_1262 ();
 sg13g2_decap_8 FILLER_59_1304 ();
 sg13g2_decap_8 FILLER_59_1311 ();
 sg13g2_decap_8 FILLER_59_1318 ();
 sg13g2_fill_1 FILLER_59_1325 ();
 sg13g2_decap_8 FILLER_59_1330 ();
 sg13g2_fill_1 FILLER_59_1337 ();
 sg13g2_fill_1 FILLER_59_1357 ();
 sg13g2_fill_2 FILLER_59_1371 ();
 sg13g2_fill_2 FILLER_59_1383 ();
 sg13g2_fill_1 FILLER_59_1385 ();
 sg13g2_decap_8 FILLER_59_1391 ();
 sg13g2_decap_8 FILLER_59_1398 ();
 sg13g2_decap_8 FILLER_59_1405 ();
 sg13g2_decap_8 FILLER_59_1412 ();
 sg13g2_decap_8 FILLER_59_1419 ();
 sg13g2_decap_4 FILLER_59_1426 ();
 sg13g2_decap_8 FILLER_59_1434 ();
 sg13g2_decap_8 FILLER_59_1441 ();
 sg13g2_decap_4 FILLER_59_1448 ();
 sg13g2_fill_1 FILLER_59_1452 ();
 sg13g2_fill_2 FILLER_59_1463 ();
 sg13g2_decap_8 FILLER_59_1480 ();
 sg13g2_decap_8 FILLER_59_1487 ();
 sg13g2_decap_8 FILLER_59_1494 ();
 sg13g2_fill_2 FILLER_59_1501 ();
 sg13g2_decap_8 FILLER_59_1507 ();
 sg13g2_decap_8 FILLER_59_1514 ();
 sg13g2_fill_1 FILLER_59_1521 ();
 sg13g2_decap_8 FILLER_59_1536 ();
 sg13g2_decap_4 FILLER_59_1548 ();
 sg13g2_fill_2 FILLER_59_1552 ();
 sg13g2_decap_8 FILLER_59_1577 ();
 sg13g2_decap_8 FILLER_59_1584 ();
 sg13g2_decap_8 FILLER_59_1591 ();
 sg13g2_fill_2 FILLER_59_1598 ();
 sg13g2_fill_1 FILLER_59_1605 ();
 sg13g2_fill_2 FILLER_59_1611 ();
 sg13g2_fill_1 FILLER_59_1613 ();
 sg13g2_decap_4 FILLER_59_1629 ();
 sg13g2_fill_1 FILLER_59_1633 ();
 sg13g2_decap_8 FILLER_59_1651 ();
 sg13g2_decap_8 FILLER_59_1658 ();
 sg13g2_decap_4 FILLER_59_1665 ();
 sg13g2_fill_1 FILLER_59_1669 ();
 sg13g2_decap_8 FILLER_59_1677 ();
 sg13g2_decap_8 FILLER_59_1684 ();
 sg13g2_decap_4 FILLER_59_1691 ();
 sg13g2_fill_1 FILLER_59_1695 ();
 sg13g2_decap_8 FILLER_59_1711 ();
 sg13g2_decap_8 FILLER_59_1718 ();
 sg13g2_decap_8 FILLER_59_1725 ();
 sg13g2_decap_8 FILLER_59_1732 ();
 sg13g2_decap_8 FILLER_59_1739 ();
 sg13g2_decap_8 FILLER_59_1750 ();
 sg13g2_decap_8 FILLER_59_1757 ();
 sg13g2_decap_8 FILLER_59_1764 ();
 sg13g2_decap_8 FILLER_59_1771 ();
 sg13g2_decap_8 FILLER_59_1786 ();
 sg13g2_decap_8 FILLER_59_1793 ();
 sg13g2_fill_1 FILLER_59_1800 ();
 sg13g2_decap_8 FILLER_59_1805 ();
 sg13g2_decap_8 FILLER_59_1812 ();
 sg13g2_decap_8 FILLER_59_1819 ();
 sg13g2_decap_8 FILLER_59_1826 ();
 sg13g2_decap_8 FILLER_59_1833 ();
 sg13g2_decap_8 FILLER_59_1840 ();
 sg13g2_decap_8 FILLER_59_1847 ();
 sg13g2_decap_8 FILLER_59_1854 ();
 sg13g2_decap_8 FILLER_59_1861 ();
 sg13g2_decap_8 FILLER_59_1868 ();
 sg13g2_decap_8 FILLER_59_1875 ();
 sg13g2_decap_8 FILLER_59_1882 ();
 sg13g2_decap_8 FILLER_59_1889 ();
 sg13g2_decap_8 FILLER_59_1896 ();
 sg13g2_decap_8 FILLER_59_1903 ();
 sg13g2_decap_8 FILLER_59_1910 ();
 sg13g2_decap_8 FILLER_59_1917 ();
 sg13g2_decap_8 FILLER_59_1924 ();
 sg13g2_fill_2 FILLER_59_1931 ();
 sg13g2_fill_1 FILLER_59_1933 ();
 sg13g2_decap_8 FILLER_59_1939 ();
 sg13g2_decap_8 FILLER_59_1946 ();
 sg13g2_decap_8 FILLER_59_1953 ();
 sg13g2_decap_8 FILLER_59_1960 ();
 sg13g2_decap_8 FILLER_59_1967 ();
 sg13g2_decap_8 FILLER_59_1974 ();
 sg13g2_decap_8 FILLER_59_1981 ();
 sg13g2_decap_8 FILLER_59_1988 ();
 sg13g2_decap_8 FILLER_59_1995 ();
 sg13g2_decap_8 FILLER_59_2002 ();
 sg13g2_decap_8 FILLER_59_2009 ();
 sg13g2_decap_8 FILLER_59_2016 ();
 sg13g2_decap_8 FILLER_59_2023 ();
 sg13g2_decap_8 FILLER_59_2030 ();
 sg13g2_decap_8 FILLER_59_2037 ();
 sg13g2_decap_4 FILLER_59_2044 ();
 sg13g2_fill_2 FILLER_59_2048 ();
 sg13g2_decap_8 FILLER_59_2053 ();
 sg13g2_decap_8 FILLER_59_2060 ();
 sg13g2_decap_8 FILLER_59_2067 ();
 sg13g2_decap_8 FILLER_59_2074 ();
 sg13g2_decap_8 FILLER_59_2081 ();
 sg13g2_decap_8 FILLER_59_2088 ();
 sg13g2_decap_8 FILLER_59_2095 ();
 sg13g2_decap_8 FILLER_59_2102 ();
 sg13g2_decap_8 FILLER_59_2109 ();
 sg13g2_decap_8 FILLER_59_2116 ();
 sg13g2_decap_8 FILLER_59_2123 ();
 sg13g2_decap_8 FILLER_59_2130 ();
 sg13g2_decap_8 FILLER_59_2137 ();
 sg13g2_decap_8 FILLER_59_2144 ();
 sg13g2_decap_8 FILLER_59_2151 ();
 sg13g2_decap_4 FILLER_59_2158 ();
 sg13g2_decap_8 FILLER_59_2166 ();
 sg13g2_decap_8 FILLER_59_2173 ();
 sg13g2_decap_8 FILLER_59_2180 ();
 sg13g2_fill_1 FILLER_59_2187 ();
 sg13g2_decap_8 FILLER_59_2191 ();
 sg13g2_decap_4 FILLER_59_2198 ();
 sg13g2_fill_2 FILLER_59_2202 ();
 sg13g2_decap_8 FILLER_59_2212 ();
 sg13g2_fill_2 FILLER_59_2219 ();
 sg13g2_decap_4 FILLER_59_2225 ();
 sg13g2_decap_8 FILLER_59_2255 ();
 sg13g2_decap_8 FILLER_59_2262 ();
 sg13g2_decap_8 FILLER_59_2269 ();
 sg13g2_decap_8 FILLER_59_2276 ();
 sg13g2_decap_8 FILLER_59_2283 ();
 sg13g2_decap_8 FILLER_59_2290 ();
 sg13g2_decap_8 FILLER_59_2297 ();
 sg13g2_decap_8 FILLER_59_2304 ();
 sg13g2_decap_8 FILLER_59_2311 ();
 sg13g2_decap_8 FILLER_59_2318 ();
 sg13g2_decap_8 FILLER_59_2325 ();
 sg13g2_decap_8 FILLER_59_2332 ();
 sg13g2_decap_8 FILLER_59_2339 ();
 sg13g2_decap_8 FILLER_59_2346 ();
 sg13g2_decap_8 FILLER_59_2353 ();
 sg13g2_decap_8 FILLER_59_2360 ();
 sg13g2_decap_8 FILLER_59_2367 ();
 sg13g2_decap_8 FILLER_59_2374 ();
 sg13g2_decap_8 FILLER_59_2381 ();
 sg13g2_decap_8 FILLER_59_2388 ();
 sg13g2_decap_8 FILLER_59_2395 ();
 sg13g2_decap_8 FILLER_59_2402 ();
 sg13g2_decap_8 FILLER_59_2409 ();
 sg13g2_decap_8 FILLER_59_2416 ();
 sg13g2_decap_8 FILLER_59_2423 ();
 sg13g2_decap_8 FILLER_59_2430 ();
 sg13g2_decap_8 FILLER_59_2437 ();
 sg13g2_decap_8 FILLER_59_2444 ();
 sg13g2_decap_8 FILLER_59_2451 ();
 sg13g2_decap_8 FILLER_59_2458 ();
 sg13g2_decap_8 FILLER_59_2465 ();
 sg13g2_decap_8 FILLER_59_2472 ();
 sg13g2_decap_8 FILLER_59_2479 ();
 sg13g2_decap_8 FILLER_59_2486 ();
 sg13g2_decap_8 FILLER_59_2493 ();
 sg13g2_decap_8 FILLER_59_2500 ();
 sg13g2_decap_8 FILLER_59_2507 ();
 sg13g2_decap_8 FILLER_59_2514 ();
 sg13g2_decap_8 FILLER_59_2521 ();
 sg13g2_decap_8 FILLER_59_2528 ();
 sg13g2_decap_8 FILLER_59_2535 ();
 sg13g2_decap_8 FILLER_59_2542 ();
 sg13g2_decap_8 FILLER_59_2549 ();
 sg13g2_decap_8 FILLER_59_2556 ();
 sg13g2_decap_8 FILLER_59_2563 ();
 sg13g2_decap_8 FILLER_59_2570 ();
 sg13g2_decap_8 FILLER_59_2577 ();
 sg13g2_decap_8 FILLER_59_2584 ();
 sg13g2_decap_8 FILLER_59_2591 ();
 sg13g2_decap_8 FILLER_59_2598 ();
 sg13g2_decap_8 FILLER_59_2605 ();
 sg13g2_decap_8 FILLER_59_2612 ();
 sg13g2_decap_8 FILLER_59_2619 ();
 sg13g2_decap_8 FILLER_59_2626 ();
 sg13g2_decap_8 FILLER_59_2633 ();
 sg13g2_decap_8 FILLER_59_2640 ();
 sg13g2_decap_8 FILLER_59_2647 ();
 sg13g2_decap_8 FILLER_59_2654 ();
 sg13g2_decap_8 FILLER_59_2661 ();
 sg13g2_fill_2 FILLER_59_2668 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_61 ();
 sg13g2_decap_8 FILLER_60_68 ();
 sg13g2_decap_8 FILLER_60_75 ();
 sg13g2_decap_8 FILLER_60_82 ();
 sg13g2_fill_2 FILLER_60_89 ();
 sg13g2_decap_8 FILLER_60_95 ();
 sg13g2_decap_8 FILLER_60_102 ();
 sg13g2_decap_8 FILLER_60_109 ();
 sg13g2_fill_1 FILLER_60_116 ();
 sg13g2_decap_8 FILLER_60_121 ();
 sg13g2_decap_4 FILLER_60_128 ();
 sg13g2_decap_4 FILLER_60_137 ();
 sg13g2_fill_2 FILLER_60_141 ();
 sg13g2_decap_4 FILLER_60_148 ();
 sg13g2_fill_1 FILLER_60_152 ();
 sg13g2_decap_8 FILLER_60_158 ();
 sg13g2_fill_1 FILLER_60_165 ();
 sg13g2_fill_1 FILLER_60_170 ();
 sg13g2_decap_8 FILLER_60_176 ();
 sg13g2_decap_4 FILLER_60_183 ();
 sg13g2_fill_2 FILLER_60_195 ();
 sg13g2_decap_8 FILLER_60_201 ();
 sg13g2_decap_8 FILLER_60_208 ();
 sg13g2_decap_8 FILLER_60_215 ();
 sg13g2_decap_8 FILLER_60_222 ();
 sg13g2_decap_8 FILLER_60_229 ();
 sg13g2_decap_8 FILLER_60_236 ();
 sg13g2_decap_8 FILLER_60_243 ();
 sg13g2_decap_8 FILLER_60_250 ();
 sg13g2_decap_8 FILLER_60_257 ();
 sg13g2_decap_8 FILLER_60_264 ();
 sg13g2_decap_8 FILLER_60_271 ();
 sg13g2_decap_8 FILLER_60_278 ();
 sg13g2_decap_8 FILLER_60_285 ();
 sg13g2_decap_8 FILLER_60_292 ();
 sg13g2_decap_8 FILLER_60_299 ();
 sg13g2_decap_8 FILLER_60_306 ();
 sg13g2_fill_2 FILLER_60_313 ();
 sg13g2_fill_1 FILLER_60_315 ();
 sg13g2_fill_1 FILLER_60_337 ();
 sg13g2_decap_8 FILLER_60_344 ();
 sg13g2_decap_8 FILLER_60_351 ();
 sg13g2_decap_8 FILLER_60_358 ();
 sg13g2_decap_8 FILLER_60_365 ();
 sg13g2_decap_8 FILLER_60_372 ();
 sg13g2_decap_8 FILLER_60_379 ();
 sg13g2_decap_8 FILLER_60_386 ();
 sg13g2_decap_8 FILLER_60_393 ();
 sg13g2_decap_8 FILLER_60_400 ();
 sg13g2_decap_8 FILLER_60_407 ();
 sg13g2_decap_8 FILLER_60_414 ();
 sg13g2_decap_4 FILLER_60_421 ();
 sg13g2_decap_8 FILLER_60_444 ();
 sg13g2_decap_8 FILLER_60_451 ();
 sg13g2_decap_8 FILLER_60_458 ();
 sg13g2_decap_8 FILLER_60_465 ();
 sg13g2_decap_4 FILLER_60_472 ();
 sg13g2_decap_8 FILLER_60_489 ();
 sg13g2_decap_8 FILLER_60_496 ();
 sg13g2_fill_2 FILLER_60_503 ();
 sg13g2_fill_1 FILLER_60_517 ();
 sg13g2_decap_8 FILLER_60_530 ();
 sg13g2_decap_8 FILLER_60_537 ();
 sg13g2_decap_4 FILLER_60_544 ();
 sg13g2_fill_2 FILLER_60_548 ();
 sg13g2_decap_8 FILLER_60_555 ();
 sg13g2_fill_1 FILLER_60_562 ();
 sg13g2_decap_8 FILLER_60_566 ();
 sg13g2_decap_8 FILLER_60_573 ();
 sg13g2_decap_8 FILLER_60_580 ();
 sg13g2_decap_8 FILLER_60_587 ();
 sg13g2_decap_8 FILLER_60_594 ();
 sg13g2_decap_8 FILLER_60_601 ();
 sg13g2_decap_8 FILLER_60_608 ();
 sg13g2_decap_8 FILLER_60_615 ();
 sg13g2_decap_4 FILLER_60_622 ();
 sg13g2_fill_1 FILLER_60_626 ();
 sg13g2_decap_8 FILLER_60_630 ();
 sg13g2_decap_8 FILLER_60_637 ();
 sg13g2_decap_8 FILLER_60_644 ();
 sg13g2_decap_8 FILLER_60_651 ();
 sg13g2_decap_8 FILLER_60_658 ();
 sg13g2_decap_4 FILLER_60_665 ();
 sg13g2_decap_8 FILLER_60_675 ();
 sg13g2_decap_8 FILLER_60_682 ();
 sg13g2_decap_8 FILLER_60_689 ();
 sg13g2_decap_8 FILLER_60_696 ();
 sg13g2_fill_1 FILLER_60_712 ();
 sg13g2_decap_8 FILLER_60_718 ();
 sg13g2_decap_8 FILLER_60_725 ();
 sg13g2_fill_1 FILLER_60_732 ();
 sg13g2_decap_8 FILLER_60_753 ();
 sg13g2_decap_8 FILLER_60_760 ();
 sg13g2_decap_8 FILLER_60_767 ();
 sg13g2_decap_8 FILLER_60_774 ();
 sg13g2_decap_8 FILLER_60_781 ();
 sg13g2_decap_8 FILLER_60_788 ();
 sg13g2_decap_8 FILLER_60_795 ();
 sg13g2_fill_1 FILLER_60_817 ();
 sg13g2_decap_8 FILLER_60_821 ();
 sg13g2_decap_8 FILLER_60_828 ();
 sg13g2_decap_8 FILLER_60_835 ();
 sg13g2_decap_8 FILLER_60_842 ();
 sg13g2_decap_8 FILLER_60_849 ();
 sg13g2_decap_8 FILLER_60_856 ();
 sg13g2_fill_2 FILLER_60_863 ();
 sg13g2_fill_1 FILLER_60_865 ();
 sg13g2_decap_4 FILLER_60_876 ();
 sg13g2_fill_1 FILLER_60_880 ();
 sg13g2_decap_8 FILLER_60_886 ();
 sg13g2_decap_8 FILLER_60_893 ();
 sg13g2_decap_4 FILLER_60_900 ();
 sg13g2_fill_1 FILLER_60_904 ();
 sg13g2_decap_8 FILLER_60_910 ();
 sg13g2_decap_8 FILLER_60_917 ();
 sg13g2_decap_8 FILLER_60_924 ();
 sg13g2_decap_8 FILLER_60_931 ();
 sg13g2_decap_8 FILLER_60_938 ();
 sg13g2_decap_8 FILLER_60_945 ();
 sg13g2_decap_8 FILLER_60_952 ();
 sg13g2_decap_8 FILLER_60_959 ();
 sg13g2_decap_8 FILLER_60_966 ();
 sg13g2_decap_4 FILLER_60_973 ();
 sg13g2_decap_8 FILLER_60_983 ();
 sg13g2_decap_8 FILLER_60_990 ();
 sg13g2_decap_8 FILLER_60_997 ();
 sg13g2_decap_8 FILLER_60_1004 ();
 sg13g2_decap_8 FILLER_60_1011 ();
 sg13g2_decap_8 FILLER_60_1018 ();
 sg13g2_decap_8 FILLER_60_1025 ();
 sg13g2_decap_8 FILLER_60_1032 ();
 sg13g2_decap_8 FILLER_60_1039 ();
 sg13g2_decap_8 FILLER_60_1046 ();
 sg13g2_decap_8 FILLER_60_1053 ();
 sg13g2_fill_2 FILLER_60_1060 ();
 sg13g2_fill_1 FILLER_60_1062 ();
 sg13g2_decap_8 FILLER_60_1067 ();
 sg13g2_decap_4 FILLER_60_1074 ();
 sg13g2_fill_2 FILLER_60_1078 ();
 sg13g2_decap_8 FILLER_60_1083 ();
 sg13g2_fill_2 FILLER_60_1090 ();
 sg13g2_fill_1 FILLER_60_1092 ();
 sg13g2_fill_2 FILLER_60_1098 ();
 sg13g2_decap_4 FILLER_60_1106 ();
 sg13g2_fill_1 FILLER_60_1110 ();
 sg13g2_decap_8 FILLER_60_1115 ();
 sg13g2_decap_8 FILLER_60_1122 ();
 sg13g2_decap_8 FILLER_60_1129 ();
 sg13g2_decap_8 FILLER_60_1136 ();
 sg13g2_decap_8 FILLER_60_1143 ();
 sg13g2_decap_8 FILLER_60_1150 ();
 sg13g2_fill_1 FILLER_60_1157 ();
 sg13g2_decap_4 FILLER_60_1162 ();
 sg13g2_fill_2 FILLER_60_1166 ();
 sg13g2_decap_8 FILLER_60_1172 ();
 sg13g2_decap_8 FILLER_60_1179 ();
 sg13g2_decap_8 FILLER_60_1186 ();
 sg13g2_decap_8 FILLER_60_1193 ();
 sg13g2_decap_8 FILLER_60_1205 ();
 sg13g2_decap_8 FILLER_60_1212 ();
 sg13g2_decap_8 FILLER_60_1219 ();
 sg13g2_decap_8 FILLER_60_1226 ();
 sg13g2_decap_8 FILLER_60_1233 ();
 sg13g2_decap_8 FILLER_60_1240 ();
 sg13g2_fill_2 FILLER_60_1247 ();
 sg13g2_decap_8 FILLER_60_1254 ();
 sg13g2_decap_8 FILLER_60_1261 ();
 sg13g2_decap_8 FILLER_60_1268 ();
 sg13g2_decap_8 FILLER_60_1275 ();
 sg13g2_decap_4 FILLER_60_1282 ();
 sg13g2_fill_2 FILLER_60_1289 ();
 sg13g2_decap_8 FILLER_60_1297 ();
 sg13g2_decap_8 FILLER_60_1304 ();
 sg13g2_decap_8 FILLER_60_1311 ();
 sg13g2_decap_8 FILLER_60_1318 ();
 sg13g2_fill_1 FILLER_60_1325 ();
 sg13g2_decap_8 FILLER_60_1331 ();
 sg13g2_decap_4 FILLER_60_1338 ();
 sg13g2_fill_2 FILLER_60_1342 ();
 sg13g2_decap_8 FILLER_60_1367 ();
 sg13g2_decap_8 FILLER_60_1374 ();
 sg13g2_decap_8 FILLER_60_1381 ();
 sg13g2_decap_8 FILLER_60_1388 ();
 sg13g2_fill_1 FILLER_60_1395 ();
 sg13g2_decap_8 FILLER_60_1404 ();
 sg13g2_decap_8 FILLER_60_1411 ();
 sg13g2_decap_8 FILLER_60_1418 ();
 sg13g2_decap_8 FILLER_60_1425 ();
 sg13g2_fill_2 FILLER_60_1432 ();
 sg13g2_decap_8 FILLER_60_1439 ();
 sg13g2_decap_8 FILLER_60_1446 ();
 sg13g2_decap_8 FILLER_60_1453 ();
 sg13g2_decap_8 FILLER_60_1460 ();
 sg13g2_decap_8 FILLER_60_1467 ();
 sg13g2_decap_8 FILLER_60_1474 ();
 sg13g2_fill_2 FILLER_60_1481 ();
 sg13g2_fill_1 FILLER_60_1491 ();
 sg13g2_decap_8 FILLER_60_1497 ();
 sg13g2_decap_8 FILLER_60_1504 ();
 sg13g2_decap_8 FILLER_60_1511 ();
 sg13g2_decap_8 FILLER_60_1518 ();
 sg13g2_decap_8 FILLER_60_1525 ();
 sg13g2_decap_8 FILLER_60_1532 ();
 sg13g2_decap_8 FILLER_60_1539 ();
 sg13g2_decap_8 FILLER_60_1546 ();
 sg13g2_decap_8 FILLER_60_1553 ();
 sg13g2_decap_8 FILLER_60_1560 ();
 sg13g2_decap_8 FILLER_60_1567 ();
 sg13g2_decap_8 FILLER_60_1574 ();
 sg13g2_decap_8 FILLER_60_1581 ();
 sg13g2_decap_8 FILLER_60_1588 ();
 sg13g2_decap_8 FILLER_60_1595 ();
 sg13g2_decap_8 FILLER_60_1602 ();
 sg13g2_decap_8 FILLER_60_1609 ();
 sg13g2_decap_8 FILLER_60_1616 ();
 sg13g2_decap_8 FILLER_60_1623 ();
 sg13g2_decap_8 FILLER_60_1630 ();
 sg13g2_decap_8 FILLER_60_1637 ();
 sg13g2_decap_8 FILLER_60_1644 ();
 sg13g2_decap_8 FILLER_60_1651 ();
 sg13g2_decap_8 FILLER_60_1658 ();
 sg13g2_decap_8 FILLER_60_1665 ();
 sg13g2_decap_8 FILLER_60_1672 ();
 sg13g2_decap_8 FILLER_60_1679 ();
 sg13g2_decap_8 FILLER_60_1686 ();
 sg13g2_fill_2 FILLER_60_1693 ();
 sg13g2_fill_1 FILLER_60_1695 ();
 sg13g2_decap_8 FILLER_60_1708 ();
 sg13g2_decap_8 FILLER_60_1715 ();
 sg13g2_decap_8 FILLER_60_1722 ();
 sg13g2_decap_8 FILLER_60_1729 ();
 sg13g2_fill_2 FILLER_60_1736 ();
 sg13g2_fill_1 FILLER_60_1738 ();
 sg13g2_decap_8 FILLER_60_1747 ();
 sg13g2_decap_8 FILLER_60_1754 ();
 sg13g2_decap_8 FILLER_60_1761 ();
 sg13g2_decap_8 FILLER_60_1768 ();
 sg13g2_decap_8 FILLER_60_1775 ();
 sg13g2_decap_8 FILLER_60_1782 ();
 sg13g2_decap_8 FILLER_60_1789 ();
 sg13g2_decap_8 FILLER_60_1796 ();
 sg13g2_fill_2 FILLER_60_1803 ();
 sg13g2_fill_1 FILLER_60_1805 ();
 sg13g2_decap_8 FILLER_60_1819 ();
 sg13g2_decap_8 FILLER_60_1826 ();
 sg13g2_decap_8 FILLER_60_1833 ();
 sg13g2_decap_8 FILLER_60_1840 ();
 sg13g2_decap_8 FILLER_60_1847 ();
 sg13g2_decap_8 FILLER_60_1854 ();
 sg13g2_decap_4 FILLER_60_1861 ();
 sg13g2_decap_8 FILLER_60_1886 ();
 sg13g2_decap_8 FILLER_60_1893 ();
 sg13g2_decap_8 FILLER_60_1900 ();
 sg13g2_decap_8 FILLER_60_1907 ();
 sg13g2_decap_8 FILLER_60_1914 ();
 sg13g2_decap_8 FILLER_60_1921 ();
 sg13g2_decap_8 FILLER_60_1928 ();
 sg13g2_decap_8 FILLER_60_1935 ();
 sg13g2_decap_8 FILLER_60_1942 ();
 sg13g2_decap_8 FILLER_60_1949 ();
 sg13g2_decap_8 FILLER_60_1956 ();
 sg13g2_decap_8 FILLER_60_1963 ();
 sg13g2_decap_8 FILLER_60_1970 ();
 sg13g2_decap_8 FILLER_60_1977 ();
 sg13g2_decap_8 FILLER_60_1984 ();
 sg13g2_decap_8 FILLER_60_1991 ();
 sg13g2_decap_8 FILLER_60_1998 ();
 sg13g2_decap_8 FILLER_60_2005 ();
 sg13g2_decap_8 FILLER_60_2012 ();
 sg13g2_decap_8 FILLER_60_2019 ();
 sg13g2_decap_8 FILLER_60_2026 ();
 sg13g2_decap_8 FILLER_60_2033 ();
 sg13g2_decap_4 FILLER_60_2040 ();
 sg13g2_fill_2 FILLER_60_2044 ();
 sg13g2_decap_4 FILLER_60_2080 ();
 sg13g2_fill_2 FILLER_60_2084 ();
 sg13g2_decap_8 FILLER_60_2098 ();
 sg13g2_decap_8 FILLER_60_2105 ();
 sg13g2_decap_8 FILLER_60_2112 ();
 sg13g2_decap_8 FILLER_60_2119 ();
 sg13g2_decap_8 FILLER_60_2126 ();
 sg13g2_decap_8 FILLER_60_2133 ();
 sg13g2_decap_8 FILLER_60_2140 ();
 sg13g2_decap_8 FILLER_60_2147 ();
 sg13g2_decap_8 FILLER_60_2154 ();
 sg13g2_decap_8 FILLER_60_2161 ();
 sg13g2_decap_8 FILLER_60_2168 ();
 sg13g2_decap_8 FILLER_60_2175 ();
 sg13g2_decap_8 FILLER_60_2188 ();
 sg13g2_decap_8 FILLER_60_2195 ();
 sg13g2_decap_8 FILLER_60_2202 ();
 sg13g2_decap_8 FILLER_60_2209 ();
 sg13g2_decap_8 FILLER_60_2216 ();
 sg13g2_decap_8 FILLER_60_2223 ();
 sg13g2_decap_8 FILLER_60_2230 ();
 sg13g2_fill_1 FILLER_60_2237 ();
 sg13g2_decap_8 FILLER_60_2242 ();
 sg13g2_decap_8 FILLER_60_2249 ();
 sg13g2_decap_8 FILLER_60_2256 ();
 sg13g2_decap_8 FILLER_60_2263 ();
 sg13g2_decap_8 FILLER_60_2270 ();
 sg13g2_decap_8 FILLER_60_2277 ();
 sg13g2_decap_8 FILLER_60_2284 ();
 sg13g2_decap_8 FILLER_60_2291 ();
 sg13g2_decap_8 FILLER_60_2298 ();
 sg13g2_decap_8 FILLER_60_2305 ();
 sg13g2_decap_8 FILLER_60_2312 ();
 sg13g2_decap_8 FILLER_60_2319 ();
 sg13g2_decap_8 FILLER_60_2326 ();
 sg13g2_decap_8 FILLER_60_2333 ();
 sg13g2_decap_8 FILLER_60_2340 ();
 sg13g2_decap_8 FILLER_60_2347 ();
 sg13g2_decap_8 FILLER_60_2354 ();
 sg13g2_decap_8 FILLER_60_2361 ();
 sg13g2_decap_8 FILLER_60_2368 ();
 sg13g2_decap_8 FILLER_60_2375 ();
 sg13g2_decap_8 FILLER_60_2382 ();
 sg13g2_decap_8 FILLER_60_2389 ();
 sg13g2_decap_8 FILLER_60_2396 ();
 sg13g2_decap_8 FILLER_60_2403 ();
 sg13g2_decap_8 FILLER_60_2410 ();
 sg13g2_decap_8 FILLER_60_2417 ();
 sg13g2_decap_8 FILLER_60_2424 ();
 sg13g2_decap_8 FILLER_60_2431 ();
 sg13g2_decap_8 FILLER_60_2438 ();
 sg13g2_decap_8 FILLER_60_2445 ();
 sg13g2_decap_8 FILLER_60_2452 ();
 sg13g2_decap_8 FILLER_60_2459 ();
 sg13g2_decap_8 FILLER_60_2466 ();
 sg13g2_decap_8 FILLER_60_2473 ();
 sg13g2_decap_8 FILLER_60_2480 ();
 sg13g2_decap_8 FILLER_60_2487 ();
 sg13g2_decap_8 FILLER_60_2494 ();
 sg13g2_decap_8 FILLER_60_2501 ();
 sg13g2_decap_8 FILLER_60_2508 ();
 sg13g2_decap_8 FILLER_60_2515 ();
 sg13g2_decap_8 FILLER_60_2522 ();
 sg13g2_decap_8 FILLER_60_2529 ();
 sg13g2_decap_8 FILLER_60_2536 ();
 sg13g2_decap_8 FILLER_60_2543 ();
 sg13g2_decap_8 FILLER_60_2550 ();
 sg13g2_decap_8 FILLER_60_2557 ();
 sg13g2_decap_8 FILLER_60_2564 ();
 sg13g2_decap_8 FILLER_60_2571 ();
 sg13g2_decap_8 FILLER_60_2578 ();
 sg13g2_decap_8 FILLER_60_2585 ();
 sg13g2_decap_8 FILLER_60_2592 ();
 sg13g2_decap_8 FILLER_60_2599 ();
 sg13g2_decap_8 FILLER_60_2606 ();
 sg13g2_decap_8 FILLER_60_2613 ();
 sg13g2_decap_8 FILLER_60_2620 ();
 sg13g2_decap_8 FILLER_60_2627 ();
 sg13g2_decap_8 FILLER_60_2634 ();
 sg13g2_decap_8 FILLER_60_2641 ();
 sg13g2_decap_8 FILLER_60_2648 ();
 sg13g2_decap_8 FILLER_60_2655 ();
 sg13g2_decap_8 FILLER_60_2662 ();
 sg13g2_fill_1 FILLER_60_2669 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_fill_1 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_62 ();
 sg13g2_decap_8 FILLER_61_69 ();
 sg13g2_fill_2 FILLER_61_76 ();
 sg13g2_fill_1 FILLER_61_78 ();
 sg13g2_decap_8 FILLER_61_83 ();
 sg13g2_decap_8 FILLER_61_90 ();
 sg13g2_decap_8 FILLER_61_97 ();
 sg13g2_decap_8 FILLER_61_104 ();
 sg13g2_decap_8 FILLER_61_120 ();
 sg13g2_decap_8 FILLER_61_127 ();
 sg13g2_decap_8 FILLER_61_134 ();
 sg13g2_decap_8 FILLER_61_141 ();
 sg13g2_decap_4 FILLER_61_148 ();
 sg13g2_decap_8 FILLER_61_157 ();
 sg13g2_decap_8 FILLER_61_164 ();
 sg13g2_decap_8 FILLER_61_171 ();
 sg13g2_decap_8 FILLER_61_178 ();
 sg13g2_decap_8 FILLER_61_185 ();
 sg13g2_decap_8 FILLER_61_192 ();
 sg13g2_decap_8 FILLER_61_199 ();
 sg13g2_decap_8 FILLER_61_206 ();
 sg13g2_decap_8 FILLER_61_213 ();
 sg13g2_decap_8 FILLER_61_220 ();
 sg13g2_decap_8 FILLER_61_227 ();
 sg13g2_decap_8 FILLER_61_234 ();
 sg13g2_decap_8 FILLER_61_241 ();
 sg13g2_decap_8 FILLER_61_248 ();
 sg13g2_decap_8 FILLER_61_255 ();
 sg13g2_decap_8 FILLER_61_262 ();
 sg13g2_decap_8 FILLER_61_269 ();
 sg13g2_decap_8 FILLER_61_276 ();
 sg13g2_decap_8 FILLER_61_283 ();
 sg13g2_decap_8 FILLER_61_290 ();
 sg13g2_decap_8 FILLER_61_297 ();
 sg13g2_fill_2 FILLER_61_304 ();
 sg13g2_fill_2 FILLER_61_317 ();
 sg13g2_decap_8 FILLER_61_353 ();
 sg13g2_decap_8 FILLER_61_360 ();
 sg13g2_decap_8 FILLER_61_367 ();
 sg13g2_decap_8 FILLER_61_374 ();
 sg13g2_decap_8 FILLER_61_381 ();
 sg13g2_decap_8 FILLER_61_388 ();
 sg13g2_decap_8 FILLER_61_395 ();
 sg13g2_decap_8 FILLER_61_402 ();
 sg13g2_decap_8 FILLER_61_409 ();
 sg13g2_fill_1 FILLER_61_416 ();
 sg13g2_decap_8 FILLER_61_421 ();
 sg13g2_decap_8 FILLER_61_428 ();
 sg13g2_decap_8 FILLER_61_435 ();
 sg13g2_decap_8 FILLER_61_442 ();
 sg13g2_decap_8 FILLER_61_449 ();
 sg13g2_fill_1 FILLER_61_456 ();
 sg13g2_decap_8 FILLER_61_463 ();
 sg13g2_fill_2 FILLER_61_470 ();
 sg13g2_fill_1 FILLER_61_472 ();
 sg13g2_fill_2 FILLER_61_488 ();
 sg13g2_decap_8 FILLER_61_494 ();
 sg13g2_decap_4 FILLER_61_501 ();
 sg13g2_decap_8 FILLER_61_516 ();
 sg13g2_fill_2 FILLER_61_523 ();
 sg13g2_decap_8 FILLER_61_529 ();
 sg13g2_decap_4 FILLER_61_536 ();
 sg13g2_fill_1 FILLER_61_545 ();
 sg13g2_decap_8 FILLER_61_551 ();
 sg13g2_decap_8 FILLER_61_558 ();
 sg13g2_decap_8 FILLER_61_565 ();
 sg13g2_decap_8 FILLER_61_572 ();
 sg13g2_decap_8 FILLER_61_579 ();
 sg13g2_fill_2 FILLER_61_586 ();
 sg13g2_fill_1 FILLER_61_588 ();
 sg13g2_decap_4 FILLER_61_594 ();
 sg13g2_fill_1 FILLER_61_598 ();
 sg13g2_decap_8 FILLER_61_604 ();
 sg13g2_decap_8 FILLER_61_611 ();
 sg13g2_fill_2 FILLER_61_618 ();
 sg13g2_fill_2 FILLER_61_625 ();
 sg13g2_decap_8 FILLER_61_639 ();
 sg13g2_decap_8 FILLER_61_646 ();
 sg13g2_decap_4 FILLER_61_656 ();
 sg13g2_decap_8 FILLER_61_681 ();
 sg13g2_decap_8 FILLER_61_688 ();
 sg13g2_decap_8 FILLER_61_695 ();
 sg13g2_decap_8 FILLER_61_702 ();
 sg13g2_decap_8 FILLER_61_709 ();
 sg13g2_decap_8 FILLER_61_716 ();
 sg13g2_decap_4 FILLER_61_723 ();
 sg13g2_fill_1 FILLER_61_727 ();
 sg13g2_fill_1 FILLER_61_755 ();
 sg13g2_decap_8 FILLER_61_768 ();
 sg13g2_decap_8 FILLER_61_775 ();
 sg13g2_decap_8 FILLER_61_782 ();
 sg13g2_decap_8 FILLER_61_789 ();
 sg13g2_decap_8 FILLER_61_811 ();
 sg13g2_decap_8 FILLER_61_818 ();
 sg13g2_fill_1 FILLER_61_825 ();
 sg13g2_decap_8 FILLER_61_830 ();
 sg13g2_decap_8 FILLER_61_837 ();
 sg13g2_decap_8 FILLER_61_844 ();
 sg13g2_decap_8 FILLER_61_851 ();
 sg13g2_decap_8 FILLER_61_858 ();
 sg13g2_decap_4 FILLER_61_865 ();
 sg13g2_fill_1 FILLER_61_869 ();
 sg13g2_decap_8 FILLER_61_875 ();
 sg13g2_decap_8 FILLER_61_882 ();
 sg13g2_decap_8 FILLER_61_889 ();
 sg13g2_decap_4 FILLER_61_896 ();
 sg13g2_fill_2 FILLER_61_900 ();
 sg13g2_fill_2 FILLER_61_917 ();
 sg13g2_fill_1 FILLER_61_919 ();
 sg13g2_decap_8 FILLER_61_926 ();
 sg13g2_decap_8 FILLER_61_933 ();
 sg13g2_decap_8 FILLER_61_940 ();
 sg13g2_fill_2 FILLER_61_947 ();
 sg13g2_fill_1 FILLER_61_949 ();
 sg13g2_decap_8 FILLER_61_954 ();
 sg13g2_decap_8 FILLER_61_961 ();
 sg13g2_decap_8 FILLER_61_968 ();
 sg13g2_decap_8 FILLER_61_975 ();
 sg13g2_decap_8 FILLER_61_982 ();
 sg13g2_decap_8 FILLER_61_989 ();
 sg13g2_decap_4 FILLER_61_996 ();
 sg13g2_decap_8 FILLER_61_1013 ();
 sg13g2_decap_8 FILLER_61_1020 ();
 sg13g2_decap_8 FILLER_61_1027 ();
 sg13g2_decap_8 FILLER_61_1034 ();
 sg13g2_fill_2 FILLER_61_1041 ();
 sg13g2_decap_8 FILLER_61_1058 ();
 sg13g2_decap_8 FILLER_61_1065 ();
 sg13g2_fill_2 FILLER_61_1072 ();
 sg13g2_fill_1 FILLER_61_1074 ();
 sg13g2_fill_1 FILLER_61_1079 ();
 sg13g2_fill_2 FILLER_61_1098 ();
 sg13g2_decap_8 FILLER_61_1104 ();
 sg13g2_decap_8 FILLER_61_1111 ();
 sg13g2_decap_8 FILLER_61_1118 ();
 sg13g2_decap_8 FILLER_61_1125 ();
 sg13g2_decap_8 FILLER_61_1132 ();
 sg13g2_decap_8 FILLER_61_1139 ();
 sg13g2_decap_8 FILLER_61_1146 ();
 sg13g2_decap_8 FILLER_61_1153 ();
 sg13g2_decap_8 FILLER_61_1160 ();
 sg13g2_decap_8 FILLER_61_1167 ();
 sg13g2_decap_8 FILLER_61_1174 ();
 sg13g2_decap_8 FILLER_61_1181 ();
 sg13g2_decap_8 FILLER_61_1188 ();
 sg13g2_decap_8 FILLER_61_1195 ();
 sg13g2_decap_8 FILLER_61_1202 ();
 sg13g2_decap_8 FILLER_61_1209 ();
 sg13g2_decap_8 FILLER_61_1216 ();
 sg13g2_decap_8 FILLER_61_1223 ();
 sg13g2_decap_4 FILLER_61_1230 ();
 sg13g2_decap_8 FILLER_61_1246 ();
 sg13g2_decap_8 FILLER_61_1253 ();
 sg13g2_decap_8 FILLER_61_1260 ();
 sg13g2_decap_8 FILLER_61_1267 ();
 sg13g2_fill_2 FILLER_61_1274 ();
 sg13g2_fill_1 FILLER_61_1276 ();
 sg13g2_decap_8 FILLER_61_1281 ();
 sg13g2_decap_8 FILLER_61_1288 ();
 sg13g2_decap_4 FILLER_61_1295 ();
 sg13g2_fill_2 FILLER_61_1299 ();
 sg13g2_decap_8 FILLER_61_1313 ();
 sg13g2_decap_8 FILLER_61_1320 ();
 sg13g2_decap_8 FILLER_61_1327 ();
 sg13g2_decap_8 FILLER_61_1334 ();
 sg13g2_decap_4 FILLER_61_1341 ();
 sg13g2_fill_2 FILLER_61_1345 ();
 sg13g2_decap_4 FILLER_61_1355 ();
 sg13g2_decap_8 FILLER_61_1374 ();
 sg13g2_decap_8 FILLER_61_1381 ();
 sg13g2_decap_8 FILLER_61_1388 ();
 sg13g2_decap_8 FILLER_61_1395 ();
 sg13g2_decap_8 FILLER_61_1402 ();
 sg13g2_decap_8 FILLER_61_1409 ();
 sg13g2_decap_8 FILLER_61_1416 ();
 sg13g2_decap_8 FILLER_61_1423 ();
 sg13g2_decap_4 FILLER_61_1430 ();
 sg13g2_decap_8 FILLER_61_1439 ();
 sg13g2_decap_8 FILLER_61_1446 ();
 sg13g2_decap_8 FILLER_61_1453 ();
 sg13g2_decap_8 FILLER_61_1460 ();
 sg13g2_decap_4 FILLER_61_1467 ();
 sg13g2_fill_2 FILLER_61_1471 ();
 sg13g2_decap_8 FILLER_61_1485 ();
 sg13g2_decap_8 FILLER_61_1492 ();
 sg13g2_decap_8 FILLER_61_1499 ();
 sg13g2_decap_8 FILLER_61_1506 ();
 sg13g2_decap_8 FILLER_61_1513 ();
 sg13g2_decap_8 FILLER_61_1520 ();
 sg13g2_fill_2 FILLER_61_1527 ();
 sg13g2_fill_1 FILLER_61_1529 ();
 sg13g2_decap_8 FILLER_61_1533 ();
 sg13g2_decap_8 FILLER_61_1540 ();
 sg13g2_decap_8 FILLER_61_1547 ();
 sg13g2_decap_8 FILLER_61_1554 ();
 sg13g2_decap_8 FILLER_61_1561 ();
 sg13g2_decap_8 FILLER_61_1568 ();
 sg13g2_decap_8 FILLER_61_1575 ();
 sg13g2_decap_8 FILLER_61_1582 ();
 sg13g2_decap_8 FILLER_61_1589 ();
 sg13g2_decap_8 FILLER_61_1596 ();
 sg13g2_decap_8 FILLER_61_1603 ();
 sg13g2_decap_8 FILLER_61_1610 ();
 sg13g2_decap_8 FILLER_61_1617 ();
 sg13g2_decap_4 FILLER_61_1624 ();
 sg13g2_fill_1 FILLER_61_1628 ();
 sg13g2_decap_8 FILLER_61_1635 ();
 sg13g2_decap_8 FILLER_61_1642 ();
 sg13g2_decap_8 FILLER_61_1649 ();
 sg13g2_decap_8 FILLER_61_1656 ();
 sg13g2_decap_4 FILLER_61_1663 ();
 sg13g2_decap_8 FILLER_61_1675 ();
 sg13g2_decap_4 FILLER_61_1682 ();
 sg13g2_fill_2 FILLER_61_1686 ();
 sg13g2_fill_2 FILLER_61_1694 ();
 sg13g2_decap_8 FILLER_61_1711 ();
 sg13g2_decap_8 FILLER_61_1718 ();
 sg13g2_decap_8 FILLER_61_1725 ();
 sg13g2_decap_8 FILLER_61_1732 ();
 sg13g2_decap_8 FILLER_61_1739 ();
 sg13g2_decap_8 FILLER_61_1746 ();
 sg13g2_decap_8 FILLER_61_1753 ();
 sg13g2_decap_8 FILLER_61_1760 ();
 sg13g2_decap_8 FILLER_61_1767 ();
 sg13g2_decap_8 FILLER_61_1774 ();
 sg13g2_decap_8 FILLER_61_1781 ();
 sg13g2_decap_8 FILLER_61_1788 ();
 sg13g2_decap_8 FILLER_61_1795 ();
 sg13g2_decap_8 FILLER_61_1806 ();
 sg13g2_decap_8 FILLER_61_1813 ();
 sg13g2_decap_8 FILLER_61_1820 ();
 sg13g2_decap_8 FILLER_61_1827 ();
 sg13g2_decap_8 FILLER_61_1834 ();
 sg13g2_decap_8 FILLER_61_1841 ();
 sg13g2_decap_8 FILLER_61_1848 ();
 sg13g2_decap_4 FILLER_61_1855 ();
 sg13g2_decap_8 FILLER_61_1912 ();
 sg13g2_decap_8 FILLER_61_1919 ();
 sg13g2_decap_8 FILLER_61_1926 ();
 sg13g2_decap_8 FILLER_61_1933 ();
 sg13g2_decap_8 FILLER_61_1940 ();
 sg13g2_fill_2 FILLER_61_1947 ();
 sg13g2_decap_4 FILLER_61_1952 ();
 sg13g2_decap_8 FILLER_61_1960 ();
 sg13g2_decap_8 FILLER_61_1967 ();
 sg13g2_decap_8 FILLER_61_1974 ();
 sg13g2_decap_4 FILLER_61_1981 ();
 sg13g2_fill_2 FILLER_61_1988 ();
 sg13g2_fill_1 FILLER_61_1990 ();
 sg13g2_decap_8 FILLER_61_1995 ();
 sg13g2_decap_8 FILLER_61_2002 ();
 sg13g2_decap_8 FILLER_61_2009 ();
 sg13g2_decap_8 FILLER_61_2016 ();
 sg13g2_decap_8 FILLER_61_2023 ();
 sg13g2_decap_8 FILLER_61_2030 ();
 sg13g2_decap_8 FILLER_61_2037 ();
 sg13g2_decap_8 FILLER_61_2044 ();
 sg13g2_decap_8 FILLER_61_2051 ();
 sg13g2_decap_8 FILLER_61_2058 ();
 sg13g2_decap_8 FILLER_61_2065 ();
 sg13g2_decap_8 FILLER_61_2072 ();
 sg13g2_decap_8 FILLER_61_2079 ();
 sg13g2_decap_8 FILLER_61_2086 ();
 sg13g2_decap_4 FILLER_61_2093 ();
 sg13g2_decap_4 FILLER_61_2101 ();
 sg13g2_fill_1 FILLER_61_2105 ();
 sg13g2_decap_8 FILLER_61_2114 ();
 sg13g2_decap_8 FILLER_61_2121 ();
 sg13g2_decap_8 FILLER_61_2128 ();
 sg13g2_decap_8 FILLER_61_2135 ();
 sg13g2_decap_8 FILLER_61_2142 ();
 sg13g2_decap_8 FILLER_61_2149 ();
 sg13g2_decap_4 FILLER_61_2156 ();
 sg13g2_fill_1 FILLER_61_2160 ();
 sg13g2_decap_4 FILLER_61_2164 ();
 sg13g2_fill_1 FILLER_61_2168 ();
 sg13g2_decap_8 FILLER_61_2174 ();
 sg13g2_decap_4 FILLER_61_2181 ();
 sg13g2_decap_8 FILLER_61_2189 ();
 sg13g2_decap_8 FILLER_61_2196 ();
 sg13g2_decap_8 FILLER_61_2203 ();
 sg13g2_decap_8 FILLER_61_2210 ();
 sg13g2_decap_8 FILLER_61_2217 ();
 sg13g2_decap_8 FILLER_61_2224 ();
 sg13g2_decap_8 FILLER_61_2231 ();
 sg13g2_decap_8 FILLER_61_2238 ();
 sg13g2_decap_8 FILLER_61_2245 ();
 sg13g2_decap_8 FILLER_61_2252 ();
 sg13g2_decap_8 FILLER_61_2259 ();
 sg13g2_decap_8 FILLER_61_2266 ();
 sg13g2_decap_8 FILLER_61_2273 ();
 sg13g2_decap_8 FILLER_61_2280 ();
 sg13g2_decap_8 FILLER_61_2287 ();
 sg13g2_decap_8 FILLER_61_2294 ();
 sg13g2_decap_8 FILLER_61_2301 ();
 sg13g2_decap_8 FILLER_61_2308 ();
 sg13g2_decap_8 FILLER_61_2315 ();
 sg13g2_decap_8 FILLER_61_2322 ();
 sg13g2_decap_8 FILLER_61_2329 ();
 sg13g2_decap_8 FILLER_61_2336 ();
 sg13g2_decap_8 FILLER_61_2343 ();
 sg13g2_decap_8 FILLER_61_2350 ();
 sg13g2_decap_8 FILLER_61_2357 ();
 sg13g2_decap_8 FILLER_61_2364 ();
 sg13g2_decap_8 FILLER_61_2371 ();
 sg13g2_decap_8 FILLER_61_2378 ();
 sg13g2_decap_8 FILLER_61_2385 ();
 sg13g2_decap_8 FILLER_61_2392 ();
 sg13g2_decap_8 FILLER_61_2399 ();
 sg13g2_decap_8 FILLER_61_2406 ();
 sg13g2_decap_8 FILLER_61_2413 ();
 sg13g2_decap_8 FILLER_61_2420 ();
 sg13g2_decap_8 FILLER_61_2427 ();
 sg13g2_decap_8 FILLER_61_2434 ();
 sg13g2_decap_8 FILLER_61_2441 ();
 sg13g2_decap_8 FILLER_61_2448 ();
 sg13g2_decap_8 FILLER_61_2455 ();
 sg13g2_decap_8 FILLER_61_2462 ();
 sg13g2_decap_8 FILLER_61_2469 ();
 sg13g2_decap_8 FILLER_61_2476 ();
 sg13g2_decap_8 FILLER_61_2483 ();
 sg13g2_decap_8 FILLER_61_2490 ();
 sg13g2_decap_8 FILLER_61_2497 ();
 sg13g2_decap_8 FILLER_61_2504 ();
 sg13g2_decap_8 FILLER_61_2511 ();
 sg13g2_decap_8 FILLER_61_2518 ();
 sg13g2_decap_8 FILLER_61_2525 ();
 sg13g2_decap_8 FILLER_61_2532 ();
 sg13g2_decap_8 FILLER_61_2539 ();
 sg13g2_decap_8 FILLER_61_2546 ();
 sg13g2_decap_8 FILLER_61_2553 ();
 sg13g2_decap_8 FILLER_61_2560 ();
 sg13g2_decap_8 FILLER_61_2567 ();
 sg13g2_decap_8 FILLER_61_2574 ();
 sg13g2_decap_8 FILLER_61_2581 ();
 sg13g2_decap_8 FILLER_61_2588 ();
 sg13g2_decap_8 FILLER_61_2595 ();
 sg13g2_decap_8 FILLER_61_2602 ();
 sg13g2_decap_8 FILLER_61_2609 ();
 sg13g2_decap_8 FILLER_61_2616 ();
 sg13g2_decap_8 FILLER_61_2623 ();
 sg13g2_decap_8 FILLER_61_2630 ();
 sg13g2_decap_8 FILLER_61_2637 ();
 sg13g2_decap_8 FILLER_61_2644 ();
 sg13g2_decap_8 FILLER_61_2651 ();
 sg13g2_decap_8 FILLER_61_2658 ();
 sg13g2_decap_4 FILLER_61_2665 ();
 sg13g2_fill_1 FILLER_61_2669 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_4 FILLER_62_49 ();
 sg13g2_fill_1 FILLER_62_53 ();
 sg13g2_fill_1 FILLER_62_59 ();
 sg13g2_decap_8 FILLER_62_65 ();
 sg13g2_fill_2 FILLER_62_72 ();
 sg13g2_fill_1 FILLER_62_74 ();
 sg13g2_decap_4 FILLER_62_79 ();
 sg13g2_fill_2 FILLER_62_83 ();
 sg13g2_decap_8 FILLER_62_90 ();
 sg13g2_decap_4 FILLER_62_97 ();
 sg13g2_fill_2 FILLER_62_101 ();
 sg13g2_fill_2 FILLER_62_115 ();
 sg13g2_decap_8 FILLER_62_121 ();
 sg13g2_decap_4 FILLER_62_128 ();
 sg13g2_fill_2 FILLER_62_132 ();
 sg13g2_decap_8 FILLER_62_139 ();
 sg13g2_decap_8 FILLER_62_146 ();
 sg13g2_decap_8 FILLER_62_153 ();
 sg13g2_decap_8 FILLER_62_160 ();
 sg13g2_decap_8 FILLER_62_167 ();
 sg13g2_decap_8 FILLER_62_174 ();
 sg13g2_decap_8 FILLER_62_181 ();
 sg13g2_decap_8 FILLER_62_188 ();
 sg13g2_decap_8 FILLER_62_195 ();
 sg13g2_decap_8 FILLER_62_202 ();
 sg13g2_decap_8 FILLER_62_209 ();
 sg13g2_decap_8 FILLER_62_216 ();
 sg13g2_decap_8 FILLER_62_223 ();
 sg13g2_decap_4 FILLER_62_230 ();
 sg13g2_fill_1 FILLER_62_249 ();
 sg13g2_decap_8 FILLER_62_254 ();
 sg13g2_decap_8 FILLER_62_261 ();
 sg13g2_decap_8 FILLER_62_268 ();
 sg13g2_decap_8 FILLER_62_275 ();
 sg13g2_decap_8 FILLER_62_282 ();
 sg13g2_decap_8 FILLER_62_289 ();
 sg13g2_decap_8 FILLER_62_296 ();
 sg13g2_decap_8 FILLER_62_303 ();
 sg13g2_fill_2 FILLER_62_310 ();
 sg13g2_fill_1 FILLER_62_312 ();
 sg13g2_decap_8 FILLER_62_350 ();
 sg13g2_decap_8 FILLER_62_357 ();
 sg13g2_decap_8 FILLER_62_364 ();
 sg13g2_decap_8 FILLER_62_371 ();
 sg13g2_decap_8 FILLER_62_378 ();
 sg13g2_decap_4 FILLER_62_385 ();
 sg13g2_fill_2 FILLER_62_389 ();
 sg13g2_fill_2 FILLER_62_403 ();
 sg13g2_decap_8 FILLER_62_415 ();
 sg13g2_decap_8 FILLER_62_422 ();
 sg13g2_decap_8 FILLER_62_429 ();
 sg13g2_decap_8 FILLER_62_436 ();
 sg13g2_decap_8 FILLER_62_443 ();
 sg13g2_decap_8 FILLER_62_450 ();
 sg13g2_decap_8 FILLER_62_467 ();
 sg13g2_fill_2 FILLER_62_474 ();
 sg13g2_decap_8 FILLER_62_481 ();
 sg13g2_fill_1 FILLER_62_488 ();
 sg13g2_decap_8 FILLER_62_493 ();
 sg13g2_decap_8 FILLER_62_500 ();
 sg13g2_decap_8 FILLER_62_507 ();
 sg13g2_decap_8 FILLER_62_514 ();
 sg13g2_decap_8 FILLER_62_521 ();
 sg13g2_decap_8 FILLER_62_528 ();
 sg13g2_decap_8 FILLER_62_535 ();
 sg13g2_decap_8 FILLER_62_542 ();
 sg13g2_decap_8 FILLER_62_549 ();
 sg13g2_decap_8 FILLER_62_556 ();
 sg13g2_decap_8 FILLER_62_563 ();
 sg13g2_decap_8 FILLER_62_570 ();
 sg13g2_decap_8 FILLER_62_577 ();
 sg13g2_decap_8 FILLER_62_584 ();
 sg13g2_decap_8 FILLER_62_591 ();
 sg13g2_decap_8 FILLER_62_598 ();
 sg13g2_decap_8 FILLER_62_605 ();
 sg13g2_decap_8 FILLER_62_612 ();
 sg13g2_decap_8 FILLER_62_619 ();
 sg13g2_fill_1 FILLER_62_626 ();
 sg13g2_decap_4 FILLER_62_631 ();
 sg13g2_decap_8 FILLER_62_639 ();
 sg13g2_decap_4 FILLER_62_646 ();
 sg13g2_decap_8 FILLER_62_665 ();
 sg13g2_decap_8 FILLER_62_672 ();
 sg13g2_decap_4 FILLER_62_679 ();
 sg13g2_decap_4 FILLER_62_686 ();
 sg13g2_decap_8 FILLER_62_693 ();
 sg13g2_fill_1 FILLER_62_700 ();
 sg13g2_decap_8 FILLER_62_713 ();
 sg13g2_decap_8 FILLER_62_720 ();
 sg13g2_fill_2 FILLER_62_727 ();
 sg13g2_decap_8 FILLER_62_737 ();
 sg13g2_decap_4 FILLER_62_744 ();
 sg13g2_fill_1 FILLER_62_748 ();
 sg13g2_decap_8 FILLER_62_760 ();
 sg13g2_decap_8 FILLER_62_767 ();
 sg13g2_fill_2 FILLER_62_774 ();
 sg13g2_fill_2 FILLER_62_780 ();
 sg13g2_fill_1 FILLER_62_782 ();
 sg13g2_decap_8 FILLER_62_786 ();
 sg13g2_decap_4 FILLER_62_793 ();
 sg13g2_fill_2 FILLER_62_797 ();
 sg13g2_decap_8 FILLER_62_804 ();
 sg13g2_decap_8 FILLER_62_811 ();
 sg13g2_decap_8 FILLER_62_818 ();
 sg13g2_decap_8 FILLER_62_825 ();
 sg13g2_decap_8 FILLER_62_832 ();
 sg13g2_decap_8 FILLER_62_839 ();
 sg13g2_decap_8 FILLER_62_846 ();
 sg13g2_decap_8 FILLER_62_857 ();
 sg13g2_fill_2 FILLER_62_864 ();
 sg13g2_fill_1 FILLER_62_866 ();
 sg13g2_decap_8 FILLER_62_873 ();
 sg13g2_decap_8 FILLER_62_880 ();
 sg13g2_decap_8 FILLER_62_887 ();
 sg13g2_decap_8 FILLER_62_894 ();
 sg13g2_decap_8 FILLER_62_901 ();
 sg13g2_decap_8 FILLER_62_908 ();
 sg13g2_decap_8 FILLER_62_915 ();
 sg13g2_decap_8 FILLER_62_922 ();
 sg13g2_decap_8 FILLER_62_929 ();
 sg13g2_decap_8 FILLER_62_936 ();
 sg13g2_fill_2 FILLER_62_943 ();
 sg13g2_fill_2 FILLER_62_963 ();
 sg13g2_decap_8 FILLER_62_970 ();
 sg13g2_decap_4 FILLER_62_977 ();
 sg13g2_decap_8 FILLER_62_985 ();
 sg13g2_decap_8 FILLER_62_992 ();
 sg13g2_fill_1 FILLER_62_999 ();
 sg13g2_decap_8 FILLER_62_1009 ();
 sg13g2_decap_8 FILLER_62_1016 ();
 sg13g2_fill_2 FILLER_62_1034 ();
 sg13g2_fill_1 FILLER_62_1036 ();
 sg13g2_decap_4 FILLER_62_1042 ();
 sg13g2_decap_8 FILLER_62_1052 ();
 sg13g2_decap_8 FILLER_62_1059 ();
 sg13g2_decap_8 FILLER_62_1066 ();
 sg13g2_decap_8 FILLER_62_1073 ();
 sg13g2_fill_2 FILLER_62_1080 ();
 sg13g2_fill_1 FILLER_62_1082 ();
 sg13g2_fill_1 FILLER_62_1088 ();
 sg13g2_decap_8 FILLER_62_1093 ();
 sg13g2_decap_8 FILLER_62_1100 ();
 sg13g2_decap_8 FILLER_62_1107 ();
 sg13g2_decap_4 FILLER_62_1114 ();
 sg13g2_fill_1 FILLER_62_1133 ();
 sg13g2_decap_8 FILLER_62_1138 ();
 sg13g2_decap_8 FILLER_62_1145 ();
 sg13g2_decap_8 FILLER_62_1152 ();
 sg13g2_decap_8 FILLER_62_1159 ();
 sg13g2_decap_8 FILLER_62_1166 ();
 sg13g2_decap_8 FILLER_62_1173 ();
 sg13g2_decap_4 FILLER_62_1180 ();
 sg13g2_decap_8 FILLER_62_1187 ();
 sg13g2_decap_8 FILLER_62_1194 ();
 sg13g2_decap_8 FILLER_62_1201 ();
 sg13g2_decap_8 FILLER_62_1208 ();
 sg13g2_decap_8 FILLER_62_1215 ();
 sg13g2_decap_4 FILLER_62_1222 ();
 sg13g2_fill_2 FILLER_62_1226 ();
 sg13g2_decap_8 FILLER_62_1239 ();
 sg13g2_decap_8 FILLER_62_1246 ();
 sg13g2_decap_8 FILLER_62_1253 ();
 sg13g2_decap_8 FILLER_62_1260 ();
 sg13g2_decap_8 FILLER_62_1267 ();
 sg13g2_decap_8 FILLER_62_1289 ();
 sg13g2_decap_4 FILLER_62_1296 ();
 sg13g2_fill_1 FILLER_62_1300 ();
 sg13g2_decap_8 FILLER_62_1306 ();
 sg13g2_fill_2 FILLER_62_1313 ();
 sg13g2_fill_1 FILLER_62_1315 ();
 sg13g2_fill_2 FILLER_62_1322 ();
 sg13g2_fill_1 FILLER_62_1324 ();
 sg13g2_decap_8 FILLER_62_1335 ();
 sg13g2_decap_8 FILLER_62_1342 ();
 sg13g2_fill_1 FILLER_62_1349 ();
 sg13g2_decap_8 FILLER_62_1364 ();
 sg13g2_decap_8 FILLER_62_1371 ();
 sg13g2_decap_8 FILLER_62_1378 ();
 sg13g2_decap_8 FILLER_62_1385 ();
 sg13g2_decap_8 FILLER_62_1392 ();
 sg13g2_fill_1 FILLER_62_1399 ();
 sg13g2_decap_8 FILLER_62_1403 ();
 sg13g2_decap_8 FILLER_62_1410 ();
 sg13g2_decap_8 FILLER_62_1417 ();
 sg13g2_decap_8 FILLER_62_1424 ();
 sg13g2_decap_8 FILLER_62_1431 ();
 sg13g2_decap_8 FILLER_62_1438 ();
 sg13g2_decap_8 FILLER_62_1445 ();
 sg13g2_decap_8 FILLER_62_1452 ();
 sg13g2_decap_8 FILLER_62_1459 ();
 sg13g2_decap_8 FILLER_62_1466 ();
 sg13g2_decap_8 FILLER_62_1473 ();
 sg13g2_decap_8 FILLER_62_1480 ();
 sg13g2_fill_2 FILLER_62_1487 ();
 sg13g2_decap_8 FILLER_62_1497 ();
 sg13g2_decap_8 FILLER_62_1504 ();
 sg13g2_fill_1 FILLER_62_1511 ();
 sg13g2_fill_2 FILLER_62_1527 ();
 sg13g2_fill_1 FILLER_62_1529 ();
 sg13g2_fill_1 FILLER_62_1535 ();
 sg13g2_decap_8 FILLER_62_1542 ();
 sg13g2_decap_8 FILLER_62_1549 ();
 sg13g2_decap_8 FILLER_62_1556 ();
 sg13g2_decap_8 FILLER_62_1563 ();
 sg13g2_decap_4 FILLER_62_1570 ();
 sg13g2_fill_1 FILLER_62_1574 ();
 sg13g2_decap_8 FILLER_62_1578 ();
 sg13g2_decap_8 FILLER_62_1585 ();
 sg13g2_decap_8 FILLER_62_1592 ();
 sg13g2_decap_8 FILLER_62_1599 ();
 sg13g2_decap_8 FILLER_62_1606 ();
 sg13g2_decap_8 FILLER_62_1613 ();
 sg13g2_decap_4 FILLER_62_1620 ();
 sg13g2_fill_2 FILLER_62_1624 ();
 sg13g2_decap_8 FILLER_62_1639 ();
 sg13g2_decap_8 FILLER_62_1646 ();
 sg13g2_fill_1 FILLER_62_1653 ();
 sg13g2_decap_8 FILLER_62_1657 ();
 sg13g2_decap_4 FILLER_62_1664 ();
 sg13g2_fill_2 FILLER_62_1668 ();
 sg13g2_decap_8 FILLER_62_1674 ();
 sg13g2_decap_8 FILLER_62_1681 ();
 sg13g2_decap_8 FILLER_62_1688 ();
 sg13g2_decap_8 FILLER_62_1695 ();
 sg13g2_fill_2 FILLER_62_1702 ();
 sg13g2_decap_8 FILLER_62_1713 ();
 sg13g2_decap_8 FILLER_62_1720 ();
 sg13g2_decap_8 FILLER_62_1727 ();
 sg13g2_decap_8 FILLER_62_1734 ();
 sg13g2_decap_8 FILLER_62_1741 ();
 sg13g2_decap_8 FILLER_62_1748 ();
 sg13g2_decap_8 FILLER_62_1755 ();
 sg13g2_decap_8 FILLER_62_1762 ();
 sg13g2_decap_8 FILLER_62_1769 ();
 sg13g2_decap_8 FILLER_62_1776 ();
 sg13g2_decap_8 FILLER_62_1783 ();
 sg13g2_decap_8 FILLER_62_1803 ();
 sg13g2_fill_2 FILLER_62_1810 ();
 sg13g2_decap_8 FILLER_62_1828 ();
 sg13g2_decap_8 FILLER_62_1835 ();
 sg13g2_decap_8 FILLER_62_1842 ();
 sg13g2_decap_8 FILLER_62_1849 ();
 sg13g2_decap_8 FILLER_62_1856 ();
 sg13g2_fill_2 FILLER_62_1863 ();
 sg13g2_decap_8 FILLER_62_1898 ();
 sg13g2_decap_8 FILLER_62_1905 ();
 sg13g2_decap_8 FILLER_62_1912 ();
 sg13g2_decap_8 FILLER_62_1919 ();
 sg13g2_decap_8 FILLER_62_1926 ();
 sg13g2_decap_8 FILLER_62_1933 ();
 sg13g2_decap_8 FILLER_62_1940 ();
 sg13g2_fill_2 FILLER_62_1947 ();
 sg13g2_decap_8 FILLER_62_1975 ();
 sg13g2_fill_2 FILLER_62_1982 ();
 sg13g2_fill_1 FILLER_62_1984 ();
 sg13g2_decap_8 FILLER_62_2014 ();
 sg13g2_decap_8 FILLER_62_2021 ();
 sg13g2_decap_8 FILLER_62_2028 ();
 sg13g2_decap_8 FILLER_62_2035 ();
 sg13g2_decap_8 FILLER_62_2042 ();
 sg13g2_decap_8 FILLER_62_2049 ();
 sg13g2_decap_8 FILLER_62_2056 ();
 sg13g2_decap_8 FILLER_62_2063 ();
 sg13g2_decap_8 FILLER_62_2070 ();
 sg13g2_decap_8 FILLER_62_2077 ();
 sg13g2_decap_8 FILLER_62_2084 ();
 sg13g2_decap_8 FILLER_62_2091 ();
 sg13g2_decap_8 FILLER_62_2098 ();
 sg13g2_decap_8 FILLER_62_2105 ();
 sg13g2_decap_8 FILLER_62_2112 ();
 sg13g2_decap_8 FILLER_62_2119 ();
 sg13g2_decap_8 FILLER_62_2126 ();
 sg13g2_decap_8 FILLER_62_2133 ();
 sg13g2_decap_8 FILLER_62_2140 ();
 sg13g2_decap_8 FILLER_62_2147 ();
 sg13g2_decap_8 FILLER_62_2154 ();
 sg13g2_decap_8 FILLER_62_2161 ();
 sg13g2_decap_8 FILLER_62_2168 ();
 sg13g2_decap_8 FILLER_62_2175 ();
 sg13g2_decap_8 FILLER_62_2182 ();
 sg13g2_decap_8 FILLER_62_2189 ();
 sg13g2_decap_8 FILLER_62_2196 ();
 sg13g2_decap_8 FILLER_62_2203 ();
 sg13g2_decap_8 FILLER_62_2210 ();
 sg13g2_decap_8 FILLER_62_2217 ();
 sg13g2_decap_8 FILLER_62_2224 ();
 sg13g2_decap_8 FILLER_62_2231 ();
 sg13g2_decap_8 FILLER_62_2238 ();
 sg13g2_decap_8 FILLER_62_2245 ();
 sg13g2_decap_8 FILLER_62_2252 ();
 sg13g2_decap_8 FILLER_62_2259 ();
 sg13g2_decap_8 FILLER_62_2266 ();
 sg13g2_decap_8 FILLER_62_2273 ();
 sg13g2_decap_8 FILLER_62_2280 ();
 sg13g2_decap_8 FILLER_62_2287 ();
 sg13g2_decap_8 FILLER_62_2294 ();
 sg13g2_decap_8 FILLER_62_2301 ();
 sg13g2_decap_8 FILLER_62_2308 ();
 sg13g2_decap_8 FILLER_62_2315 ();
 sg13g2_decap_8 FILLER_62_2322 ();
 sg13g2_decap_8 FILLER_62_2329 ();
 sg13g2_decap_8 FILLER_62_2336 ();
 sg13g2_decap_8 FILLER_62_2343 ();
 sg13g2_decap_8 FILLER_62_2350 ();
 sg13g2_decap_8 FILLER_62_2357 ();
 sg13g2_decap_8 FILLER_62_2364 ();
 sg13g2_decap_8 FILLER_62_2371 ();
 sg13g2_decap_8 FILLER_62_2378 ();
 sg13g2_decap_8 FILLER_62_2385 ();
 sg13g2_decap_8 FILLER_62_2392 ();
 sg13g2_decap_8 FILLER_62_2399 ();
 sg13g2_decap_8 FILLER_62_2406 ();
 sg13g2_decap_8 FILLER_62_2413 ();
 sg13g2_decap_8 FILLER_62_2420 ();
 sg13g2_decap_8 FILLER_62_2427 ();
 sg13g2_decap_8 FILLER_62_2434 ();
 sg13g2_decap_8 FILLER_62_2441 ();
 sg13g2_decap_8 FILLER_62_2448 ();
 sg13g2_decap_8 FILLER_62_2455 ();
 sg13g2_decap_8 FILLER_62_2462 ();
 sg13g2_decap_8 FILLER_62_2469 ();
 sg13g2_decap_8 FILLER_62_2476 ();
 sg13g2_decap_8 FILLER_62_2483 ();
 sg13g2_decap_8 FILLER_62_2490 ();
 sg13g2_decap_8 FILLER_62_2497 ();
 sg13g2_decap_8 FILLER_62_2504 ();
 sg13g2_decap_8 FILLER_62_2511 ();
 sg13g2_decap_8 FILLER_62_2518 ();
 sg13g2_decap_8 FILLER_62_2525 ();
 sg13g2_decap_8 FILLER_62_2532 ();
 sg13g2_decap_8 FILLER_62_2539 ();
 sg13g2_decap_8 FILLER_62_2546 ();
 sg13g2_decap_8 FILLER_62_2553 ();
 sg13g2_decap_8 FILLER_62_2560 ();
 sg13g2_decap_8 FILLER_62_2567 ();
 sg13g2_decap_8 FILLER_62_2574 ();
 sg13g2_decap_8 FILLER_62_2581 ();
 sg13g2_decap_8 FILLER_62_2588 ();
 sg13g2_decap_8 FILLER_62_2595 ();
 sg13g2_decap_8 FILLER_62_2602 ();
 sg13g2_decap_8 FILLER_62_2609 ();
 sg13g2_decap_8 FILLER_62_2616 ();
 sg13g2_decap_8 FILLER_62_2623 ();
 sg13g2_decap_8 FILLER_62_2630 ();
 sg13g2_decap_8 FILLER_62_2637 ();
 sg13g2_decap_8 FILLER_62_2644 ();
 sg13g2_decap_8 FILLER_62_2651 ();
 sg13g2_decap_8 FILLER_62_2658 ();
 sg13g2_decap_4 FILLER_62_2665 ();
 sg13g2_fill_1 FILLER_62_2669 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_fill_1 FILLER_63_56 ();
 sg13g2_decap_4 FILLER_63_63 ();
 sg13g2_fill_2 FILLER_63_67 ();
 sg13g2_decap_8 FILLER_63_73 ();
 sg13g2_decap_8 FILLER_63_80 ();
 sg13g2_decap_8 FILLER_63_87 ();
 sg13g2_decap_8 FILLER_63_94 ();
 sg13g2_decap_8 FILLER_63_101 ();
 sg13g2_decap_8 FILLER_63_108 ();
 sg13g2_decap_8 FILLER_63_115 ();
 sg13g2_decap_8 FILLER_63_122 ();
 sg13g2_fill_1 FILLER_63_129 ();
 sg13g2_decap_8 FILLER_63_137 ();
 sg13g2_decap_8 FILLER_63_144 ();
 sg13g2_decap_8 FILLER_63_151 ();
 sg13g2_decap_8 FILLER_63_158 ();
 sg13g2_decap_8 FILLER_63_165 ();
 sg13g2_fill_2 FILLER_63_172 ();
 sg13g2_decap_8 FILLER_63_178 ();
 sg13g2_decap_8 FILLER_63_185 ();
 sg13g2_decap_8 FILLER_63_192 ();
 sg13g2_decap_8 FILLER_63_199 ();
 sg13g2_decap_8 FILLER_63_206 ();
 sg13g2_decap_8 FILLER_63_213 ();
 sg13g2_decap_8 FILLER_63_220 ();
 sg13g2_decap_8 FILLER_63_227 ();
 sg13g2_decap_8 FILLER_63_234 ();
 sg13g2_fill_2 FILLER_63_241 ();
 sg13g2_decap_8 FILLER_63_269 ();
 sg13g2_decap_8 FILLER_63_276 ();
 sg13g2_decap_8 FILLER_63_283 ();
 sg13g2_decap_8 FILLER_63_290 ();
 sg13g2_decap_4 FILLER_63_297 ();
 sg13g2_fill_1 FILLER_63_301 ();
 sg13g2_fill_1 FILLER_63_325 ();
 sg13g2_decap_8 FILLER_63_352 ();
 sg13g2_decap_8 FILLER_63_359 ();
 sg13g2_decap_8 FILLER_63_366 ();
 sg13g2_decap_8 FILLER_63_373 ();
 sg13g2_decap_8 FILLER_63_380 ();
 sg13g2_decap_8 FILLER_63_387 ();
 sg13g2_fill_2 FILLER_63_399 ();
 sg13g2_decap_8 FILLER_63_406 ();
 sg13g2_decap_8 FILLER_63_413 ();
 sg13g2_decap_8 FILLER_63_420 ();
 sg13g2_decap_8 FILLER_63_427 ();
 sg13g2_decap_4 FILLER_63_434 ();
 sg13g2_fill_2 FILLER_63_438 ();
 sg13g2_decap_8 FILLER_63_444 ();
 sg13g2_decap_8 FILLER_63_451 ();
 sg13g2_decap_8 FILLER_63_458 ();
 sg13g2_decap_8 FILLER_63_465 ();
 sg13g2_fill_1 FILLER_63_472 ();
 sg13g2_decap_8 FILLER_63_478 ();
 sg13g2_decap_8 FILLER_63_485 ();
 sg13g2_decap_8 FILLER_63_492 ();
 sg13g2_decap_8 FILLER_63_499 ();
 sg13g2_decap_8 FILLER_63_506 ();
 sg13g2_decap_8 FILLER_63_517 ();
 sg13g2_decap_8 FILLER_63_524 ();
 sg13g2_decap_8 FILLER_63_531 ();
 sg13g2_decap_4 FILLER_63_538 ();
 sg13g2_fill_2 FILLER_63_542 ();
 sg13g2_decap_8 FILLER_63_548 ();
 sg13g2_decap_8 FILLER_63_555 ();
 sg13g2_decap_8 FILLER_63_562 ();
 sg13g2_decap_4 FILLER_63_569 ();
 sg13g2_fill_1 FILLER_63_573 ();
 sg13g2_decap_8 FILLER_63_577 ();
 sg13g2_decap_8 FILLER_63_584 ();
 sg13g2_decap_8 FILLER_63_591 ();
 sg13g2_decap_8 FILLER_63_598 ();
 sg13g2_decap_8 FILLER_63_605 ();
 sg13g2_decap_8 FILLER_63_612 ();
 sg13g2_decap_8 FILLER_63_619 ();
 sg13g2_decap_8 FILLER_63_626 ();
 sg13g2_decap_8 FILLER_63_633 ();
 sg13g2_decap_8 FILLER_63_640 ();
 sg13g2_decap_4 FILLER_63_647 ();
 sg13g2_fill_2 FILLER_63_651 ();
 sg13g2_decap_8 FILLER_63_657 ();
 sg13g2_decap_8 FILLER_63_664 ();
 sg13g2_decap_4 FILLER_63_671 ();
 sg13g2_fill_2 FILLER_63_675 ();
 sg13g2_fill_1 FILLER_63_682 ();
 sg13g2_fill_1 FILLER_63_688 ();
 sg13g2_decap_8 FILLER_63_706 ();
 sg13g2_decap_8 FILLER_63_713 ();
 sg13g2_decap_8 FILLER_63_720 ();
 sg13g2_decap_8 FILLER_63_727 ();
 sg13g2_decap_8 FILLER_63_734 ();
 sg13g2_decap_8 FILLER_63_741 ();
 sg13g2_decap_4 FILLER_63_748 ();
 sg13g2_decap_8 FILLER_63_755 ();
 sg13g2_decap_8 FILLER_63_762 ();
 sg13g2_decap_8 FILLER_63_769 ();
 sg13g2_decap_8 FILLER_63_776 ();
 sg13g2_decap_8 FILLER_63_789 ();
 sg13g2_decap_8 FILLER_63_796 ();
 sg13g2_decap_8 FILLER_63_803 ();
 sg13g2_decap_8 FILLER_63_810 ();
 sg13g2_decap_8 FILLER_63_817 ();
 sg13g2_decap_8 FILLER_63_824 ();
 sg13g2_decap_8 FILLER_63_831 ();
 sg13g2_decap_8 FILLER_63_838 ();
 sg13g2_decap_8 FILLER_63_845 ();
 sg13g2_decap_8 FILLER_63_852 ();
 sg13g2_decap_8 FILLER_63_859 ();
 sg13g2_fill_2 FILLER_63_866 ();
 sg13g2_decap_8 FILLER_63_872 ();
 sg13g2_decap_8 FILLER_63_879 ();
 sg13g2_decap_8 FILLER_63_886 ();
 sg13g2_decap_8 FILLER_63_893 ();
 sg13g2_decap_8 FILLER_63_900 ();
 sg13g2_decap_8 FILLER_63_907 ();
 sg13g2_decap_8 FILLER_63_914 ();
 sg13g2_decap_8 FILLER_63_921 ();
 sg13g2_decap_8 FILLER_63_928 ();
 sg13g2_fill_1 FILLER_63_935 ();
 sg13g2_decap_8 FILLER_63_939 ();
 sg13g2_decap_8 FILLER_63_946 ();
 sg13g2_decap_4 FILLER_63_953 ();
 sg13g2_decap_8 FILLER_63_961 ();
 sg13g2_decap_8 FILLER_63_968 ();
 sg13g2_decap_8 FILLER_63_975 ();
 sg13g2_decap_8 FILLER_63_982 ();
 sg13g2_decap_8 FILLER_63_989 ();
 sg13g2_decap_8 FILLER_63_996 ();
 sg13g2_decap_8 FILLER_63_1006 ();
 sg13g2_decap_8 FILLER_63_1013 ();
 sg13g2_decap_8 FILLER_63_1020 ();
 sg13g2_decap_8 FILLER_63_1027 ();
 sg13g2_decap_8 FILLER_63_1034 ();
 sg13g2_decap_8 FILLER_63_1041 ();
 sg13g2_decap_8 FILLER_63_1048 ();
 sg13g2_decap_8 FILLER_63_1055 ();
 sg13g2_decap_8 FILLER_63_1062 ();
 sg13g2_decap_8 FILLER_63_1069 ();
 sg13g2_decap_8 FILLER_63_1076 ();
 sg13g2_fill_2 FILLER_63_1083 ();
 sg13g2_fill_1 FILLER_63_1085 ();
 sg13g2_fill_2 FILLER_63_1089 ();
 sg13g2_fill_1 FILLER_63_1091 ();
 sg13g2_decap_8 FILLER_63_1098 ();
 sg13g2_decap_8 FILLER_63_1105 ();
 sg13g2_decap_4 FILLER_63_1112 ();
 sg13g2_fill_2 FILLER_63_1116 ();
 sg13g2_decap_8 FILLER_63_1130 ();
 sg13g2_decap_8 FILLER_63_1137 ();
 sg13g2_decap_8 FILLER_63_1144 ();
 sg13g2_decap_8 FILLER_63_1151 ();
 sg13g2_decap_8 FILLER_63_1158 ();
 sg13g2_decap_8 FILLER_63_1165 ();
 sg13g2_fill_1 FILLER_63_1190 ();
 sg13g2_fill_2 FILLER_63_1196 ();
 sg13g2_decap_8 FILLER_63_1203 ();
 sg13g2_decap_8 FILLER_63_1210 ();
 sg13g2_decap_8 FILLER_63_1217 ();
 sg13g2_decap_8 FILLER_63_1224 ();
 sg13g2_fill_2 FILLER_63_1231 ();
 sg13g2_fill_1 FILLER_63_1233 ();
 sg13g2_fill_1 FILLER_63_1237 ();
 sg13g2_decap_8 FILLER_63_1247 ();
 sg13g2_decap_8 FILLER_63_1254 ();
 sg13g2_decap_8 FILLER_63_1261 ();
 sg13g2_decap_8 FILLER_63_1268 ();
 sg13g2_fill_2 FILLER_63_1275 ();
 sg13g2_decap_8 FILLER_63_1283 ();
 sg13g2_decap_8 FILLER_63_1290 ();
 sg13g2_decap_8 FILLER_63_1297 ();
 sg13g2_decap_8 FILLER_63_1308 ();
 sg13g2_decap_8 FILLER_63_1315 ();
 sg13g2_decap_8 FILLER_63_1322 ();
 sg13g2_decap_8 FILLER_63_1329 ();
 sg13g2_decap_8 FILLER_63_1336 ();
 sg13g2_decap_8 FILLER_63_1343 ();
 sg13g2_decap_8 FILLER_63_1350 ();
 sg13g2_decap_8 FILLER_63_1357 ();
 sg13g2_decap_8 FILLER_63_1364 ();
 sg13g2_decap_8 FILLER_63_1371 ();
 sg13g2_decap_8 FILLER_63_1378 ();
 sg13g2_decap_8 FILLER_63_1385 ();
 sg13g2_decap_8 FILLER_63_1392 ();
 sg13g2_fill_1 FILLER_63_1399 ();
 sg13g2_decap_8 FILLER_63_1405 ();
 sg13g2_decap_8 FILLER_63_1412 ();
 sg13g2_decap_8 FILLER_63_1419 ();
 sg13g2_decap_8 FILLER_63_1426 ();
 sg13g2_decap_8 FILLER_63_1433 ();
 sg13g2_decap_8 FILLER_63_1440 ();
 sg13g2_decap_8 FILLER_63_1447 ();
 sg13g2_decap_4 FILLER_63_1454 ();
 sg13g2_decap_8 FILLER_63_1463 ();
 sg13g2_decap_8 FILLER_63_1470 ();
 sg13g2_decap_8 FILLER_63_1477 ();
 sg13g2_decap_8 FILLER_63_1484 ();
 sg13g2_decap_8 FILLER_63_1491 ();
 sg13g2_decap_8 FILLER_63_1498 ();
 sg13g2_decap_4 FILLER_63_1505 ();
 sg13g2_decap_8 FILLER_63_1526 ();
 sg13g2_fill_2 FILLER_63_1533 ();
 sg13g2_fill_1 FILLER_63_1535 ();
 sg13g2_decap_8 FILLER_63_1540 ();
 sg13g2_decap_4 FILLER_63_1553 ();
 sg13g2_fill_2 FILLER_63_1557 ();
 sg13g2_decap_8 FILLER_63_1564 ();
 sg13g2_decap_4 FILLER_63_1571 ();
 sg13g2_fill_1 FILLER_63_1579 ();
 sg13g2_decap_8 FILLER_63_1588 ();
 sg13g2_fill_1 FILLER_63_1595 ();
 sg13g2_decap_8 FILLER_63_1602 ();
 sg13g2_decap_8 FILLER_63_1609 ();
 sg13g2_decap_4 FILLER_63_1616 ();
 sg13g2_fill_1 FILLER_63_1620 ();
 sg13g2_fill_1 FILLER_63_1626 ();
 sg13g2_fill_1 FILLER_63_1641 ();
 sg13g2_fill_1 FILLER_63_1657 ();
 sg13g2_decap_8 FILLER_63_1668 ();
 sg13g2_decap_8 FILLER_63_1675 ();
 sg13g2_fill_2 FILLER_63_1682 ();
 sg13g2_decap_4 FILLER_63_1689 ();
 sg13g2_fill_1 FILLER_63_1693 ();
 sg13g2_decap_8 FILLER_63_1702 ();
 sg13g2_decap_8 FILLER_63_1709 ();
 sg13g2_decap_8 FILLER_63_1716 ();
 sg13g2_decap_8 FILLER_63_1723 ();
 sg13g2_decap_8 FILLER_63_1730 ();
 sg13g2_fill_1 FILLER_63_1737 ();
 sg13g2_decap_8 FILLER_63_1742 ();
 sg13g2_decap_8 FILLER_63_1753 ();
 sg13g2_decap_8 FILLER_63_1760 ();
 sg13g2_decap_8 FILLER_63_1767 ();
 sg13g2_decap_8 FILLER_63_1774 ();
 sg13g2_decap_8 FILLER_63_1781 ();
 sg13g2_decap_8 FILLER_63_1788 ();
 sg13g2_decap_8 FILLER_63_1795 ();
 sg13g2_decap_8 FILLER_63_1802 ();
 sg13g2_decap_8 FILLER_63_1809 ();
 sg13g2_decap_8 FILLER_63_1816 ();
 sg13g2_decap_8 FILLER_63_1823 ();
 sg13g2_decap_8 FILLER_63_1830 ();
 sg13g2_decap_8 FILLER_63_1837 ();
 sg13g2_decap_8 FILLER_63_1844 ();
 sg13g2_decap_8 FILLER_63_1851 ();
 sg13g2_decap_8 FILLER_63_1858 ();
 sg13g2_decap_8 FILLER_63_1865 ();
 sg13g2_decap_8 FILLER_63_1872 ();
 sg13g2_decap_8 FILLER_63_1879 ();
 sg13g2_decap_8 FILLER_63_1886 ();
 sg13g2_decap_8 FILLER_63_1893 ();
 sg13g2_decap_8 FILLER_63_1900 ();
 sg13g2_decap_8 FILLER_63_1907 ();
 sg13g2_decap_8 FILLER_63_1914 ();
 sg13g2_decap_8 FILLER_63_1921 ();
 sg13g2_decap_8 FILLER_63_1928 ();
 sg13g2_decap_8 FILLER_63_1935 ();
 sg13g2_decap_8 FILLER_63_1942 ();
 sg13g2_decap_8 FILLER_63_1949 ();
 sg13g2_decap_8 FILLER_63_1956 ();
 sg13g2_decap_8 FILLER_63_1963 ();
 sg13g2_decap_8 FILLER_63_1970 ();
 sg13g2_decap_8 FILLER_63_1977 ();
 sg13g2_decap_8 FILLER_63_1984 ();
 sg13g2_decap_8 FILLER_63_1991 ();
 sg13g2_decap_4 FILLER_63_1998 ();
 sg13g2_decap_4 FILLER_63_2006 ();
 sg13g2_fill_1 FILLER_63_2010 ();
 sg13g2_decap_8 FILLER_63_2019 ();
 sg13g2_decap_8 FILLER_63_2026 ();
 sg13g2_decap_8 FILLER_63_2033 ();
 sg13g2_decap_8 FILLER_63_2040 ();
 sg13g2_decap_8 FILLER_63_2047 ();
 sg13g2_decap_8 FILLER_63_2054 ();
 sg13g2_decap_8 FILLER_63_2061 ();
 sg13g2_decap_8 FILLER_63_2068 ();
 sg13g2_decap_8 FILLER_63_2075 ();
 sg13g2_decap_8 FILLER_63_2082 ();
 sg13g2_decap_8 FILLER_63_2089 ();
 sg13g2_fill_2 FILLER_63_2096 ();
 sg13g2_fill_1 FILLER_63_2098 ();
 sg13g2_decap_4 FILLER_63_2102 ();
 sg13g2_decap_8 FILLER_63_2110 ();
 sg13g2_decap_8 FILLER_63_2117 ();
 sg13g2_decap_8 FILLER_63_2124 ();
 sg13g2_decap_8 FILLER_63_2131 ();
 sg13g2_decap_8 FILLER_63_2138 ();
 sg13g2_decap_8 FILLER_63_2145 ();
 sg13g2_decap_8 FILLER_63_2152 ();
 sg13g2_decap_8 FILLER_63_2159 ();
 sg13g2_decap_8 FILLER_63_2166 ();
 sg13g2_decap_8 FILLER_63_2173 ();
 sg13g2_decap_4 FILLER_63_2180 ();
 sg13g2_decap_8 FILLER_63_2190 ();
 sg13g2_decap_8 FILLER_63_2197 ();
 sg13g2_decap_8 FILLER_63_2204 ();
 sg13g2_decap_8 FILLER_63_2211 ();
 sg13g2_decap_8 FILLER_63_2218 ();
 sg13g2_decap_8 FILLER_63_2225 ();
 sg13g2_decap_8 FILLER_63_2232 ();
 sg13g2_decap_8 FILLER_63_2239 ();
 sg13g2_decap_8 FILLER_63_2246 ();
 sg13g2_decap_8 FILLER_63_2253 ();
 sg13g2_decap_8 FILLER_63_2260 ();
 sg13g2_decap_8 FILLER_63_2267 ();
 sg13g2_decap_8 FILLER_63_2274 ();
 sg13g2_decap_8 FILLER_63_2281 ();
 sg13g2_decap_8 FILLER_63_2288 ();
 sg13g2_decap_8 FILLER_63_2295 ();
 sg13g2_decap_8 FILLER_63_2302 ();
 sg13g2_decap_8 FILLER_63_2309 ();
 sg13g2_decap_8 FILLER_63_2316 ();
 sg13g2_decap_8 FILLER_63_2323 ();
 sg13g2_decap_8 FILLER_63_2330 ();
 sg13g2_decap_8 FILLER_63_2337 ();
 sg13g2_decap_8 FILLER_63_2344 ();
 sg13g2_decap_8 FILLER_63_2351 ();
 sg13g2_decap_8 FILLER_63_2358 ();
 sg13g2_decap_8 FILLER_63_2365 ();
 sg13g2_decap_8 FILLER_63_2372 ();
 sg13g2_decap_8 FILLER_63_2379 ();
 sg13g2_decap_8 FILLER_63_2386 ();
 sg13g2_decap_8 FILLER_63_2393 ();
 sg13g2_decap_8 FILLER_63_2400 ();
 sg13g2_decap_8 FILLER_63_2407 ();
 sg13g2_decap_8 FILLER_63_2414 ();
 sg13g2_decap_8 FILLER_63_2421 ();
 sg13g2_decap_8 FILLER_63_2428 ();
 sg13g2_decap_8 FILLER_63_2435 ();
 sg13g2_decap_8 FILLER_63_2442 ();
 sg13g2_decap_8 FILLER_63_2449 ();
 sg13g2_decap_8 FILLER_63_2456 ();
 sg13g2_decap_8 FILLER_63_2463 ();
 sg13g2_decap_8 FILLER_63_2470 ();
 sg13g2_decap_8 FILLER_63_2477 ();
 sg13g2_decap_8 FILLER_63_2484 ();
 sg13g2_decap_8 FILLER_63_2491 ();
 sg13g2_decap_8 FILLER_63_2498 ();
 sg13g2_decap_8 FILLER_63_2505 ();
 sg13g2_decap_8 FILLER_63_2512 ();
 sg13g2_decap_8 FILLER_63_2519 ();
 sg13g2_decap_8 FILLER_63_2526 ();
 sg13g2_decap_8 FILLER_63_2533 ();
 sg13g2_decap_8 FILLER_63_2540 ();
 sg13g2_decap_8 FILLER_63_2547 ();
 sg13g2_decap_8 FILLER_63_2554 ();
 sg13g2_decap_8 FILLER_63_2561 ();
 sg13g2_decap_8 FILLER_63_2568 ();
 sg13g2_decap_8 FILLER_63_2575 ();
 sg13g2_decap_8 FILLER_63_2582 ();
 sg13g2_decap_8 FILLER_63_2589 ();
 sg13g2_decap_8 FILLER_63_2596 ();
 sg13g2_decap_8 FILLER_63_2603 ();
 sg13g2_decap_8 FILLER_63_2610 ();
 sg13g2_decap_8 FILLER_63_2617 ();
 sg13g2_decap_8 FILLER_63_2624 ();
 sg13g2_decap_8 FILLER_63_2631 ();
 sg13g2_decap_8 FILLER_63_2638 ();
 sg13g2_decap_8 FILLER_63_2645 ();
 sg13g2_decap_8 FILLER_63_2652 ();
 sg13g2_decap_8 FILLER_63_2659 ();
 sg13g2_decap_4 FILLER_63_2666 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_91 ();
 sg13g2_decap_8 FILLER_64_98 ();
 sg13g2_decap_8 FILLER_64_105 ();
 sg13g2_decap_8 FILLER_64_112 ();
 sg13g2_decap_8 FILLER_64_119 ();
 sg13g2_decap_8 FILLER_64_126 ();
 sg13g2_decap_8 FILLER_64_133 ();
 sg13g2_decap_8 FILLER_64_140 ();
 sg13g2_decap_8 FILLER_64_147 ();
 sg13g2_decap_8 FILLER_64_154 ();
 sg13g2_decap_8 FILLER_64_161 ();
 sg13g2_decap_8 FILLER_64_173 ();
 sg13g2_decap_8 FILLER_64_180 ();
 sg13g2_decap_8 FILLER_64_187 ();
 sg13g2_decap_8 FILLER_64_194 ();
 sg13g2_decap_8 FILLER_64_201 ();
 sg13g2_decap_8 FILLER_64_208 ();
 sg13g2_decap_8 FILLER_64_215 ();
 sg13g2_decap_8 FILLER_64_222 ();
 sg13g2_decap_8 FILLER_64_229 ();
 sg13g2_decap_8 FILLER_64_236 ();
 sg13g2_decap_8 FILLER_64_243 ();
 sg13g2_decap_8 FILLER_64_250 ();
 sg13g2_decap_8 FILLER_64_257 ();
 sg13g2_decap_8 FILLER_64_264 ();
 sg13g2_decap_8 FILLER_64_271 ();
 sg13g2_decap_8 FILLER_64_278 ();
 sg13g2_decap_8 FILLER_64_285 ();
 sg13g2_decap_8 FILLER_64_292 ();
 sg13g2_decap_8 FILLER_64_299 ();
 sg13g2_fill_2 FILLER_64_306 ();
 sg13g2_fill_1 FILLER_64_308 ();
 sg13g2_fill_1 FILLER_64_328 ();
 sg13g2_fill_2 FILLER_64_335 ();
 sg13g2_decap_8 FILLER_64_352 ();
 sg13g2_decap_8 FILLER_64_359 ();
 sg13g2_decap_8 FILLER_64_366 ();
 sg13g2_decap_8 FILLER_64_373 ();
 sg13g2_decap_8 FILLER_64_380 ();
 sg13g2_decap_8 FILLER_64_387 ();
 sg13g2_decap_8 FILLER_64_394 ();
 sg13g2_decap_8 FILLER_64_401 ();
 sg13g2_decap_8 FILLER_64_408 ();
 sg13g2_decap_8 FILLER_64_415 ();
 sg13g2_decap_8 FILLER_64_422 ();
 sg13g2_decap_8 FILLER_64_429 ();
 sg13g2_decap_8 FILLER_64_436 ();
 sg13g2_decap_8 FILLER_64_443 ();
 sg13g2_decap_8 FILLER_64_450 ();
 sg13g2_decap_8 FILLER_64_457 ();
 sg13g2_fill_2 FILLER_64_464 ();
 sg13g2_decap_8 FILLER_64_469 ();
 sg13g2_decap_8 FILLER_64_476 ();
 sg13g2_decap_8 FILLER_64_483 ();
 sg13g2_decap_8 FILLER_64_490 ();
 sg13g2_decap_8 FILLER_64_497 ();
 sg13g2_decap_8 FILLER_64_504 ();
 sg13g2_decap_8 FILLER_64_511 ();
 sg13g2_decap_8 FILLER_64_518 ();
 sg13g2_decap_8 FILLER_64_525 ();
 sg13g2_decap_8 FILLER_64_532 ();
 sg13g2_decap_8 FILLER_64_539 ();
 sg13g2_decap_8 FILLER_64_546 ();
 sg13g2_decap_8 FILLER_64_553 ();
 sg13g2_decap_4 FILLER_64_560 ();
 sg13g2_fill_2 FILLER_64_564 ();
 sg13g2_decap_8 FILLER_64_580 ();
 sg13g2_decap_8 FILLER_64_587 ();
 sg13g2_decap_8 FILLER_64_594 ();
 sg13g2_decap_8 FILLER_64_601 ();
 sg13g2_decap_4 FILLER_64_608 ();
 sg13g2_fill_2 FILLER_64_612 ();
 sg13g2_decap_4 FILLER_64_618 ();
 sg13g2_decap_8 FILLER_64_628 ();
 sg13g2_decap_8 FILLER_64_635 ();
 sg13g2_fill_2 FILLER_64_642 ();
 sg13g2_fill_1 FILLER_64_644 ();
 sg13g2_decap_8 FILLER_64_664 ();
 sg13g2_fill_2 FILLER_64_671 ();
 sg13g2_fill_1 FILLER_64_692 ();
 sg13g2_decap_8 FILLER_64_698 ();
 sg13g2_decap_8 FILLER_64_705 ();
 sg13g2_decap_8 FILLER_64_712 ();
 sg13g2_decap_8 FILLER_64_719 ();
 sg13g2_decap_4 FILLER_64_726 ();
 sg13g2_decap_8 FILLER_64_735 ();
 sg13g2_decap_8 FILLER_64_742 ();
 sg13g2_decap_8 FILLER_64_749 ();
 sg13g2_decap_8 FILLER_64_756 ();
 sg13g2_decap_8 FILLER_64_763 ();
 sg13g2_decap_4 FILLER_64_770 ();
 sg13g2_fill_1 FILLER_64_774 ();
 sg13g2_decap_8 FILLER_64_779 ();
 sg13g2_decap_8 FILLER_64_786 ();
 sg13g2_decap_4 FILLER_64_793 ();
 sg13g2_fill_1 FILLER_64_797 ();
 sg13g2_decap_8 FILLER_64_803 ();
 sg13g2_decap_8 FILLER_64_810 ();
 sg13g2_decap_8 FILLER_64_817 ();
 sg13g2_decap_8 FILLER_64_824 ();
 sg13g2_fill_2 FILLER_64_831 ();
 sg13g2_decap_8 FILLER_64_838 ();
 sg13g2_decap_8 FILLER_64_845 ();
 sg13g2_decap_8 FILLER_64_852 ();
 sg13g2_decap_8 FILLER_64_859 ();
 sg13g2_decap_8 FILLER_64_870 ();
 sg13g2_decap_4 FILLER_64_877 ();
 sg13g2_fill_1 FILLER_64_881 ();
 sg13g2_decap_8 FILLER_64_888 ();
 sg13g2_decap_8 FILLER_64_895 ();
 sg13g2_fill_1 FILLER_64_902 ();
 sg13g2_decap_8 FILLER_64_908 ();
 sg13g2_decap_8 FILLER_64_915 ();
 sg13g2_decap_8 FILLER_64_922 ();
 sg13g2_decap_4 FILLER_64_929 ();
 sg13g2_decap_8 FILLER_64_936 ();
 sg13g2_decap_8 FILLER_64_943 ();
 sg13g2_decap_8 FILLER_64_950 ();
 sg13g2_decap_8 FILLER_64_957 ();
 sg13g2_decap_8 FILLER_64_964 ();
 sg13g2_decap_4 FILLER_64_971 ();
 sg13g2_decap_8 FILLER_64_980 ();
 sg13g2_decap_8 FILLER_64_987 ();
 sg13g2_decap_8 FILLER_64_994 ();
 sg13g2_decap_8 FILLER_64_1001 ();
 sg13g2_decap_8 FILLER_64_1008 ();
 sg13g2_decap_8 FILLER_64_1015 ();
 sg13g2_decap_8 FILLER_64_1022 ();
 sg13g2_decap_8 FILLER_64_1029 ();
 sg13g2_decap_4 FILLER_64_1036 ();
 sg13g2_fill_1 FILLER_64_1040 ();
 sg13g2_decap_8 FILLER_64_1056 ();
 sg13g2_decap_8 FILLER_64_1063 ();
 sg13g2_decap_8 FILLER_64_1070 ();
 sg13g2_fill_2 FILLER_64_1077 ();
 sg13g2_fill_2 FILLER_64_1084 ();
 sg13g2_decap_8 FILLER_64_1101 ();
 sg13g2_decap_8 FILLER_64_1108 ();
 sg13g2_decap_4 FILLER_64_1115 ();
 sg13g2_fill_2 FILLER_64_1119 ();
 sg13g2_decap_8 FILLER_64_1124 ();
 sg13g2_decap_8 FILLER_64_1131 ();
 sg13g2_decap_8 FILLER_64_1138 ();
 sg13g2_fill_1 FILLER_64_1145 ();
 sg13g2_decap_8 FILLER_64_1152 ();
 sg13g2_decap_8 FILLER_64_1159 ();
 sg13g2_decap_8 FILLER_64_1166 ();
 sg13g2_decap_8 FILLER_64_1173 ();
 sg13g2_decap_8 FILLER_64_1180 ();
 sg13g2_decap_8 FILLER_64_1187 ();
 sg13g2_decap_8 FILLER_64_1194 ();
 sg13g2_decap_8 FILLER_64_1201 ();
 sg13g2_decap_8 FILLER_64_1214 ();
 sg13g2_decap_8 FILLER_64_1221 ();
 sg13g2_fill_2 FILLER_64_1228 ();
 sg13g2_decap_8 FILLER_64_1243 ();
 sg13g2_decap_8 FILLER_64_1250 ();
 sg13g2_decap_8 FILLER_64_1257 ();
 sg13g2_decap_8 FILLER_64_1264 ();
 sg13g2_decap_8 FILLER_64_1271 ();
 sg13g2_decap_8 FILLER_64_1278 ();
 sg13g2_decap_8 FILLER_64_1285 ();
 sg13g2_decap_8 FILLER_64_1292 ();
 sg13g2_decap_8 FILLER_64_1299 ();
 sg13g2_decap_8 FILLER_64_1306 ();
 sg13g2_decap_8 FILLER_64_1313 ();
 sg13g2_decap_8 FILLER_64_1323 ();
 sg13g2_decap_8 FILLER_64_1330 ();
 sg13g2_decap_8 FILLER_64_1337 ();
 sg13g2_decap_8 FILLER_64_1344 ();
 sg13g2_decap_8 FILLER_64_1351 ();
 sg13g2_decap_8 FILLER_64_1358 ();
 sg13g2_decap_8 FILLER_64_1365 ();
 sg13g2_decap_8 FILLER_64_1372 ();
 sg13g2_decap_8 FILLER_64_1379 ();
 sg13g2_decap_8 FILLER_64_1386 ();
 sg13g2_decap_8 FILLER_64_1393 ();
 sg13g2_decap_8 FILLER_64_1400 ();
 sg13g2_decap_8 FILLER_64_1415 ();
 sg13g2_decap_8 FILLER_64_1422 ();
 sg13g2_decap_8 FILLER_64_1429 ();
 sg13g2_decap_8 FILLER_64_1436 ();
 sg13g2_decap_8 FILLER_64_1443 ();
 sg13g2_decap_8 FILLER_64_1450 ();
 sg13g2_decap_8 FILLER_64_1457 ();
 sg13g2_decap_8 FILLER_64_1464 ();
 sg13g2_decap_8 FILLER_64_1471 ();
 sg13g2_decap_8 FILLER_64_1478 ();
 sg13g2_fill_2 FILLER_64_1485 ();
 sg13g2_decap_4 FILLER_64_1493 ();
 sg13g2_fill_2 FILLER_64_1497 ();
 sg13g2_fill_1 FILLER_64_1511 ();
 sg13g2_decap_8 FILLER_64_1525 ();
 sg13g2_decap_8 FILLER_64_1532 ();
 sg13g2_decap_8 FILLER_64_1539 ();
 sg13g2_decap_8 FILLER_64_1546 ();
 sg13g2_decap_8 FILLER_64_1553 ();
 sg13g2_decap_8 FILLER_64_1560 ();
 sg13g2_decap_8 FILLER_64_1567 ();
 sg13g2_fill_1 FILLER_64_1574 ();
 sg13g2_decap_8 FILLER_64_1578 ();
 sg13g2_decap_8 FILLER_64_1585 ();
 sg13g2_decap_8 FILLER_64_1592 ();
 sg13g2_decap_8 FILLER_64_1599 ();
 sg13g2_decap_8 FILLER_64_1606 ();
 sg13g2_decap_8 FILLER_64_1613 ();
 sg13g2_decap_8 FILLER_64_1620 ();
 sg13g2_decap_8 FILLER_64_1627 ();
 sg13g2_decap_8 FILLER_64_1634 ();
 sg13g2_fill_1 FILLER_64_1641 ();
 sg13g2_decap_8 FILLER_64_1650 ();
 sg13g2_decap_8 FILLER_64_1657 ();
 sg13g2_decap_8 FILLER_64_1664 ();
 sg13g2_decap_8 FILLER_64_1671 ();
 sg13g2_decap_8 FILLER_64_1678 ();
 sg13g2_decap_8 FILLER_64_1685 ();
 sg13g2_decap_8 FILLER_64_1692 ();
 sg13g2_decap_8 FILLER_64_1699 ();
 sg13g2_decap_8 FILLER_64_1706 ();
 sg13g2_decap_8 FILLER_64_1713 ();
 sg13g2_decap_8 FILLER_64_1720 ();
 sg13g2_decap_8 FILLER_64_1727 ();
 sg13g2_decap_8 FILLER_64_1734 ();
 sg13g2_decap_4 FILLER_64_1741 ();
 sg13g2_fill_2 FILLER_64_1745 ();
 sg13g2_decap_8 FILLER_64_1762 ();
 sg13g2_decap_8 FILLER_64_1769 ();
 sg13g2_decap_8 FILLER_64_1776 ();
 sg13g2_decap_8 FILLER_64_1783 ();
 sg13g2_decap_8 FILLER_64_1790 ();
 sg13g2_decap_8 FILLER_64_1797 ();
 sg13g2_decap_8 FILLER_64_1804 ();
 sg13g2_decap_8 FILLER_64_1811 ();
 sg13g2_decap_8 FILLER_64_1818 ();
 sg13g2_decap_8 FILLER_64_1825 ();
 sg13g2_decap_8 FILLER_64_1832 ();
 sg13g2_decap_8 FILLER_64_1839 ();
 sg13g2_decap_8 FILLER_64_1846 ();
 sg13g2_decap_8 FILLER_64_1853 ();
 sg13g2_decap_8 FILLER_64_1860 ();
 sg13g2_decap_8 FILLER_64_1867 ();
 sg13g2_decap_8 FILLER_64_1874 ();
 sg13g2_decap_8 FILLER_64_1881 ();
 sg13g2_decap_8 FILLER_64_1888 ();
 sg13g2_decap_8 FILLER_64_1895 ();
 sg13g2_decap_8 FILLER_64_1902 ();
 sg13g2_decap_8 FILLER_64_1909 ();
 sg13g2_decap_8 FILLER_64_1916 ();
 sg13g2_decap_8 FILLER_64_1923 ();
 sg13g2_decap_8 FILLER_64_1930 ();
 sg13g2_decap_8 FILLER_64_1937 ();
 sg13g2_decap_8 FILLER_64_1944 ();
 sg13g2_decap_8 FILLER_64_1951 ();
 sg13g2_decap_4 FILLER_64_1958 ();
 sg13g2_fill_2 FILLER_64_1962 ();
 sg13g2_decap_8 FILLER_64_1974 ();
 sg13g2_decap_8 FILLER_64_1981 ();
 sg13g2_decap_8 FILLER_64_1988 ();
 sg13g2_decap_8 FILLER_64_1995 ();
 sg13g2_decap_8 FILLER_64_2002 ();
 sg13g2_decap_8 FILLER_64_2009 ();
 sg13g2_decap_8 FILLER_64_2016 ();
 sg13g2_decap_8 FILLER_64_2023 ();
 sg13g2_decap_8 FILLER_64_2030 ();
 sg13g2_decap_8 FILLER_64_2037 ();
 sg13g2_decap_8 FILLER_64_2044 ();
 sg13g2_decap_8 FILLER_64_2051 ();
 sg13g2_decap_8 FILLER_64_2058 ();
 sg13g2_fill_2 FILLER_64_2065 ();
 sg13g2_decap_8 FILLER_64_2070 ();
 sg13g2_decap_8 FILLER_64_2077 ();
 sg13g2_decap_8 FILLER_64_2084 ();
 sg13g2_decap_8 FILLER_64_2091 ();
 sg13g2_fill_1 FILLER_64_2098 ();
 sg13g2_decap_8 FILLER_64_2125 ();
 sg13g2_decap_8 FILLER_64_2132 ();
 sg13g2_decap_8 FILLER_64_2139 ();
 sg13g2_decap_8 FILLER_64_2146 ();
 sg13g2_decap_8 FILLER_64_2153 ();
 sg13g2_decap_8 FILLER_64_2160 ();
 sg13g2_decap_8 FILLER_64_2167 ();
 sg13g2_decap_8 FILLER_64_2174 ();
 sg13g2_decap_4 FILLER_64_2181 ();
 sg13g2_fill_1 FILLER_64_2185 ();
 sg13g2_decap_8 FILLER_64_2190 ();
 sg13g2_decap_8 FILLER_64_2197 ();
 sg13g2_decap_8 FILLER_64_2204 ();
 sg13g2_decap_8 FILLER_64_2211 ();
 sg13g2_decap_8 FILLER_64_2218 ();
 sg13g2_decap_8 FILLER_64_2225 ();
 sg13g2_decap_8 FILLER_64_2232 ();
 sg13g2_decap_8 FILLER_64_2239 ();
 sg13g2_decap_8 FILLER_64_2246 ();
 sg13g2_decap_8 FILLER_64_2253 ();
 sg13g2_decap_8 FILLER_64_2260 ();
 sg13g2_decap_8 FILLER_64_2267 ();
 sg13g2_decap_8 FILLER_64_2274 ();
 sg13g2_decap_8 FILLER_64_2281 ();
 sg13g2_decap_8 FILLER_64_2288 ();
 sg13g2_decap_8 FILLER_64_2295 ();
 sg13g2_decap_8 FILLER_64_2302 ();
 sg13g2_decap_8 FILLER_64_2309 ();
 sg13g2_decap_8 FILLER_64_2316 ();
 sg13g2_decap_8 FILLER_64_2323 ();
 sg13g2_decap_8 FILLER_64_2330 ();
 sg13g2_decap_8 FILLER_64_2337 ();
 sg13g2_decap_8 FILLER_64_2344 ();
 sg13g2_decap_8 FILLER_64_2351 ();
 sg13g2_decap_8 FILLER_64_2358 ();
 sg13g2_decap_8 FILLER_64_2365 ();
 sg13g2_decap_8 FILLER_64_2372 ();
 sg13g2_decap_8 FILLER_64_2379 ();
 sg13g2_decap_8 FILLER_64_2386 ();
 sg13g2_decap_8 FILLER_64_2393 ();
 sg13g2_decap_8 FILLER_64_2400 ();
 sg13g2_decap_8 FILLER_64_2407 ();
 sg13g2_decap_8 FILLER_64_2414 ();
 sg13g2_decap_8 FILLER_64_2421 ();
 sg13g2_decap_8 FILLER_64_2428 ();
 sg13g2_decap_8 FILLER_64_2435 ();
 sg13g2_decap_8 FILLER_64_2442 ();
 sg13g2_decap_8 FILLER_64_2449 ();
 sg13g2_decap_8 FILLER_64_2456 ();
 sg13g2_decap_8 FILLER_64_2463 ();
 sg13g2_decap_8 FILLER_64_2470 ();
 sg13g2_decap_8 FILLER_64_2477 ();
 sg13g2_decap_8 FILLER_64_2484 ();
 sg13g2_decap_8 FILLER_64_2491 ();
 sg13g2_decap_8 FILLER_64_2498 ();
 sg13g2_decap_8 FILLER_64_2505 ();
 sg13g2_decap_8 FILLER_64_2512 ();
 sg13g2_decap_8 FILLER_64_2519 ();
 sg13g2_decap_8 FILLER_64_2526 ();
 sg13g2_decap_8 FILLER_64_2533 ();
 sg13g2_decap_8 FILLER_64_2540 ();
 sg13g2_decap_8 FILLER_64_2547 ();
 sg13g2_decap_8 FILLER_64_2554 ();
 sg13g2_decap_8 FILLER_64_2561 ();
 sg13g2_decap_8 FILLER_64_2568 ();
 sg13g2_decap_8 FILLER_64_2575 ();
 sg13g2_decap_8 FILLER_64_2582 ();
 sg13g2_decap_8 FILLER_64_2589 ();
 sg13g2_decap_8 FILLER_64_2596 ();
 sg13g2_decap_8 FILLER_64_2603 ();
 sg13g2_decap_8 FILLER_64_2610 ();
 sg13g2_decap_8 FILLER_64_2617 ();
 sg13g2_decap_8 FILLER_64_2624 ();
 sg13g2_decap_8 FILLER_64_2631 ();
 sg13g2_decap_8 FILLER_64_2638 ();
 sg13g2_decap_8 FILLER_64_2645 ();
 sg13g2_decap_8 FILLER_64_2652 ();
 sg13g2_decap_8 FILLER_64_2659 ();
 sg13g2_decap_4 FILLER_64_2666 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_64 ();
 sg13g2_decap_4 FILLER_65_71 ();
 sg13g2_fill_1 FILLER_65_79 ();
 sg13g2_decap_8 FILLER_65_85 ();
 sg13g2_decap_8 FILLER_65_92 ();
 sg13g2_decap_8 FILLER_65_99 ();
 sg13g2_decap_8 FILLER_65_106 ();
 sg13g2_decap_4 FILLER_65_113 ();
 sg13g2_fill_1 FILLER_65_117 ();
 sg13g2_decap_8 FILLER_65_122 ();
 sg13g2_decap_8 FILLER_65_129 ();
 sg13g2_decap_8 FILLER_65_136 ();
 sg13g2_decap_8 FILLER_65_143 ();
 sg13g2_decap_8 FILLER_65_150 ();
 sg13g2_decap_8 FILLER_65_157 ();
 sg13g2_decap_4 FILLER_65_164 ();
 sg13g2_fill_1 FILLER_65_168 ();
 sg13g2_decap_8 FILLER_65_173 ();
 sg13g2_decap_4 FILLER_65_180 ();
 sg13g2_fill_2 FILLER_65_184 ();
 sg13g2_fill_2 FILLER_65_191 ();
 sg13g2_fill_1 FILLER_65_193 ();
 sg13g2_decap_8 FILLER_65_198 ();
 sg13g2_decap_8 FILLER_65_205 ();
 sg13g2_decap_8 FILLER_65_212 ();
 sg13g2_decap_8 FILLER_65_219 ();
 sg13g2_decap_8 FILLER_65_226 ();
 sg13g2_decap_8 FILLER_65_233 ();
 sg13g2_decap_8 FILLER_65_240 ();
 sg13g2_decap_8 FILLER_65_247 ();
 sg13g2_decap_8 FILLER_65_254 ();
 sg13g2_decap_8 FILLER_65_261 ();
 sg13g2_decap_8 FILLER_65_268 ();
 sg13g2_decap_8 FILLER_65_275 ();
 sg13g2_decap_8 FILLER_65_282 ();
 sg13g2_decap_8 FILLER_65_289 ();
 sg13g2_decap_8 FILLER_65_296 ();
 sg13g2_decap_8 FILLER_65_303 ();
 sg13g2_decap_4 FILLER_65_310 ();
 sg13g2_decap_8 FILLER_65_343 ();
 sg13g2_decap_8 FILLER_65_350 ();
 sg13g2_decap_8 FILLER_65_357 ();
 sg13g2_decap_8 FILLER_65_364 ();
 sg13g2_decap_8 FILLER_65_371 ();
 sg13g2_decap_8 FILLER_65_378 ();
 sg13g2_fill_1 FILLER_65_385 ();
 sg13g2_decap_8 FILLER_65_404 ();
 sg13g2_decap_8 FILLER_65_411 ();
 sg13g2_decap_8 FILLER_65_418 ();
 sg13g2_decap_8 FILLER_65_425 ();
 sg13g2_decap_8 FILLER_65_432 ();
 sg13g2_decap_8 FILLER_65_439 ();
 sg13g2_fill_2 FILLER_65_446 ();
 sg13g2_fill_1 FILLER_65_448 ();
 sg13g2_decap_8 FILLER_65_473 ();
 sg13g2_decap_8 FILLER_65_480 ();
 sg13g2_fill_1 FILLER_65_487 ();
 sg13g2_decap_8 FILLER_65_493 ();
 sg13g2_decap_8 FILLER_65_500 ();
 sg13g2_decap_8 FILLER_65_507 ();
 sg13g2_decap_8 FILLER_65_514 ();
 sg13g2_decap_8 FILLER_65_521 ();
 sg13g2_decap_8 FILLER_65_528 ();
 sg13g2_decap_8 FILLER_65_535 ();
 sg13g2_fill_2 FILLER_65_542 ();
 sg13g2_fill_1 FILLER_65_544 ();
 sg13g2_decap_4 FILLER_65_549 ();
 sg13g2_decap_8 FILLER_65_557 ();
 sg13g2_decap_8 FILLER_65_564 ();
 sg13g2_fill_2 FILLER_65_571 ();
 sg13g2_decap_4 FILLER_65_578 ();
 sg13g2_decap_8 FILLER_65_587 ();
 sg13g2_decap_8 FILLER_65_594 ();
 sg13g2_decap_8 FILLER_65_601 ();
 sg13g2_decap_8 FILLER_65_608 ();
 sg13g2_decap_8 FILLER_65_615 ();
 sg13g2_decap_8 FILLER_65_622 ();
 sg13g2_decap_8 FILLER_65_629 ();
 sg13g2_decap_8 FILLER_65_636 ();
 sg13g2_decap_8 FILLER_65_643 ();
 sg13g2_decap_8 FILLER_65_650 ();
 sg13g2_fill_1 FILLER_65_657 ();
 sg13g2_decap_8 FILLER_65_661 ();
 sg13g2_decap_8 FILLER_65_668 ();
 sg13g2_decap_8 FILLER_65_675 ();
 sg13g2_decap_8 FILLER_65_690 ();
 sg13g2_decap_8 FILLER_65_697 ();
 sg13g2_decap_8 FILLER_65_704 ();
 sg13g2_decap_8 FILLER_65_711 ();
 sg13g2_decap_8 FILLER_65_718 ();
 sg13g2_decap_8 FILLER_65_725 ();
 sg13g2_decap_8 FILLER_65_732 ();
 sg13g2_decap_8 FILLER_65_739 ();
 sg13g2_decap_8 FILLER_65_746 ();
 sg13g2_decap_8 FILLER_65_753 ();
 sg13g2_decap_8 FILLER_65_760 ();
 sg13g2_decap_8 FILLER_65_767 ();
 sg13g2_decap_8 FILLER_65_774 ();
 sg13g2_decap_8 FILLER_65_781 ();
 sg13g2_decap_8 FILLER_65_788 ();
 sg13g2_decap_8 FILLER_65_795 ();
 sg13g2_decap_8 FILLER_65_802 ();
 sg13g2_fill_2 FILLER_65_809 ();
 sg13g2_decap_8 FILLER_65_815 ();
 sg13g2_decap_8 FILLER_65_822 ();
 sg13g2_decap_8 FILLER_65_829 ();
 sg13g2_decap_8 FILLER_65_836 ();
 sg13g2_decap_8 FILLER_65_843 ();
 sg13g2_decap_8 FILLER_65_850 ();
 sg13g2_decap_8 FILLER_65_857 ();
 sg13g2_decap_8 FILLER_65_864 ();
 sg13g2_decap_8 FILLER_65_871 ();
 sg13g2_decap_8 FILLER_65_878 ();
 sg13g2_decap_8 FILLER_65_885 ();
 sg13g2_decap_8 FILLER_65_892 ();
 sg13g2_fill_1 FILLER_65_899 ();
 sg13g2_decap_4 FILLER_65_905 ();
 sg13g2_fill_1 FILLER_65_909 ();
 sg13g2_decap_8 FILLER_65_914 ();
 sg13g2_decap_8 FILLER_65_921 ();
 sg13g2_decap_8 FILLER_65_928 ();
 sg13g2_decap_8 FILLER_65_935 ();
 sg13g2_decap_8 FILLER_65_942 ();
 sg13g2_decap_8 FILLER_65_949 ();
 sg13g2_decap_8 FILLER_65_956 ();
 sg13g2_decap_8 FILLER_65_963 ();
 sg13g2_decap_8 FILLER_65_970 ();
 sg13g2_decap_8 FILLER_65_977 ();
 sg13g2_decap_8 FILLER_65_984 ();
 sg13g2_decap_8 FILLER_65_991 ();
 sg13g2_decap_8 FILLER_65_998 ();
 sg13g2_decap_8 FILLER_65_1005 ();
 sg13g2_decap_8 FILLER_65_1012 ();
 sg13g2_decap_8 FILLER_65_1019 ();
 sg13g2_decap_8 FILLER_65_1026 ();
 sg13g2_decap_8 FILLER_65_1033 ();
 sg13g2_fill_1 FILLER_65_1040 ();
 sg13g2_decap_8 FILLER_65_1049 ();
 sg13g2_decap_8 FILLER_65_1056 ();
 sg13g2_decap_8 FILLER_65_1063 ();
 sg13g2_decap_8 FILLER_65_1070 ();
 sg13g2_decap_8 FILLER_65_1077 ();
 sg13g2_fill_2 FILLER_65_1084 ();
 sg13g2_decap_8 FILLER_65_1089 ();
 sg13g2_fill_2 FILLER_65_1096 ();
 sg13g2_decap_8 FILLER_65_1113 ();
 sg13g2_decap_8 FILLER_65_1120 ();
 sg13g2_decap_8 FILLER_65_1127 ();
 sg13g2_decap_8 FILLER_65_1134 ();
 sg13g2_decap_4 FILLER_65_1141 ();
 sg13g2_fill_2 FILLER_65_1145 ();
 sg13g2_decap_8 FILLER_65_1150 ();
 sg13g2_decap_8 FILLER_65_1157 ();
 sg13g2_decap_8 FILLER_65_1164 ();
 sg13g2_decap_8 FILLER_65_1171 ();
 sg13g2_decap_8 FILLER_65_1178 ();
 sg13g2_decap_8 FILLER_65_1185 ();
 sg13g2_decap_8 FILLER_65_1192 ();
 sg13g2_decap_8 FILLER_65_1199 ();
 sg13g2_decap_8 FILLER_65_1206 ();
 sg13g2_decap_8 FILLER_65_1213 ();
 sg13g2_decap_8 FILLER_65_1220 ();
 sg13g2_decap_8 FILLER_65_1227 ();
 sg13g2_decap_4 FILLER_65_1234 ();
 sg13g2_decap_8 FILLER_65_1241 ();
 sg13g2_fill_1 FILLER_65_1248 ();
 sg13g2_decap_4 FILLER_65_1254 ();
 sg13g2_fill_2 FILLER_65_1258 ();
 sg13g2_decap_8 FILLER_65_1279 ();
 sg13g2_decap_8 FILLER_65_1286 ();
 sg13g2_decap_8 FILLER_65_1293 ();
 sg13g2_decap_4 FILLER_65_1300 ();
 sg13g2_fill_2 FILLER_65_1304 ();
 sg13g2_decap_8 FILLER_65_1311 ();
 sg13g2_fill_2 FILLER_65_1318 ();
 sg13g2_fill_1 FILLER_65_1324 ();
 sg13g2_decap_8 FILLER_65_1336 ();
 sg13g2_decap_8 FILLER_65_1343 ();
 sg13g2_decap_4 FILLER_65_1350 ();
 sg13g2_decap_8 FILLER_65_1374 ();
 sg13g2_decap_8 FILLER_65_1381 ();
 sg13g2_decap_8 FILLER_65_1392 ();
 sg13g2_decap_4 FILLER_65_1399 ();
 sg13g2_decap_4 FILLER_65_1408 ();
 sg13g2_fill_2 FILLER_65_1412 ();
 sg13g2_decap_8 FILLER_65_1418 ();
 sg13g2_decap_4 FILLER_65_1425 ();
 sg13g2_fill_2 FILLER_65_1429 ();
 sg13g2_decap_8 FILLER_65_1435 ();
 sg13g2_decap_8 FILLER_65_1442 ();
 sg13g2_decap_4 FILLER_65_1449 ();
 sg13g2_fill_2 FILLER_65_1453 ();
 sg13g2_fill_2 FILLER_65_1458 ();
 sg13g2_decap_4 FILLER_65_1466 ();
 sg13g2_fill_2 FILLER_65_1470 ();
 sg13g2_decap_8 FILLER_65_1478 ();
 sg13g2_decap_8 FILLER_65_1485 ();
 sg13g2_decap_8 FILLER_65_1492 ();
 sg13g2_decap_4 FILLER_65_1499 ();
 sg13g2_fill_2 FILLER_65_1503 ();
 sg13g2_decap_8 FILLER_65_1525 ();
 sg13g2_decap_8 FILLER_65_1532 ();
 sg13g2_decap_8 FILLER_65_1539 ();
 sg13g2_decap_8 FILLER_65_1546 ();
 sg13g2_fill_1 FILLER_65_1553 ();
 sg13g2_decap_8 FILLER_65_1559 ();
 sg13g2_decap_4 FILLER_65_1566 ();
 sg13g2_decap_8 FILLER_65_1574 ();
 sg13g2_decap_4 FILLER_65_1581 ();
 sg13g2_fill_2 FILLER_65_1585 ();
 sg13g2_decap_8 FILLER_65_1591 ();
 sg13g2_decap_8 FILLER_65_1598 ();
 sg13g2_decap_4 FILLER_65_1605 ();
 sg13g2_decap_8 FILLER_65_1624 ();
 sg13g2_decap_8 FILLER_65_1631 ();
 sg13g2_decap_8 FILLER_65_1638 ();
 sg13g2_fill_1 FILLER_65_1645 ();
 sg13g2_decap_8 FILLER_65_1650 ();
 sg13g2_decap_8 FILLER_65_1657 ();
 sg13g2_decap_8 FILLER_65_1664 ();
 sg13g2_decap_8 FILLER_65_1671 ();
 sg13g2_decap_8 FILLER_65_1678 ();
 sg13g2_decap_8 FILLER_65_1685 ();
 sg13g2_fill_2 FILLER_65_1692 ();
 sg13g2_fill_1 FILLER_65_1694 ();
 sg13g2_decap_4 FILLER_65_1700 ();
 sg13g2_fill_2 FILLER_65_1704 ();
 sg13g2_decap_8 FILLER_65_1710 ();
 sg13g2_decap_8 FILLER_65_1717 ();
 sg13g2_decap_8 FILLER_65_1724 ();
 sg13g2_decap_4 FILLER_65_1731 ();
 sg13g2_fill_1 FILLER_65_1735 ();
 sg13g2_decap_4 FILLER_65_1741 ();
 sg13g2_fill_2 FILLER_65_1745 ();
 sg13g2_decap_8 FILLER_65_1751 ();
 sg13g2_decap_8 FILLER_65_1758 ();
 sg13g2_decap_4 FILLER_65_1765 ();
 sg13g2_decap_8 FILLER_65_1808 ();
 sg13g2_decap_8 FILLER_65_1815 ();
 sg13g2_decap_8 FILLER_65_1822 ();
 sg13g2_decap_8 FILLER_65_1829 ();
 sg13g2_decap_8 FILLER_65_1836 ();
 sg13g2_decap_8 FILLER_65_1843 ();
 sg13g2_decap_8 FILLER_65_1850 ();
 sg13g2_decap_8 FILLER_65_1857 ();
 sg13g2_decap_8 FILLER_65_1864 ();
 sg13g2_decap_8 FILLER_65_1871 ();
 sg13g2_decap_8 FILLER_65_1878 ();
 sg13g2_decap_8 FILLER_65_1885 ();
 sg13g2_decap_8 FILLER_65_1892 ();
 sg13g2_decap_8 FILLER_65_1899 ();
 sg13g2_decap_8 FILLER_65_1906 ();
 sg13g2_decap_8 FILLER_65_1913 ();
 sg13g2_decap_8 FILLER_65_1920 ();
 sg13g2_decap_8 FILLER_65_1927 ();
 sg13g2_decap_8 FILLER_65_1934 ();
 sg13g2_decap_8 FILLER_65_1941 ();
 sg13g2_decap_8 FILLER_65_1948 ();
 sg13g2_decap_8 FILLER_65_1955 ();
 sg13g2_decap_8 FILLER_65_1962 ();
 sg13g2_decap_4 FILLER_65_1969 ();
 sg13g2_decap_8 FILLER_65_1976 ();
 sg13g2_decap_8 FILLER_65_1983 ();
 sg13g2_decap_8 FILLER_65_1990 ();
 sg13g2_decap_8 FILLER_65_1997 ();
 sg13g2_decap_8 FILLER_65_2004 ();
 sg13g2_decap_8 FILLER_65_2011 ();
 sg13g2_fill_1 FILLER_65_2018 ();
 sg13g2_decap_8 FILLER_65_2023 ();
 sg13g2_decap_8 FILLER_65_2030 ();
 sg13g2_decap_8 FILLER_65_2037 ();
 sg13g2_decap_8 FILLER_65_2044 ();
 sg13g2_decap_8 FILLER_65_2051 ();
 sg13g2_fill_2 FILLER_65_2058 ();
 sg13g2_fill_1 FILLER_65_2060 ();
 sg13g2_decap_8 FILLER_65_2065 ();
 sg13g2_decap_8 FILLER_65_2072 ();
 sg13g2_decap_8 FILLER_65_2079 ();
 sg13g2_decap_8 FILLER_65_2086 ();
 sg13g2_decap_8 FILLER_65_2093 ();
 sg13g2_decap_8 FILLER_65_2100 ();
 sg13g2_decap_8 FILLER_65_2107 ();
 sg13g2_decap_8 FILLER_65_2114 ();
 sg13g2_decap_8 FILLER_65_2121 ();
 sg13g2_decap_8 FILLER_65_2128 ();
 sg13g2_decap_8 FILLER_65_2135 ();
 sg13g2_fill_1 FILLER_65_2142 ();
 sg13g2_fill_1 FILLER_65_2157 ();
 sg13g2_decap_8 FILLER_65_2161 ();
 sg13g2_decap_8 FILLER_65_2168 ();
 sg13g2_decap_8 FILLER_65_2175 ();
 sg13g2_fill_1 FILLER_65_2182 ();
 sg13g2_decap_8 FILLER_65_2191 ();
 sg13g2_decap_8 FILLER_65_2198 ();
 sg13g2_decap_8 FILLER_65_2205 ();
 sg13g2_decap_8 FILLER_65_2212 ();
 sg13g2_decap_8 FILLER_65_2219 ();
 sg13g2_fill_1 FILLER_65_2226 ();
 sg13g2_decap_8 FILLER_65_2230 ();
 sg13g2_decap_8 FILLER_65_2237 ();
 sg13g2_decap_8 FILLER_65_2244 ();
 sg13g2_decap_8 FILLER_65_2251 ();
 sg13g2_decap_8 FILLER_65_2258 ();
 sg13g2_decap_8 FILLER_65_2265 ();
 sg13g2_decap_8 FILLER_65_2272 ();
 sg13g2_decap_8 FILLER_65_2279 ();
 sg13g2_decap_8 FILLER_65_2286 ();
 sg13g2_decap_8 FILLER_65_2293 ();
 sg13g2_decap_8 FILLER_65_2300 ();
 sg13g2_decap_8 FILLER_65_2307 ();
 sg13g2_decap_8 FILLER_65_2314 ();
 sg13g2_decap_8 FILLER_65_2321 ();
 sg13g2_decap_8 FILLER_65_2328 ();
 sg13g2_decap_8 FILLER_65_2335 ();
 sg13g2_decap_8 FILLER_65_2342 ();
 sg13g2_decap_8 FILLER_65_2349 ();
 sg13g2_decap_8 FILLER_65_2356 ();
 sg13g2_decap_8 FILLER_65_2363 ();
 sg13g2_decap_8 FILLER_65_2370 ();
 sg13g2_decap_8 FILLER_65_2377 ();
 sg13g2_decap_8 FILLER_65_2384 ();
 sg13g2_decap_8 FILLER_65_2391 ();
 sg13g2_decap_8 FILLER_65_2398 ();
 sg13g2_decap_8 FILLER_65_2405 ();
 sg13g2_decap_8 FILLER_65_2412 ();
 sg13g2_decap_8 FILLER_65_2419 ();
 sg13g2_decap_8 FILLER_65_2426 ();
 sg13g2_decap_8 FILLER_65_2433 ();
 sg13g2_decap_8 FILLER_65_2440 ();
 sg13g2_decap_8 FILLER_65_2447 ();
 sg13g2_decap_8 FILLER_65_2454 ();
 sg13g2_decap_8 FILLER_65_2461 ();
 sg13g2_decap_8 FILLER_65_2468 ();
 sg13g2_decap_8 FILLER_65_2475 ();
 sg13g2_decap_8 FILLER_65_2482 ();
 sg13g2_decap_8 FILLER_65_2489 ();
 sg13g2_decap_8 FILLER_65_2496 ();
 sg13g2_decap_8 FILLER_65_2503 ();
 sg13g2_decap_8 FILLER_65_2510 ();
 sg13g2_decap_8 FILLER_65_2517 ();
 sg13g2_decap_8 FILLER_65_2524 ();
 sg13g2_decap_8 FILLER_65_2531 ();
 sg13g2_decap_8 FILLER_65_2538 ();
 sg13g2_decap_8 FILLER_65_2545 ();
 sg13g2_decap_8 FILLER_65_2552 ();
 sg13g2_decap_8 FILLER_65_2559 ();
 sg13g2_decap_8 FILLER_65_2566 ();
 sg13g2_decap_8 FILLER_65_2573 ();
 sg13g2_decap_8 FILLER_65_2580 ();
 sg13g2_decap_8 FILLER_65_2587 ();
 sg13g2_decap_8 FILLER_65_2594 ();
 sg13g2_decap_8 FILLER_65_2601 ();
 sg13g2_decap_8 FILLER_65_2608 ();
 sg13g2_decap_8 FILLER_65_2615 ();
 sg13g2_decap_8 FILLER_65_2622 ();
 sg13g2_decap_8 FILLER_65_2629 ();
 sg13g2_decap_8 FILLER_65_2636 ();
 sg13g2_decap_8 FILLER_65_2643 ();
 sg13g2_decap_8 FILLER_65_2650 ();
 sg13g2_decap_8 FILLER_65_2657 ();
 sg13g2_decap_4 FILLER_65_2664 ();
 sg13g2_fill_2 FILLER_65_2668 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_4 FILLER_66_70 ();
 sg13g2_fill_1 FILLER_66_74 ();
 sg13g2_decap_8 FILLER_66_86 ();
 sg13g2_decap_8 FILLER_66_93 ();
 sg13g2_decap_8 FILLER_66_100 ();
 sg13g2_decap_8 FILLER_66_107 ();
 sg13g2_decap_8 FILLER_66_124 ();
 sg13g2_decap_8 FILLER_66_131 ();
 sg13g2_decap_8 FILLER_66_138 ();
 sg13g2_decap_4 FILLER_66_145 ();
 sg13g2_fill_1 FILLER_66_149 ();
 sg13g2_decap_4 FILLER_66_155 ();
 sg13g2_decap_4 FILLER_66_168 ();
 sg13g2_fill_1 FILLER_66_172 ();
 sg13g2_decap_8 FILLER_66_177 ();
 sg13g2_decap_8 FILLER_66_184 ();
 sg13g2_decap_8 FILLER_66_191 ();
 sg13g2_decap_8 FILLER_66_198 ();
 sg13g2_decap_8 FILLER_66_205 ();
 sg13g2_decap_8 FILLER_66_212 ();
 sg13g2_decap_8 FILLER_66_219 ();
 sg13g2_decap_8 FILLER_66_226 ();
 sg13g2_decap_8 FILLER_66_233 ();
 sg13g2_decap_8 FILLER_66_240 ();
 sg13g2_decap_8 FILLER_66_247 ();
 sg13g2_fill_1 FILLER_66_266 ();
 sg13g2_decap_8 FILLER_66_274 ();
 sg13g2_decap_8 FILLER_66_281 ();
 sg13g2_decap_8 FILLER_66_288 ();
 sg13g2_decap_8 FILLER_66_295 ();
 sg13g2_decap_8 FILLER_66_302 ();
 sg13g2_decap_8 FILLER_66_309 ();
 sg13g2_decap_8 FILLER_66_316 ();
 sg13g2_decap_8 FILLER_66_323 ();
 sg13g2_decap_8 FILLER_66_330 ();
 sg13g2_decap_8 FILLER_66_337 ();
 sg13g2_decap_8 FILLER_66_344 ();
 sg13g2_decap_8 FILLER_66_351 ();
 sg13g2_decap_8 FILLER_66_358 ();
 sg13g2_decap_8 FILLER_66_365 ();
 sg13g2_fill_2 FILLER_66_372 ();
 sg13g2_fill_1 FILLER_66_397 ();
 sg13g2_decap_8 FILLER_66_410 ();
 sg13g2_decap_8 FILLER_66_417 ();
 sg13g2_decap_4 FILLER_66_424 ();
 sg13g2_decap_8 FILLER_66_452 ();
 sg13g2_decap_8 FILLER_66_459 ();
 sg13g2_decap_8 FILLER_66_466 ();
 sg13g2_decap_8 FILLER_66_473 ();
 sg13g2_decap_8 FILLER_66_480 ();
 sg13g2_decap_8 FILLER_66_491 ();
 sg13g2_decap_8 FILLER_66_498 ();
 sg13g2_decap_8 FILLER_66_505 ();
 sg13g2_decap_4 FILLER_66_512 ();
 sg13g2_decap_8 FILLER_66_521 ();
 sg13g2_decap_8 FILLER_66_528 ();
 sg13g2_decap_8 FILLER_66_535 ();
 sg13g2_decap_8 FILLER_66_542 ();
 sg13g2_decap_4 FILLER_66_549 ();
 sg13g2_fill_2 FILLER_66_553 ();
 sg13g2_decap_8 FILLER_66_560 ();
 sg13g2_decap_4 FILLER_66_567 ();
 sg13g2_fill_2 FILLER_66_571 ();
 sg13g2_decap_8 FILLER_66_576 ();
 sg13g2_decap_8 FILLER_66_583 ();
 sg13g2_decap_8 FILLER_66_590 ();
 sg13g2_decap_8 FILLER_66_597 ();
 sg13g2_decap_8 FILLER_66_604 ();
 sg13g2_fill_2 FILLER_66_611 ();
 sg13g2_decap_8 FILLER_66_631 ();
 sg13g2_decap_8 FILLER_66_638 ();
 sg13g2_decap_8 FILLER_66_645 ();
 sg13g2_decap_8 FILLER_66_670 ();
 sg13g2_decap_4 FILLER_66_677 ();
 sg13g2_fill_1 FILLER_66_681 ();
 sg13g2_decap_8 FILLER_66_693 ();
 sg13g2_decap_8 FILLER_66_700 ();
 sg13g2_decap_8 FILLER_66_707 ();
 sg13g2_decap_8 FILLER_66_714 ();
 sg13g2_decap_4 FILLER_66_721 ();
 sg13g2_fill_2 FILLER_66_725 ();
 sg13g2_fill_2 FILLER_66_731 ();
 sg13g2_decap_8 FILLER_66_737 ();
 sg13g2_decap_8 FILLER_66_744 ();
 sg13g2_decap_8 FILLER_66_751 ();
 sg13g2_decap_8 FILLER_66_758 ();
 sg13g2_decap_8 FILLER_66_765 ();
 sg13g2_decap_8 FILLER_66_772 ();
 sg13g2_decap_8 FILLER_66_787 ();
 sg13g2_decap_8 FILLER_66_794 ();
 sg13g2_decap_8 FILLER_66_801 ();
 sg13g2_fill_2 FILLER_66_808 ();
 sg13g2_decap_8 FILLER_66_815 ();
 sg13g2_decap_8 FILLER_66_822 ();
 sg13g2_decap_8 FILLER_66_829 ();
 sg13g2_decap_8 FILLER_66_836 ();
 sg13g2_decap_8 FILLER_66_843 ();
 sg13g2_decap_8 FILLER_66_850 ();
 sg13g2_decap_8 FILLER_66_857 ();
 sg13g2_decap_8 FILLER_66_864 ();
 sg13g2_decap_8 FILLER_66_871 ();
 sg13g2_decap_8 FILLER_66_878 ();
 sg13g2_decap_8 FILLER_66_885 ();
 sg13g2_decap_8 FILLER_66_892 ();
 sg13g2_decap_8 FILLER_66_899 ();
 sg13g2_decap_8 FILLER_66_906 ();
 sg13g2_decap_8 FILLER_66_913 ();
 sg13g2_decap_8 FILLER_66_920 ();
 sg13g2_decap_4 FILLER_66_927 ();
 sg13g2_fill_1 FILLER_66_931 ();
 sg13g2_decap_8 FILLER_66_935 ();
 sg13g2_decap_8 FILLER_66_942 ();
 sg13g2_decap_8 FILLER_66_949 ();
 sg13g2_decap_8 FILLER_66_956 ();
 sg13g2_decap_8 FILLER_66_963 ();
 sg13g2_decap_8 FILLER_66_970 ();
 sg13g2_decap_8 FILLER_66_977 ();
 sg13g2_decap_8 FILLER_66_984 ();
 sg13g2_decap_8 FILLER_66_991 ();
 sg13g2_decap_8 FILLER_66_998 ();
 sg13g2_fill_2 FILLER_66_1005 ();
 sg13g2_decap_8 FILLER_66_1020 ();
 sg13g2_decap_8 FILLER_66_1027 ();
 sg13g2_fill_1 FILLER_66_1034 ();
 sg13g2_fill_2 FILLER_66_1039 ();
 sg13g2_decap_8 FILLER_66_1053 ();
 sg13g2_decap_8 FILLER_66_1060 ();
 sg13g2_decap_8 FILLER_66_1067 ();
 sg13g2_decap_8 FILLER_66_1074 ();
 sg13g2_decap_8 FILLER_66_1081 ();
 sg13g2_decap_8 FILLER_66_1088 ();
 sg13g2_fill_1 FILLER_66_1095 ();
 sg13g2_decap_8 FILLER_66_1106 ();
 sg13g2_decap_8 FILLER_66_1113 ();
 sg13g2_decap_8 FILLER_66_1120 ();
 sg13g2_decap_8 FILLER_66_1127 ();
 sg13g2_decap_8 FILLER_66_1134 ();
 sg13g2_decap_4 FILLER_66_1141 ();
 sg13g2_fill_2 FILLER_66_1145 ();
 sg13g2_decap_8 FILLER_66_1153 ();
 sg13g2_decap_8 FILLER_66_1160 ();
 sg13g2_decap_8 FILLER_66_1167 ();
 sg13g2_decap_8 FILLER_66_1174 ();
 sg13g2_fill_2 FILLER_66_1181 ();
 sg13g2_fill_1 FILLER_66_1183 ();
 sg13g2_decap_8 FILLER_66_1189 ();
 sg13g2_decap_8 FILLER_66_1196 ();
 sg13g2_decap_8 FILLER_66_1203 ();
 sg13g2_fill_2 FILLER_66_1210 ();
 sg13g2_fill_1 FILLER_66_1212 ();
 sg13g2_decap_8 FILLER_66_1219 ();
 sg13g2_decap_8 FILLER_66_1226 ();
 sg13g2_decap_8 FILLER_66_1233 ();
 sg13g2_decap_8 FILLER_66_1240 ();
 sg13g2_decap_8 FILLER_66_1247 ();
 sg13g2_decap_8 FILLER_66_1254 ();
 sg13g2_decap_8 FILLER_66_1261 ();
 sg13g2_fill_1 FILLER_66_1268 ();
 sg13g2_decap_8 FILLER_66_1276 ();
 sg13g2_decap_4 FILLER_66_1292 ();
 sg13g2_fill_1 FILLER_66_1296 ();
 sg13g2_fill_2 FILLER_66_1301 ();
 sg13g2_fill_1 FILLER_66_1303 ();
 sg13g2_decap_8 FILLER_66_1308 ();
 sg13g2_decap_4 FILLER_66_1315 ();
 sg13g2_fill_1 FILLER_66_1319 ();
 sg13g2_decap_8 FILLER_66_1323 ();
 sg13g2_decap_8 FILLER_66_1330 ();
 sg13g2_fill_2 FILLER_66_1337 ();
 sg13g2_fill_2 FILLER_66_1351 ();
 sg13g2_fill_1 FILLER_66_1353 ();
 sg13g2_decap_8 FILLER_66_1358 ();
 sg13g2_decap_8 FILLER_66_1365 ();
 sg13g2_decap_8 FILLER_66_1372 ();
 sg13g2_decap_8 FILLER_66_1379 ();
 sg13g2_decap_8 FILLER_66_1386 ();
 sg13g2_decap_8 FILLER_66_1393 ();
 sg13g2_decap_8 FILLER_66_1400 ();
 sg13g2_fill_2 FILLER_66_1407 ();
 sg13g2_fill_1 FILLER_66_1409 ();
 sg13g2_decap_8 FILLER_66_1416 ();
 sg13g2_decap_8 FILLER_66_1423 ();
 sg13g2_decap_8 FILLER_66_1430 ();
 sg13g2_decap_8 FILLER_66_1437 ();
 sg13g2_fill_2 FILLER_66_1444 ();
 sg13g2_decap_8 FILLER_66_1477 ();
 sg13g2_decap_8 FILLER_66_1484 ();
 sg13g2_decap_4 FILLER_66_1491 ();
 sg13g2_decap_8 FILLER_66_1503 ();
 sg13g2_decap_8 FILLER_66_1510 ();
 sg13g2_decap_8 FILLER_66_1517 ();
 sg13g2_decap_8 FILLER_66_1524 ();
 sg13g2_decap_8 FILLER_66_1531 ();
 sg13g2_decap_4 FILLER_66_1538 ();
 sg13g2_decap_8 FILLER_66_1545 ();
 sg13g2_decap_8 FILLER_66_1552 ();
 sg13g2_decap_8 FILLER_66_1559 ();
 sg13g2_decap_8 FILLER_66_1566 ();
 sg13g2_decap_8 FILLER_66_1573 ();
 sg13g2_decap_8 FILLER_66_1580 ();
 sg13g2_decap_4 FILLER_66_1587 ();
 sg13g2_decap_8 FILLER_66_1596 ();
 sg13g2_decap_4 FILLER_66_1603 ();
 sg13g2_fill_2 FILLER_66_1607 ();
 sg13g2_decap_8 FILLER_66_1613 ();
 sg13g2_fill_2 FILLER_66_1620 ();
 sg13g2_decap_8 FILLER_66_1625 ();
 sg13g2_decap_8 FILLER_66_1632 ();
 sg13g2_decap_8 FILLER_66_1639 ();
 sg13g2_decap_8 FILLER_66_1646 ();
 sg13g2_decap_8 FILLER_66_1653 ();
 sg13g2_fill_2 FILLER_66_1660 ();
 sg13g2_decap_8 FILLER_66_1665 ();
 sg13g2_decap_8 FILLER_66_1672 ();
 sg13g2_decap_8 FILLER_66_1679 ();
 sg13g2_decap_8 FILLER_66_1686 ();
 sg13g2_decap_8 FILLER_66_1693 ();
 sg13g2_decap_8 FILLER_66_1700 ();
 sg13g2_decap_8 FILLER_66_1707 ();
 sg13g2_decap_8 FILLER_66_1714 ();
 sg13g2_decap_8 FILLER_66_1721 ();
 sg13g2_decap_8 FILLER_66_1728 ();
 sg13g2_decap_8 FILLER_66_1735 ();
 sg13g2_decap_8 FILLER_66_1742 ();
 sg13g2_decap_8 FILLER_66_1749 ();
 sg13g2_decap_8 FILLER_66_1772 ();
 sg13g2_decap_8 FILLER_66_1779 ();
 sg13g2_decap_8 FILLER_66_1786 ();
 sg13g2_decap_8 FILLER_66_1793 ();
 sg13g2_decap_8 FILLER_66_1800 ();
 sg13g2_decap_8 FILLER_66_1807 ();
 sg13g2_decap_8 FILLER_66_1814 ();
 sg13g2_decap_8 FILLER_66_1821 ();
 sg13g2_decap_8 FILLER_66_1828 ();
 sg13g2_decap_8 FILLER_66_1835 ();
 sg13g2_decap_8 FILLER_66_1842 ();
 sg13g2_decap_8 FILLER_66_1849 ();
 sg13g2_decap_8 FILLER_66_1856 ();
 sg13g2_decap_8 FILLER_66_1863 ();
 sg13g2_decap_8 FILLER_66_1870 ();
 sg13g2_decap_8 FILLER_66_1877 ();
 sg13g2_decap_8 FILLER_66_1884 ();
 sg13g2_decap_8 FILLER_66_1891 ();
 sg13g2_decap_8 FILLER_66_1898 ();
 sg13g2_decap_8 FILLER_66_1905 ();
 sg13g2_decap_8 FILLER_66_1912 ();
 sg13g2_decap_8 FILLER_66_1919 ();
 sg13g2_decap_8 FILLER_66_1926 ();
 sg13g2_decap_8 FILLER_66_1933 ();
 sg13g2_decap_8 FILLER_66_1940 ();
 sg13g2_decap_8 FILLER_66_1947 ();
 sg13g2_decap_8 FILLER_66_1954 ();
 sg13g2_decap_8 FILLER_66_1961 ();
 sg13g2_decap_8 FILLER_66_1968 ();
 sg13g2_decap_8 FILLER_66_1975 ();
 sg13g2_decap_8 FILLER_66_1982 ();
 sg13g2_decap_8 FILLER_66_1989 ();
 sg13g2_fill_2 FILLER_66_1996 ();
 sg13g2_fill_1 FILLER_66_1998 ();
 sg13g2_decap_8 FILLER_66_2007 ();
 sg13g2_decap_4 FILLER_66_2014 ();
 sg13g2_fill_1 FILLER_66_2018 ();
 sg13g2_decap_8 FILLER_66_2030 ();
 sg13g2_decap_8 FILLER_66_2037 ();
 sg13g2_decap_8 FILLER_66_2044 ();
 sg13g2_decap_8 FILLER_66_2051 ();
 sg13g2_fill_2 FILLER_66_2058 ();
 sg13g2_decap_8 FILLER_66_2064 ();
 sg13g2_decap_8 FILLER_66_2071 ();
 sg13g2_decap_8 FILLER_66_2078 ();
 sg13g2_decap_4 FILLER_66_2085 ();
 sg13g2_fill_1 FILLER_66_2089 ();
 sg13g2_decap_8 FILLER_66_2099 ();
 sg13g2_decap_8 FILLER_66_2106 ();
 sg13g2_decap_8 FILLER_66_2113 ();
 sg13g2_decap_8 FILLER_66_2120 ();
 sg13g2_decap_8 FILLER_66_2127 ();
 sg13g2_decap_8 FILLER_66_2134 ();
 sg13g2_decap_4 FILLER_66_2141 ();
 sg13g2_fill_1 FILLER_66_2145 ();
 sg13g2_decap_8 FILLER_66_2149 ();
 sg13g2_decap_8 FILLER_66_2156 ();
 sg13g2_decap_8 FILLER_66_2163 ();
 sg13g2_decap_8 FILLER_66_2170 ();
 sg13g2_decap_8 FILLER_66_2177 ();
 sg13g2_fill_1 FILLER_66_2184 ();
 sg13g2_decap_8 FILLER_66_2192 ();
 sg13g2_fill_1 FILLER_66_2199 ();
 sg13g2_decap_8 FILLER_66_2204 ();
 sg13g2_decap_8 FILLER_66_2211 ();
 sg13g2_decap_8 FILLER_66_2218 ();
 sg13g2_fill_2 FILLER_66_2225 ();
 sg13g2_decap_8 FILLER_66_2257 ();
 sg13g2_decap_8 FILLER_66_2264 ();
 sg13g2_decap_8 FILLER_66_2271 ();
 sg13g2_decap_8 FILLER_66_2278 ();
 sg13g2_decap_8 FILLER_66_2285 ();
 sg13g2_decap_8 FILLER_66_2292 ();
 sg13g2_decap_8 FILLER_66_2299 ();
 sg13g2_decap_8 FILLER_66_2306 ();
 sg13g2_decap_8 FILLER_66_2313 ();
 sg13g2_decap_8 FILLER_66_2320 ();
 sg13g2_decap_8 FILLER_66_2327 ();
 sg13g2_decap_8 FILLER_66_2334 ();
 sg13g2_decap_8 FILLER_66_2341 ();
 sg13g2_decap_8 FILLER_66_2348 ();
 sg13g2_decap_8 FILLER_66_2355 ();
 sg13g2_decap_8 FILLER_66_2362 ();
 sg13g2_decap_8 FILLER_66_2369 ();
 sg13g2_decap_8 FILLER_66_2376 ();
 sg13g2_decap_8 FILLER_66_2383 ();
 sg13g2_decap_8 FILLER_66_2390 ();
 sg13g2_decap_8 FILLER_66_2397 ();
 sg13g2_decap_8 FILLER_66_2404 ();
 sg13g2_decap_8 FILLER_66_2411 ();
 sg13g2_decap_8 FILLER_66_2418 ();
 sg13g2_decap_8 FILLER_66_2425 ();
 sg13g2_decap_8 FILLER_66_2432 ();
 sg13g2_decap_8 FILLER_66_2439 ();
 sg13g2_decap_8 FILLER_66_2446 ();
 sg13g2_decap_8 FILLER_66_2453 ();
 sg13g2_decap_8 FILLER_66_2460 ();
 sg13g2_decap_8 FILLER_66_2467 ();
 sg13g2_decap_8 FILLER_66_2474 ();
 sg13g2_decap_8 FILLER_66_2481 ();
 sg13g2_decap_8 FILLER_66_2488 ();
 sg13g2_decap_8 FILLER_66_2495 ();
 sg13g2_decap_8 FILLER_66_2502 ();
 sg13g2_decap_8 FILLER_66_2509 ();
 sg13g2_decap_8 FILLER_66_2516 ();
 sg13g2_decap_8 FILLER_66_2523 ();
 sg13g2_decap_8 FILLER_66_2530 ();
 sg13g2_decap_8 FILLER_66_2537 ();
 sg13g2_decap_8 FILLER_66_2544 ();
 sg13g2_decap_8 FILLER_66_2551 ();
 sg13g2_decap_8 FILLER_66_2558 ();
 sg13g2_decap_8 FILLER_66_2565 ();
 sg13g2_decap_8 FILLER_66_2572 ();
 sg13g2_decap_8 FILLER_66_2579 ();
 sg13g2_decap_8 FILLER_66_2586 ();
 sg13g2_decap_8 FILLER_66_2593 ();
 sg13g2_decap_8 FILLER_66_2600 ();
 sg13g2_decap_8 FILLER_66_2607 ();
 sg13g2_decap_8 FILLER_66_2614 ();
 sg13g2_decap_8 FILLER_66_2621 ();
 sg13g2_decap_8 FILLER_66_2628 ();
 sg13g2_decap_8 FILLER_66_2635 ();
 sg13g2_decap_8 FILLER_66_2642 ();
 sg13g2_decap_8 FILLER_66_2649 ();
 sg13g2_decap_8 FILLER_66_2656 ();
 sg13g2_decap_8 FILLER_66_2663 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_4 FILLER_67_70 ();
 sg13g2_fill_1 FILLER_67_74 ();
 sg13g2_decap_8 FILLER_67_79 ();
 sg13g2_decap_8 FILLER_67_86 ();
 sg13g2_decap_8 FILLER_67_93 ();
 sg13g2_decap_8 FILLER_67_100 ();
 sg13g2_decap_4 FILLER_67_107 ();
 sg13g2_decap_8 FILLER_67_119 ();
 sg13g2_decap_8 FILLER_67_126 ();
 sg13g2_decap_8 FILLER_67_133 ();
 sg13g2_decap_8 FILLER_67_140 ();
 sg13g2_decap_8 FILLER_67_147 ();
 sg13g2_decap_8 FILLER_67_154 ();
 sg13g2_decap_8 FILLER_67_161 ();
 sg13g2_decap_8 FILLER_67_168 ();
 sg13g2_decap_8 FILLER_67_175 ();
 sg13g2_decap_8 FILLER_67_182 ();
 sg13g2_decap_8 FILLER_67_189 ();
 sg13g2_decap_8 FILLER_67_196 ();
 sg13g2_decap_8 FILLER_67_203 ();
 sg13g2_decap_8 FILLER_67_210 ();
 sg13g2_decap_8 FILLER_67_217 ();
 sg13g2_decap_8 FILLER_67_224 ();
 sg13g2_decap_8 FILLER_67_231 ();
 sg13g2_decap_8 FILLER_67_238 ();
 sg13g2_decap_8 FILLER_67_245 ();
 sg13g2_decap_8 FILLER_67_252 ();
 sg13g2_decap_4 FILLER_67_259 ();
 sg13g2_decap_8 FILLER_67_289 ();
 sg13g2_decap_8 FILLER_67_296 ();
 sg13g2_decap_8 FILLER_67_303 ();
 sg13g2_decap_8 FILLER_67_310 ();
 sg13g2_decap_8 FILLER_67_317 ();
 sg13g2_decap_8 FILLER_67_324 ();
 sg13g2_decap_8 FILLER_67_331 ();
 sg13g2_decap_8 FILLER_67_338 ();
 sg13g2_decap_8 FILLER_67_345 ();
 sg13g2_decap_8 FILLER_67_352 ();
 sg13g2_decap_8 FILLER_67_359 ();
 sg13g2_decap_8 FILLER_67_366 ();
 sg13g2_decap_8 FILLER_67_373 ();
 sg13g2_decap_8 FILLER_67_380 ();
 sg13g2_decap_4 FILLER_67_387 ();
 sg13g2_fill_2 FILLER_67_391 ();
 sg13g2_decap_8 FILLER_67_402 ();
 sg13g2_decap_8 FILLER_67_409 ();
 sg13g2_decap_8 FILLER_67_416 ();
 sg13g2_decap_8 FILLER_67_423 ();
 sg13g2_decap_8 FILLER_67_430 ();
 sg13g2_fill_2 FILLER_67_437 ();
 sg13g2_fill_1 FILLER_67_439 ();
 sg13g2_decap_8 FILLER_67_445 ();
 sg13g2_decap_8 FILLER_67_452 ();
 sg13g2_decap_8 FILLER_67_459 ();
 sg13g2_decap_8 FILLER_67_466 ();
 sg13g2_fill_2 FILLER_67_473 ();
 sg13g2_fill_1 FILLER_67_475 ();
 sg13g2_fill_2 FILLER_67_480 ();
 sg13g2_fill_1 FILLER_67_482 ();
 sg13g2_decap_8 FILLER_67_488 ();
 sg13g2_decap_8 FILLER_67_495 ();
 sg13g2_decap_8 FILLER_67_502 ();
 sg13g2_fill_2 FILLER_67_509 ();
 sg13g2_fill_1 FILLER_67_511 ();
 sg13g2_decap_8 FILLER_67_520 ();
 sg13g2_decap_8 FILLER_67_527 ();
 sg13g2_decap_8 FILLER_67_534 ();
 sg13g2_decap_4 FILLER_67_549 ();
 sg13g2_fill_1 FILLER_67_553 ();
 sg13g2_decap_8 FILLER_67_562 ();
 sg13g2_decap_8 FILLER_67_569 ();
 sg13g2_decap_8 FILLER_67_576 ();
 sg13g2_decap_8 FILLER_67_583 ();
 sg13g2_decap_8 FILLER_67_590 ();
 sg13g2_decap_8 FILLER_67_597 ();
 sg13g2_decap_8 FILLER_67_604 ();
 sg13g2_decap_8 FILLER_67_611 ();
 sg13g2_fill_1 FILLER_67_618 ();
 sg13g2_decap_8 FILLER_67_624 ();
 sg13g2_decap_8 FILLER_67_631 ();
 sg13g2_decap_8 FILLER_67_638 ();
 sg13g2_fill_2 FILLER_67_645 ();
 sg13g2_decap_8 FILLER_67_688 ();
 sg13g2_decap_8 FILLER_67_695 ();
 sg13g2_decap_8 FILLER_67_702 ();
 sg13g2_decap_8 FILLER_67_709 ();
 sg13g2_decap_8 FILLER_67_716 ();
 sg13g2_decap_8 FILLER_67_723 ();
 sg13g2_fill_1 FILLER_67_730 ();
 sg13g2_decap_8 FILLER_67_739 ();
 sg13g2_decap_8 FILLER_67_746 ();
 sg13g2_decap_8 FILLER_67_753 ();
 sg13g2_decap_4 FILLER_67_760 ();
 sg13g2_fill_2 FILLER_67_764 ();
 sg13g2_decap_8 FILLER_67_778 ();
 sg13g2_decap_8 FILLER_67_785 ();
 sg13g2_fill_2 FILLER_67_792 ();
 sg13g2_decap_8 FILLER_67_799 ();
 sg13g2_decap_4 FILLER_67_806 ();
 sg13g2_fill_1 FILLER_67_810 ();
 sg13g2_decap_8 FILLER_67_815 ();
 sg13g2_decap_8 FILLER_67_822 ();
 sg13g2_decap_8 FILLER_67_829 ();
 sg13g2_decap_8 FILLER_67_836 ();
 sg13g2_decap_8 FILLER_67_843 ();
 sg13g2_fill_1 FILLER_67_869 ();
 sg13g2_decap_8 FILLER_67_876 ();
 sg13g2_decap_8 FILLER_67_883 ();
 sg13g2_decap_8 FILLER_67_890 ();
 sg13g2_decap_8 FILLER_67_897 ();
 sg13g2_decap_8 FILLER_67_904 ();
 sg13g2_decap_4 FILLER_67_911 ();
 sg13g2_decap_8 FILLER_67_918 ();
 sg13g2_decap_4 FILLER_67_925 ();
 sg13g2_decap_8 FILLER_67_936 ();
 sg13g2_decap_8 FILLER_67_943 ();
 sg13g2_decap_8 FILLER_67_950 ();
 sg13g2_fill_1 FILLER_67_957 ();
 sg13g2_fill_2 FILLER_67_966 ();
 sg13g2_fill_1 FILLER_67_968 ();
 sg13g2_decap_8 FILLER_67_985 ();
 sg13g2_fill_2 FILLER_67_992 ();
 sg13g2_fill_1 FILLER_67_1009 ();
 sg13g2_decap_8 FILLER_67_1015 ();
 sg13g2_decap_8 FILLER_67_1022 ();
 sg13g2_fill_2 FILLER_67_1029 ();
 sg13g2_fill_1 FILLER_67_1031 ();
 sg13g2_decap_8 FILLER_67_1056 ();
 sg13g2_decap_8 FILLER_67_1063 ();
 sg13g2_decap_8 FILLER_67_1070 ();
 sg13g2_decap_4 FILLER_67_1077 ();
 sg13g2_fill_2 FILLER_67_1081 ();
 sg13g2_decap_8 FILLER_67_1088 ();
 sg13g2_decap_8 FILLER_67_1095 ();
 sg13g2_fill_1 FILLER_67_1102 ();
 sg13g2_decap_8 FILLER_67_1107 ();
 sg13g2_decap_8 FILLER_67_1114 ();
 sg13g2_decap_8 FILLER_67_1121 ();
 sg13g2_decap_8 FILLER_67_1128 ();
 sg13g2_decap_8 FILLER_67_1135 ();
 sg13g2_decap_8 FILLER_67_1142 ();
 sg13g2_decap_8 FILLER_67_1149 ();
 sg13g2_fill_1 FILLER_67_1156 ();
 sg13g2_decap_8 FILLER_67_1160 ();
 sg13g2_decap_8 FILLER_67_1167 ();
 sg13g2_decap_8 FILLER_67_1174 ();
 sg13g2_decap_8 FILLER_67_1181 ();
 sg13g2_decap_8 FILLER_67_1188 ();
 sg13g2_decap_8 FILLER_67_1195 ();
 sg13g2_decap_8 FILLER_67_1202 ();
 sg13g2_fill_1 FILLER_67_1209 ();
 sg13g2_decap_8 FILLER_67_1215 ();
 sg13g2_decap_8 FILLER_67_1222 ();
 sg13g2_decap_8 FILLER_67_1229 ();
 sg13g2_decap_8 FILLER_67_1236 ();
 sg13g2_decap_8 FILLER_67_1243 ();
 sg13g2_decap_8 FILLER_67_1250 ();
 sg13g2_decap_8 FILLER_67_1257 ();
 sg13g2_decap_4 FILLER_67_1264 ();
 sg13g2_fill_1 FILLER_67_1268 ();
 sg13g2_decap_8 FILLER_67_1281 ();
 sg13g2_decap_8 FILLER_67_1288 ();
 sg13g2_decap_8 FILLER_67_1295 ();
 sg13g2_decap_8 FILLER_67_1302 ();
 sg13g2_decap_8 FILLER_67_1309 ();
 sg13g2_decap_8 FILLER_67_1316 ();
 sg13g2_decap_8 FILLER_67_1323 ();
 sg13g2_decap_8 FILLER_67_1330 ();
 sg13g2_fill_2 FILLER_67_1337 ();
 sg13g2_decap_8 FILLER_67_1349 ();
 sg13g2_decap_4 FILLER_67_1356 ();
 sg13g2_fill_1 FILLER_67_1360 ();
 sg13g2_decap_8 FILLER_67_1366 ();
 sg13g2_decap_8 FILLER_67_1373 ();
 sg13g2_decap_8 FILLER_67_1380 ();
 sg13g2_decap_8 FILLER_67_1387 ();
 sg13g2_decap_8 FILLER_67_1394 ();
 sg13g2_decap_8 FILLER_67_1401 ();
 sg13g2_decap_8 FILLER_67_1413 ();
 sg13g2_decap_8 FILLER_67_1420 ();
 sg13g2_decap_8 FILLER_67_1427 ();
 sg13g2_decap_8 FILLER_67_1434 ();
 sg13g2_decap_8 FILLER_67_1441 ();
 sg13g2_decap_4 FILLER_67_1448 ();
 sg13g2_decap_8 FILLER_67_1462 ();
 sg13g2_decap_8 FILLER_67_1469 ();
 sg13g2_fill_2 FILLER_67_1476 ();
 sg13g2_fill_1 FILLER_67_1478 ();
 sg13g2_decap_8 FILLER_67_1482 ();
 sg13g2_decap_8 FILLER_67_1489 ();
 sg13g2_decap_4 FILLER_67_1496 ();
 sg13g2_decap_8 FILLER_67_1503 ();
 sg13g2_decap_8 FILLER_67_1510 ();
 sg13g2_decap_8 FILLER_67_1517 ();
 sg13g2_decap_8 FILLER_67_1524 ();
 sg13g2_decap_8 FILLER_67_1531 ();
 sg13g2_fill_2 FILLER_67_1538 ();
 sg13g2_fill_1 FILLER_67_1540 ();
 sg13g2_decap_8 FILLER_67_1548 ();
 sg13g2_decap_8 FILLER_67_1555 ();
 sg13g2_decap_4 FILLER_67_1562 ();
 sg13g2_fill_1 FILLER_67_1566 ();
 sg13g2_decap_8 FILLER_67_1570 ();
 sg13g2_decap_8 FILLER_67_1577 ();
 sg13g2_decap_4 FILLER_67_1584 ();
 sg13g2_fill_2 FILLER_67_1588 ();
 sg13g2_decap_8 FILLER_67_1594 ();
 sg13g2_decap_4 FILLER_67_1601 ();
 sg13g2_fill_2 FILLER_67_1605 ();
 sg13g2_fill_2 FILLER_67_1611 ();
 sg13g2_decap_8 FILLER_67_1635 ();
 sg13g2_fill_2 FILLER_67_1642 ();
 sg13g2_fill_2 FILLER_67_1668 ();
 sg13g2_decap_8 FILLER_67_1677 ();
 sg13g2_decap_8 FILLER_67_1684 ();
 sg13g2_decap_8 FILLER_67_1691 ();
 sg13g2_decap_8 FILLER_67_1713 ();
 sg13g2_decap_8 FILLER_67_1720 ();
 sg13g2_decap_8 FILLER_67_1727 ();
 sg13g2_decap_8 FILLER_67_1734 ();
 sg13g2_decap_8 FILLER_67_1741 ();
 sg13g2_decap_8 FILLER_67_1748 ();
 sg13g2_decap_8 FILLER_67_1755 ();
 sg13g2_decap_8 FILLER_67_1762 ();
 sg13g2_decap_8 FILLER_67_1769 ();
 sg13g2_decap_4 FILLER_67_1776 ();
 sg13g2_decap_8 FILLER_67_1784 ();
 sg13g2_decap_8 FILLER_67_1791 ();
 sg13g2_fill_2 FILLER_67_1798 ();
 sg13g2_fill_1 FILLER_67_1800 ();
 sg13g2_decap_8 FILLER_67_1805 ();
 sg13g2_decap_8 FILLER_67_1812 ();
 sg13g2_decap_8 FILLER_67_1819 ();
 sg13g2_decap_8 FILLER_67_1826 ();
 sg13g2_decap_8 FILLER_67_1833 ();
 sg13g2_decap_8 FILLER_67_1840 ();
 sg13g2_decap_8 FILLER_67_1847 ();
 sg13g2_decap_8 FILLER_67_1854 ();
 sg13g2_decap_8 FILLER_67_1861 ();
 sg13g2_decap_8 FILLER_67_1868 ();
 sg13g2_decap_8 FILLER_67_1875 ();
 sg13g2_decap_8 FILLER_67_1882 ();
 sg13g2_decap_8 FILLER_67_1889 ();
 sg13g2_decap_8 FILLER_67_1896 ();
 sg13g2_decap_8 FILLER_67_1903 ();
 sg13g2_decap_8 FILLER_67_1910 ();
 sg13g2_decap_8 FILLER_67_1917 ();
 sg13g2_decap_8 FILLER_67_1924 ();
 sg13g2_decap_8 FILLER_67_1931 ();
 sg13g2_decap_8 FILLER_67_1938 ();
 sg13g2_decap_8 FILLER_67_1945 ();
 sg13g2_decap_8 FILLER_67_1952 ();
 sg13g2_decap_8 FILLER_67_1959 ();
 sg13g2_fill_1 FILLER_67_1966 ();
 sg13g2_decap_8 FILLER_67_1974 ();
 sg13g2_decap_8 FILLER_67_1981 ();
 sg13g2_decap_8 FILLER_67_1988 ();
 sg13g2_decap_8 FILLER_67_1995 ();
 sg13g2_decap_8 FILLER_67_2002 ();
 sg13g2_decap_8 FILLER_67_2009 ();
 sg13g2_decap_4 FILLER_67_2016 ();
 sg13g2_fill_1 FILLER_67_2020 ();
 sg13g2_decap_8 FILLER_67_2026 ();
 sg13g2_decap_8 FILLER_67_2033 ();
 sg13g2_decap_8 FILLER_67_2040 ();
 sg13g2_decap_8 FILLER_67_2047 ();
 sg13g2_decap_8 FILLER_67_2054 ();
 sg13g2_decap_8 FILLER_67_2061 ();
 sg13g2_decap_8 FILLER_67_2068 ();
 sg13g2_decap_8 FILLER_67_2075 ();
 sg13g2_decap_8 FILLER_67_2082 ();
 sg13g2_decap_8 FILLER_67_2089 ();
 sg13g2_fill_2 FILLER_67_2096 ();
 sg13g2_fill_1 FILLER_67_2098 ();
 sg13g2_decap_8 FILLER_67_2103 ();
 sg13g2_decap_8 FILLER_67_2110 ();
 sg13g2_decap_8 FILLER_67_2117 ();
 sg13g2_decap_8 FILLER_67_2124 ();
 sg13g2_decap_8 FILLER_67_2131 ();
 sg13g2_decap_4 FILLER_67_2138 ();
 sg13g2_fill_2 FILLER_67_2142 ();
 sg13g2_decap_8 FILLER_67_2148 ();
 sg13g2_decap_8 FILLER_67_2158 ();
 sg13g2_decap_8 FILLER_67_2165 ();
 sg13g2_decap_8 FILLER_67_2172 ();
 sg13g2_decap_8 FILLER_67_2179 ();
 sg13g2_decap_8 FILLER_67_2186 ();
 sg13g2_decap_8 FILLER_67_2193 ();
 sg13g2_decap_8 FILLER_67_2200 ();
 sg13g2_decap_8 FILLER_67_2207 ();
 sg13g2_decap_8 FILLER_67_2214 ();
 sg13g2_decap_8 FILLER_67_2221 ();
 sg13g2_decap_8 FILLER_67_2228 ();
 sg13g2_decap_8 FILLER_67_2235 ();
 sg13g2_decap_8 FILLER_67_2242 ();
 sg13g2_decap_8 FILLER_67_2249 ();
 sg13g2_decap_8 FILLER_67_2256 ();
 sg13g2_decap_8 FILLER_67_2263 ();
 sg13g2_decap_8 FILLER_67_2270 ();
 sg13g2_decap_8 FILLER_67_2277 ();
 sg13g2_decap_8 FILLER_67_2284 ();
 sg13g2_decap_8 FILLER_67_2291 ();
 sg13g2_decap_8 FILLER_67_2298 ();
 sg13g2_decap_8 FILLER_67_2305 ();
 sg13g2_decap_8 FILLER_67_2312 ();
 sg13g2_decap_8 FILLER_67_2319 ();
 sg13g2_decap_8 FILLER_67_2326 ();
 sg13g2_decap_8 FILLER_67_2333 ();
 sg13g2_decap_8 FILLER_67_2340 ();
 sg13g2_decap_8 FILLER_67_2347 ();
 sg13g2_decap_8 FILLER_67_2354 ();
 sg13g2_decap_8 FILLER_67_2361 ();
 sg13g2_decap_8 FILLER_67_2368 ();
 sg13g2_decap_8 FILLER_67_2375 ();
 sg13g2_decap_8 FILLER_67_2382 ();
 sg13g2_decap_8 FILLER_67_2389 ();
 sg13g2_decap_8 FILLER_67_2396 ();
 sg13g2_decap_8 FILLER_67_2403 ();
 sg13g2_decap_8 FILLER_67_2410 ();
 sg13g2_decap_8 FILLER_67_2417 ();
 sg13g2_decap_8 FILLER_67_2424 ();
 sg13g2_decap_8 FILLER_67_2431 ();
 sg13g2_decap_8 FILLER_67_2438 ();
 sg13g2_decap_8 FILLER_67_2445 ();
 sg13g2_decap_8 FILLER_67_2452 ();
 sg13g2_decap_8 FILLER_67_2459 ();
 sg13g2_decap_8 FILLER_67_2466 ();
 sg13g2_decap_8 FILLER_67_2473 ();
 sg13g2_decap_8 FILLER_67_2480 ();
 sg13g2_decap_8 FILLER_67_2487 ();
 sg13g2_decap_8 FILLER_67_2494 ();
 sg13g2_decap_8 FILLER_67_2501 ();
 sg13g2_decap_8 FILLER_67_2508 ();
 sg13g2_decap_8 FILLER_67_2515 ();
 sg13g2_decap_8 FILLER_67_2522 ();
 sg13g2_decap_8 FILLER_67_2529 ();
 sg13g2_decap_8 FILLER_67_2536 ();
 sg13g2_decap_8 FILLER_67_2543 ();
 sg13g2_decap_8 FILLER_67_2550 ();
 sg13g2_decap_8 FILLER_67_2557 ();
 sg13g2_decap_8 FILLER_67_2564 ();
 sg13g2_decap_8 FILLER_67_2571 ();
 sg13g2_decap_8 FILLER_67_2578 ();
 sg13g2_decap_8 FILLER_67_2585 ();
 sg13g2_decap_8 FILLER_67_2592 ();
 sg13g2_decap_8 FILLER_67_2599 ();
 sg13g2_decap_8 FILLER_67_2606 ();
 sg13g2_decap_8 FILLER_67_2613 ();
 sg13g2_decap_8 FILLER_67_2620 ();
 sg13g2_decap_8 FILLER_67_2627 ();
 sg13g2_decap_8 FILLER_67_2634 ();
 sg13g2_decap_8 FILLER_67_2641 ();
 sg13g2_decap_8 FILLER_67_2648 ();
 sg13g2_decap_8 FILLER_67_2655 ();
 sg13g2_decap_8 FILLER_67_2662 ();
 sg13g2_fill_1 FILLER_67_2669 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_4 FILLER_68_35 ();
 sg13g2_fill_1 FILLER_68_39 ();
 sg13g2_decap_8 FILLER_68_66 ();
 sg13g2_fill_1 FILLER_68_73 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_4 FILLER_68_105 ();
 sg13g2_fill_2 FILLER_68_109 ();
 sg13g2_decap_4 FILLER_68_114 ();
 sg13g2_fill_1 FILLER_68_118 ();
 sg13g2_decap_8 FILLER_68_124 ();
 sg13g2_decap_8 FILLER_68_131 ();
 sg13g2_decap_4 FILLER_68_138 ();
 sg13g2_fill_1 FILLER_68_142 ();
 sg13g2_decap_8 FILLER_68_154 ();
 sg13g2_decap_8 FILLER_68_161 ();
 sg13g2_decap_8 FILLER_68_168 ();
 sg13g2_decap_8 FILLER_68_175 ();
 sg13g2_decap_8 FILLER_68_182 ();
 sg13g2_decap_8 FILLER_68_189 ();
 sg13g2_decap_8 FILLER_68_196 ();
 sg13g2_decap_8 FILLER_68_203 ();
 sg13g2_decap_8 FILLER_68_210 ();
 sg13g2_decap_8 FILLER_68_217 ();
 sg13g2_decap_8 FILLER_68_224 ();
 sg13g2_decap_8 FILLER_68_231 ();
 sg13g2_decap_8 FILLER_68_238 ();
 sg13g2_decap_8 FILLER_68_245 ();
 sg13g2_decap_8 FILLER_68_257 ();
 sg13g2_fill_2 FILLER_68_264 ();
 sg13g2_fill_1 FILLER_68_266 ();
 sg13g2_decap_8 FILLER_68_271 ();
 sg13g2_decap_8 FILLER_68_278 ();
 sg13g2_decap_8 FILLER_68_285 ();
 sg13g2_decap_8 FILLER_68_292 ();
 sg13g2_decap_8 FILLER_68_299 ();
 sg13g2_decap_8 FILLER_68_306 ();
 sg13g2_decap_8 FILLER_68_313 ();
 sg13g2_decap_8 FILLER_68_320 ();
 sg13g2_decap_8 FILLER_68_327 ();
 sg13g2_decap_8 FILLER_68_334 ();
 sg13g2_decap_8 FILLER_68_341 ();
 sg13g2_decap_8 FILLER_68_348 ();
 sg13g2_decap_4 FILLER_68_355 ();
 sg13g2_fill_2 FILLER_68_359 ();
 sg13g2_decap_8 FILLER_68_365 ();
 sg13g2_decap_8 FILLER_68_372 ();
 sg13g2_decap_8 FILLER_68_379 ();
 sg13g2_decap_8 FILLER_68_386 ();
 sg13g2_decap_8 FILLER_68_393 ();
 sg13g2_decap_8 FILLER_68_400 ();
 sg13g2_decap_8 FILLER_68_407 ();
 sg13g2_decap_8 FILLER_68_414 ();
 sg13g2_decap_8 FILLER_68_421 ();
 sg13g2_decap_4 FILLER_68_428 ();
 sg13g2_decap_8 FILLER_68_436 ();
 sg13g2_decap_8 FILLER_68_443 ();
 sg13g2_decap_8 FILLER_68_450 ();
 sg13g2_decap_8 FILLER_68_460 ();
 sg13g2_decap_8 FILLER_68_467 ();
 sg13g2_decap_8 FILLER_68_474 ();
 sg13g2_decap_8 FILLER_68_481 ();
 sg13g2_decap_8 FILLER_68_488 ();
 sg13g2_decap_8 FILLER_68_495 ();
 sg13g2_decap_8 FILLER_68_502 ();
 sg13g2_decap_4 FILLER_68_509 ();
 sg13g2_fill_1 FILLER_68_513 ();
 sg13g2_decap_8 FILLER_68_518 ();
 sg13g2_decap_8 FILLER_68_525 ();
 sg13g2_decap_8 FILLER_68_532 ();
 sg13g2_decap_8 FILLER_68_539 ();
 sg13g2_decap_8 FILLER_68_546 ();
 sg13g2_decap_4 FILLER_68_553 ();
 sg13g2_fill_1 FILLER_68_557 ();
 sg13g2_decap_8 FILLER_68_561 ();
 sg13g2_decap_8 FILLER_68_568 ();
 sg13g2_decap_8 FILLER_68_575 ();
 sg13g2_decap_8 FILLER_68_582 ();
 sg13g2_decap_8 FILLER_68_593 ();
 sg13g2_decap_8 FILLER_68_600 ();
 sg13g2_decap_8 FILLER_68_607 ();
 sg13g2_decap_8 FILLER_68_614 ();
 sg13g2_decap_8 FILLER_68_621 ();
 sg13g2_decap_8 FILLER_68_628 ();
 sg13g2_decap_8 FILLER_68_635 ();
 sg13g2_decap_8 FILLER_68_642 ();
 sg13g2_decap_4 FILLER_68_649 ();
 sg13g2_decap_8 FILLER_68_657 ();
 sg13g2_fill_2 FILLER_68_672 ();
 sg13g2_decap_8 FILLER_68_690 ();
 sg13g2_decap_8 FILLER_68_697 ();
 sg13g2_fill_2 FILLER_68_704 ();
 sg13g2_decap_8 FILLER_68_712 ();
 sg13g2_decap_4 FILLER_68_719 ();
 sg13g2_fill_1 FILLER_68_723 ();
 sg13g2_decap_4 FILLER_68_729 ();
 sg13g2_fill_1 FILLER_68_733 ();
 sg13g2_decap_8 FILLER_68_738 ();
 sg13g2_decap_8 FILLER_68_745 ();
 sg13g2_decap_4 FILLER_68_752 ();
 sg13g2_fill_1 FILLER_68_756 ();
 sg13g2_decap_8 FILLER_68_773 ();
 sg13g2_decap_8 FILLER_68_780 ();
 sg13g2_decap_8 FILLER_68_787 ();
 sg13g2_decap_8 FILLER_68_794 ();
 sg13g2_decap_8 FILLER_68_801 ();
 sg13g2_decap_8 FILLER_68_808 ();
 sg13g2_decap_8 FILLER_68_815 ();
 sg13g2_decap_8 FILLER_68_822 ();
 sg13g2_fill_2 FILLER_68_829 ();
 sg13g2_fill_1 FILLER_68_831 ();
 sg13g2_fill_1 FILLER_68_859 ();
 sg13g2_decap_8 FILLER_68_883 ();
 sg13g2_decap_8 FILLER_68_896 ();
 sg13g2_decap_8 FILLER_68_903 ();
 sg13g2_fill_2 FILLER_68_910 ();
 sg13g2_decap_8 FILLER_68_925 ();
 sg13g2_decap_8 FILLER_68_932 ();
 sg13g2_decap_8 FILLER_68_939 ();
 sg13g2_decap_8 FILLER_68_946 ();
 sg13g2_decap_8 FILLER_68_953 ();
 sg13g2_decap_8 FILLER_68_960 ();
 sg13g2_decap_8 FILLER_68_967 ();
 sg13g2_decap_8 FILLER_68_974 ();
 sg13g2_decap_8 FILLER_68_981 ();
 sg13g2_decap_8 FILLER_68_988 ();
 sg13g2_decap_4 FILLER_68_995 ();
 sg13g2_fill_1 FILLER_68_999 ();
 sg13g2_decap_8 FILLER_68_1011 ();
 sg13g2_decap_8 FILLER_68_1018 ();
 sg13g2_decap_8 FILLER_68_1025 ();
 sg13g2_decap_4 FILLER_68_1032 ();
 sg13g2_decap_8 FILLER_68_1040 ();
 sg13g2_decap_8 FILLER_68_1047 ();
 sg13g2_decap_8 FILLER_68_1054 ();
 sg13g2_decap_8 FILLER_68_1061 ();
 sg13g2_decap_8 FILLER_68_1068 ();
 sg13g2_decap_8 FILLER_68_1075 ();
 sg13g2_decap_8 FILLER_68_1082 ();
 sg13g2_decap_8 FILLER_68_1089 ();
 sg13g2_decap_8 FILLER_68_1096 ();
 sg13g2_decap_8 FILLER_68_1103 ();
 sg13g2_decap_8 FILLER_68_1110 ();
 sg13g2_decap_8 FILLER_68_1117 ();
 sg13g2_decap_8 FILLER_68_1124 ();
 sg13g2_decap_8 FILLER_68_1131 ();
 sg13g2_fill_2 FILLER_68_1138 ();
 sg13g2_fill_2 FILLER_68_1155 ();
 sg13g2_decap_8 FILLER_68_1169 ();
 sg13g2_decap_8 FILLER_68_1176 ();
 sg13g2_decap_8 FILLER_68_1183 ();
 sg13g2_decap_8 FILLER_68_1190 ();
 sg13g2_decap_8 FILLER_68_1197 ();
 sg13g2_decap_8 FILLER_68_1204 ();
 sg13g2_decap_4 FILLER_68_1211 ();
 sg13g2_fill_2 FILLER_68_1215 ();
 sg13g2_decap_8 FILLER_68_1222 ();
 sg13g2_decap_8 FILLER_68_1229 ();
 sg13g2_decap_8 FILLER_68_1236 ();
 sg13g2_decap_8 FILLER_68_1243 ();
 sg13g2_decap_8 FILLER_68_1250 ();
 sg13g2_decap_8 FILLER_68_1257 ();
 sg13g2_decap_8 FILLER_68_1264 ();
 sg13g2_decap_8 FILLER_68_1271 ();
 sg13g2_fill_2 FILLER_68_1278 ();
 sg13g2_decap_8 FILLER_68_1285 ();
 sg13g2_decap_8 FILLER_68_1292 ();
 sg13g2_decap_8 FILLER_68_1299 ();
 sg13g2_decap_4 FILLER_68_1306 ();
 sg13g2_fill_2 FILLER_68_1310 ();
 sg13g2_decap_8 FILLER_68_1327 ();
 sg13g2_decap_8 FILLER_68_1334 ();
 sg13g2_decap_8 FILLER_68_1341 ();
 sg13g2_decap_8 FILLER_68_1363 ();
 sg13g2_decap_8 FILLER_68_1370 ();
 sg13g2_decap_4 FILLER_68_1377 ();
 sg13g2_decap_8 FILLER_68_1385 ();
 sg13g2_decap_4 FILLER_68_1392 ();
 sg13g2_fill_1 FILLER_68_1396 ();
 sg13g2_decap_8 FILLER_68_1401 ();
 sg13g2_decap_8 FILLER_68_1408 ();
 sg13g2_decap_8 FILLER_68_1415 ();
 sg13g2_decap_8 FILLER_68_1422 ();
 sg13g2_decap_8 FILLER_68_1429 ();
 sg13g2_decap_8 FILLER_68_1436 ();
 sg13g2_fill_1 FILLER_68_1443 ();
 sg13g2_decap_8 FILLER_68_1449 ();
 sg13g2_decap_8 FILLER_68_1456 ();
 sg13g2_fill_2 FILLER_68_1463 ();
 sg13g2_decap_8 FILLER_68_1470 ();
 sg13g2_fill_2 FILLER_68_1477 ();
 sg13g2_decap_8 FILLER_68_1483 ();
 sg13g2_fill_2 FILLER_68_1490 ();
 sg13g2_fill_2 FILLER_68_1498 ();
 sg13g2_fill_1 FILLER_68_1506 ();
 sg13g2_decap_4 FILLER_68_1536 ();
 sg13g2_fill_1 FILLER_68_1540 ();
 sg13g2_decap_8 FILLER_68_1546 ();
 sg13g2_decap_8 FILLER_68_1553 ();
 sg13g2_decap_8 FILLER_68_1560 ();
 sg13g2_decap_8 FILLER_68_1571 ();
 sg13g2_decap_8 FILLER_68_1578 ();
 sg13g2_decap_8 FILLER_68_1585 ();
 sg13g2_decap_8 FILLER_68_1592 ();
 sg13g2_decap_8 FILLER_68_1599 ();
 sg13g2_decap_4 FILLER_68_1606 ();
 sg13g2_decap_8 FILLER_68_1614 ();
 sg13g2_fill_1 FILLER_68_1621 ();
 sg13g2_decap_8 FILLER_68_1626 ();
 sg13g2_decap_4 FILLER_68_1633 ();
 sg13g2_fill_1 FILLER_68_1637 ();
 sg13g2_fill_2 FILLER_68_1651 ();
 sg13g2_decap_8 FILLER_68_1657 ();
 sg13g2_decap_4 FILLER_68_1664 ();
 sg13g2_fill_2 FILLER_68_1668 ();
 sg13g2_decap_8 FILLER_68_1674 ();
 sg13g2_decap_8 FILLER_68_1681 ();
 sg13g2_decap_8 FILLER_68_1688 ();
 sg13g2_fill_2 FILLER_68_1695 ();
 sg13g2_fill_1 FILLER_68_1697 ();
 sg13g2_decap_8 FILLER_68_1718 ();
 sg13g2_fill_1 FILLER_68_1725 ();
 sg13g2_decap_8 FILLER_68_1747 ();
 sg13g2_decap_8 FILLER_68_1754 ();
 sg13g2_decap_8 FILLER_68_1761 ();
 sg13g2_decap_8 FILLER_68_1768 ();
 sg13g2_decap_8 FILLER_68_1775 ();
 sg13g2_decap_8 FILLER_68_1782 ();
 sg13g2_decap_8 FILLER_68_1789 ();
 sg13g2_decap_8 FILLER_68_1796 ();
 sg13g2_decap_8 FILLER_68_1803 ();
 sg13g2_decap_8 FILLER_68_1810 ();
 sg13g2_decap_8 FILLER_68_1817 ();
 sg13g2_decap_8 FILLER_68_1824 ();
 sg13g2_decap_8 FILLER_68_1831 ();
 sg13g2_decap_8 FILLER_68_1838 ();
 sg13g2_decap_8 FILLER_68_1845 ();
 sg13g2_decap_8 FILLER_68_1852 ();
 sg13g2_decap_8 FILLER_68_1859 ();
 sg13g2_decap_8 FILLER_68_1866 ();
 sg13g2_decap_8 FILLER_68_1873 ();
 sg13g2_decap_8 FILLER_68_1880 ();
 sg13g2_decap_8 FILLER_68_1887 ();
 sg13g2_decap_8 FILLER_68_1894 ();
 sg13g2_decap_8 FILLER_68_1901 ();
 sg13g2_decap_8 FILLER_68_1908 ();
 sg13g2_decap_8 FILLER_68_1915 ();
 sg13g2_decap_8 FILLER_68_1922 ();
 sg13g2_decap_8 FILLER_68_1929 ();
 sg13g2_decap_8 FILLER_68_1936 ();
 sg13g2_decap_8 FILLER_68_1943 ();
 sg13g2_decap_8 FILLER_68_1950 ();
 sg13g2_decap_8 FILLER_68_1957 ();
 sg13g2_fill_2 FILLER_68_1964 ();
 sg13g2_fill_1 FILLER_68_1966 ();
 sg13g2_decap_8 FILLER_68_2001 ();
 sg13g2_fill_1 FILLER_68_2008 ();
 sg13g2_decap_8 FILLER_68_2012 ();
 sg13g2_decap_8 FILLER_68_2019 ();
 sg13g2_decap_8 FILLER_68_2026 ();
 sg13g2_decap_8 FILLER_68_2033 ();
 sg13g2_decap_8 FILLER_68_2040 ();
 sg13g2_decap_8 FILLER_68_2047 ();
 sg13g2_decap_8 FILLER_68_2054 ();
 sg13g2_decap_8 FILLER_68_2061 ();
 sg13g2_decap_8 FILLER_68_2068 ();
 sg13g2_decap_8 FILLER_68_2075 ();
 sg13g2_decap_8 FILLER_68_2082 ();
 sg13g2_decap_8 FILLER_68_2089 ();
 sg13g2_decap_8 FILLER_68_2096 ();
 sg13g2_decap_8 FILLER_68_2103 ();
 sg13g2_decap_8 FILLER_68_2110 ();
 sg13g2_decap_8 FILLER_68_2117 ();
 sg13g2_decap_8 FILLER_68_2124 ();
 sg13g2_decap_8 FILLER_68_2131 ();
 sg13g2_decap_8 FILLER_68_2138 ();
 sg13g2_decap_8 FILLER_68_2145 ();
 sg13g2_decap_8 FILLER_68_2152 ();
 sg13g2_decap_8 FILLER_68_2159 ();
 sg13g2_decap_8 FILLER_68_2166 ();
 sg13g2_decap_8 FILLER_68_2173 ();
 sg13g2_decap_8 FILLER_68_2180 ();
 sg13g2_decap_8 FILLER_68_2187 ();
 sg13g2_decap_8 FILLER_68_2194 ();
 sg13g2_decap_8 FILLER_68_2201 ();
 sg13g2_decap_8 FILLER_68_2208 ();
 sg13g2_decap_8 FILLER_68_2215 ();
 sg13g2_decap_8 FILLER_68_2222 ();
 sg13g2_decap_8 FILLER_68_2229 ();
 sg13g2_decap_8 FILLER_68_2236 ();
 sg13g2_decap_8 FILLER_68_2243 ();
 sg13g2_decap_8 FILLER_68_2250 ();
 sg13g2_decap_8 FILLER_68_2257 ();
 sg13g2_decap_8 FILLER_68_2264 ();
 sg13g2_decap_8 FILLER_68_2271 ();
 sg13g2_decap_8 FILLER_68_2278 ();
 sg13g2_decap_8 FILLER_68_2285 ();
 sg13g2_decap_8 FILLER_68_2292 ();
 sg13g2_decap_8 FILLER_68_2299 ();
 sg13g2_decap_8 FILLER_68_2306 ();
 sg13g2_decap_8 FILLER_68_2313 ();
 sg13g2_decap_8 FILLER_68_2320 ();
 sg13g2_decap_8 FILLER_68_2327 ();
 sg13g2_decap_8 FILLER_68_2334 ();
 sg13g2_decap_8 FILLER_68_2341 ();
 sg13g2_decap_8 FILLER_68_2348 ();
 sg13g2_decap_8 FILLER_68_2355 ();
 sg13g2_decap_8 FILLER_68_2362 ();
 sg13g2_decap_8 FILLER_68_2369 ();
 sg13g2_decap_8 FILLER_68_2376 ();
 sg13g2_decap_8 FILLER_68_2383 ();
 sg13g2_decap_8 FILLER_68_2390 ();
 sg13g2_decap_8 FILLER_68_2397 ();
 sg13g2_decap_8 FILLER_68_2404 ();
 sg13g2_decap_8 FILLER_68_2411 ();
 sg13g2_decap_8 FILLER_68_2418 ();
 sg13g2_decap_8 FILLER_68_2425 ();
 sg13g2_decap_8 FILLER_68_2432 ();
 sg13g2_decap_8 FILLER_68_2439 ();
 sg13g2_decap_8 FILLER_68_2446 ();
 sg13g2_decap_8 FILLER_68_2453 ();
 sg13g2_decap_8 FILLER_68_2460 ();
 sg13g2_decap_8 FILLER_68_2467 ();
 sg13g2_decap_8 FILLER_68_2474 ();
 sg13g2_decap_8 FILLER_68_2481 ();
 sg13g2_decap_8 FILLER_68_2488 ();
 sg13g2_decap_8 FILLER_68_2495 ();
 sg13g2_decap_8 FILLER_68_2502 ();
 sg13g2_decap_8 FILLER_68_2509 ();
 sg13g2_decap_8 FILLER_68_2516 ();
 sg13g2_decap_8 FILLER_68_2523 ();
 sg13g2_decap_8 FILLER_68_2530 ();
 sg13g2_decap_8 FILLER_68_2537 ();
 sg13g2_decap_8 FILLER_68_2544 ();
 sg13g2_decap_8 FILLER_68_2551 ();
 sg13g2_decap_8 FILLER_68_2558 ();
 sg13g2_decap_8 FILLER_68_2565 ();
 sg13g2_decap_8 FILLER_68_2572 ();
 sg13g2_decap_8 FILLER_68_2579 ();
 sg13g2_decap_8 FILLER_68_2586 ();
 sg13g2_decap_8 FILLER_68_2593 ();
 sg13g2_decap_8 FILLER_68_2600 ();
 sg13g2_decap_8 FILLER_68_2607 ();
 sg13g2_decap_8 FILLER_68_2614 ();
 sg13g2_decap_8 FILLER_68_2621 ();
 sg13g2_decap_8 FILLER_68_2628 ();
 sg13g2_decap_8 FILLER_68_2635 ();
 sg13g2_decap_8 FILLER_68_2642 ();
 sg13g2_decap_8 FILLER_68_2649 ();
 sg13g2_decap_8 FILLER_68_2656 ();
 sg13g2_decap_8 FILLER_68_2663 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_46 ();
 sg13g2_decap_8 FILLER_69_53 ();
 sg13g2_decap_8 FILLER_69_60 ();
 sg13g2_decap_8 FILLER_69_67 ();
 sg13g2_decap_8 FILLER_69_74 ();
 sg13g2_decap_8 FILLER_69_81 ();
 sg13g2_decap_8 FILLER_69_88 ();
 sg13g2_decap_8 FILLER_69_95 ();
 sg13g2_decap_8 FILLER_69_102 ();
 sg13g2_decap_8 FILLER_69_109 ();
 sg13g2_decap_8 FILLER_69_116 ();
 sg13g2_decap_8 FILLER_69_123 ();
 sg13g2_decap_8 FILLER_69_130 ();
 sg13g2_decap_8 FILLER_69_137 ();
 sg13g2_decap_8 FILLER_69_144 ();
 sg13g2_decap_8 FILLER_69_151 ();
 sg13g2_decap_4 FILLER_69_158 ();
 sg13g2_decap_8 FILLER_69_166 ();
 sg13g2_decap_8 FILLER_69_173 ();
 sg13g2_decap_8 FILLER_69_180 ();
 sg13g2_decap_8 FILLER_69_187 ();
 sg13g2_decap_8 FILLER_69_194 ();
 sg13g2_decap_8 FILLER_69_201 ();
 sg13g2_decap_8 FILLER_69_208 ();
 sg13g2_decap_8 FILLER_69_219 ();
 sg13g2_decap_8 FILLER_69_226 ();
 sg13g2_decap_8 FILLER_69_233 ();
 sg13g2_decap_8 FILLER_69_240 ();
 sg13g2_decap_8 FILLER_69_247 ();
 sg13g2_decap_8 FILLER_69_254 ();
 sg13g2_decap_8 FILLER_69_261 ();
 sg13g2_fill_1 FILLER_69_268 ();
 sg13g2_decap_8 FILLER_69_273 ();
 sg13g2_decap_8 FILLER_69_280 ();
 sg13g2_decap_8 FILLER_69_287 ();
 sg13g2_decap_8 FILLER_69_294 ();
 sg13g2_fill_1 FILLER_69_301 ();
 sg13g2_decap_8 FILLER_69_313 ();
 sg13g2_decap_8 FILLER_69_320 ();
 sg13g2_decap_8 FILLER_69_327 ();
 sg13g2_decap_8 FILLER_69_334 ();
 sg13g2_decap_8 FILLER_69_341 ();
 sg13g2_decap_8 FILLER_69_348 ();
 sg13g2_decap_8 FILLER_69_355 ();
 sg13g2_decap_8 FILLER_69_362 ();
 sg13g2_decap_8 FILLER_69_369 ();
 sg13g2_decap_8 FILLER_69_376 ();
 sg13g2_decap_8 FILLER_69_383 ();
 sg13g2_decap_8 FILLER_69_390 ();
 sg13g2_decap_8 FILLER_69_397 ();
 sg13g2_decap_8 FILLER_69_404 ();
 sg13g2_decap_8 FILLER_69_411 ();
 sg13g2_decap_8 FILLER_69_418 ();
 sg13g2_decap_8 FILLER_69_425 ();
 sg13g2_fill_1 FILLER_69_432 ();
 sg13g2_decap_4 FILLER_69_438 ();
 sg13g2_decap_8 FILLER_69_465 ();
 sg13g2_decap_8 FILLER_69_472 ();
 sg13g2_fill_2 FILLER_69_479 ();
 sg13g2_decap_8 FILLER_69_485 ();
 sg13g2_decap_8 FILLER_69_492 ();
 sg13g2_decap_8 FILLER_69_499 ();
 sg13g2_decap_8 FILLER_69_506 ();
 sg13g2_decap_8 FILLER_69_513 ();
 sg13g2_decap_8 FILLER_69_520 ();
 sg13g2_decap_8 FILLER_69_527 ();
 sg13g2_decap_4 FILLER_69_534 ();
 sg13g2_fill_2 FILLER_69_538 ();
 sg13g2_fill_2 FILLER_69_544 ();
 sg13g2_fill_1 FILLER_69_546 ();
 sg13g2_fill_2 FILLER_69_556 ();
 sg13g2_decap_8 FILLER_69_570 ();
 sg13g2_decap_4 FILLER_69_577 ();
 sg13g2_fill_2 FILLER_69_581 ();
 sg13g2_decap_4 FILLER_69_587 ();
 sg13g2_decap_8 FILLER_69_595 ();
 sg13g2_decap_8 FILLER_69_602 ();
 sg13g2_decap_8 FILLER_69_609 ();
 sg13g2_decap_4 FILLER_69_616 ();
 sg13g2_fill_1 FILLER_69_620 ();
 sg13g2_decap_8 FILLER_69_626 ();
 sg13g2_decap_8 FILLER_69_633 ();
 sg13g2_decap_8 FILLER_69_640 ();
 sg13g2_decap_4 FILLER_69_647 ();
 sg13g2_fill_2 FILLER_69_651 ();
 sg13g2_decap_4 FILLER_69_656 ();
 sg13g2_fill_2 FILLER_69_660 ();
 sg13g2_decap_8 FILLER_69_695 ();
 sg13g2_decap_8 FILLER_69_702 ();
 sg13g2_decap_8 FILLER_69_709 ();
 sg13g2_fill_1 FILLER_69_716 ();
 sg13g2_decap_8 FILLER_69_726 ();
 sg13g2_decap_8 FILLER_69_733 ();
 sg13g2_decap_8 FILLER_69_740 ();
 sg13g2_decap_8 FILLER_69_747 ();
 sg13g2_decap_8 FILLER_69_754 ();
 sg13g2_decap_8 FILLER_69_761 ();
 sg13g2_decap_8 FILLER_69_768 ();
 sg13g2_decap_4 FILLER_69_775 ();
 sg13g2_fill_2 FILLER_69_779 ();
 sg13g2_decap_8 FILLER_69_791 ();
 sg13g2_decap_8 FILLER_69_798 ();
 sg13g2_decap_8 FILLER_69_805 ();
 sg13g2_decap_8 FILLER_69_812 ();
 sg13g2_decap_8 FILLER_69_819 ();
 sg13g2_decap_4 FILLER_69_832 ();
 sg13g2_fill_2 FILLER_69_836 ();
 sg13g2_decap_8 FILLER_69_875 ();
 sg13g2_decap_8 FILLER_69_882 ();
 sg13g2_decap_8 FILLER_69_889 ();
 sg13g2_decap_8 FILLER_69_896 ();
 sg13g2_decap_8 FILLER_69_903 ();
 sg13g2_decap_4 FILLER_69_910 ();
 sg13g2_fill_1 FILLER_69_914 ();
 sg13g2_decap_8 FILLER_69_920 ();
 sg13g2_decap_8 FILLER_69_927 ();
 sg13g2_decap_8 FILLER_69_934 ();
 sg13g2_fill_1 FILLER_69_941 ();
 sg13g2_decap_8 FILLER_69_948 ();
 sg13g2_decap_8 FILLER_69_955 ();
 sg13g2_decap_8 FILLER_69_962 ();
 sg13g2_decap_4 FILLER_69_969 ();
 sg13g2_decap_8 FILLER_69_985 ();
 sg13g2_decap_8 FILLER_69_992 ();
 sg13g2_decap_8 FILLER_69_1008 ();
 sg13g2_decap_8 FILLER_69_1015 ();
 sg13g2_decap_8 FILLER_69_1022 ();
 sg13g2_decap_4 FILLER_69_1029 ();
 sg13g2_fill_2 FILLER_69_1033 ();
 sg13g2_decap_8 FILLER_69_1040 ();
 sg13g2_decap_8 FILLER_69_1047 ();
 sg13g2_decap_8 FILLER_69_1054 ();
 sg13g2_decap_8 FILLER_69_1061 ();
 sg13g2_decap_8 FILLER_69_1068 ();
 sg13g2_decap_8 FILLER_69_1075 ();
 sg13g2_decap_8 FILLER_69_1082 ();
 sg13g2_decap_8 FILLER_69_1089 ();
 sg13g2_decap_8 FILLER_69_1100 ();
 sg13g2_decap_8 FILLER_69_1107 ();
 sg13g2_decap_8 FILLER_69_1114 ();
 sg13g2_decap_8 FILLER_69_1121 ();
 sg13g2_fill_1 FILLER_69_1128 ();
 sg13g2_decap_8 FILLER_69_1139 ();
 sg13g2_decap_4 FILLER_69_1146 ();
 sg13g2_fill_2 FILLER_69_1150 ();
 sg13g2_decap_8 FILLER_69_1174 ();
 sg13g2_decap_8 FILLER_69_1181 ();
 sg13g2_decap_8 FILLER_69_1188 ();
 sg13g2_decap_8 FILLER_69_1195 ();
 sg13g2_decap_8 FILLER_69_1207 ();
 sg13g2_decap_8 FILLER_69_1214 ();
 sg13g2_decap_8 FILLER_69_1221 ();
 sg13g2_fill_1 FILLER_69_1228 ();
 sg13g2_decap_8 FILLER_69_1233 ();
 sg13g2_decap_8 FILLER_69_1240 ();
 sg13g2_decap_8 FILLER_69_1247 ();
 sg13g2_decap_8 FILLER_69_1254 ();
 sg13g2_decap_8 FILLER_69_1261 ();
 sg13g2_decap_8 FILLER_69_1268 ();
 sg13g2_decap_8 FILLER_69_1275 ();
 sg13g2_fill_2 FILLER_69_1282 ();
 sg13g2_decap_8 FILLER_69_1287 ();
 sg13g2_decap_8 FILLER_69_1294 ();
 sg13g2_decap_8 FILLER_69_1301 ();
 sg13g2_fill_2 FILLER_69_1313 ();
 sg13g2_decap_8 FILLER_69_1320 ();
 sg13g2_decap_8 FILLER_69_1327 ();
 sg13g2_decap_8 FILLER_69_1334 ();
 sg13g2_decap_8 FILLER_69_1341 ();
 sg13g2_decap_8 FILLER_69_1356 ();
 sg13g2_decap_8 FILLER_69_1363 ();
 sg13g2_decap_4 FILLER_69_1370 ();
 sg13g2_fill_1 FILLER_69_1374 ();
 sg13g2_decap_4 FILLER_69_1379 ();
 sg13g2_fill_2 FILLER_69_1383 ();
 sg13g2_decap_4 FILLER_69_1389 ();
 sg13g2_fill_1 FILLER_69_1393 ();
 sg13g2_decap_8 FILLER_69_1409 ();
 sg13g2_decap_8 FILLER_69_1416 ();
 sg13g2_decap_8 FILLER_69_1423 ();
 sg13g2_decap_8 FILLER_69_1430 ();
 sg13g2_decap_8 FILLER_69_1437 ();
 sg13g2_decap_8 FILLER_69_1444 ();
 sg13g2_decap_8 FILLER_69_1451 ();
 sg13g2_decap_8 FILLER_69_1458 ();
 sg13g2_decap_8 FILLER_69_1465 ();
 sg13g2_decap_4 FILLER_69_1472 ();
 sg13g2_fill_2 FILLER_69_1476 ();
 sg13g2_decap_8 FILLER_69_1483 ();
 sg13g2_decap_4 FILLER_69_1490 ();
 sg13g2_fill_1 FILLER_69_1494 ();
 sg13g2_decap_4 FILLER_69_1514 ();
 sg13g2_fill_2 FILLER_69_1518 ();
 sg13g2_decap_4 FILLER_69_1535 ();
 sg13g2_fill_2 FILLER_69_1539 ();
 sg13g2_decap_8 FILLER_69_1544 ();
 sg13g2_decap_8 FILLER_69_1551 ();
 sg13g2_decap_8 FILLER_69_1558 ();
 sg13g2_decap_8 FILLER_69_1565 ();
 sg13g2_decap_8 FILLER_69_1577 ();
 sg13g2_decap_8 FILLER_69_1584 ();
 sg13g2_decap_8 FILLER_69_1591 ();
 sg13g2_decap_8 FILLER_69_1598 ();
 sg13g2_decap_8 FILLER_69_1605 ();
 sg13g2_decap_8 FILLER_69_1612 ();
 sg13g2_fill_2 FILLER_69_1619 ();
 sg13g2_fill_1 FILLER_69_1621 ();
 sg13g2_decap_8 FILLER_69_1637 ();
 sg13g2_decap_8 FILLER_69_1647 ();
 sg13g2_decap_8 FILLER_69_1654 ();
 sg13g2_decap_8 FILLER_69_1661 ();
 sg13g2_decap_8 FILLER_69_1668 ();
 sg13g2_decap_8 FILLER_69_1675 ();
 sg13g2_decap_8 FILLER_69_1682 ();
 sg13g2_decap_8 FILLER_69_1689 ();
 sg13g2_decap_8 FILLER_69_1696 ();
 sg13g2_decap_8 FILLER_69_1703 ();
 sg13g2_decap_8 FILLER_69_1710 ();
 sg13g2_decap_8 FILLER_69_1717 ();
 sg13g2_decap_8 FILLER_69_1724 ();
 sg13g2_decap_8 FILLER_69_1731 ();
 sg13g2_decap_8 FILLER_69_1738 ();
 sg13g2_decap_8 FILLER_69_1745 ();
 sg13g2_decap_8 FILLER_69_1752 ();
 sg13g2_fill_2 FILLER_69_1759 ();
 sg13g2_decap_8 FILLER_69_1765 ();
 sg13g2_decap_8 FILLER_69_1772 ();
 sg13g2_decap_8 FILLER_69_1779 ();
 sg13g2_decap_8 FILLER_69_1786 ();
 sg13g2_decap_8 FILLER_69_1793 ();
 sg13g2_decap_8 FILLER_69_1800 ();
 sg13g2_decap_8 FILLER_69_1807 ();
 sg13g2_decap_8 FILLER_69_1814 ();
 sg13g2_decap_8 FILLER_69_1821 ();
 sg13g2_decap_8 FILLER_69_1828 ();
 sg13g2_decap_8 FILLER_69_1835 ();
 sg13g2_decap_8 FILLER_69_1842 ();
 sg13g2_decap_8 FILLER_69_1849 ();
 sg13g2_decap_8 FILLER_69_1856 ();
 sg13g2_decap_8 FILLER_69_1863 ();
 sg13g2_decap_8 FILLER_69_1870 ();
 sg13g2_decap_8 FILLER_69_1877 ();
 sg13g2_decap_8 FILLER_69_1884 ();
 sg13g2_decap_8 FILLER_69_1891 ();
 sg13g2_decap_8 FILLER_69_1898 ();
 sg13g2_decap_8 FILLER_69_1905 ();
 sg13g2_decap_8 FILLER_69_1912 ();
 sg13g2_decap_8 FILLER_69_1919 ();
 sg13g2_decap_8 FILLER_69_1926 ();
 sg13g2_decap_8 FILLER_69_1933 ();
 sg13g2_decap_8 FILLER_69_1940 ();
 sg13g2_decap_8 FILLER_69_1947 ();
 sg13g2_decap_8 FILLER_69_1954 ();
 sg13g2_decap_4 FILLER_69_1961 ();
 sg13g2_decap_8 FILLER_69_1969 ();
 sg13g2_decap_8 FILLER_69_1976 ();
 sg13g2_decap_8 FILLER_69_1983 ();
 sg13g2_decap_8 FILLER_69_1990 ();
 sg13g2_decap_8 FILLER_69_1997 ();
 sg13g2_decap_8 FILLER_69_2004 ();
 sg13g2_decap_8 FILLER_69_2011 ();
 sg13g2_fill_2 FILLER_69_2018 ();
 sg13g2_decap_8 FILLER_69_2034 ();
 sg13g2_decap_8 FILLER_69_2041 ();
 sg13g2_decap_8 FILLER_69_2048 ();
 sg13g2_decap_4 FILLER_69_2055 ();
 sg13g2_decap_8 FILLER_69_2065 ();
 sg13g2_decap_8 FILLER_69_2072 ();
 sg13g2_decap_8 FILLER_69_2079 ();
 sg13g2_decap_8 FILLER_69_2086 ();
 sg13g2_decap_8 FILLER_69_2093 ();
 sg13g2_fill_2 FILLER_69_2100 ();
 sg13g2_fill_1 FILLER_69_2102 ();
 sg13g2_decap_8 FILLER_69_2106 ();
 sg13g2_decap_8 FILLER_69_2113 ();
 sg13g2_decap_8 FILLER_69_2120 ();
 sg13g2_decap_8 FILLER_69_2127 ();
 sg13g2_decap_8 FILLER_69_2134 ();
 sg13g2_decap_8 FILLER_69_2141 ();
 sg13g2_decap_8 FILLER_69_2148 ();
 sg13g2_fill_1 FILLER_69_2155 ();
 sg13g2_decap_8 FILLER_69_2162 ();
 sg13g2_decap_8 FILLER_69_2169 ();
 sg13g2_decap_8 FILLER_69_2176 ();
 sg13g2_decap_4 FILLER_69_2183 ();
 sg13g2_fill_2 FILLER_69_2187 ();
 sg13g2_decap_8 FILLER_69_2192 ();
 sg13g2_decap_8 FILLER_69_2199 ();
 sg13g2_decap_8 FILLER_69_2206 ();
 sg13g2_decap_8 FILLER_69_2213 ();
 sg13g2_decap_8 FILLER_69_2220 ();
 sg13g2_decap_8 FILLER_69_2227 ();
 sg13g2_decap_8 FILLER_69_2234 ();
 sg13g2_decap_8 FILLER_69_2241 ();
 sg13g2_decap_8 FILLER_69_2248 ();
 sg13g2_decap_8 FILLER_69_2255 ();
 sg13g2_decap_8 FILLER_69_2262 ();
 sg13g2_decap_8 FILLER_69_2269 ();
 sg13g2_decap_8 FILLER_69_2276 ();
 sg13g2_decap_8 FILLER_69_2283 ();
 sg13g2_decap_8 FILLER_69_2290 ();
 sg13g2_decap_8 FILLER_69_2297 ();
 sg13g2_decap_8 FILLER_69_2304 ();
 sg13g2_decap_8 FILLER_69_2311 ();
 sg13g2_decap_8 FILLER_69_2318 ();
 sg13g2_decap_8 FILLER_69_2325 ();
 sg13g2_decap_8 FILLER_69_2332 ();
 sg13g2_decap_8 FILLER_69_2339 ();
 sg13g2_decap_8 FILLER_69_2346 ();
 sg13g2_decap_8 FILLER_69_2353 ();
 sg13g2_decap_8 FILLER_69_2360 ();
 sg13g2_decap_8 FILLER_69_2367 ();
 sg13g2_decap_8 FILLER_69_2374 ();
 sg13g2_decap_8 FILLER_69_2381 ();
 sg13g2_decap_8 FILLER_69_2388 ();
 sg13g2_decap_8 FILLER_69_2395 ();
 sg13g2_decap_8 FILLER_69_2402 ();
 sg13g2_decap_8 FILLER_69_2409 ();
 sg13g2_decap_8 FILLER_69_2416 ();
 sg13g2_decap_8 FILLER_69_2423 ();
 sg13g2_decap_8 FILLER_69_2430 ();
 sg13g2_decap_8 FILLER_69_2437 ();
 sg13g2_decap_8 FILLER_69_2444 ();
 sg13g2_decap_8 FILLER_69_2451 ();
 sg13g2_decap_8 FILLER_69_2458 ();
 sg13g2_decap_8 FILLER_69_2465 ();
 sg13g2_decap_8 FILLER_69_2472 ();
 sg13g2_decap_8 FILLER_69_2479 ();
 sg13g2_decap_8 FILLER_69_2486 ();
 sg13g2_decap_8 FILLER_69_2493 ();
 sg13g2_decap_8 FILLER_69_2500 ();
 sg13g2_decap_8 FILLER_69_2507 ();
 sg13g2_decap_8 FILLER_69_2514 ();
 sg13g2_decap_8 FILLER_69_2521 ();
 sg13g2_decap_8 FILLER_69_2528 ();
 sg13g2_decap_8 FILLER_69_2535 ();
 sg13g2_decap_8 FILLER_69_2542 ();
 sg13g2_decap_8 FILLER_69_2549 ();
 sg13g2_decap_8 FILLER_69_2556 ();
 sg13g2_decap_8 FILLER_69_2563 ();
 sg13g2_decap_8 FILLER_69_2570 ();
 sg13g2_decap_8 FILLER_69_2577 ();
 sg13g2_decap_8 FILLER_69_2584 ();
 sg13g2_decap_8 FILLER_69_2591 ();
 sg13g2_decap_8 FILLER_69_2598 ();
 sg13g2_decap_8 FILLER_69_2605 ();
 sg13g2_decap_8 FILLER_69_2612 ();
 sg13g2_decap_8 FILLER_69_2619 ();
 sg13g2_decap_8 FILLER_69_2626 ();
 sg13g2_decap_8 FILLER_69_2633 ();
 sg13g2_decap_8 FILLER_69_2640 ();
 sg13g2_decap_8 FILLER_69_2647 ();
 sg13g2_decap_8 FILLER_69_2654 ();
 sg13g2_decap_8 FILLER_69_2661 ();
 sg13g2_fill_2 FILLER_69_2668 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_8 FILLER_70_105 ();
 sg13g2_decap_8 FILLER_70_112 ();
 sg13g2_decap_8 FILLER_70_119 ();
 sg13g2_decap_8 FILLER_70_126 ();
 sg13g2_decap_8 FILLER_70_133 ();
 sg13g2_decap_8 FILLER_70_140 ();
 sg13g2_decap_8 FILLER_70_147 ();
 sg13g2_decap_8 FILLER_70_154 ();
 sg13g2_decap_8 FILLER_70_161 ();
 sg13g2_decap_8 FILLER_70_168 ();
 sg13g2_decap_8 FILLER_70_175 ();
 sg13g2_decap_8 FILLER_70_182 ();
 sg13g2_decap_8 FILLER_70_189 ();
 sg13g2_decap_8 FILLER_70_196 ();
 sg13g2_decap_8 FILLER_70_203 ();
 sg13g2_decap_8 FILLER_70_210 ();
 sg13g2_decap_8 FILLER_70_217 ();
 sg13g2_decap_8 FILLER_70_224 ();
 sg13g2_decap_8 FILLER_70_231 ();
 sg13g2_decap_8 FILLER_70_238 ();
 sg13g2_decap_8 FILLER_70_245 ();
 sg13g2_decap_8 FILLER_70_252 ();
 sg13g2_decap_8 FILLER_70_259 ();
 sg13g2_decap_8 FILLER_70_266 ();
 sg13g2_decap_8 FILLER_70_273 ();
 sg13g2_decap_8 FILLER_70_280 ();
 sg13g2_decap_8 FILLER_70_287 ();
 sg13g2_decap_8 FILLER_70_294 ();
 sg13g2_decap_8 FILLER_70_301 ();
 sg13g2_decap_8 FILLER_70_308 ();
 sg13g2_decap_8 FILLER_70_315 ();
 sg13g2_decap_8 FILLER_70_322 ();
 sg13g2_decap_8 FILLER_70_329 ();
 sg13g2_decap_8 FILLER_70_336 ();
 sg13g2_decap_8 FILLER_70_343 ();
 sg13g2_decap_8 FILLER_70_350 ();
 sg13g2_decap_8 FILLER_70_357 ();
 sg13g2_decap_8 FILLER_70_364 ();
 sg13g2_decap_4 FILLER_70_371 ();
 sg13g2_fill_1 FILLER_70_375 ();
 sg13g2_fill_2 FILLER_70_381 ();
 sg13g2_fill_1 FILLER_70_383 ();
 sg13g2_decap_8 FILLER_70_388 ();
 sg13g2_decap_8 FILLER_70_395 ();
 sg13g2_decap_8 FILLER_70_402 ();
 sg13g2_decap_8 FILLER_70_409 ();
 sg13g2_decap_8 FILLER_70_416 ();
 sg13g2_decap_8 FILLER_70_423 ();
 sg13g2_decap_8 FILLER_70_430 ();
 sg13g2_decap_8 FILLER_70_437 ();
 sg13g2_decap_8 FILLER_70_444 ();
 sg13g2_decap_8 FILLER_70_451 ();
 sg13g2_decap_4 FILLER_70_458 ();
 sg13g2_fill_2 FILLER_70_462 ();
 sg13g2_decap_8 FILLER_70_468 ();
 sg13g2_decap_8 FILLER_70_475 ();
 sg13g2_decap_8 FILLER_70_482 ();
 sg13g2_fill_2 FILLER_70_489 ();
 sg13g2_decap_8 FILLER_70_506 ();
 sg13g2_decap_8 FILLER_70_513 ();
 sg13g2_decap_8 FILLER_70_520 ();
 sg13g2_decap_8 FILLER_70_527 ();
 sg13g2_decap_4 FILLER_70_534 ();
 sg13g2_fill_2 FILLER_70_538 ();
 sg13g2_decap_4 FILLER_70_544 ();
 sg13g2_fill_1 FILLER_70_548 ();
 sg13g2_fill_1 FILLER_70_554 ();
 sg13g2_decap_8 FILLER_70_565 ();
 sg13g2_decap_8 FILLER_70_572 ();
 sg13g2_decap_8 FILLER_70_579 ();
 sg13g2_decap_8 FILLER_70_586 ();
 sg13g2_fill_1 FILLER_70_593 ();
 sg13g2_decap_8 FILLER_70_598 ();
 sg13g2_decap_8 FILLER_70_605 ();
 sg13g2_decap_8 FILLER_70_612 ();
 sg13g2_fill_2 FILLER_70_619 ();
 sg13g2_decap_8 FILLER_70_636 ();
 sg13g2_decap_8 FILLER_70_643 ();
 sg13g2_decap_8 FILLER_70_650 ();
 sg13g2_decap_8 FILLER_70_657 ();
 sg13g2_decap_8 FILLER_70_664 ();
 sg13g2_decap_8 FILLER_70_671 ();
 sg13g2_decap_4 FILLER_70_678 ();
 sg13g2_fill_1 FILLER_70_682 ();
 sg13g2_decap_8 FILLER_70_689 ();
 sg13g2_decap_8 FILLER_70_696 ();
 sg13g2_decap_8 FILLER_70_703 ();
 sg13g2_decap_8 FILLER_70_710 ();
 sg13g2_decap_8 FILLER_70_722 ();
 sg13g2_decap_8 FILLER_70_729 ();
 sg13g2_decap_8 FILLER_70_736 ();
 sg13g2_decap_8 FILLER_70_743 ();
 sg13g2_decap_8 FILLER_70_750 ();
 sg13g2_decap_8 FILLER_70_757 ();
 sg13g2_decap_8 FILLER_70_764 ();
 sg13g2_decap_8 FILLER_70_771 ();
 sg13g2_decap_8 FILLER_70_778 ();
 sg13g2_decap_8 FILLER_70_785 ();
 sg13g2_decap_8 FILLER_70_792 ();
 sg13g2_decap_8 FILLER_70_799 ();
 sg13g2_fill_1 FILLER_70_806 ();
 sg13g2_decap_8 FILLER_70_822 ();
 sg13g2_decap_8 FILLER_70_829 ();
 sg13g2_decap_8 FILLER_70_836 ();
 sg13g2_decap_8 FILLER_70_843 ();
 sg13g2_decap_4 FILLER_70_850 ();
 sg13g2_fill_2 FILLER_70_854 ();
 sg13g2_decap_8 FILLER_70_862 ();
 sg13g2_decap_8 FILLER_70_869 ();
 sg13g2_decap_8 FILLER_70_876 ();
 sg13g2_decap_8 FILLER_70_883 ();
 sg13g2_decap_8 FILLER_70_890 ();
 sg13g2_decap_8 FILLER_70_897 ();
 sg13g2_decap_8 FILLER_70_904 ();
 sg13g2_decap_4 FILLER_70_911 ();
 sg13g2_decap_8 FILLER_70_924 ();
 sg13g2_decap_8 FILLER_70_931 ();
 sg13g2_decap_8 FILLER_70_938 ();
 sg13g2_fill_1 FILLER_70_945 ();
 sg13g2_decap_8 FILLER_70_949 ();
 sg13g2_decap_8 FILLER_70_956 ();
 sg13g2_decap_8 FILLER_70_963 ();
 sg13g2_decap_8 FILLER_70_979 ();
 sg13g2_decap_8 FILLER_70_986 ();
 sg13g2_decap_4 FILLER_70_993 ();
 sg13g2_fill_2 FILLER_70_997 ();
 sg13g2_fill_1 FILLER_70_1002 ();
 sg13g2_decap_8 FILLER_70_1018 ();
 sg13g2_decap_8 FILLER_70_1025 ();
 sg13g2_decap_8 FILLER_70_1032 ();
 sg13g2_fill_2 FILLER_70_1039 ();
 sg13g2_decap_8 FILLER_70_1045 ();
 sg13g2_decap_8 FILLER_70_1052 ();
 sg13g2_decap_8 FILLER_70_1059 ();
 sg13g2_fill_2 FILLER_70_1066 ();
 sg13g2_fill_1 FILLER_70_1068 ();
 sg13g2_decap_8 FILLER_70_1084 ();
 sg13g2_decap_8 FILLER_70_1091 ();
 sg13g2_fill_1 FILLER_70_1098 ();
 sg13g2_decap_8 FILLER_70_1104 ();
 sg13g2_decap_8 FILLER_70_1111 ();
 sg13g2_decap_8 FILLER_70_1118 ();
 sg13g2_decap_8 FILLER_70_1125 ();
 sg13g2_decap_8 FILLER_70_1132 ();
 sg13g2_fill_2 FILLER_70_1139 ();
 sg13g2_fill_2 FILLER_70_1160 ();
 sg13g2_decap_8 FILLER_70_1165 ();
 sg13g2_decap_8 FILLER_70_1172 ();
 sg13g2_decap_8 FILLER_70_1179 ();
 sg13g2_decap_8 FILLER_70_1186 ();
 sg13g2_decap_8 FILLER_70_1193 ();
 sg13g2_decap_8 FILLER_70_1200 ();
 sg13g2_decap_8 FILLER_70_1207 ();
 sg13g2_decap_8 FILLER_70_1214 ();
 sg13g2_decap_8 FILLER_70_1221 ();
 sg13g2_decap_4 FILLER_70_1228 ();
 sg13g2_fill_2 FILLER_70_1232 ();
 sg13g2_decap_8 FILLER_70_1249 ();
 sg13g2_decap_8 FILLER_70_1256 ();
 sg13g2_decap_4 FILLER_70_1263 ();
 sg13g2_decap_8 FILLER_70_1272 ();
 sg13g2_decap_4 FILLER_70_1279 ();
 sg13g2_fill_1 FILLER_70_1283 ();
 sg13g2_decap_8 FILLER_70_1288 ();
 sg13g2_decap_8 FILLER_70_1295 ();
 sg13g2_decap_8 FILLER_70_1302 ();
 sg13g2_decap_4 FILLER_70_1309 ();
 sg13g2_fill_1 FILLER_70_1313 ();
 sg13g2_decap_8 FILLER_70_1319 ();
 sg13g2_decap_8 FILLER_70_1326 ();
 sg13g2_decap_4 FILLER_70_1333 ();
 sg13g2_fill_2 FILLER_70_1337 ();
 sg13g2_decap_4 FILLER_70_1344 ();
 sg13g2_decap_8 FILLER_70_1367 ();
 sg13g2_decap_8 FILLER_70_1374 ();
 sg13g2_decap_8 FILLER_70_1381 ();
 sg13g2_decap_4 FILLER_70_1388 ();
 sg13g2_fill_2 FILLER_70_1392 ();
 sg13g2_decap_8 FILLER_70_1398 ();
 sg13g2_decap_8 FILLER_70_1405 ();
 sg13g2_decap_8 FILLER_70_1412 ();
 sg13g2_fill_2 FILLER_70_1419 ();
 sg13g2_decap_8 FILLER_70_1426 ();
 sg13g2_decap_8 FILLER_70_1433 ();
 sg13g2_decap_8 FILLER_70_1440 ();
 sg13g2_decap_8 FILLER_70_1447 ();
 sg13g2_decap_8 FILLER_70_1454 ();
 sg13g2_decap_8 FILLER_70_1461 ();
 sg13g2_decap_8 FILLER_70_1468 ();
 sg13g2_fill_2 FILLER_70_1475 ();
 sg13g2_fill_1 FILLER_70_1477 ();
 sg13g2_decap_4 FILLER_70_1481 ();
 sg13g2_fill_1 FILLER_70_1485 ();
 sg13g2_fill_2 FILLER_70_1498 ();
 sg13g2_fill_2 FILLER_70_1505 ();
 sg13g2_fill_1 FILLER_70_1507 ();
 sg13g2_decap_4 FILLER_70_1513 ();
 sg13g2_decap_8 FILLER_70_1524 ();
 sg13g2_fill_2 FILLER_70_1531 ();
 sg13g2_decap_8 FILLER_70_1538 ();
 sg13g2_decap_8 FILLER_70_1545 ();
 sg13g2_decap_8 FILLER_70_1552 ();
 sg13g2_decap_8 FILLER_70_1559 ();
 sg13g2_decap_8 FILLER_70_1566 ();
 sg13g2_decap_8 FILLER_70_1573 ();
 sg13g2_decap_8 FILLER_70_1580 ();
 sg13g2_decap_8 FILLER_70_1587 ();
 sg13g2_decap_8 FILLER_70_1594 ();
 sg13g2_decap_8 FILLER_70_1601 ();
 sg13g2_decap_8 FILLER_70_1608 ();
 sg13g2_decap_8 FILLER_70_1615 ();
 sg13g2_decap_8 FILLER_70_1622 ();
 sg13g2_decap_8 FILLER_70_1629 ();
 sg13g2_decap_8 FILLER_70_1636 ();
 sg13g2_decap_8 FILLER_70_1643 ();
 sg13g2_decap_8 FILLER_70_1650 ();
 sg13g2_decap_8 FILLER_70_1665 ();
 sg13g2_decap_8 FILLER_70_1672 ();
 sg13g2_decap_8 FILLER_70_1679 ();
 sg13g2_decap_8 FILLER_70_1686 ();
 sg13g2_decap_4 FILLER_70_1693 ();
 sg13g2_fill_2 FILLER_70_1697 ();
 sg13g2_decap_8 FILLER_70_1702 ();
 sg13g2_decap_8 FILLER_70_1709 ();
 sg13g2_decap_8 FILLER_70_1716 ();
 sg13g2_decap_8 FILLER_70_1723 ();
 sg13g2_decap_8 FILLER_70_1730 ();
 sg13g2_decap_8 FILLER_70_1737 ();
 sg13g2_fill_2 FILLER_70_1744 ();
 sg13g2_fill_1 FILLER_70_1746 ();
 sg13g2_decap_8 FILLER_70_1759 ();
 sg13g2_decap_8 FILLER_70_1766 ();
 sg13g2_decap_8 FILLER_70_1773 ();
 sg13g2_decap_8 FILLER_70_1780 ();
 sg13g2_decap_8 FILLER_70_1787 ();
 sg13g2_decap_8 FILLER_70_1794 ();
 sg13g2_decap_8 FILLER_70_1801 ();
 sg13g2_decap_8 FILLER_70_1808 ();
 sg13g2_decap_8 FILLER_70_1815 ();
 sg13g2_decap_8 FILLER_70_1822 ();
 sg13g2_decap_8 FILLER_70_1829 ();
 sg13g2_decap_8 FILLER_70_1836 ();
 sg13g2_decap_8 FILLER_70_1843 ();
 sg13g2_decap_8 FILLER_70_1850 ();
 sg13g2_decap_8 FILLER_70_1857 ();
 sg13g2_decap_8 FILLER_70_1864 ();
 sg13g2_decap_8 FILLER_70_1871 ();
 sg13g2_decap_8 FILLER_70_1878 ();
 sg13g2_decap_8 FILLER_70_1885 ();
 sg13g2_decap_8 FILLER_70_1892 ();
 sg13g2_decap_8 FILLER_70_1899 ();
 sg13g2_decap_8 FILLER_70_1906 ();
 sg13g2_decap_8 FILLER_70_1913 ();
 sg13g2_decap_8 FILLER_70_1920 ();
 sg13g2_decap_8 FILLER_70_1927 ();
 sg13g2_decap_8 FILLER_70_1934 ();
 sg13g2_decap_8 FILLER_70_1941 ();
 sg13g2_decap_8 FILLER_70_1948 ();
 sg13g2_decap_8 FILLER_70_1955 ();
 sg13g2_decap_8 FILLER_70_1962 ();
 sg13g2_decap_8 FILLER_70_1969 ();
 sg13g2_decap_8 FILLER_70_1976 ();
 sg13g2_decap_8 FILLER_70_1983 ();
 sg13g2_decap_8 FILLER_70_1990 ();
 sg13g2_decap_8 FILLER_70_1997 ();
 sg13g2_decap_8 FILLER_70_2004 ();
 sg13g2_decap_8 FILLER_70_2011 ();
 sg13g2_decap_8 FILLER_70_2018 ();
 sg13g2_decap_8 FILLER_70_2025 ();
 sg13g2_decap_8 FILLER_70_2032 ();
 sg13g2_decap_8 FILLER_70_2039 ();
 sg13g2_decap_8 FILLER_70_2046 ();
 sg13g2_decap_4 FILLER_70_2053 ();
 sg13g2_fill_2 FILLER_70_2057 ();
 sg13g2_decap_8 FILLER_70_2062 ();
 sg13g2_decap_8 FILLER_70_2069 ();
 sg13g2_decap_8 FILLER_70_2076 ();
 sg13g2_decap_8 FILLER_70_2083 ();
 sg13g2_decap_4 FILLER_70_2090 ();
 sg13g2_fill_2 FILLER_70_2094 ();
 sg13g2_fill_2 FILLER_70_2108 ();
 sg13g2_fill_1 FILLER_70_2110 ();
 sg13g2_decap_8 FILLER_70_2120 ();
 sg13g2_decap_8 FILLER_70_2127 ();
 sg13g2_decap_8 FILLER_70_2134 ();
 sg13g2_decap_8 FILLER_70_2141 ();
 sg13g2_decap_8 FILLER_70_2148 ();
 sg13g2_fill_1 FILLER_70_2155 ();
 sg13g2_decap_8 FILLER_70_2167 ();
 sg13g2_decap_8 FILLER_70_2174 ();
 sg13g2_decap_8 FILLER_70_2181 ();
 sg13g2_decap_4 FILLER_70_2200 ();
 sg13g2_fill_1 FILLER_70_2204 ();
 sg13g2_decap_8 FILLER_70_2231 ();
 sg13g2_decap_8 FILLER_70_2238 ();
 sg13g2_decap_8 FILLER_70_2245 ();
 sg13g2_decap_8 FILLER_70_2252 ();
 sg13g2_decap_8 FILLER_70_2259 ();
 sg13g2_decap_8 FILLER_70_2266 ();
 sg13g2_decap_8 FILLER_70_2273 ();
 sg13g2_decap_8 FILLER_70_2280 ();
 sg13g2_decap_8 FILLER_70_2287 ();
 sg13g2_decap_8 FILLER_70_2294 ();
 sg13g2_decap_8 FILLER_70_2301 ();
 sg13g2_decap_8 FILLER_70_2308 ();
 sg13g2_decap_8 FILLER_70_2315 ();
 sg13g2_decap_8 FILLER_70_2322 ();
 sg13g2_decap_8 FILLER_70_2329 ();
 sg13g2_decap_8 FILLER_70_2336 ();
 sg13g2_decap_8 FILLER_70_2343 ();
 sg13g2_decap_8 FILLER_70_2350 ();
 sg13g2_decap_8 FILLER_70_2357 ();
 sg13g2_decap_8 FILLER_70_2364 ();
 sg13g2_decap_8 FILLER_70_2371 ();
 sg13g2_decap_8 FILLER_70_2378 ();
 sg13g2_decap_8 FILLER_70_2385 ();
 sg13g2_decap_8 FILLER_70_2392 ();
 sg13g2_decap_8 FILLER_70_2399 ();
 sg13g2_decap_8 FILLER_70_2406 ();
 sg13g2_decap_8 FILLER_70_2413 ();
 sg13g2_decap_8 FILLER_70_2420 ();
 sg13g2_decap_8 FILLER_70_2427 ();
 sg13g2_decap_8 FILLER_70_2434 ();
 sg13g2_decap_8 FILLER_70_2441 ();
 sg13g2_decap_8 FILLER_70_2448 ();
 sg13g2_decap_8 FILLER_70_2455 ();
 sg13g2_decap_8 FILLER_70_2462 ();
 sg13g2_decap_8 FILLER_70_2469 ();
 sg13g2_decap_8 FILLER_70_2476 ();
 sg13g2_decap_8 FILLER_70_2483 ();
 sg13g2_decap_8 FILLER_70_2490 ();
 sg13g2_decap_8 FILLER_70_2497 ();
 sg13g2_decap_8 FILLER_70_2504 ();
 sg13g2_decap_8 FILLER_70_2511 ();
 sg13g2_decap_8 FILLER_70_2518 ();
 sg13g2_decap_8 FILLER_70_2525 ();
 sg13g2_decap_8 FILLER_70_2532 ();
 sg13g2_decap_8 FILLER_70_2539 ();
 sg13g2_decap_8 FILLER_70_2546 ();
 sg13g2_decap_8 FILLER_70_2553 ();
 sg13g2_decap_8 FILLER_70_2560 ();
 sg13g2_decap_8 FILLER_70_2567 ();
 sg13g2_decap_8 FILLER_70_2574 ();
 sg13g2_decap_8 FILLER_70_2581 ();
 sg13g2_decap_8 FILLER_70_2588 ();
 sg13g2_decap_8 FILLER_70_2595 ();
 sg13g2_decap_8 FILLER_70_2602 ();
 sg13g2_decap_8 FILLER_70_2609 ();
 sg13g2_decap_8 FILLER_70_2616 ();
 sg13g2_decap_8 FILLER_70_2623 ();
 sg13g2_decap_8 FILLER_70_2630 ();
 sg13g2_decap_8 FILLER_70_2637 ();
 sg13g2_decap_8 FILLER_70_2644 ();
 sg13g2_decap_8 FILLER_70_2651 ();
 sg13g2_decap_8 FILLER_70_2658 ();
 sg13g2_decap_4 FILLER_70_2665 ();
 sg13g2_fill_1 FILLER_70_2669 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_112 ();
 sg13g2_decap_8 FILLER_71_119 ();
 sg13g2_decap_8 FILLER_71_126 ();
 sg13g2_decap_8 FILLER_71_133 ();
 sg13g2_decap_8 FILLER_71_140 ();
 sg13g2_decap_8 FILLER_71_147 ();
 sg13g2_decap_4 FILLER_71_154 ();
 sg13g2_decap_8 FILLER_71_162 ();
 sg13g2_decap_8 FILLER_71_169 ();
 sg13g2_decap_8 FILLER_71_176 ();
 sg13g2_decap_8 FILLER_71_183 ();
 sg13g2_decap_8 FILLER_71_190 ();
 sg13g2_decap_8 FILLER_71_197 ();
 sg13g2_decap_8 FILLER_71_204 ();
 sg13g2_decap_8 FILLER_71_211 ();
 sg13g2_decap_8 FILLER_71_218 ();
 sg13g2_decap_8 FILLER_71_225 ();
 sg13g2_decap_8 FILLER_71_232 ();
 sg13g2_decap_8 FILLER_71_239 ();
 sg13g2_decap_8 FILLER_71_246 ();
 sg13g2_decap_8 FILLER_71_253 ();
 sg13g2_decap_8 FILLER_71_260 ();
 sg13g2_decap_8 FILLER_71_267 ();
 sg13g2_decap_8 FILLER_71_274 ();
 sg13g2_decap_8 FILLER_71_281 ();
 sg13g2_decap_8 FILLER_71_288 ();
 sg13g2_decap_8 FILLER_71_295 ();
 sg13g2_decap_8 FILLER_71_302 ();
 sg13g2_decap_8 FILLER_71_309 ();
 sg13g2_decap_8 FILLER_71_316 ();
 sg13g2_decap_8 FILLER_71_323 ();
 sg13g2_decap_8 FILLER_71_330 ();
 sg13g2_decap_8 FILLER_71_347 ();
 sg13g2_decap_8 FILLER_71_354 ();
 sg13g2_decap_8 FILLER_71_361 ();
 sg13g2_decap_8 FILLER_71_368 ();
 sg13g2_decap_8 FILLER_71_375 ();
 sg13g2_decap_8 FILLER_71_382 ();
 sg13g2_fill_2 FILLER_71_389 ();
 sg13g2_fill_1 FILLER_71_391 ();
 sg13g2_decap_4 FILLER_71_407 ();
 sg13g2_fill_2 FILLER_71_411 ();
 sg13g2_fill_2 FILLER_71_417 ();
 sg13g2_fill_1 FILLER_71_419 ();
 sg13g2_decap_8 FILLER_71_425 ();
 sg13g2_decap_4 FILLER_71_432 ();
 sg13g2_decap_8 FILLER_71_440 ();
 sg13g2_decap_8 FILLER_71_447 ();
 sg13g2_decap_8 FILLER_71_454 ();
 sg13g2_decap_8 FILLER_71_461 ();
 sg13g2_decap_8 FILLER_71_468 ();
 sg13g2_decap_8 FILLER_71_475 ();
 sg13g2_decap_8 FILLER_71_482 ();
 sg13g2_decap_4 FILLER_71_489 ();
 sg13g2_fill_1 FILLER_71_493 ();
 sg13g2_decap_8 FILLER_71_498 ();
 sg13g2_decap_4 FILLER_71_505 ();
 sg13g2_fill_2 FILLER_71_509 ();
 sg13g2_decap_8 FILLER_71_514 ();
 sg13g2_fill_2 FILLER_71_521 ();
 sg13g2_decap_8 FILLER_71_528 ();
 sg13g2_decap_8 FILLER_71_535 ();
 sg13g2_decap_8 FILLER_71_542 ();
 sg13g2_decap_4 FILLER_71_549 ();
 sg13g2_fill_2 FILLER_71_553 ();
 sg13g2_decap_8 FILLER_71_564 ();
 sg13g2_decap_8 FILLER_71_571 ();
 sg13g2_decap_8 FILLER_71_578 ();
 sg13g2_decap_8 FILLER_71_585 ();
 sg13g2_decap_8 FILLER_71_592 ();
 sg13g2_decap_8 FILLER_71_599 ();
 sg13g2_decap_8 FILLER_71_606 ();
 sg13g2_fill_2 FILLER_71_613 ();
 sg13g2_fill_1 FILLER_71_615 ();
 sg13g2_decap_4 FILLER_71_619 ();
 sg13g2_fill_1 FILLER_71_623 ();
 sg13g2_decap_4 FILLER_71_628 ();
 sg13g2_fill_1 FILLER_71_632 ();
 sg13g2_decap_8 FILLER_71_636 ();
 sg13g2_decap_8 FILLER_71_643 ();
 sg13g2_decap_8 FILLER_71_650 ();
 sg13g2_decap_8 FILLER_71_657 ();
 sg13g2_decap_8 FILLER_71_664 ();
 sg13g2_decap_8 FILLER_71_671 ();
 sg13g2_decap_8 FILLER_71_678 ();
 sg13g2_decap_8 FILLER_71_685 ();
 sg13g2_fill_2 FILLER_71_692 ();
 sg13g2_fill_1 FILLER_71_694 ();
 sg13g2_fill_2 FILLER_71_702 ();
 sg13g2_decap_8 FILLER_71_708 ();
 sg13g2_decap_8 FILLER_71_715 ();
 sg13g2_decap_4 FILLER_71_722 ();
 sg13g2_fill_1 FILLER_71_726 ();
 sg13g2_decap_8 FILLER_71_742 ();
 sg13g2_decap_8 FILLER_71_749 ();
 sg13g2_decap_8 FILLER_71_756 ();
 sg13g2_decap_8 FILLER_71_763 ();
 sg13g2_decap_4 FILLER_71_770 ();
 sg13g2_fill_1 FILLER_71_774 ();
 sg13g2_decap_8 FILLER_71_794 ();
 sg13g2_decap_8 FILLER_71_801 ();
 sg13g2_fill_2 FILLER_71_808 ();
 sg13g2_decap_8 FILLER_71_815 ();
 sg13g2_decap_8 FILLER_71_822 ();
 sg13g2_decap_8 FILLER_71_835 ();
 sg13g2_decap_8 FILLER_71_842 ();
 sg13g2_fill_2 FILLER_71_849 ();
 sg13g2_fill_1 FILLER_71_851 ();
 sg13g2_decap_8 FILLER_71_867 ();
 sg13g2_decap_8 FILLER_71_874 ();
 sg13g2_decap_8 FILLER_71_881 ();
 sg13g2_decap_4 FILLER_71_888 ();
 sg13g2_fill_2 FILLER_71_892 ();
 sg13g2_decap_8 FILLER_71_898 ();
 sg13g2_decap_8 FILLER_71_905 ();
 sg13g2_decap_8 FILLER_71_912 ();
 sg13g2_decap_8 FILLER_71_919 ();
 sg13g2_decap_4 FILLER_71_926 ();
 sg13g2_fill_2 FILLER_71_930 ();
 sg13g2_fill_2 FILLER_71_944 ();
 sg13g2_decap_8 FILLER_71_965 ();
 sg13g2_decap_4 FILLER_71_972 ();
 sg13g2_decap_8 FILLER_71_991 ();
 sg13g2_fill_1 FILLER_71_998 ();
 sg13g2_fill_1 FILLER_71_1005 ();
 sg13g2_decap_8 FILLER_71_1011 ();
 sg13g2_decap_8 FILLER_71_1018 ();
 sg13g2_decap_8 FILLER_71_1025 ();
 sg13g2_decap_8 FILLER_71_1032 ();
 sg13g2_decap_8 FILLER_71_1039 ();
 sg13g2_decap_8 FILLER_71_1046 ();
 sg13g2_decap_8 FILLER_71_1053 ();
 sg13g2_decap_8 FILLER_71_1060 ();
 sg13g2_decap_4 FILLER_71_1067 ();
 sg13g2_fill_1 FILLER_71_1071 ();
 sg13g2_decap_8 FILLER_71_1076 ();
 sg13g2_decap_8 FILLER_71_1083 ();
 sg13g2_decap_8 FILLER_71_1090 ();
 sg13g2_decap_4 FILLER_71_1097 ();
 sg13g2_fill_2 FILLER_71_1106 ();
 sg13g2_fill_1 FILLER_71_1108 ();
 sg13g2_decap_8 FILLER_71_1114 ();
 sg13g2_decap_8 FILLER_71_1121 ();
 sg13g2_decap_8 FILLER_71_1128 ();
 sg13g2_decap_8 FILLER_71_1135 ();
 sg13g2_decap_8 FILLER_71_1142 ();
 sg13g2_fill_1 FILLER_71_1149 ();
 sg13g2_decap_8 FILLER_71_1165 ();
 sg13g2_decap_8 FILLER_71_1172 ();
 sg13g2_decap_8 FILLER_71_1179 ();
 sg13g2_decap_8 FILLER_71_1186 ();
 sg13g2_decap_8 FILLER_71_1193 ();
 sg13g2_decap_8 FILLER_71_1200 ();
 sg13g2_decap_8 FILLER_71_1207 ();
 sg13g2_decap_8 FILLER_71_1214 ();
 sg13g2_decap_8 FILLER_71_1221 ();
 sg13g2_decap_4 FILLER_71_1228 ();
 sg13g2_fill_1 FILLER_71_1232 ();
 sg13g2_decap_8 FILLER_71_1246 ();
 sg13g2_decap_8 FILLER_71_1253 ();
 sg13g2_decap_8 FILLER_71_1260 ();
 sg13g2_decap_8 FILLER_71_1267 ();
 sg13g2_decap_8 FILLER_71_1274 ();
 sg13g2_fill_2 FILLER_71_1281 ();
 sg13g2_fill_1 FILLER_71_1283 ();
 sg13g2_decap_8 FILLER_71_1287 ();
 sg13g2_decap_4 FILLER_71_1294 ();
 sg13g2_fill_2 FILLER_71_1298 ();
 sg13g2_decap_8 FILLER_71_1306 ();
 sg13g2_fill_1 FILLER_71_1313 ();
 sg13g2_decap_8 FILLER_71_1317 ();
 sg13g2_decap_8 FILLER_71_1324 ();
 sg13g2_decap_8 FILLER_71_1331 ();
 sg13g2_decap_8 FILLER_71_1338 ();
 sg13g2_decap_8 FILLER_71_1345 ();
 sg13g2_fill_1 FILLER_71_1352 ();
 sg13g2_decap_8 FILLER_71_1356 ();
 sg13g2_decap_8 FILLER_71_1363 ();
 sg13g2_decap_8 FILLER_71_1370 ();
 sg13g2_decap_8 FILLER_71_1377 ();
 sg13g2_decap_8 FILLER_71_1384 ();
 sg13g2_fill_2 FILLER_71_1391 ();
 sg13g2_decap_8 FILLER_71_1397 ();
 sg13g2_decap_8 FILLER_71_1404 ();
 sg13g2_decap_8 FILLER_71_1411 ();
 sg13g2_decap_8 FILLER_71_1418 ();
 sg13g2_decap_8 FILLER_71_1425 ();
 sg13g2_decap_4 FILLER_71_1432 ();
 sg13g2_decap_8 FILLER_71_1440 ();
 sg13g2_decap_8 FILLER_71_1447 ();
 sg13g2_decap_8 FILLER_71_1454 ();
 sg13g2_decap_8 FILLER_71_1461 ();
 sg13g2_decap_8 FILLER_71_1468 ();
 sg13g2_decap_8 FILLER_71_1475 ();
 sg13g2_decap_8 FILLER_71_1482 ();
 sg13g2_decap_8 FILLER_71_1489 ();
 sg13g2_decap_8 FILLER_71_1496 ();
 sg13g2_decap_8 FILLER_71_1503 ();
 sg13g2_decap_8 FILLER_71_1510 ();
 sg13g2_fill_2 FILLER_71_1517 ();
 sg13g2_fill_1 FILLER_71_1519 ();
 sg13g2_decap_8 FILLER_71_1523 ();
 sg13g2_decap_8 FILLER_71_1530 ();
 sg13g2_decap_4 FILLER_71_1537 ();
 sg13g2_fill_2 FILLER_71_1541 ();
 sg13g2_decap_8 FILLER_71_1547 ();
 sg13g2_decap_8 FILLER_71_1554 ();
 sg13g2_decap_8 FILLER_71_1561 ();
 sg13g2_fill_2 FILLER_71_1568 ();
 sg13g2_fill_1 FILLER_71_1570 ();
 sg13g2_decap_8 FILLER_71_1586 ();
 sg13g2_decap_8 FILLER_71_1593 ();
 sg13g2_decap_8 FILLER_71_1600 ();
 sg13g2_fill_1 FILLER_71_1607 ();
 sg13g2_decap_8 FILLER_71_1623 ();
 sg13g2_decap_8 FILLER_71_1633 ();
 sg13g2_decap_8 FILLER_71_1640 ();
 sg13g2_decap_8 FILLER_71_1651 ();
 sg13g2_decap_4 FILLER_71_1658 ();
 sg13g2_fill_1 FILLER_71_1662 ();
 sg13g2_decap_8 FILLER_71_1666 ();
 sg13g2_decap_8 FILLER_71_1673 ();
 sg13g2_decap_8 FILLER_71_1680 ();
 sg13g2_decap_8 FILLER_71_1687 ();
 sg13g2_decap_4 FILLER_71_1694 ();
 sg13g2_fill_1 FILLER_71_1698 ();
 sg13g2_decap_8 FILLER_71_1702 ();
 sg13g2_decap_8 FILLER_71_1709 ();
 sg13g2_decap_8 FILLER_71_1716 ();
 sg13g2_decap_8 FILLER_71_1723 ();
 sg13g2_fill_2 FILLER_71_1730 ();
 sg13g2_fill_1 FILLER_71_1732 ();
 sg13g2_decap_8 FILLER_71_1736 ();
 sg13g2_decap_8 FILLER_71_1743 ();
 sg13g2_decap_8 FILLER_71_1750 ();
 sg13g2_decap_8 FILLER_71_1757 ();
 sg13g2_decap_8 FILLER_71_1764 ();
 sg13g2_decap_8 FILLER_71_1771 ();
 sg13g2_decap_8 FILLER_71_1778 ();
 sg13g2_decap_8 FILLER_71_1785 ();
 sg13g2_decap_8 FILLER_71_1792 ();
 sg13g2_decap_8 FILLER_71_1799 ();
 sg13g2_decap_8 FILLER_71_1806 ();
 sg13g2_decap_8 FILLER_71_1813 ();
 sg13g2_decap_8 FILLER_71_1820 ();
 sg13g2_decap_8 FILLER_71_1827 ();
 sg13g2_decap_4 FILLER_71_1834 ();
 sg13g2_decap_8 FILLER_71_1851 ();
 sg13g2_decap_8 FILLER_71_1858 ();
 sg13g2_decap_8 FILLER_71_1865 ();
 sg13g2_decap_8 FILLER_71_1872 ();
 sg13g2_decap_8 FILLER_71_1879 ();
 sg13g2_decap_8 FILLER_71_1886 ();
 sg13g2_decap_8 FILLER_71_1893 ();
 sg13g2_decap_8 FILLER_71_1900 ();
 sg13g2_decap_8 FILLER_71_1907 ();
 sg13g2_decap_8 FILLER_71_1914 ();
 sg13g2_decap_8 FILLER_71_1921 ();
 sg13g2_decap_8 FILLER_71_1928 ();
 sg13g2_decap_8 FILLER_71_1935 ();
 sg13g2_decap_8 FILLER_71_1942 ();
 sg13g2_decap_8 FILLER_71_1949 ();
 sg13g2_decap_8 FILLER_71_1956 ();
 sg13g2_decap_8 FILLER_71_1963 ();
 sg13g2_decap_8 FILLER_71_1970 ();
 sg13g2_decap_8 FILLER_71_1977 ();
 sg13g2_decap_8 FILLER_71_1984 ();
 sg13g2_decap_8 FILLER_71_1991 ();
 sg13g2_decap_8 FILLER_71_1998 ();
 sg13g2_decap_8 FILLER_71_2005 ();
 sg13g2_decap_8 FILLER_71_2012 ();
 sg13g2_decap_4 FILLER_71_2019 ();
 sg13g2_fill_2 FILLER_71_2023 ();
 sg13g2_decap_8 FILLER_71_2030 ();
 sg13g2_decap_8 FILLER_71_2037 ();
 sg13g2_decap_8 FILLER_71_2044 ();
 sg13g2_decap_4 FILLER_71_2051 ();
 sg13g2_fill_2 FILLER_71_2055 ();
 sg13g2_decap_8 FILLER_71_2065 ();
 sg13g2_decap_8 FILLER_71_2072 ();
 sg13g2_decap_8 FILLER_71_2079 ();
 sg13g2_decap_8 FILLER_71_2086 ();
 sg13g2_decap_4 FILLER_71_2093 ();
 sg13g2_fill_1 FILLER_71_2097 ();
 sg13g2_decap_8 FILLER_71_2101 ();
 sg13g2_decap_8 FILLER_71_2108 ();
 sg13g2_decap_8 FILLER_71_2115 ();
 sg13g2_decap_8 FILLER_71_2122 ();
 sg13g2_decap_8 FILLER_71_2129 ();
 sg13g2_decap_8 FILLER_71_2136 ();
 sg13g2_fill_2 FILLER_71_2143 ();
 sg13g2_fill_1 FILLER_71_2145 ();
 sg13g2_decap_8 FILLER_71_2149 ();
 sg13g2_decap_8 FILLER_71_2156 ();
 sg13g2_decap_8 FILLER_71_2163 ();
 sg13g2_decap_8 FILLER_71_2170 ();
 sg13g2_decap_8 FILLER_71_2177 ();
 sg13g2_decap_8 FILLER_71_2184 ();
 sg13g2_decap_8 FILLER_71_2191 ();
 sg13g2_decap_8 FILLER_71_2198 ();
 sg13g2_decap_8 FILLER_71_2205 ();
 sg13g2_fill_1 FILLER_71_2212 ();
 sg13g2_decap_8 FILLER_71_2217 ();
 sg13g2_decap_8 FILLER_71_2224 ();
 sg13g2_decap_8 FILLER_71_2231 ();
 sg13g2_decap_8 FILLER_71_2238 ();
 sg13g2_decap_8 FILLER_71_2245 ();
 sg13g2_decap_8 FILLER_71_2252 ();
 sg13g2_decap_8 FILLER_71_2259 ();
 sg13g2_decap_8 FILLER_71_2266 ();
 sg13g2_decap_8 FILLER_71_2273 ();
 sg13g2_decap_8 FILLER_71_2280 ();
 sg13g2_decap_8 FILLER_71_2287 ();
 sg13g2_decap_8 FILLER_71_2294 ();
 sg13g2_decap_8 FILLER_71_2301 ();
 sg13g2_decap_8 FILLER_71_2308 ();
 sg13g2_decap_8 FILLER_71_2315 ();
 sg13g2_decap_8 FILLER_71_2322 ();
 sg13g2_decap_8 FILLER_71_2329 ();
 sg13g2_decap_8 FILLER_71_2336 ();
 sg13g2_decap_8 FILLER_71_2343 ();
 sg13g2_decap_8 FILLER_71_2350 ();
 sg13g2_decap_8 FILLER_71_2357 ();
 sg13g2_decap_8 FILLER_71_2364 ();
 sg13g2_decap_8 FILLER_71_2371 ();
 sg13g2_decap_8 FILLER_71_2378 ();
 sg13g2_decap_8 FILLER_71_2385 ();
 sg13g2_decap_8 FILLER_71_2392 ();
 sg13g2_decap_8 FILLER_71_2399 ();
 sg13g2_decap_8 FILLER_71_2406 ();
 sg13g2_decap_8 FILLER_71_2413 ();
 sg13g2_decap_8 FILLER_71_2420 ();
 sg13g2_decap_8 FILLER_71_2427 ();
 sg13g2_decap_8 FILLER_71_2434 ();
 sg13g2_decap_8 FILLER_71_2441 ();
 sg13g2_decap_8 FILLER_71_2448 ();
 sg13g2_decap_8 FILLER_71_2455 ();
 sg13g2_decap_8 FILLER_71_2462 ();
 sg13g2_decap_8 FILLER_71_2469 ();
 sg13g2_decap_8 FILLER_71_2476 ();
 sg13g2_decap_8 FILLER_71_2483 ();
 sg13g2_decap_8 FILLER_71_2490 ();
 sg13g2_decap_8 FILLER_71_2497 ();
 sg13g2_decap_8 FILLER_71_2504 ();
 sg13g2_decap_8 FILLER_71_2511 ();
 sg13g2_decap_8 FILLER_71_2518 ();
 sg13g2_decap_8 FILLER_71_2525 ();
 sg13g2_decap_8 FILLER_71_2532 ();
 sg13g2_decap_8 FILLER_71_2539 ();
 sg13g2_decap_8 FILLER_71_2546 ();
 sg13g2_decap_8 FILLER_71_2553 ();
 sg13g2_decap_8 FILLER_71_2560 ();
 sg13g2_decap_8 FILLER_71_2567 ();
 sg13g2_decap_8 FILLER_71_2574 ();
 sg13g2_decap_8 FILLER_71_2581 ();
 sg13g2_decap_8 FILLER_71_2588 ();
 sg13g2_decap_8 FILLER_71_2595 ();
 sg13g2_decap_8 FILLER_71_2602 ();
 sg13g2_decap_8 FILLER_71_2609 ();
 sg13g2_decap_8 FILLER_71_2616 ();
 sg13g2_decap_8 FILLER_71_2623 ();
 sg13g2_decap_8 FILLER_71_2630 ();
 sg13g2_decap_8 FILLER_71_2637 ();
 sg13g2_decap_8 FILLER_71_2644 ();
 sg13g2_decap_8 FILLER_71_2651 ();
 sg13g2_decap_8 FILLER_71_2658 ();
 sg13g2_decap_4 FILLER_71_2665 ();
 sg13g2_fill_1 FILLER_71_2669 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_fill_1 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_83 ();
 sg13g2_decap_8 FILLER_72_90 ();
 sg13g2_decap_8 FILLER_72_97 ();
 sg13g2_decap_4 FILLER_72_104 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_119 ();
 sg13g2_decap_8 FILLER_72_126 ();
 sg13g2_decap_8 FILLER_72_133 ();
 sg13g2_decap_8 FILLER_72_140 ();
 sg13g2_decap_4 FILLER_72_147 ();
 sg13g2_fill_1 FILLER_72_151 ();
 sg13g2_decap_8 FILLER_72_178 ();
 sg13g2_decap_8 FILLER_72_185 ();
 sg13g2_fill_2 FILLER_72_192 ();
 sg13g2_fill_1 FILLER_72_194 ();
 sg13g2_decap_4 FILLER_72_198 ();
 sg13g2_decap_8 FILLER_72_206 ();
 sg13g2_decap_8 FILLER_72_213 ();
 sg13g2_decap_8 FILLER_72_220 ();
 sg13g2_decap_8 FILLER_72_227 ();
 sg13g2_decap_4 FILLER_72_234 ();
 sg13g2_fill_1 FILLER_72_238 ();
 sg13g2_decap_8 FILLER_72_254 ();
 sg13g2_decap_8 FILLER_72_261 ();
 sg13g2_decap_8 FILLER_72_268 ();
 sg13g2_decap_8 FILLER_72_275 ();
 sg13g2_fill_1 FILLER_72_282 ();
 sg13g2_fill_1 FILLER_72_298 ();
 sg13g2_decap_8 FILLER_72_303 ();
 sg13g2_decap_8 FILLER_72_310 ();
 sg13g2_decap_8 FILLER_72_317 ();
 sg13g2_decap_8 FILLER_72_324 ();
 sg13g2_decap_8 FILLER_72_331 ();
 sg13g2_decap_8 FILLER_72_338 ();
 sg13g2_decap_8 FILLER_72_345 ();
 sg13g2_decap_8 FILLER_72_352 ();
 sg13g2_decap_8 FILLER_72_359 ();
 sg13g2_decap_8 FILLER_72_366 ();
 sg13g2_fill_1 FILLER_72_373 ();
 sg13g2_decap_8 FILLER_72_377 ();
 sg13g2_decap_8 FILLER_72_384 ();
 sg13g2_decap_4 FILLER_72_391 ();
 sg13g2_decap_8 FILLER_72_402 ();
 sg13g2_decap_8 FILLER_72_409 ();
 sg13g2_decap_8 FILLER_72_416 ();
 sg13g2_decap_8 FILLER_72_423 ();
 sg13g2_decap_8 FILLER_72_430 ();
 sg13g2_fill_2 FILLER_72_437 ();
 sg13g2_fill_1 FILLER_72_439 ();
 sg13g2_decap_8 FILLER_72_444 ();
 sg13g2_decap_8 FILLER_72_451 ();
 sg13g2_decap_8 FILLER_72_458 ();
 sg13g2_decap_8 FILLER_72_465 ();
 sg13g2_decap_8 FILLER_72_472 ();
 sg13g2_decap_8 FILLER_72_479 ();
 sg13g2_fill_1 FILLER_72_486 ();
 sg13g2_decap_8 FILLER_72_502 ();
 sg13g2_decap_8 FILLER_72_509 ();
 sg13g2_decap_8 FILLER_72_516 ();
 sg13g2_decap_8 FILLER_72_523 ();
 sg13g2_fill_1 FILLER_72_530 ();
 sg13g2_decap_8 FILLER_72_536 ();
 sg13g2_decap_8 FILLER_72_543 ();
 sg13g2_decap_8 FILLER_72_550 ();
 sg13g2_fill_2 FILLER_72_557 ();
 sg13g2_decap_8 FILLER_72_564 ();
 sg13g2_decap_8 FILLER_72_571 ();
 sg13g2_decap_8 FILLER_72_578 ();
 sg13g2_decap_8 FILLER_72_585 ();
 sg13g2_decap_8 FILLER_72_592 ();
 sg13g2_fill_2 FILLER_72_599 ();
 sg13g2_fill_1 FILLER_72_601 ();
 sg13g2_fill_1 FILLER_72_612 ();
 sg13g2_fill_1 FILLER_72_622 ();
 sg13g2_decap_8 FILLER_72_641 ();
 sg13g2_decap_8 FILLER_72_648 ();
 sg13g2_decap_8 FILLER_72_655 ();
 sg13g2_fill_1 FILLER_72_662 ();
 sg13g2_fill_2 FILLER_72_669 ();
 sg13g2_fill_1 FILLER_72_671 ();
 sg13g2_decap_8 FILLER_72_676 ();
 sg13g2_fill_2 FILLER_72_683 ();
 sg13g2_fill_1 FILLER_72_685 ();
 sg13g2_decap_4 FILLER_72_689 ();
 sg13g2_fill_2 FILLER_72_693 ();
 sg13g2_fill_2 FILLER_72_700 ();
 sg13g2_fill_1 FILLER_72_702 ();
 sg13g2_decap_8 FILLER_72_709 ();
 sg13g2_decap_4 FILLER_72_716 ();
 sg13g2_decap_8 FILLER_72_738 ();
 sg13g2_decap_8 FILLER_72_745 ();
 sg13g2_decap_8 FILLER_72_752 ();
 sg13g2_decap_8 FILLER_72_759 ();
 sg13g2_decap_8 FILLER_72_766 ();
 sg13g2_decap_4 FILLER_72_773 ();
 sg13g2_decap_8 FILLER_72_786 ();
 sg13g2_decap_8 FILLER_72_793 ();
 sg13g2_decap_8 FILLER_72_800 ();
 sg13g2_fill_2 FILLER_72_807 ();
 sg13g2_fill_1 FILLER_72_809 ();
 sg13g2_decap_4 FILLER_72_816 ();
 sg13g2_fill_1 FILLER_72_820 ();
 sg13g2_fill_1 FILLER_72_828 ();
 sg13g2_decap_8 FILLER_72_839 ();
 sg13g2_decap_8 FILLER_72_846 ();
 sg13g2_fill_2 FILLER_72_853 ();
 sg13g2_decap_8 FILLER_72_860 ();
 sg13g2_decap_8 FILLER_72_867 ();
 sg13g2_decap_8 FILLER_72_874 ();
 sg13g2_decap_8 FILLER_72_881 ();
 sg13g2_fill_2 FILLER_72_888 ();
 sg13g2_decap_8 FILLER_72_895 ();
 sg13g2_decap_8 FILLER_72_902 ();
 sg13g2_decap_8 FILLER_72_909 ();
 sg13g2_decap_8 FILLER_72_916 ();
 sg13g2_decap_4 FILLER_72_923 ();
 sg13g2_fill_2 FILLER_72_927 ();
 sg13g2_decap_8 FILLER_72_933 ();
 sg13g2_fill_1 FILLER_72_940 ();
 sg13g2_fill_1 FILLER_72_945 ();
 sg13g2_fill_2 FILLER_72_962 ();
 sg13g2_decap_8 FILLER_72_990 ();
 sg13g2_decap_8 FILLER_72_997 ();
 sg13g2_fill_2 FILLER_72_1004 ();
 sg13g2_fill_1 FILLER_72_1009 ();
 sg13g2_decap_8 FILLER_72_1015 ();
 sg13g2_decap_8 FILLER_72_1022 ();
 sg13g2_decap_4 FILLER_72_1039 ();
 sg13g2_decap_8 FILLER_72_1048 ();
 sg13g2_decap_8 FILLER_72_1055 ();
 sg13g2_decap_8 FILLER_72_1062 ();
 sg13g2_fill_2 FILLER_72_1069 ();
 sg13g2_fill_1 FILLER_72_1071 ();
 sg13g2_decap_8 FILLER_72_1084 ();
 sg13g2_decap_8 FILLER_72_1091 ();
 sg13g2_decap_4 FILLER_72_1103 ();
 sg13g2_fill_2 FILLER_72_1107 ();
 sg13g2_decap_8 FILLER_72_1113 ();
 sg13g2_decap_8 FILLER_72_1120 ();
 sg13g2_decap_8 FILLER_72_1127 ();
 sg13g2_fill_1 FILLER_72_1134 ();
 sg13g2_decap_8 FILLER_72_1150 ();
 sg13g2_decap_8 FILLER_72_1157 ();
 sg13g2_fill_2 FILLER_72_1169 ();
 sg13g2_fill_1 FILLER_72_1171 ();
 sg13g2_decap_8 FILLER_72_1176 ();
 sg13g2_decap_8 FILLER_72_1187 ();
 sg13g2_fill_2 FILLER_72_1194 ();
 sg13g2_decap_8 FILLER_72_1227 ();
 sg13g2_decap_8 FILLER_72_1238 ();
 sg13g2_decap_8 FILLER_72_1245 ();
 sg13g2_decap_8 FILLER_72_1252 ();
 sg13g2_decap_8 FILLER_72_1259 ();
 sg13g2_decap_8 FILLER_72_1266 ();
 sg13g2_decap_8 FILLER_72_1273 ();
 sg13g2_decap_8 FILLER_72_1280 ();
 sg13g2_decap_8 FILLER_72_1287 ();
 sg13g2_decap_8 FILLER_72_1294 ();
 sg13g2_decap_8 FILLER_72_1301 ();
 sg13g2_decap_8 FILLER_72_1308 ();
 sg13g2_fill_1 FILLER_72_1315 ();
 sg13g2_decap_8 FILLER_72_1320 ();
 sg13g2_decap_8 FILLER_72_1327 ();
 sg13g2_decap_8 FILLER_72_1334 ();
 sg13g2_decap_8 FILLER_72_1341 ();
 sg13g2_fill_1 FILLER_72_1352 ();
 sg13g2_decap_8 FILLER_72_1358 ();
 sg13g2_decap_8 FILLER_72_1365 ();
 sg13g2_decap_8 FILLER_72_1372 ();
 sg13g2_decap_4 FILLER_72_1379 ();
 sg13g2_fill_2 FILLER_72_1391 ();
 sg13g2_decap_4 FILLER_72_1428 ();
 sg13g2_fill_1 FILLER_72_1432 ();
 sg13g2_decap_8 FILLER_72_1448 ();
 sg13g2_decap_4 FILLER_72_1455 ();
 sg13g2_fill_2 FILLER_72_1459 ();
 sg13g2_decap_8 FILLER_72_1467 ();
 sg13g2_decap_8 FILLER_72_1474 ();
 sg13g2_decap_8 FILLER_72_1481 ();
 sg13g2_decap_8 FILLER_72_1488 ();
 sg13g2_decap_8 FILLER_72_1495 ();
 sg13g2_decap_8 FILLER_72_1502 ();
 sg13g2_decap_8 FILLER_72_1509 ();
 sg13g2_decap_8 FILLER_72_1516 ();
 sg13g2_decap_8 FILLER_72_1523 ();
 sg13g2_decap_4 FILLER_72_1530 ();
 sg13g2_decap_8 FILLER_72_1539 ();
 sg13g2_decap_8 FILLER_72_1546 ();
 sg13g2_decap_8 FILLER_72_1553 ();
 sg13g2_fill_2 FILLER_72_1560 ();
 sg13g2_decap_4 FILLER_72_1566 ();
 sg13g2_fill_1 FILLER_72_1570 ();
 sg13g2_decap_8 FILLER_72_1575 ();
 sg13g2_decap_8 FILLER_72_1582 ();
 sg13g2_decap_8 FILLER_72_1589 ();
 sg13g2_decap_8 FILLER_72_1596 ();
 sg13g2_fill_2 FILLER_72_1603 ();
 sg13g2_fill_1 FILLER_72_1624 ();
 sg13g2_decap_4 FILLER_72_1649 ();
 sg13g2_fill_1 FILLER_72_1653 ();
 sg13g2_decap_8 FILLER_72_1674 ();
 sg13g2_decap_8 FILLER_72_1681 ();
 sg13g2_decap_8 FILLER_72_1688 ();
 sg13g2_fill_1 FILLER_72_1695 ();
 sg13g2_decap_8 FILLER_72_1708 ();
 sg13g2_decap_8 FILLER_72_1715 ();
 sg13g2_decap_8 FILLER_72_1722 ();
 sg13g2_fill_1 FILLER_72_1729 ();
 sg13g2_decap_8 FILLER_72_1746 ();
 sg13g2_decap_8 FILLER_72_1753 ();
 sg13g2_decap_8 FILLER_72_1760 ();
 sg13g2_decap_8 FILLER_72_1767 ();
 sg13g2_decap_8 FILLER_72_1774 ();
 sg13g2_decap_8 FILLER_72_1781 ();
 sg13g2_decap_8 FILLER_72_1788 ();
 sg13g2_decap_8 FILLER_72_1795 ();
 sg13g2_decap_8 FILLER_72_1802 ();
 sg13g2_decap_8 FILLER_72_1809 ();
 sg13g2_decap_8 FILLER_72_1816 ();
 sg13g2_decap_8 FILLER_72_1823 ();
 sg13g2_decap_8 FILLER_72_1830 ();
 sg13g2_decap_8 FILLER_72_1837 ();
 sg13g2_decap_8 FILLER_72_1844 ();
 sg13g2_decap_8 FILLER_72_1851 ();
 sg13g2_decap_8 FILLER_72_1858 ();
 sg13g2_decap_8 FILLER_72_1865 ();
 sg13g2_decap_8 FILLER_72_1872 ();
 sg13g2_decap_8 FILLER_72_1879 ();
 sg13g2_decap_8 FILLER_72_1886 ();
 sg13g2_decap_8 FILLER_72_1893 ();
 sg13g2_decap_8 FILLER_72_1900 ();
 sg13g2_decap_8 FILLER_72_1907 ();
 sg13g2_decap_8 FILLER_72_1914 ();
 sg13g2_decap_8 FILLER_72_1921 ();
 sg13g2_decap_8 FILLER_72_1928 ();
 sg13g2_decap_8 FILLER_72_1935 ();
 sg13g2_decap_8 FILLER_72_1942 ();
 sg13g2_decap_8 FILLER_72_1949 ();
 sg13g2_decap_8 FILLER_72_1956 ();
 sg13g2_decap_8 FILLER_72_1963 ();
 sg13g2_decap_8 FILLER_72_1970 ();
 sg13g2_decap_8 FILLER_72_1977 ();
 sg13g2_decap_8 FILLER_72_2010 ();
 sg13g2_decap_8 FILLER_72_2017 ();
 sg13g2_fill_1 FILLER_72_2024 ();
 sg13g2_decap_8 FILLER_72_2029 ();
 sg13g2_decap_8 FILLER_72_2036 ();
 sg13g2_decap_8 FILLER_72_2043 ();
 sg13g2_decap_8 FILLER_72_2050 ();
 sg13g2_decap_8 FILLER_72_2057 ();
 sg13g2_decap_8 FILLER_72_2064 ();
 sg13g2_decap_8 FILLER_72_2071 ();
 sg13g2_decap_4 FILLER_72_2078 ();
 sg13g2_fill_1 FILLER_72_2082 ();
 sg13g2_decap_8 FILLER_72_2091 ();
 sg13g2_decap_8 FILLER_72_2098 ();
 sg13g2_decap_8 FILLER_72_2105 ();
 sg13g2_decap_4 FILLER_72_2112 ();
 sg13g2_fill_1 FILLER_72_2116 ();
 sg13g2_decap_8 FILLER_72_2125 ();
 sg13g2_decap_8 FILLER_72_2132 ();
 sg13g2_decap_8 FILLER_72_2139 ();
 sg13g2_decap_8 FILLER_72_2146 ();
 sg13g2_decap_8 FILLER_72_2153 ();
 sg13g2_decap_8 FILLER_72_2160 ();
 sg13g2_decap_8 FILLER_72_2167 ();
 sg13g2_decap_8 FILLER_72_2174 ();
 sg13g2_decap_8 FILLER_72_2181 ();
 sg13g2_decap_8 FILLER_72_2188 ();
 sg13g2_decap_8 FILLER_72_2195 ();
 sg13g2_decap_8 FILLER_72_2202 ();
 sg13g2_decap_8 FILLER_72_2209 ();
 sg13g2_decap_8 FILLER_72_2216 ();
 sg13g2_decap_8 FILLER_72_2223 ();
 sg13g2_decap_8 FILLER_72_2230 ();
 sg13g2_decap_8 FILLER_72_2237 ();
 sg13g2_decap_8 FILLER_72_2244 ();
 sg13g2_decap_8 FILLER_72_2251 ();
 sg13g2_decap_8 FILLER_72_2258 ();
 sg13g2_decap_8 FILLER_72_2265 ();
 sg13g2_decap_8 FILLER_72_2272 ();
 sg13g2_decap_8 FILLER_72_2279 ();
 sg13g2_decap_8 FILLER_72_2286 ();
 sg13g2_decap_8 FILLER_72_2293 ();
 sg13g2_decap_8 FILLER_72_2300 ();
 sg13g2_decap_8 FILLER_72_2307 ();
 sg13g2_decap_8 FILLER_72_2314 ();
 sg13g2_decap_8 FILLER_72_2321 ();
 sg13g2_decap_8 FILLER_72_2328 ();
 sg13g2_decap_8 FILLER_72_2335 ();
 sg13g2_decap_8 FILLER_72_2342 ();
 sg13g2_decap_8 FILLER_72_2349 ();
 sg13g2_decap_8 FILLER_72_2356 ();
 sg13g2_decap_8 FILLER_72_2363 ();
 sg13g2_decap_8 FILLER_72_2370 ();
 sg13g2_decap_8 FILLER_72_2377 ();
 sg13g2_decap_8 FILLER_72_2384 ();
 sg13g2_decap_8 FILLER_72_2391 ();
 sg13g2_decap_8 FILLER_72_2398 ();
 sg13g2_decap_8 FILLER_72_2405 ();
 sg13g2_decap_8 FILLER_72_2412 ();
 sg13g2_decap_8 FILLER_72_2419 ();
 sg13g2_decap_8 FILLER_72_2426 ();
 sg13g2_decap_8 FILLER_72_2433 ();
 sg13g2_decap_8 FILLER_72_2440 ();
 sg13g2_decap_8 FILLER_72_2447 ();
 sg13g2_decap_8 FILLER_72_2454 ();
 sg13g2_decap_8 FILLER_72_2461 ();
 sg13g2_decap_8 FILLER_72_2468 ();
 sg13g2_decap_8 FILLER_72_2475 ();
 sg13g2_decap_8 FILLER_72_2482 ();
 sg13g2_decap_8 FILLER_72_2489 ();
 sg13g2_decap_8 FILLER_72_2496 ();
 sg13g2_decap_8 FILLER_72_2503 ();
 sg13g2_decap_8 FILLER_72_2510 ();
 sg13g2_decap_8 FILLER_72_2517 ();
 sg13g2_decap_8 FILLER_72_2524 ();
 sg13g2_decap_8 FILLER_72_2531 ();
 sg13g2_decap_8 FILLER_72_2538 ();
 sg13g2_decap_8 FILLER_72_2545 ();
 sg13g2_decap_8 FILLER_72_2552 ();
 sg13g2_decap_8 FILLER_72_2559 ();
 sg13g2_decap_8 FILLER_72_2566 ();
 sg13g2_decap_8 FILLER_72_2573 ();
 sg13g2_decap_8 FILLER_72_2580 ();
 sg13g2_decap_8 FILLER_72_2587 ();
 sg13g2_decap_8 FILLER_72_2594 ();
 sg13g2_decap_8 FILLER_72_2601 ();
 sg13g2_decap_8 FILLER_72_2608 ();
 sg13g2_decap_8 FILLER_72_2615 ();
 sg13g2_decap_8 FILLER_72_2622 ();
 sg13g2_decap_8 FILLER_72_2629 ();
 sg13g2_decap_8 FILLER_72_2636 ();
 sg13g2_decap_8 FILLER_72_2643 ();
 sg13g2_decap_8 FILLER_72_2650 ();
 sg13g2_decap_8 FILLER_72_2657 ();
 sg13g2_decap_4 FILLER_72_2664 ();
 sg13g2_fill_2 FILLER_72_2668 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_fill_2 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_69 ();
 sg13g2_decap_8 FILLER_73_76 ();
 sg13g2_decap_8 FILLER_73_83 ();
 sg13g2_decap_8 FILLER_73_90 ();
 sg13g2_decap_4 FILLER_73_97 ();
 sg13g2_fill_1 FILLER_73_101 ();
 sg13g2_decap_8 FILLER_73_128 ();
 sg13g2_decap_8 FILLER_73_135 ();
 sg13g2_decap_8 FILLER_73_142 ();
 sg13g2_decap_8 FILLER_73_149 ();
 sg13g2_decap_8 FILLER_73_156 ();
 sg13g2_decap_8 FILLER_73_163 ();
 sg13g2_decap_8 FILLER_73_170 ();
 sg13g2_decap_8 FILLER_73_177 ();
 sg13g2_decap_8 FILLER_73_184 ();
 sg13g2_fill_1 FILLER_73_191 ();
 sg13g2_decap_8 FILLER_73_221 ();
 sg13g2_decap_8 FILLER_73_228 ();
 sg13g2_decap_8 FILLER_73_235 ();
 sg13g2_decap_8 FILLER_73_268 ();
 sg13g2_decap_8 FILLER_73_275 ();
 sg13g2_decap_8 FILLER_73_282 ();
 sg13g2_fill_2 FILLER_73_289 ();
 sg13g2_fill_1 FILLER_73_291 ();
 sg13g2_decap_8 FILLER_73_318 ();
 sg13g2_decap_8 FILLER_73_325 ();
 sg13g2_decap_8 FILLER_73_332 ();
 sg13g2_decap_8 FILLER_73_339 ();
 sg13g2_decap_8 FILLER_73_346 ();
 sg13g2_decap_8 FILLER_73_353 ();
 sg13g2_decap_8 FILLER_73_360 ();
 sg13g2_decap_8 FILLER_73_367 ();
 sg13g2_decap_8 FILLER_73_374 ();
 sg13g2_decap_8 FILLER_73_381 ();
 sg13g2_decap_8 FILLER_73_388 ();
 sg13g2_fill_2 FILLER_73_395 ();
 sg13g2_decap_4 FILLER_73_401 ();
 sg13g2_fill_1 FILLER_73_405 ();
 sg13g2_decap_8 FILLER_73_411 ();
 sg13g2_decap_8 FILLER_73_418 ();
 sg13g2_fill_2 FILLER_73_425 ();
 sg13g2_fill_1 FILLER_73_427 ();
 sg13g2_decap_8 FILLER_73_433 ();
 sg13g2_decap_8 FILLER_73_440 ();
 sg13g2_decap_4 FILLER_73_447 ();
 sg13g2_decap_8 FILLER_73_466 ();
 sg13g2_decap_8 FILLER_73_473 ();
 sg13g2_decap_8 FILLER_73_480 ();
 sg13g2_fill_2 FILLER_73_487 ();
 sg13g2_fill_1 FILLER_73_489 ();
 sg13g2_decap_8 FILLER_73_495 ();
 sg13g2_decap_8 FILLER_73_502 ();
 sg13g2_decap_8 FILLER_73_509 ();
 sg13g2_decap_8 FILLER_73_520 ();
 sg13g2_decap_8 FILLER_73_527 ();
 sg13g2_decap_8 FILLER_73_534 ();
 sg13g2_decap_8 FILLER_73_541 ();
 sg13g2_decap_8 FILLER_73_548 ();
 sg13g2_decap_8 FILLER_73_555 ();
 sg13g2_decap_4 FILLER_73_562 ();
 sg13g2_decap_8 FILLER_73_571 ();
 sg13g2_decap_8 FILLER_73_578 ();
 sg13g2_decap_8 FILLER_73_585 ();
 sg13g2_decap_8 FILLER_73_592 ();
 sg13g2_decap_8 FILLER_73_599 ();
 sg13g2_decap_8 FILLER_73_606 ();
 sg13g2_decap_4 FILLER_73_613 ();
 sg13g2_fill_2 FILLER_73_617 ();
 sg13g2_decap_8 FILLER_73_633 ();
 sg13g2_decap_8 FILLER_73_640 ();
 sg13g2_decap_8 FILLER_73_647 ();
 sg13g2_decap_8 FILLER_73_654 ();
 sg13g2_fill_2 FILLER_73_661 ();
 sg13g2_decap_8 FILLER_73_667 ();
 sg13g2_decap_8 FILLER_73_674 ();
 sg13g2_fill_2 FILLER_73_681 ();
 sg13g2_decap_8 FILLER_73_691 ();
 sg13g2_decap_4 FILLER_73_698 ();
 sg13g2_fill_1 FILLER_73_702 ();
 sg13g2_decap_8 FILLER_73_708 ();
 sg13g2_decap_8 FILLER_73_715 ();
 sg13g2_decap_8 FILLER_73_722 ();
 sg13g2_decap_8 FILLER_73_729 ();
 sg13g2_decap_8 FILLER_73_736 ();
 sg13g2_decap_8 FILLER_73_743 ();
 sg13g2_decap_8 FILLER_73_750 ();
 sg13g2_decap_8 FILLER_73_757 ();
 sg13g2_decap_8 FILLER_73_764 ();
 sg13g2_decap_4 FILLER_73_771 ();
 sg13g2_decap_8 FILLER_73_780 ();
 sg13g2_decap_8 FILLER_73_787 ();
 sg13g2_decap_8 FILLER_73_794 ();
 sg13g2_decap_8 FILLER_73_801 ();
 sg13g2_decap_8 FILLER_73_808 ();
 sg13g2_decap_4 FILLER_73_815 ();
 sg13g2_fill_2 FILLER_73_819 ();
 sg13g2_fill_2 FILLER_73_826 ();
 sg13g2_fill_1 FILLER_73_828 ();
 sg13g2_decap_8 FILLER_73_834 ();
 sg13g2_decap_8 FILLER_73_841 ();
 sg13g2_decap_8 FILLER_73_848 ();
 sg13g2_decap_8 FILLER_73_865 ();
 sg13g2_decap_8 FILLER_73_872 ();
 sg13g2_decap_8 FILLER_73_879 ();
 sg13g2_decap_8 FILLER_73_886 ();
 sg13g2_decap_8 FILLER_73_893 ();
 sg13g2_decap_8 FILLER_73_900 ();
 sg13g2_decap_8 FILLER_73_907 ();
 sg13g2_fill_2 FILLER_73_914 ();
 sg13g2_fill_1 FILLER_73_916 ();
 sg13g2_decap_8 FILLER_73_929 ();
 sg13g2_decap_4 FILLER_73_936 ();
 sg13g2_fill_1 FILLER_73_940 ();
 sg13g2_fill_2 FILLER_73_944 ();
 sg13g2_decap_8 FILLER_73_949 ();
 sg13g2_decap_8 FILLER_73_956 ();
 sg13g2_decap_8 FILLER_73_963 ();
 sg13g2_decap_8 FILLER_73_970 ();
 sg13g2_decap_4 FILLER_73_977 ();
 sg13g2_fill_1 FILLER_73_981 ();
 sg13g2_decap_8 FILLER_73_986 ();
 sg13g2_decap_8 FILLER_73_993 ();
 sg13g2_decap_8 FILLER_73_1000 ();
 sg13g2_decap_8 FILLER_73_1007 ();
 sg13g2_decap_8 FILLER_73_1014 ();
 sg13g2_decap_8 FILLER_73_1021 ();
 sg13g2_decap_8 FILLER_73_1028 ();
 sg13g2_decap_8 FILLER_73_1035 ();
 sg13g2_decap_8 FILLER_73_1042 ();
 sg13g2_decap_8 FILLER_73_1049 ();
 sg13g2_decap_8 FILLER_73_1056 ();
 sg13g2_decap_8 FILLER_73_1063 ();
 sg13g2_fill_2 FILLER_73_1070 ();
 sg13g2_fill_1 FILLER_73_1072 ();
 sg13g2_decap_8 FILLER_73_1087 ();
 sg13g2_decap_8 FILLER_73_1094 ();
 sg13g2_decap_8 FILLER_73_1101 ();
 sg13g2_decap_8 FILLER_73_1108 ();
 sg13g2_decap_8 FILLER_73_1115 ();
 sg13g2_decap_8 FILLER_73_1122 ();
 sg13g2_decap_8 FILLER_73_1129 ();
 sg13g2_fill_2 FILLER_73_1136 ();
 sg13g2_decap_8 FILLER_73_1165 ();
 sg13g2_decap_8 FILLER_73_1172 ();
 sg13g2_decap_8 FILLER_73_1179 ();
 sg13g2_decap_4 FILLER_73_1186 ();
 sg13g2_decap_4 FILLER_73_1212 ();
 sg13g2_fill_1 FILLER_73_1216 ();
 sg13g2_decap_8 FILLER_73_1222 ();
 sg13g2_decap_8 FILLER_73_1229 ();
 sg13g2_decap_8 FILLER_73_1236 ();
 sg13g2_decap_8 FILLER_73_1243 ();
 sg13g2_decap_8 FILLER_73_1250 ();
 sg13g2_decap_8 FILLER_73_1257 ();
 sg13g2_decap_4 FILLER_73_1264 ();
 sg13g2_fill_1 FILLER_73_1268 ();
 sg13g2_decap_8 FILLER_73_1273 ();
 sg13g2_decap_8 FILLER_73_1280 ();
 sg13g2_decap_8 FILLER_73_1287 ();
 sg13g2_decap_4 FILLER_73_1294 ();
 sg13g2_fill_1 FILLER_73_1298 ();
 sg13g2_decap_8 FILLER_73_1305 ();
 sg13g2_decap_4 FILLER_73_1312 ();
 sg13g2_fill_1 FILLER_73_1316 ();
 sg13g2_decap_8 FILLER_73_1321 ();
 sg13g2_decap_8 FILLER_73_1328 ();
 sg13g2_decap_8 FILLER_73_1335 ();
 sg13g2_decap_8 FILLER_73_1342 ();
 sg13g2_decap_8 FILLER_73_1349 ();
 sg13g2_fill_1 FILLER_73_1356 ();
 sg13g2_decap_8 FILLER_73_1365 ();
 sg13g2_decap_8 FILLER_73_1372 ();
 sg13g2_decap_8 FILLER_73_1379 ();
 sg13g2_decap_8 FILLER_73_1386 ();
 sg13g2_decap_8 FILLER_73_1393 ();
 sg13g2_decap_8 FILLER_73_1400 ();
 sg13g2_decap_4 FILLER_73_1407 ();
 sg13g2_fill_2 FILLER_73_1411 ();
 sg13g2_decap_8 FILLER_73_1417 ();
 sg13g2_decap_8 FILLER_73_1424 ();
 sg13g2_fill_2 FILLER_73_1431 ();
 sg13g2_decap_8 FILLER_73_1437 ();
 sg13g2_decap_8 FILLER_73_1444 ();
 sg13g2_decap_8 FILLER_73_1451 ();
 sg13g2_decap_8 FILLER_73_1474 ();
 sg13g2_decap_8 FILLER_73_1481 ();
 sg13g2_decap_8 FILLER_73_1488 ();
 sg13g2_fill_2 FILLER_73_1495 ();
 sg13g2_fill_1 FILLER_73_1497 ();
 sg13g2_decap_8 FILLER_73_1505 ();
 sg13g2_decap_8 FILLER_73_1512 ();
 sg13g2_decap_8 FILLER_73_1519 ();
 sg13g2_decap_8 FILLER_73_1526 ();
 sg13g2_fill_2 FILLER_73_1533 ();
 sg13g2_fill_1 FILLER_73_1535 ();
 sg13g2_decap_8 FILLER_73_1541 ();
 sg13g2_decap_8 FILLER_73_1548 ();
 sg13g2_decap_8 FILLER_73_1555 ();
 sg13g2_fill_2 FILLER_73_1562 ();
 sg13g2_decap_8 FILLER_73_1569 ();
 sg13g2_decap_8 FILLER_73_1576 ();
 sg13g2_decap_8 FILLER_73_1583 ();
 sg13g2_decap_8 FILLER_73_1590 ();
 sg13g2_decap_8 FILLER_73_1597 ();
 sg13g2_decap_4 FILLER_73_1604 ();
 sg13g2_decap_8 FILLER_73_1614 ();
 sg13g2_decap_8 FILLER_73_1621 ();
 sg13g2_decap_8 FILLER_73_1636 ();
 sg13g2_decap_8 FILLER_73_1643 ();
 sg13g2_decap_8 FILLER_73_1650 ();
 sg13g2_decap_4 FILLER_73_1657 ();
 sg13g2_fill_2 FILLER_73_1661 ();
 sg13g2_decap_8 FILLER_73_1666 ();
 sg13g2_decap_8 FILLER_73_1673 ();
 sg13g2_decap_8 FILLER_73_1680 ();
 sg13g2_decap_8 FILLER_73_1687 ();
 sg13g2_decap_4 FILLER_73_1694 ();
 sg13g2_fill_1 FILLER_73_1698 ();
 sg13g2_decap_8 FILLER_73_1702 ();
 sg13g2_decap_8 FILLER_73_1709 ();
 sg13g2_decap_8 FILLER_73_1716 ();
 sg13g2_decap_8 FILLER_73_1723 ();
 sg13g2_decap_8 FILLER_73_1730 ();
 sg13g2_decap_8 FILLER_73_1737 ();
 sg13g2_decap_8 FILLER_73_1744 ();
 sg13g2_decap_8 FILLER_73_1751 ();
 sg13g2_decap_8 FILLER_73_1758 ();
 sg13g2_decap_8 FILLER_73_1765 ();
 sg13g2_decap_8 FILLER_73_1772 ();
 sg13g2_decap_8 FILLER_73_1779 ();
 sg13g2_decap_8 FILLER_73_1786 ();
 sg13g2_decap_8 FILLER_73_1793 ();
 sg13g2_decap_8 FILLER_73_1800 ();
 sg13g2_decap_8 FILLER_73_1807 ();
 sg13g2_decap_8 FILLER_73_1814 ();
 sg13g2_decap_8 FILLER_73_1821 ();
 sg13g2_decap_8 FILLER_73_1828 ();
 sg13g2_decap_8 FILLER_73_1835 ();
 sg13g2_decap_8 FILLER_73_1842 ();
 sg13g2_decap_8 FILLER_73_1849 ();
 sg13g2_decap_8 FILLER_73_1856 ();
 sg13g2_decap_8 FILLER_73_1863 ();
 sg13g2_decap_8 FILLER_73_1870 ();
 sg13g2_decap_8 FILLER_73_1877 ();
 sg13g2_decap_8 FILLER_73_1884 ();
 sg13g2_decap_8 FILLER_73_1891 ();
 sg13g2_decap_8 FILLER_73_1898 ();
 sg13g2_decap_8 FILLER_73_1905 ();
 sg13g2_decap_8 FILLER_73_1912 ();
 sg13g2_decap_8 FILLER_73_1919 ();
 sg13g2_fill_2 FILLER_73_1926 ();
 sg13g2_decap_8 FILLER_73_1941 ();
 sg13g2_decap_8 FILLER_73_1948 ();
 sg13g2_decap_8 FILLER_73_1955 ();
 sg13g2_decap_8 FILLER_73_1962 ();
 sg13g2_decap_8 FILLER_73_1969 ();
 sg13g2_decap_8 FILLER_73_1976 ();
 sg13g2_decap_4 FILLER_73_1983 ();
 sg13g2_fill_2 FILLER_73_1987 ();
 sg13g2_decap_8 FILLER_73_1993 ();
 sg13g2_decap_8 FILLER_73_2000 ();
 sg13g2_decap_8 FILLER_73_2007 ();
 sg13g2_decap_8 FILLER_73_2014 ();
 sg13g2_decap_8 FILLER_73_2021 ();
 sg13g2_decap_8 FILLER_73_2028 ();
 sg13g2_decap_8 FILLER_73_2035 ();
 sg13g2_decap_8 FILLER_73_2042 ();
 sg13g2_decap_8 FILLER_73_2049 ();
 sg13g2_decap_8 FILLER_73_2056 ();
 sg13g2_decap_8 FILLER_73_2063 ();
 sg13g2_decap_8 FILLER_73_2070 ();
 sg13g2_decap_8 FILLER_73_2077 ();
 sg13g2_decap_8 FILLER_73_2084 ();
 sg13g2_decap_8 FILLER_73_2091 ();
 sg13g2_decap_8 FILLER_73_2098 ();
 sg13g2_decap_8 FILLER_73_2105 ();
 sg13g2_decap_8 FILLER_73_2112 ();
 sg13g2_decap_8 FILLER_73_2119 ();
 sg13g2_decap_8 FILLER_73_2126 ();
 sg13g2_decap_8 FILLER_73_2133 ();
 sg13g2_decap_8 FILLER_73_2140 ();
 sg13g2_decap_8 FILLER_73_2147 ();
 sg13g2_decap_8 FILLER_73_2154 ();
 sg13g2_decap_4 FILLER_73_2161 ();
 sg13g2_fill_1 FILLER_73_2165 ();
 sg13g2_decap_8 FILLER_73_2174 ();
 sg13g2_decap_8 FILLER_73_2181 ();
 sg13g2_decap_8 FILLER_73_2188 ();
 sg13g2_decap_8 FILLER_73_2195 ();
 sg13g2_decap_8 FILLER_73_2202 ();
 sg13g2_decap_8 FILLER_73_2209 ();
 sg13g2_decap_8 FILLER_73_2216 ();
 sg13g2_decap_8 FILLER_73_2223 ();
 sg13g2_decap_8 FILLER_73_2230 ();
 sg13g2_decap_8 FILLER_73_2237 ();
 sg13g2_decap_8 FILLER_73_2244 ();
 sg13g2_decap_8 FILLER_73_2251 ();
 sg13g2_decap_8 FILLER_73_2258 ();
 sg13g2_decap_8 FILLER_73_2265 ();
 sg13g2_decap_8 FILLER_73_2272 ();
 sg13g2_decap_8 FILLER_73_2279 ();
 sg13g2_decap_8 FILLER_73_2286 ();
 sg13g2_decap_8 FILLER_73_2293 ();
 sg13g2_decap_8 FILLER_73_2300 ();
 sg13g2_decap_8 FILLER_73_2307 ();
 sg13g2_decap_8 FILLER_73_2314 ();
 sg13g2_decap_8 FILLER_73_2321 ();
 sg13g2_decap_8 FILLER_73_2328 ();
 sg13g2_decap_8 FILLER_73_2335 ();
 sg13g2_decap_8 FILLER_73_2342 ();
 sg13g2_decap_8 FILLER_73_2349 ();
 sg13g2_decap_8 FILLER_73_2356 ();
 sg13g2_decap_8 FILLER_73_2363 ();
 sg13g2_decap_8 FILLER_73_2370 ();
 sg13g2_decap_8 FILLER_73_2377 ();
 sg13g2_decap_8 FILLER_73_2384 ();
 sg13g2_decap_8 FILLER_73_2391 ();
 sg13g2_decap_8 FILLER_73_2398 ();
 sg13g2_decap_8 FILLER_73_2405 ();
 sg13g2_decap_8 FILLER_73_2412 ();
 sg13g2_decap_8 FILLER_73_2419 ();
 sg13g2_decap_8 FILLER_73_2426 ();
 sg13g2_decap_8 FILLER_73_2433 ();
 sg13g2_decap_8 FILLER_73_2440 ();
 sg13g2_decap_8 FILLER_73_2447 ();
 sg13g2_decap_8 FILLER_73_2454 ();
 sg13g2_decap_8 FILLER_73_2461 ();
 sg13g2_decap_8 FILLER_73_2468 ();
 sg13g2_decap_8 FILLER_73_2475 ();
 sg13g2_decap_8 FILLER_73_2482 ();
 sg13g2_decap_8 FILLER_73_2489 ();
 sg13g2_decap_8 FILLER_73_2496 ();
 sg13g2_decap_8 FILLER_73_2503 ();
 sg13g2_decap_8 FILLER_73_2510 ();
 sg13g2_decap_8 FILLER_73_2517 ();
 sg13g2_decap_8 FILLER_73_2524 ();
 sg13g2_decap_8 FILLER_73_2531 ();
 sg13g2_decap_8 FILLER_73_2538 ();
 sg13g2_decap_8 FILLER_73_2545 ();
 sg13g2_decap_8 FILLER_73_2552 ();
 sg13g2_decap_8 FILLER_73_2559 ();
 sg13g2_decap_8 FILLER_73_2566 ();
 sg13g2_decap_8 FILLER_73_2573 ();
 sg13g2_decap_8 FILLER_73_2580 ();
 sg13g2_decap_8 FILLER_73_2587 ();
 sg13g2_decap_8 FILLER_73_2594 ();
 sg13g2_decap_8 FILLER_73_2601 ();
 sg13g2_decap_8 FILLER_73_2608 ();
 sg13g2_decap_8 FILLER_73_2615 ();
 sg13g2_decap_8 FILLER_73_2622 ();
 sg13g2_decap_8 FILLER_73_2629 ();
 sg13g2_decap_8 FILLER_73_2636 ();
 sg13g2_decap_8 FILLER_73_2643 ();
 sg13g2_decap_8 FILLER_73_2650 ();
 sg13g2_decap_8 FILLER_73_2657 ();
 sg13g2_decap_4 FILLER_73_2664 ();
 sg13g2_fill_2 FILLER_73_2668 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_decap_8 FILLER_74_119 ();
 sg13g2_fill_2 FILLER_74_126 ();
 sg13g2_fill_1 FILLER_74_128 ();
 sg13g2_fill_1 FILLER_74_144 ();
 sg13g2_decap_8 FILLER_74_149 ();
 sg13g2_decap_8 FILLER_74_156 ();
 sg13g2_decap_8 FILLER_74_163 ();
 sg13g2_decap_8 FILLER_74_170 ();
 sg13g2_decap_8 FILLER_74_177 ();
 sg13g2_decap_8 FILLER_74_184 ();
 sg13g2_decap_8 FILLER_74_191 ();
 sg13g2_decap_8 FILLER_74_198 ();
 sg13g2_decap_8 FILLER_74_205 ();
 sg13g2_decap_8 FILLER_74_212 ();
 sg13g2_decap_8 FILLER_74_219 ();
 sg13g2_decap_8 FILLER_74_226 ();
 sg13g2_decap_8 FILLER_74_233 ();
 sg13g2_decap_8 FILLER_74_240 ();
 sg13g2_fill_2 FILLER_74_247 ();
 sg13g2_decap_8 FILLER_74_253 ();
 sg13g2_decap_8 FILLER_74_260 ();
 sg13g2_decap_8 FILLER_74_267 ();
 sg13g2_decap_8 FILLER_74_274 ();
 sg13g2_decap_8 FILLER_74_281 ();
 sg13g2_decap_8 FILLER_74_288 ();
 sg13g2_decap_8 FILLER_74_295 ();
 sg13g2_decap_8 FILLER_74_302 ();
 sg13g2_decap_8 FILLER_74_309 ();
 sg13g2_decap_8 FILLER_74_316 ();
 sg13g2_decap_8 FILLER_74_323 ();
 sg13g2_decap_8 FILLER_74_330 ();
 sg13g2_decap_8 FILLER_74_337 ();
 sg13g2_decap_8 FILLER_74_344 ();
 sg13g2_decap_8 FILLER_74_351 ();
 sg13g2_decap_8 FILLER_74_358 ();
 sg13g2_decap_8 FILLER_74_365 ();
 sg13g2_decap_8 FILLER_74_372 ();
 sg13g2_decap_8 FILLER_74_379 ();
 sg13g2_decap_8 FILLER_74_386 ();
 sg13g2_decap_8 FILLER_74_393 ();
 sg13g2_decap_8 FILLER_74_400 ();
 sg13g2_decap_8 FILLER_74_407 ();
 sg13g2_decap_8 FILLER_74_414 ();
 sg13g2_decap_4 FILLER_74_421 ();
 sg13g2_fill_1 FILLER_74_425 ();
 sg13g2_fill_1 FILLER_74_444 ();
 sg13g2_decap_8 FILLER_74_461 ();
 sg13g2_decap_8 FILLER_74_468 ();
 sg13g2_decap_8 FILLER_74_475 ();
 sg13g2_decap_8 FILLER_74_482 ();
 sg13g2_decap_8 FILLER_74_489 ();
 sg13g2_decap_8 FILLER_74_496 ();
 sg13g2_decap_8 FILLER_74_503 ();
 sg13g2_decap_8 FILLER_74_510 ();
 sg13g2_decap_8 FILLER_74_517 ();
 sg13g2_decap_8 FILLER_74_524 ();
 sg13g2_decap_8 FILLER_74_531 ();
 sg13g2_decap_8 FILLER_74_538 ();
 sg13g2_decap_8 FILLER_74_545 ();
 sg13g2_decap_8 FILLER_74_552 ();
 sg13g2_decap_8 FILLER_74_559 ();
 sg13g2_decap_4 FILLER_74_566 ();
 sg13g2_fill_2 FILLER_74_579 ();
 sg13g2_decap_8 FILLER_74_585 ();
 sg13g2_decap_8 FILLER_74_592 ();
 sg13g2_decap_8 FILLER_74_599 ();
 sg13g2_decap_8 FILLER_74_606 ();
 sg13g2_decap_8 FILLER_74_613 ();
 sg13g2_decap_8 FILLER_74_620 ();
 sg13g2_decap_8 FILLER_74_627 ();
 sg13g2_decap_8 FILLER_74_634 ();
 sg13g2_decap_8 FILLER_74_641 ();
 sg13g2_decap_8 FILLER_74_648 ();
 sg13g2_decap_8 FILLER_74_655 ();
 sg13g2_fill_2 FILLER_74_662 ();
 sg13g2_decap_8 FILLER_74_673 ();
 sg13g2_decap_8 FILLER_74_680 ();
 sg13g2_decap_8 FILLER_74_687 ();
 sg13g2_decap_8 FILLER_74_694 ();
 sg13g2_decap_8 FILLER_74_701 ();
 sg13g2_decap_8 FILLER_74_708 ();
 sg13g2_decap_8 FILLER_74_715 ();
 sg13g2_decap_4 FILLER_74_722 ();
 sg13g2_fill_1 FILLER_74_726 ();
 sg13g2_decap_8 FILLER_74_739 ();
 sg13g2_decap_8 FILLER_74_746 ();
 sg13g2_decap_8 FILLER_74_753 ();
 sg13g2_decap_8 FILLER_74_760 ();
 sg13g2_decap_8 FILLER_74_767 ();
 sg13g2_decap_8 FILLER_74_774 ();
 sg13g2_decap_8 FILLER_74_781 ();
 sg13g2_decap_8 FILLER_74_788 ();
 sg13g2_decap_8 FILLER_74_795 ();
 sg13g2_decap_8 FILLER_74_802 ();
 sg13g2_decap_8 FILLER_74_809 ();
 sg13g2_decap_8 FILLER_74_816 ();
 sg13g2_decap_8 FILLER_74_823 ();
 sg13g2_decap_8 FILLER_74_830 ();
 sg13g2_decap_8 FILLER_74_837 ();
 sg13g2_decap_8 FILLER_74_844 ();
 sg13g2_decap_8 FILLER_74_851 ();
 sg13g2_decap_8 FILLER_74_858 ();
 sg13g2_decap_8 FILLER_74_865 ();
 sg13g2_decap_8 FILLER_74_872 ();
 sg13g2_decap_8 FILLER_74_879 ();
 sg13g2_decap_8 FILLER_74_886 ();
 sg13g2_decap_8 FILLER_74_893 ();
 sg13g2_decap_8 FILLER_74_900 ();
 sg13g2_decap_8 FILLER_74_907 ();
 sg13g2_fill_2 FILLER_74_914 ();
 sg13g2_fill_1 FILLER_74_916 ();
 sg13g2_decap_8 FILLER_74_921 ();
 sg13g2_decap_8 FILLER_74_928 ();
 sg13g2_decap_8 FILLER_74_935 ();
 sg13g2_decap_8 FILLER_74_942 ();
 sg13g2_decap_8 FILLER_74_949 ();
 sg13g2_decap_8 FILLER_74_956 ();
 sg13g2_decap_8 FILLER_74_963 ();
 sg13g2_decap_8 FILLER_74_970 ();
 sg13g2_decap_8 FILLER_74_977 ();
 sg13g2_decap_8 FILLER_74_984 ();
 sg13g2_decap_8 FILLER_74_991 ();
 sg13g2_decap_8 FILLER_74_998 ();
 sg13g2_decap_8 FILLER_74_1005 ();
 sg13g2_decap_8 FILLER_74_1012 ();
 sg13g2_decap_8 FILLER_74_1019 ();
 sg13g2_decap_8 FILLER_74_1026 ();
 sg13g2_fill_1 FILLER_74_1033 ();
 sg13g2_decap_8 FILLER_74_1039 ();
 sg13g2_decap_8 FILLER_74_1046 ();
 sg13g2_decap_8 FILLER_74_1053 ();
 sg13g2_decap_8 FILLER_74_1060 ();
 sg13g2_decap_8 FILLER_74_1067 ();
 sg13g2_fill_2 FILLER_74_1074 ();
 sg13g2_decap_8 FILLER_74_1084 ();
 sg13g2_decap_8 FILLER_74_1091 ();
 sg13g2_decap_8 FILLER_74_1098 ();
 sg13g2_decap_8 FILLER_74_1105 ();
 sg13g2_decap_8 FILLER_74_1112 ();
 sg13g2_decap_8 FILLER_74_1119 ();
 sg13g2_decap_8 FILLER_74_1126 ();
 sg13g2_decap_8 FILLER_74_1133 ();
 sg13g2_decap_8 FILLER_74_1140 ();
 sg13g2_decap_4 FILLER_74_1147 ();
 sg13g2_decap_8 FILLER_74_1159 ();
 sg13g2_decap_8 FILLER_74_1166 ();
 sg13g2_decap_8 FILLER_74_1173 ();
 sg13g2_decap_8 FILLER_74_1180 ();
 sg13g2_decap_8 FILLER_74_1187 ();
 sg13g2_decap_8 FILLER_74_1194 ();
 sg13g2_decap_8 FILLER_74_1201 ();
 sg13g2_decap_8 FILLER_74_1208 ();
 sg13g2_decap_8 FILLER_74_1215 ();
 sg13g2_decap_8 FILLER_74_1222 ();
 sg13g2_decap_8 FILLER_74_1229 ();
 sg13g2_decap_8 FILLER_74_1236 ();
 sg13g2_decap_8 FILLER_74_1243 ();
 sg13g2_decap_8 FILLER_74_1250 ();
 sg13g2_decap_8 FILLER_74_1257 ();
 sg13g2_decap_8 FILLER_74_1264 ();
 sg13g2_decap_8 FILLER_74_1271 ();
 sg13g2_decap_8 FILLER_74_1278 ();
 sg13g2_decap_8 FILLER_74_1285 ();
 sg13g2_decap_4 FILLER_74_1292 ();
 sg13g2_fill_1 FILLER_74_1296 ();
 sg13g2_fill_2 FILLER_74_1301 ();
 sg13g2_decap_8 FILLER_74_1308 ();
 sg13g2_decap_8 FILLER_74_1315 ();
 sg13g2_decap_8 FILLER_74_1322 ();
 sg13g2_decap_8 FILLER_74_1329 ();
 sg13g2_decap_8 FILLER_74_1336 ();
 sg13g2_decap_8 FILLER_74_1343 ();
 sg13g2_decap_8 FILLER_74_1350 ();
 sg13g2_decap_8 FILLER_74_1357 ();
 sg13g2_decap_8 FILLER_74_1364 ();
 sg13g2_decap_8 FILLER_74_1371 ();
 sg13g2_decap_8 FILLER_74_1378 ();
 sg13g2_decap_8 FILLER_74_1385 ();
 sg13g2_decap_8 FILLER_74_1392 ();
 sg13g2_decap_8 FILLER_74_1399 ();
 sg13g2_decap_4 FILLER_74_1406 ();
 sg13g2_decap_8 FILLER_74_1422 ();
 sg13g2_decap_8 FILLER_74_1429 ();
 sg13g2_decap_8 FILLER_74_1436 ();
 sg13g2_decap_8 FILLER_74_1443 ();
 sg13g2_decap_8 FILLER_74_1450 ();
 sg13g2_decap_8 FILLER_74_1462 ();
 sg13g2_decap_8 FILLER_74_1469 ();
 sg13g2_decap_8 FILLER_74_1476 ();
 sg13g2_decap_8 FILLER_74_1483 ();
 sg13g2_decap_8 FILLER_74_1490 ();
 sg13g2_decap_8 FILLER_74_1497 ();
 sg13g2_decap_8 FILLER_74_1504 ();
 sg13g2_decap_8 FILLER_74_1511 ();
 sg13g2_decap_8 FILLER_74_1518 ();
 sg13g2_decap_8 FILLER_74_1525 ();
 sg13g2_decap_8 FILLER_74_1532 ();
 sg13g2_decap_8 FILLER_74_1539 ();
 sg13g2_decap_8 FILLER_74_1546 ();
 sg13g2_decap_8 FILLER_74_1553 ();
 sg13g2_decap_8 FILLER_74_1560 ();
 sg13g2_decap_8 FILLER_74_1567 ();
 sg13g2_decap_8 FILLER_74_1574 ();
 sg13g2_decap_8 FILLER_74_1581 ();
 sg13g2_decap_8 FILLER_74_1588 ();
 sg13g2_decap_8 FILLER_74_1595 ();
 sg13g2_decap_8 FILLER_74_1602 ();
 sg13g2_decap_8 FILLER_74_1609 ();
 sg13g2_decap_8 FILLER_74_1616 ();
 sg13g2_decap_4 FILLER_74_1623 ();
 sg13g2_fill_2 FILLER_74_1627 ();
 sg13g2_decap_8 FILLER_74_1634 ();
 sg13g2_decap_8 FILLER_74_1641 ();
 sg13g2_decap_8 FILLER_74_1648 ();
 sg13g2_decap_4 FILLER_74_1655 ();
 sg13g2_fill_2 FILLER_74_1659 ();
 sg13g2_decap_8 FILLER_74_1665 ();
 sg13g2_decap_8 FILLER_74_1672 ();
 sg13g2_decap_8 FILLER_74_1679 ();
 sg13g2_decap_8 FILLER_74_1686 ();
 sg13g2_decap_8 FILLER_74_1693 ();
 sg13g2_decap_8 FILLER_74_1700 ();
 sg13g2_decap_8 FILLER_74_1707 ();
 sg13g2_decap_8 FILLER_74_1714 ();
 sg13g2_decap_8 FILLER_74_1721 ();
 sg13g2_decap_8 FILLER_74_1728 ();
 sg13g2_decap_8 FILLER_74_1735 ();
 sg13g2_decap_8 FILLER_74_1742 ();
 sg13g2_decap_8 FILLER_74_1749 ();
 sg13g2_decap_8 FILLER_74_1756 ();
 sg13g2_decap_8 FILLER_74_1763 ();
 sg13g2_decap_8 FILLER_74_1770 ();
 sg13g2_decap_8 FILLER_74_1777 ();
 sg13g2_decap_8 FILLER_74_1784 ();
 sg13g2_decap_8 FILLER_74_1791 ();
 sg13g2_decap_8 FILLER_74_1798 ();
 sg13g2_decap_8 FILLER_74_1805 ();
 sg13g2_decap_8 FILLER_74_1812 ();
 sg13g2_decap_8 FILLER_74_1819 ();
 sg13g2_decap_8 FILLER_74_1826 ();
 sg13g2_decap_8 FILLER_74_1833 ();
 sg13g2_decap_8 FILLER_74_1840 ();
 sg13g2_decap_8 FILLER_74_1847 ();
 sg13g2_decap_8 FILLER_74_1854 ();
 sg13g2_decap_8 FILLER_74_1861 ();
 sg13g2_decap_8 FILLER_74_1868 ();
 sg13g2_decap_8 FILLER_74_1875 ();
 sg13g2_decap_8 FILLER_74_1882 ();
 sg13g2_decap_8 FILLER_74_1889 ();
 sg13g2_decap_8 FILLER_74_1896 ();
 sg13g2_decap_8 FILLER_74_1903 ();
 sg13g2_decap_8 FILLER_74_1910 ();
 sg13g2_decap_8 FILLER_74_1917 ();
 sg13g2_decap_8 FILLER_74_1924 ();
 sg13g2_decap_8 FILLER_74_1931 ();
 sg13g2_decap_8 FILLER_74_1938 ();
 sg13g2_decap_8 FILLER_74_1945 ();
 sg13g2_decap_8 FILLER_74_1952 ();
 sg13g2_decap_8 FILLER_74_1959 ();
 sg13g2_decap_8 FILLER_74_1966 ();
 sg13g2_decap_8 FILLER_74_1973 ();
 sg13g2_decap_8 FILLER_74_1980 ();
 sg13g2_decap_8 FILLER_74_1987 ();
 sg13g2_decap_8 FILLER_74_1994 ();
 sg13g2_decap_8 FILLER_74_2001 ();
 sg13g2_decap_8 FILLER_74_2008 ();
 sg13g2_decap_4 FILLER_74_2015 ();
 sg13g2_decap_8 FILLER_74_2032 ();
 sg13g2_decap_8 FILLER_74_2039 ();
 sg13g2_decap_8 FILLER_74_2046 ();
 sg13g2_decap_8 FILLER_74_2053 ();
 sg13g2_decap_8 FILLER_74_2060 ();
 sg13g2_decap_8 FILLER_74_2067 ();
 sg13g2_decap_8 FILLER_74_2074 ();
 sg13g2_decap_8 FILLER_74_2081 ();
 sg13g2_decap_8 FILLER_74_2088 ();
 sg13g2_decap_8 FILLER_74_2095 ();
 sg13g2_decap_8 FILLER_74_2102 ();
 sg13g2_decap_8 FILLER_74_2109 ();
 sg13g2_decap_8 FILLER_74_2116 ();
 sg13g2_decap_8 FILLER_74_2123 ();
 sg13g2_decap_8 FILLER_74_2130 ();
 sg13g2_decap_8 FILLER_74_2137 ();
 sg13g2_decap_8 FILLER_74_2144 ();
 sg13g2_decap_8 FILLER_74_2151 ();
 sg13g2_decap_8 FILLER_74_2158 ();
 sg13g2_decap_8 FILLER_74_2169 ();
 sg13g2_decap_8 FILLER_74_2176 ();
 sg13g2_decap_8 FILLER_74_2183 ();
 sg13g2_decap_8 FILLER_74_2190 ();
 sg13g2_decap_8 FILLER_74_2197 ();
 sg13g2_decap_8 FILLER_74_2204 ();
 sg13g2_decap_8 FILLER_74_2211 ();
 sg13g2_decap_8 FILLER_74_2218 ();
 sg13g2_decap_8 FILLER_74_2225 ();
 sg13g2_decap_8 FILLER_74_2232 ();
 sg13g2_decap_8 FILLER_74_2239 ();
 sg13g2_decap_8 FILLER_74_2246 ();
 sg13g2_decap_8 FILLER_74_2253 ();
 sg13g2_decap_8 FILLER_74_2260 ();
 sg13g2_decap_8 FILLER_74_2267 ();
 sg13g2_decap_8 FILLER_74_2274 ();
 sg13g2_decap_8 FILLER_74_2281 ();
 sg13g2_decap_8 FILLER_74_2288 ();
 sg13g2_decap_8 FILLER_74_2295 ();
 sg13g2_decap_8 FILLER_74_2302 ();
 sg13g2_decap_8 FILLER_74_2309 ();
 sg13g2_decap_8 FILLER_74_2316 ();
 sg13g2_decap_8 FILLER_74_2323 ();
 sg13g2_decap_8 FILLER_74_2330 ();
 sg13g2_decap_8 FILLER_74_2337 ();
 sg13g2_decap_8 FILLER_74_2344 ();
 sg13g2_decap_8 FILLER_74_2351 ();
 sg13g2_decap_8 FILLER_74_2358 ();
 sg13g2_decap_8 FILLER_74_2365 ();
 sg13g2_decap_8 FILLER_74_2372 ();
 sg13g2_decap_8 FILLER_74_2379 ();
 sg13g2_decap_8 FILLER_74_2386 ();
 sg13g2_decap_8 FILLER_74_2393 ();
 sg13g2_decap_8 FILLER_74_2400 ();
 sg13g2_decap_8 FILLER_74_2407 ();
 sg13g2_decap_8 FILLER_74_2414 ();
 sg13g2_decap_8 FILLER_74_2421 ();
 sg13g2_decap_8 FILLER_74_2428 ();
 sg13g2_decap_8 FILLER_74_2435 ();
 sg13g2_decap_8 FILLER_74_2442 ();
 sg13g2_decap_8 FILLER_74_2449 ();
 sg13g2_decap_8 FILLER_74_2456 ();
 sg13g2_decap_8 FILLER_74_2463 ();
 sg13g2_decap_8 FILLER_74_2470 ();
 sg13g2_decap_8 FILLER_74_2477 ();
 sg13g2_decap_8 FILLER_74_2484 ();
 sg13g2_decap_8 FILLER_74_2491 ();
 sg13g2_decap_8 FILLER_74_2498 ();
 sg13g2_decap_8 FILLER_74_2505 ();
 sg13g2_decap_8 FILLER_74_2512 ();
 sg13g2_decap_8 FILLER_74_2519 ();
 sg13g2_decap_8 FILLER_74_2526 ();
 sg13g2_decap_8 FILLER_74_2533 ();
 sg13g2_decap_8 FILLER_74_2540 ();
 sg13g2_decap_8 FILLER_74_2547 ();
 sg13g2_decap_8 FILLER_74_2554 ();
 sg13g2_decap_8 FILLER_74_2561 ();
 sg13g2_decap_8 FILLER_74_2568 ();
 sg13g2_decap_8 FILLER_74_2575 ();
 sg13g2_decap_8 FILLER_74_2582 ();
 sg13g2_decap_8 FILLER_74_2589 ();
 sg13g2_decap_8 FILLER_74_2596 ();
 sg13g2_decap_8 FILLER_74_2603 ();
 sg13g2_decap_8 FILLER_74_2610 ();
 sg13g2_decap_8 FILLER_74_2617 ();
 sg13g2_decap_8 FILLER_74_2624 ();
 sg13g2_decap_8 FILLER_74_2631 ();
 sg13g2_decap_8 FILLER_74_2638 ();
 sg13g2_decap_8 FILLER_74_2645 ();
 sg13g2_decap_8 FILLER_74_2652 ();
 sg13g2_decap_8 FILLER_74_2659 ();
 sg13g2_decap_4 FILLER_74_2666 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_4 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_164 ();
 sg13g2_decap_8 FILLER_75_171 ();
 sg13g2_decap_8 FILLER_75_178 ();
 sg13g2_decap_8 FILLER_75_185 ();
 sg13g2_decap_8 FILLER_75_192 ();
 sg13g2_decap_8 FILLER_75_199 ();
 sg13g2_decap_8 FILLER_75_206 ();
 sg13g2_decap_8 FILLER_75_213 ();
 sg13g2_decap_8 FILLER_75_220 ();
 sg13g2_decap_8 FILLER_75_227 ();
 sg13g2_decap_8 FILLER_75_234 ();
 sg13g2_decap_8 FILLER_75_241 ();
 sg13g2_decap_8 FILLER_75_248 ();
 sg13g2_decap_8 FILLER_75_255 ();
 sg13g2_decap_8 FILLER_75_262 ();
 sg13g2_decap_8 FILLER_75_269 ();
 sg13g2_decap_8 FILLER_75_276 ();
 sg13g2_decap_8 FILLER_75_283 ();
 sg13g2_decap_8 FILLER_75_290 ();
 sg13g2_decap_8 FILLER_75_297 ();
 sg13g2_decap_8 FILLER_75_304 ();
 sg13g2_decap_8 FILLER_75_311 ();
 sg13g2_decap_8 FILLER_75_318 ();
 sg13g2_decap_8 FILLER_75_325 ();
 sg13g2_decap_8 FILLER_75_332 ();
 sg13g2_decap_8 FILLER_75_339 ();
 sg13g2_decap_8 FILLER_75_346 ();
 sg13g2_decap_8 FILLER_75_353 ();
 sg13g2_decap_8 FILLER_75_360 ();
 sg13g2_decap_8 FILLER_75_367 ();
 sg13g2_decap_8 FILLER_75_374 ();
 sg13g2_decap_8 FILLER_75_381 ();
 sg13g2_decap_8 FILLER_75_388 ();
 sg13g2_decap_8 FILLER_75_395 ();
 sg13g2_decap_8 FILLER_75_402 ();
 sg13g2_decap_8 FILLER_75_409 ();
 sg13g2_decap_8 FILLER_75_416 ();
 sg13g2_decap_8 FILLER_75_423 ();
 sg13g2_decap_8 FILLER_75_430 ();
 sg13g2_decap_4 FILLER_75_437 ();
 sg13g2_decap_8 FILLER_75_445 ();
 sg13g2_decap_8 FILLER_75_466 ();
 sg13g2_decap_4 FILLER_75_473 ();
 sg13g2_fill_1 FILLER_75_477 ();
 sg13g2_decap_4 FILLER_75_483 ();
 sg13g2_fill_2 FILLER_75_487 ();
 sg13g2_decap_8 FILLER_75_494 ();
 sg13g2_decap_8 FILLER_75_501 ();
 sg13g2_decap_8 FILLER_75_508 ();
 sg13g2_decap_8 FILLER_75_515 ();
 sg13g2_decap_8 FILLER_75_522 ();
 sg13g2_decap_8 FILLER_75_529 ();
 sg13g2_decap_8 FILLER_75_536 ();
 sg13g2_decap_8 FILLER_75_543 ();
 sg13g2_decap_8 FILLER_75_550 ();
 sg13g2_decap_8 FILLER_75_557 ();
 sg13g2_decap_8 FILLER_75_564 ();
 sg13g2_decap_8 FILLER_75_571 ();
 sg13g2_decap_8 FILLER_75_578 ();
 sg13g2_decap_8 FILLER_75_585 ();
 sg13g2_decap_8 FILLER_75_592 ();
 sg13g2_decap_8 FILLER_75_599 ();
 sg13g2_decap_8 FILLER_75_606 ();
 sg13g2_decap_8 FILLER_75_613 ();
 sg13g2_decap_8 FILLER_75_620 ();
 sg13g2_decap_8 FILLER_75_627 ();
 sg13g2_decap_8 FILLER_75_634 ();
 sg13g2_decap_8 FILLER_75_641 ();
 sg13g2_decap_8 FILLER_75_648 ();
 sg13g2_decap_8 FILLER_75_655 ();
 sg13g2_decap_8 FILLER_75_662 ();
 sg13g2_decap_8 FILLER_75_669 ();
 sg13g2_decap_8 FILLER_75_676 ();
 sg13g2_decap_8 FILLER_75_683 ();
 sg13g2_decap_8 FILLER_75_690 ();
 sg13g2_fill_2 FILLER_75_697 ();
 sg13g2_fill_1 FILLER_75_699 ();
 sg13g2_decap_8 FILLER_75_735 ();
 sg13g2_decap_8 FILLER_75_742 ();
 sg13g2_decap_8 FILLER_75_749 ();
 sg13g2_decap_8 FILLER_75_756 ();
 sg13g2_decap_8 FILLER_75_763 ();
 sg13g2_decap_8 FILLER_75_770 ();
 sg13g2_decap_8 FILLER_75_777 ();
 sg13g2_decap_8 FILLER_75_784 ();
 sg13g2_decap_8 FILLER_75_791 ();
 sg13g2_decap_8 FILLER_75_798 ();
 sg13g2_decap_8 FILLER_75_805 ();
 sg13g2_decap_8 FILLER_75_812 ();
 sg13g2_decap_8 FILLER_75_819 ();
 sg13g2_decap_8 FILLER_75_826 ();
 sg13g2_decap_8 FILLER_75_833 ();
 sg13g2_decap_8 FILLER_75_840 ();
 sg13g2_decap_8 FILLER_75_847 ();
 sg13g2_decap_8 FILLER_75_854 ();
 sg13g2_decap_8 FILLER_75_861 ();
 sg13g2_decap_8 FILLER_75_868 ();
 sg13g2_decap_4 FILLER_75_875 ();
 sg13g2_fill_1 FILLER_75_879 ();
 sg13g2_decap_8 FILLER_75_883 ();
 sg13g2_decap_8 FILLER_75_890 ();
 sg13g2_decap_8 FILLER_75_897 ();
 sg13g2_decap_8 FILLER_75_904 ();
 sg13g2_decap_4 FILLER_75_911 ();
 sg13g2_fill_1 FILLER_75_915 ();
 sg13g2_decap_8 FILLER_75_921 ();
 sg13g2_decap_8 FILLER_75_928 ();
 sg13g2_decap_8 FILLER_75_935 ();
 sg13g2_decap_8 FILLER_75_942 ();
 sg13g2_fill_2 FILLER_75_949 ();
 sg13g2_fill_1 FILLER_75_951 ();
 sg13g2_fill_1 FILLER_75_964 ();
 sg13g2_decap_8 FILLER_75_973 ();
 sg13g2_fill_1 FILLER_75_980 ();
 sg13g2_decap_8 FILLER_75_993 ();
 sg13g2_decap_8 FILLER_75_1000 ();
 sg13g2_decap_4 FILLER_75_1007 ();
 sg13g2_decap_8 FILLER_75_1026 ();
 sg13g2_decap_8 FILLER_75_1033 ();
 sg13g2_decap_8 FILLER_75_1040 ();
 sg13g2_decap_8 FILLER_75_1047 ();
 sg13g2_decap_8 FILLER_75_1054 ();
 sg13g2_decap_8 FILLER_75_1061 ();
 sg13g2_decap_4 FILLER_75_1068 ();
 sg13g2_fill_1 FILLER_75_1072 ();
 sg13g2_decap_8 FILLER_75_1088 ();
 sg13g2_decap_8 FILLER_75_1095 ();
 sg13g2_decap_8 FILLER_75_1102 ();
 sg13g2_decap_8 FILLER_75_1109 ();
 sg13g2_decap_8 FILLER_75_1116 ();
 sg13g2_decap_8 FILLER_75_1123 ();
 sg13g2_decap_4 FILLER_75_1130 ();
 sg13g2_decap_8 FILLER_75_1138 ();
 sg13g2_decap_8 FILLER_75_1145 ();
 sg13g2_decap_8 FILLER_75_1156 ();
 sg13g2_decap_8 FILLER_75_1163 ();
 sg13g2_decap_8 FILLER_75_1170 ();
 sg13g2_decap_8 FILLER_75_1177 ();
 sg13g2_decap_8 FILLER_75_1184 ();
 sg13g2_decap_8 FILLER_75_1191 ();
 sg13g2_fill_2 FILLER_75_1198 ();
 sg13g2_fill_1 FILLER_75_1200 ();
 sg13g2_decap_8 FILLER_75_1205 ();
 sg13g2_decap_8 FILLER_75_1212 ();
 sg13g2_decap_8 FILLER_75_1219 ();
 sg13g2_decap_4 FILLER_75_1226 ();
 sg13g2_fill_2 FILLER_75_1230 ();
 sg13g2_decap_8 FILLER_75_1241 ();
 sg13g2_decap_8 FILLER_75_1248 ();
 sg13g2_decap_8 FILLER_75_1255 ();
 sg13g2_decap_8 FILLER_75_1262 ();
 sg13g2_decap_4 FILLER_75_1269 ();
 sg13g2_fill_1 FILLER_75_1282 ();
 sg13g2_decap_8 FILLER_75_1291 ();
 sg13g2_decap_8 FILLER_75_1298 ();
 sg13g2_decap_8 FILLER_75_1305 ();
 sg13g2_decap_8 FILLER_75_1312 ();
 sg13g2_decap_8 FILLER_75_1319 ();
 sg13g2_decap_8 FILLER_75_1326 ();
 sg13g2_decap_8 FILLER_75_1333 ();
 sg13g2_decap_8 FILLER_75_1340 ();
 sg13g2_decap_8 FILLER_75_1347 ();
 sg13g2_decap_8 FILLER_75_1354 ();
 sg13g2_decap_8 FILLER_75_1361 ();
 sg13g2_fill_2 FILLER_75_1368 ();
 sg13g2_fill_1 FILLER_75_1370 ();
 sg13g2_decap_4 FILLER_75_1380 ();
 sg13g2_fill_1 FILLER_75_1384 ();
 sg13g2_decap_8 FILLER_75_1400 ();
 sg13g2_fill_2 FILLER_75_1407 ();
 sg13g2_fill_1 FILLER_75_1409 ();
 sg13g2_decap_8 FILLER_75_1420 ();
 sg13g2_decap_8 FILLER_75_1427 ();
 sg13g2_decap_8 FILLER_75_1434 ();
 sg13g2_decap_8 FILLER_75_1441 ();
 sg13g2_decap_8 FILLER_75_1448 ();
 sg13g2_decap_8 FILLER_75_1455 ();
 sg13g2_decap_8 FILLER_75_1462 ();
 sg13g2_decap_8 FILLER_75_1469 ();
 sg13g2_decap_8 FILLER_75_1476 ();
 sg13g2_decap_8 FILLER_75_1483 ();
 sg13g2_decap_8 FILLER_75_1490 ();
 sg13g2_decap_8 FILLER_75_1502 ();
 sg13g2_decap_8 FILLER_75_1509 ();
 sg13g2_decap_8 FILLER_75_1516 ();
 sg13g2_decap_8 FILLER_75_1523 ();
 sg13g2_decap_8 FILLER_75_1530 ();
 sg13g2_decap_8 FILLER_75_1537 ();
 sg13g2_decap_8 FILLER_75_1544 ();
 sg13g2_decap_8 FILLER_75_1551 ();
 sg13g2_fill_2 FILLER_75_1558 ();
 sg13g2_decap_8 FILLER_75_1563 ();
 sg13g2_decap_8 FILLER_75_1570 ();
 sg13g2_decap_8 FILLER_75_1577 ();
 sg13g2_decap_8 FILLER_75_1584 ();
 sg13g2_decap_8 FILLER_75_1591 ();
 sg13g2_decap_8 FILLER_75_1598 ();
 sg13g2_decap_8 FILLER_75_1605 ();
 sg13g2_decap_8 FILLER_75_1612 ();
 sg13g2_decap_8 FILLER_75_1619 ();
 sg13g2_decap_8 FILLER_75_1626 ();
 sg13g2_decap_8 FILLER_75_1633 ();
 sg13g2_decap_8 FILLER_75_1640 ();
 sg13g2_decap_8 FILLER_75_1647 ();
 sg13g2_decap_8 FILLER_75_1654 ();
 sg13g2_decap_8 FILLER_75_1661 ();
 sg13g2_decap_8 FILLER_75_1668 ();
 sg13g2_decap_8 FILLER_75_1675 ();
 sg13g2_fill_2 FILLER_75_1682 ();
 sg13g2_decap_8 FILLER_75_1687 ();
 sg13g2_decap_8 FILLER_75_1694 ();
 sg13g2_decap_8 FILLER_75_1701 ();
 sg13g2_decap_8 FILLER_75_1708 ();
 sg13g2_decap_8 FILLER_75_1715 ();
 sg13g2_decap_8 FILLER_75_1722 ();
 sg13g2_decap_8 FILLER_75_1729 ();
 sg13g2_decap_8 FILLER_75_1736 ();
 sg13g2_decap_8 FILLER_75_1743 ();
 sg13g2_decap_8 FILLER_75_1750 ();
 sg13g2_decap_8 FILLER_75_1757 ();
 sg13g2_decap_8 FILLER_75_1764 ();
 sg13g2_decap_8 FILLER_75_1771 ();
 sg13g2_decap_8 FILLER_75_1778 ();
 sg13g2_decap_8 FILLER_75_1785 ();
 sg13g2_decap_8 FILLER_75_1792 ();
 sg13g2_decap_8 FILLER_75_1799 ();
 sg13g2_decap_8 FILLER_75_1806 ();
 sg13g2_decap_8 FILLER_75_1813 ();
 sg13g2_decap_8 FILLER_75_1820 ();
 sg13g2_decap_8 FILLER_75_1827 ();
 sg13g2_decap_8 FILLER_75_1834 ();
 sg13g2_decap_8 FILLER_75_1841 ();
 sg13g2_decap_8 FILLER_75_1848 ();
 sg13g2_decap_8 FILLER_75_1855 ();
 sg13g2_decap_8 FILLER_75_1862 ();
 sg13g2_decap_8 FILLER_75_1869 ();
 sg13g2_decap_8 FILLER_75_1876 ();
 sg13g2_decap_8 FILLER_75_1883 ();
 sg13g2_decap_8 FILLER_75_1890 ();
 sg13g2_decap_8 FILLER_75_1897 ();
 sg13g2_decap_8 FILLER_75_1904 ();
 sg13g2_decap_8 FILLER_75_1911 ();
 sg13g2_decap_8 FILLER_75_1918 ();
 sg13g2_decap_8 FILLER_75_1925 ();
 sg13g2_decap_8 FILLER_75_1932 ();
 sg13g2_decap_8 FILLER_75_1939 ();
 sg13g2_decap_8 FILLER_75_1946 ();
 sg13g2_decap_8 FILLER_75_1953 ();
 sg13g2_decap_8 FILLER_75_1960 ();
 sg13g2_decap_8 FILLER_75_1967 ();
 sg13g2_decap_8 FILLER_75_1974 ();
 sg13g2_decap_8 FILLER_75_1981 ();
 sg13g2_decap_8 FILLER_75_1988 ();
 sg13g2_decap_8 FILLER_75_1995 ();
 sg13g2_decap_8 FILLER_75_2002 ();
 sg13g2_decap_8 FILLER_75_2009 ();
 sg13g2_decap_8 FILLER_75_2016 ();
 sg13g2_decap_8 FILLER_75_2023 ();
 sg13g2_decap_8 FILLER_75_2030 ();
 sg13g2_decap_8 FILLER_75_2037 ();
 sg13g2_decap_8 FILLER_75_2044 ();
 sg13g2_decap_4 FILLER_75_2051 ();
 sg13g2_fill_2 FILLER_75_2055 ();
 sg13g2_decap_8 FILLER_75_2061 ();
 sg13g2_decap_8 FILLER_75_2068 ();
 sg13g2_decap_8 FILLER_75_2075 ();
 sg13g2_decap_4 FILLER_75_2082 ();
 sg13g2_fill_1 FILLER_75_2086 ();
 sg13g2_decap_8 FILLER_75_2091 ();
 sg13g2_decap_8 FILLER_75_2098 ();
 sg13g2_decap_8 FILLER_75_2105 ();
 sg13g2_decap_8 FILLER_75_2112 ();
 sg13g2_decap_4 FILLER_75_2119 ();
 sg13g2_decap_8 FILLER_75_2127 ();
 sg13g2_decap_8 FILLER_75_2134 ();
 sg13g2_decap_8 FILLER_75_2141 ();
 sg13g2_decap_8 FILLER_75_2148 ();
 sg13g2_decap_8 FILLER_75_2155 ();
 sg13g2_decap_4 FILLER_75_2162 ();
 sg13g2_fill_2 FILLER_75_2166 ();
 sg13g2_decap_8 FILLER_75_2172 ();
 sg13g2_decap_8 FILLER_75_2179 ();
 sg13g2_decap_8 FILLER_75_2186 ();
 sg13g2_decap_8 FILLER_75_2193 ();
 sg13g2_decap_8 FILLER_75_2200 ();
 sg13g2_decap_8 FILLER_75_2207 ();
 sg13g2_decap_8 FILLER_75_2214 ();
 sg13g2_decap_8 FILLER_75_2221 ();
 sg13g2_decap_8 FILLER_75_2228 ();
 sg13g2_decap_8 FILLER_75_2235 ();
 sg13g2_decap_8 FILLER_75_2242 ();
 sg13g2_decap_8 FILLER_75_2249 ();
 sg13g2_decap_8 FILLER_75_2256 ();
 sg13g2_decap_8 FILLER_75_2263 ();
 sg13g2_decap_8 FILLER_75_2270 ();
 sg13g2_decap_8 FILLER_75_2277 ();
 sg13g2_decap_8 FILLER_75_2284 ();
 sg13g2_decap_8 FILLER_75_2291 ();
 sg13g2_decap_8 FILLER_75_2298 ();
 sg13g2_decap_8 FILLER_75_2305 ();
 sg13g2_decap_8 FILLER_75_2312 ();
 sg13g2_decap_8 FILLER_75_2319 ();
 sg13g2_decap_8 FILLER_75_2326 ();
 sg13g2_decap_8 FILLER_75_2333 ();
 sg13g2_decap_8 FILLER_75_2340 ();
 sg13g2_decap_8 FILLER_75_2347 ();
 sg13g2_decap_8 FILLER_75_2354 ();
 sg13g2_decap_8 FILLER_75_2361 ();
 sg13g2_decap_8 FILLER_75_2368 ();
 sg13g2_decap_8 FILLER_75_2375 ();
 sg13g2_decap_8 FILLER_75_2382 ();
 sg13g2_decap_8 FILLER_75_2389 ();
 sg13g2_decap_8 FILLER_75_2396 ();
 sg13g2_decap_8 FILLER_75_2403 ();
 sg13g2_decap_8 FILLER_75_2410 ();
 sg13g2_decap_8 FILLER_75_2417 ();
 sg13g2_decap_8 FILLER_75_2424 ();
 sg13g2_decap_8 FILLER_75_2431 ();
 sg13g2_decap_8 FILLER_75_2438 ();
 sg13g2_decap_8 FILLER_75_2445 ();
 sg13g2_decap_8 FILLER_75_2452 ();
 sg13g2_decap_8 FILLER_75_2459 ();
 sg13g2_decap_8 FILLER_75_2466 ();
 sg13g2_decap_8 FILLER_75_2473 ();
 sg13g2_decap_8 FILLER_75_2480 ();
 sg13g2_decap_8 FILLER_75_2487 ();
 sg13g2_decap_8 FILLER_75_2494 ();
 sg13g2_decap_8 FILLER_75_2501 ();
 sg13g2_decap_8 FILLER_75_2508 ();
 sg13g2_decap_8 FILLER_75_2515 ();
 sg13g2_decap_8 FILLER_75_2522 ();
 sg13g2_decap_8 FILLER_75_2529 ();
 sg13g2_decap_8 FILLER_75_2536 ();
 sg13g2_decap_8 FILLER_75_2543 ();
 sg13g2_decap_8 FILLER_75_2550 ();
 sg13g2_decap_8 FILLER_75_2557 ();
 sg13g2_decap_8 FILLER_75_2564 ();
 sg13g2_decap_8 FILLER_75_2571 ();
 sg13g2_decap_8 FILLER_75_2578 ();
 sg13g2_decap_8 FILLER_75_2585 ();
 sg13g2_decap_8 FILLER_75_2592 ();
 sg13g2_decap_8 FILLER_75_2599 ();
 sg13g2_decap_8 FILLER_75_2606 ();
 sg13g2_decap_8 FILLER_75_2613 ();
 sg13g2_decap_8 FILLER_75_2620 ();
 sg13g2_decap_8 FILLER_75_2627 ();
 sg13g2_decap_8 FILLER_75_2634 ();
 sg13g2_decap_8 FILLER_75_2641 ();
 sg13g2_decap_8 FILLER_75_2648 ();
 sg13g2_decap_8 FILLER_75_2655 ();
 sg13g2_decap_8 FILLER_75_2662 ();
 sg13g2_fill_1 FILLER_75_2669 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_decap_8 FILLER_76_140 ();
 sg13g2_decap_8 FILLER_76_147 ();
 sg13g2_decap_4 FILLER_76_154 ();
 sg13g2_fill_2 FILLER_76_158 ();
 sg13g2_decap_8 FILLER_76_175 ();
 sg13g2_decap_8 FILLER_76_182 ();
 sg13g2_decap_8 FILLER_76_189 ();
 sg13g2_decap_8 FILLER_76_196 ();
 sg13g2_decap_8 FILLER_76_203 ();
 sg13g2_decap_8 FILLER_76_210 ();
 sg13g2_decap_8 FILLER_76_217 ();
 sg13g2_decap_8 FILLER_76_224 ();
 sg13g2_decap_8 FILLER_76_231 ();
 sg13g2_decap_8 FILLER_76_238 ();
 sg13g2_decap_8 FILLER_76_245 ();
 sg13g2_decap_8 FILLER_76_252 ();
 sg13g2_decap_8 FILLER_76_259 ();
 sg13g2_decap_8 FILLER_76_266 ();
 sg13g2_decap_8 FILLER_76_273 ();
 sg13g2_decap_8 FILLER_76_280 ();
 sg13g2_decap_8 FILLER_76_287 ();
 sg13g2_decap_8 FILLER_76_294 ();
 sg13g2_decap_8 FILLER_76_301 ();
 sg13g2_decap_8 FILLER_76_308 ();
 sg13g2_decap_8 FILLER_76_315 ();
 sg13g2_decap_8 FILLER_76_322 ();
 sg13g2_decap_8 FILLER_76_329 ();
 sg13g2_decap_8 FILLER_76_336 ();
 sg13g2_decap_8 FILLER_76_343 ();
 sg13g2_decap_8 FILLER_76_350 ();
 sg13g2_decap_8 FILLER_76_357 ();
 sg13g2_decap_8 FILLER_76_364 ();
 sg13g2_decap_8 FILLER_76_371 ();
 sg13g2_decap_8 FILLER_76_378 ();
 sg13g2_fill_2 FILLER_76_385 ();
 sg13g2_decap_8 FILLER_76_402 ();
 sg13g2_decap_8 FILLER_76_409 ();
 sg13g2_decap_8 FILLER_76_416 ();
 sg13g2_decap_8 FILLER_76_423 ();
 sg13g2_decap_8 FILLER_76_430 ();
 sg13g2_decap_8 FILLER_76_437 ();
 sg13g2_decap_8 FILLER_76_444 ();
 sg13g2_decap_8 FILLER_76_451 ();
 sg13g2_decap_8 FILLER_76_458 ();
 sg13g2_decap_8 FILLER_76_465 ();
 sg13g2_decap_8 FILLER_76_472 ();
 sg13g2_decap_8 FILLER_76_479 ();
 sg13g2_decap_8 FILLER_76_486 ();
 sg13g2_decap_8 FILLER_76_493 ();
 sg13g2_decap_8 FILLER_76_500 ();
 sg13g2_decap_8 FILLER_76_507 ();
 sg13g2_decap_8 FILLER_76_514 ();
 sg13g2_decap_8 FILLER_76_521 ();
 sg13g2_decap_8 FILLER_76_528 ();
 sg13g2_decap_8 FILLER_76_535 ();
 sg13g2_decap_8 FILLER_76_542 ();
 sg13g2_decap_8 FILLER_76_549 ();
 sg13g2_decap_4 FILLER_76_556 ();
 sg13g2_decap_8 FILLER_76_565 ();
 sg13g2_decap_8 FILLER_76_572 ();
 sg13g2_decap_8 FILLER_76_579 ();
 sg13g2_decap_8 FILLER_76_586 ();
 sg13g2_decap_8 FILLER_76_593 ();
 sg13g2_decap_8 FILLER_76_600 ();
 sg13g2_decap_4 FILLER_76_615 ();
 sg13g2_fill_1 FILLER_76_619 ();
 sg13g2_decap_8 FILLER_76_624 ();
 sg13g2_decap_8 FILLER_76_631 ();
 sg13g2_decap_8 FILLER_76_638 ();
 sg13g2_decap_8 FILLER_76_645 ();
 sg13g2_decap_8 FILLER_76_652 ();
 sg13g2_decap_8 FILLER_76_659 ();
 sg13g2_decap_8 FILLER_76_666 ();
 sg13g2_decap_8 FILLER_76_673 ();
 sg13g2_decap_8 FILLER_76_680 ();
 sg13g2_decap_8 FILLER_76_687 ();
 sg13g2_decap_8 FILLER_76_694 ();
 sg13g2_decap_4 FILLER_76_705 ();
 sg13g2_decap_4 FILLER_76_712 ();
 sg13g2_fill_2 FILLER_76_716 ();
 sg13g2_decap_4 FILLER_76_722 ();
 sg13g2_fill_1 FILLER_76_726 ();
 sg13g2_decap_8 FILLER_76_739 ();
 sg13g2_decap_8 FILLER_76_746 ();
 sg13g2_decap_8 FILLER_76_753 ();
 sg13g2_decap_8 FILLER_76_760 ();
 sg13g2_decap_8 FILLER_76_767 ();
 sg13g2_decap_8 FILLER_76_797 ();
 sg13g2_decap_8 FILLER_76_804 ();
 sg13g2_decap_8 FILLER_76_811 ();
 sg13g2_decap_4 FILLER_76_818 ();
 sg13g2_fill_2 FILLER_76_822 ();
 sg13g2_decap_8 FILLER_76_828 ();
 sg13g2_decap_8 FILLER_76_835 ();
 sg13g2_decap_8 FILLER_76_842 ();
 sg13g2_decap_4 FILLER_76_849 ();
 sg13g2_fill_2 FILLER_76_853 ();
 sg13g2_fill_2 FILLER_76_861 ();
 sg13g2_fill_1 FILLER_76_863 ();
 sg13g2_fill_1 FILLER_76_879 ();
 sg13g2_decap_8 FILLER_76_884 ();
 sg13g2_decap_8 FILLER_76_891 ();
 sg13g2_decap_8 FILLER_76_898 ();
 sg13g2_decap_8 FILLER_76_905 ();
 sg13g2_decap_4 FILLER_76_912 ();
 sg13g2_decap_8 FILLER_76_927 ();
 sg13g2_decap_8 FILLER_76_934 ();
 sg13g2_decap_8 FILLER_76_941 ();
 sg13g2_fill_1 FILLER_76_948 ();
 sg13g2_fill_1 FILLER_76_965 ();
 sg13g2_decap_8 FILLER_76_970 ();
 sg13g2_fill_1 FILLER_76_977 ();
 sg13g2_decap_8 FILLER_76_985 ();
 sg13g2_decap_8 FILLER_76_992 ();
 sg13g2_decap_4 FILLER_76_999 ();
 sg13g2_fill_2 FILLER_76_1003 ();
 sg13g2_decap_4 FILLER_76_1008 ();
 sg13g2_fill_2 FILLER_76_1012 ();
 sg13g2_decap_8 FILLER_76_1018 ();
 sg13g2_decap_8 FILLER_76_1025 ();
 sg13g2_decap_8 FILLER_76_1032 ();
 sg13g2_decap_8 FILLER_76_1039 ();
 sg13g2_decap_8 FILLER_76_1046 ();
 sg13g2_decap_8 FILLER_76_1053 ();
 sg13g2_decap_8 FILLER_76_1060 ();
 sg13g2_decap_8 FILLER_76_1067 ();
 sg13g2_fill_2 FILLER_76_1074 ();
 sg13g2_decap_8 FILLER_76_1081 ();
 sg13g2_decap_8 FILLER_76_1088 ();
 sg13g2_decap_8 FILLER_76_1095 ();
 sg13g2_decap_8 FILLER_76_1102 ();
 sg13g2_decap_8 FILLER_76_1109 ();
 sg13g2_decap_8 FILLER_76_1116 ();
 sg13g2_decap_8 FILLER_76_1123 ();
 sg13g2_decap_4 FILLER_76_1130 ();
 sg13g2_fill_1 FILLER_76_1134 ();
 sg13g2_decap_8 FILLER_76_1141 ();
 sg13g2_decap_8 FILLER_76_1148 ();
 sg13g2_decap_8 FILLER_76_1155 ();
 sg13g2_decap_8 FILLER_76_1162 ();
 sg13g2_decap_4 FILLER_76_1169 ();
 sg13g2_decap_8 FILLER_76_1177 ();
 sg13g2_decap_8 FILLER_76_1184 ();
 sg13g2_decap_8 FILLER_76_1191 ();
 sg13g2_decap_8 FILLER_76_1198 ();
 sg13g2_decap_8 FILLER_76_1205 ();
 sg13g2_decap_8 FILLER_76_1212 ();
 sg13g2_decap_8 FILLER_76_1219 ();
 sg13g2_decap_8 FILLER_76_1226 ();
 sg13g2_decap_8 FILLER_76_1233 ();
 sg13g2_decap_8 FILLER_76_1240 ();
 sg13g2_decap_8 FILLER_76_1247 ();
 sg13g2_decap_8 FILLER_76_1254 ();
 sg13g2_decap_8 FILLER_76_1261 ();
 sg13g2_decap_4 FILLER_76_1268 ();
 sg13g2_fill_1 FILLER_76_1272 ();
 sg13g2_decap_8 FILLER_76_1278 ();
 sg13g2_decap_8 FILLER_76_1285 ();
 sg13g2_decap_8 FILLER_76_1292 ();
 sg13g2_fill_1 FILLER_76_1299 ();
 sg13g2_decap_8 FILLER_76_1304 ();
 sg13g2_decap_8 FILLER_76_1311 ();
 sg13g2_fill_2 FILLER_76_1318 ();
 sg13g2_decap_8 FILLER_76_1332 ();
 sg13g2_decap_8 FILLER_76_1339 ();
 sg13g2_decap_8 FILLER_76_1346 ();
 sg13g2_decap_8 FILLER_76_1353 ();
 sg13g2_decap_4 FILLER_76_1360 ();
 sg13g2_fill_2 FILLER_76_1369 ();
 sg13g2_fill_2 FILLER_76_1374 ();
 sg13g2_fill_1 FILLER_76_1376 ();
 sg13g2_decap_4 FILLER_76_1381 ();
 sg13g2_decap_8 FILLER_76_1390 ();
 sg13g2_decap_8 FILLER_76_1397 ();
 sg13g2_decap_8 FILLER_76_1404 ();
 sg13g2_decap_4 FILLER_76_1411 ();
 sg13g2_fill_1 FILLER_76_1415 ();
 sg13g2_fill_1 FILLER_76_1431 ();
 sg13g2_fill_2 FILLER_76_1447 ();
 sg13g2_fill_1 FILLER_76_1455 ();
 sg13g2_decap_8 FILLER_76_1471 ();
 sg13g2_decap_8 FILLER_76_1478 ();
 sg13g2_decap_8 FILLER_76_1485 ();
 sg13g2_decap_8 FILLER_76_1492 ();
 sg13g2_decap_8 FILLER_76_1499 ();
 sg13g2_decap_8 FILLER_76_1506 ();
 sg13g2_fill_1 FILLER_76_1513 ();
 sg13g2_decap_8 FILLER_76_1519 ();
 sg13g2_decap_8 FILLER_76_1529 ();
 sg13g2_fill_2 FILLER_76_1536 ();
 sg13g2_fill_1 FILLER_76_1538 ();
 sg13g2_decap_8 FILLER_76_1545 ();
 sg13g2_decap_8 FILLER_76_1552 ();
 sg13g2_fill_1 FILLER_76_1559 ();
 sg13g2_decap_8 FILLER_76_1564 ();
 sg13g2_decap_8 FILLER_76_1571 ();
 sg13g2_decap_8 FILLER_76_1578 ();
 sg13g2_decap_8 FILLER_76_1585 ();
 sg13g2_decap_8 FILLER_76_1592 ();
 sg13g2_decap_8 FILLER_76_1599 ();
 sg13g2_decap_8 FILLER_76_1606 ();
 sg13g2_decap_8 FILLER_76_1613 ();
 sg13g2_decap_8 FILLER_76_1620 ();
 sg13g2_decap_8 FILLER_76_1627 ();
 sg13g2_fill_1 FILLER_76_1634 ();
 sg13g2_decap_8 FILLER_76_1650 ();
 sg13g2_decap_8 FILLER_76_1657 ();
 sg13g2_decap_8 FILLER_76_1664 ();
 sg13g2_decap_8 FILLER_76_1671 ();
 sg13g2_decap_4 FILLER_76_1678 ();
 sg13g2_fill_2 FILLER_76_1682 ();
 sg13g2_decap_8 FILLER_76_1688 ();
 sg13g2_decap_8 FILLER_76_1695 ();
 sg13g2_decap_8 FILLER_76_1702 ();
 sg13g2_decap_8 FILLER_76_1709 ();
 sg13g2_decap_8 FILLER_76_1716 ();
 sg13g2_decap_8 FILLER_76_1723 ();
 sg13g2_decap_8 FILLER_76_1730 ();
 sg13g2_decap_8 FILLER_76_1737 ();
 sg13g2_decap_8 FILLER_76_1744 ();
 sg13g2_decap_8 FILLER_76_1751 ();
 sg13g2_decap_8 FILLER_76_1758 ();
 sg13g2_decap_8 FILLER_76_1765 ();
 sg13g2_decap_8 FILLER_76_1772 ();
 sg13g2_decap_8 FILLER_76_1779 ();
 sg13g2_decap_8 FILLER_76_1786 ();
 sg13g2_decap_8 FILLER_76_1793 ();
 sg13g2_decap_8 FILLER_76_1800 ();
 sg13g2_decap_8 FILLER_76_1807 ();
 sg13g2_decap_8 FILLER_76_1814 ();
 sg13g2_decap_8 FILLER_76_1821 ();
 sg13g2_decap_8 FILLER_76_1828 ();
 sg13g2_decap_8 FILLER_76_1835 ();
 sg13g2_decap_8 FILLER_76_1842 ();
 sg13g2_decap_8 FILLER_76_1849 ();
 sg13g2_decap_8 FILLER_76_1856 ();
 sg13g2_decap_8 FILLER_76_1863 ();
 sg13g2_decap_8 FILLER_76_1870 ();
 sg13g2_decap_8 FILLER_76_1877 ();
 sg13g2_decap_8 FILLER_76_1884 ();
 sg13g2_decap_8 FILLER_76_1891 ();
 sg13g2_decap_8 FILLER_76_1898 ();
 sg13g2_decap_8 FILLER_76_1905 ();
 sg13g2_decap_8 FILLER_76_1912 ();
 sg13g2_decap_8 FILLER_76_1919 ();
 sg13g2_decap_8 FILLER_76_1926 ();
 sg13g2_decap_8 FILLER_76_1933 ();
 sg13g2_decap_8 FILLER_76_1940 ();
 sg13g2_decap_8 FILLER_76_1947 ();
 sg13g2_decap_8 FILLER_76_1954 ();
 sg13g2_decap_8 FILLER_76_1961 ();
 sg13g2_decap_8 FILLER_76_1968 ();
 sg13g2_decap_8 FILLER_76_1975 ();
 sg13g2_decap_8 FILLER_76_1982 ();
 sg13g2_decap_8 FILLER_76_1989 ();
 sg13g2_decap_8 FILLER_76_1996 ();
 sg13g2_decap_8 FILLER_76_2003 ();
 sg13g2_decap_8 FILLER_76_2010 ();
 sg13g2_decap_8 FILLER_76_2017 ();
 sg13g2_decap_8 FILLER_76_2024 ();
 sg13g2_decap_8 FILLER_76_2031 ();
 sg13g2_decap_8 FILLER_76_2038 ();
 sg13g2_decap_8 FILLER_76_2045 ();
 sg13g2_decap_8 FILLER_76_2052 ();
 sg13g2_decap_8 FILLER_76_2059 ();
 sg13g2_decap_8 FILLER_76_2066 ();
 sg13g2_decap_8 FILLER_76_2073 ();
 sg13g2_decap_8 FILLER_76_2080 ();
 sg13g2_decap_8 FILLER_76_2087 ();
 sg13g2_decap_8 FILLER_76_2094 ();
 sg13g2_decap_8 FILLER_76_2101 ();
 sg13g2_decap_8 FILLER_76_2108 ();
 sg13g2_decap_8 FILLER_76_2115 ();
 sg13g2_decap_8 FILLER_76_2122 ();
 sg13g2_decap_8 FILLER_76_2129 ();
 sg13g2_decap_8 FILLER_76_2136 ();
 sg13g2_decap_8 FILLER_76_2143 ();
 sg13g2_decap_8 FILLER_76_2150 ();
 sg13g2_decap_8 FILLER_76_2157 ();
 sg13g2_decap_8 FILLER_76_2164 ();
 sg13g2_decap_8 FILLER_76_2171 ();
 sg13g2_decap_8 FILLER_76_2178 ();
 sg13g2_decap_8 FILLER_76_2185 ();
 sg13g2_decap_8 FILLER_76_2192 ();
 sg13g2_decap_8 FILLER_76_2199 ();
 sg13g2_decap_8 FILLER_76_2206 ();
 sg13g2_decap_8 FILLER_76_2213 ();
 sg13g2_decap_8 FILLER_76_2220 ();
 sg13g2_decap_8 FILLER_76_2227 ();
 sg13g2_decap_8 FILLER_76_2234 ();
 sg13g2_decap_8 FILLER_76_2241 ();
 sg13g2_decap_8 FILLER_76_2248 ();
 sg13g2_decap_8 FILLER_76_2255 ();
 sg13g2_decap_8 FILLER_76_2262 ();
 sg13g2_decap_8 FILLER_76_2269 ();
 sg13g2_decap_8 FILLER_76_2276 ();
 sg13g2_decap_8 FILLER_76_2283 ();
 sg13g2_decap_8 FILLER_76_2290 ();
 sg13g2_decap_8 FILLER_76_2297 ();
 sg13g2_decap_8 FILLER_76_2304 ();
 sg13g2_decap_8 FILLER_76_2311 ();
 sg13g2_decap_8 FILLER_76_2318 ();
 sg13g2_decap_8 FILLER_76_2325 ();
 sg13g2_decap_8 FILLER_76_2332 ();
 sg13g2_decap_8 FILLER_76_2339 ();
 sg13g2_decap_8 FILLER_76_2346 ();
 sg13g2_decap_8 FILLER_76_2353 ();
 sg13g2_decap_8 FILLER_76_2360 ();
 sg13g2_decap_8 FILLER_76_2367 ();
 sg13g2_decap_8 FILLER_76_2374 ();
 sg13g2_decap_8 FILLER_76_2381 ();
 sg13g2_decap_8 FILLER_76_2388 ();
 sg13g2_decap_8 FILLER_76_2395 ();
 sg13g2_decap_8 FILLER_76_2402 ();
 sg13g2_decap_8 FILLER_76_2409 ();
 sg13g2_decap_8 FILLER_76_2416 ();
 sg13g2_decap_8 FILLER_76_2423 ();
 sg13g2_decap_8 FILLER_76_2430 ();
 sg13g2_decap_8 FILLER_76_2437 ();
 sg13g2_decap_8 FILLER_76_2444 ();
 sg13g2_decap_8 FILLER_76_2451 ();
 sg13g2_decap_8 FILLER_76_2458 ();
 sg13g2_decap_8 FILLER_76_2465 ();
 sg13g2_decap_8 FILLER_76_2472 ();
 sg13g2_decap_8 FILLER_76_2479 ();
 sg13g2_decap_8 FILLER_76_2486 ();
 sg13g2_decap_8 FILLER_76_2493 ();
 sg13g2_decap_8 FILLER_76_2500 ();
 sg13g2_decap_8 FILLER_76_2507 ();
 sg13g2_decap_8 FILLER_76_2514 ();
 sg13g2_decap_8 FILLER_76_2521 ();
 sg13g2_decap_8 FILLER_76_2528 ();
 sg13g2_decap_8 FILLER_76_2535 ();
 sg13g2_decap_8 FILLER_76_2542 ();
 sg13g2_decap_8 FILLER_76_2549 ();
 sg13g2_decap_8 FILLER_76_2556 ();
 sg13g2_decap_8 FILLER_76_2563 ();
 sg13g2_decap_8 FILLER_76_2570 ();
 sg13g2_decap_8 FILLER_76_2577 ();
 sg13g2_decap_8 FILLER_76_2584 ();
 sg13g2_decap_8 FILLER_76_2591 ();
 sg13g2_decap_8 FILLER_76_2598 ();
 sg13g2_decap_8 FILLER_76_2605 ();
 sg13g2_decap_8 FILLER_76_2612 ();
 sg13g2_decap_8 FILLER_76_2619 ();
 sg13g2_decap_8 FILLER_76_2626 ();
 sg13g2_decap_8 FILLER_76_2633 ();
 sg13g2_decap_8 FILLER_76_2640 ();
 sg13g2_decap_8 FILLER_76_2647 ();
 sg13g2_decap_8 FILLER_76_2654 ();
 sg13g2_decap_8 FILLER_76_2661 ();
 sg13g2_fill_2 FILLER_76_2668 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_fill_1 FILLER_77_147 ();
 sg13g2_decap_8 FILLER_77_189 ();
 sg13g2_decap_8 FILLER_77_196 ();
 sg13g2_decap_8 FILLER_77_203 ();
 sg13g2_decap_4 FILLER_77_210 ();
 sg13g2_fill_1 FILLER_77_214 ();
 sg13g2_decap_8 FILLER_77_230 ();
 sg13g2_decap_8 FILLER_77_237 ();
 sg13g2_decap_8 FILLER_77_244 ();
 sg13g2_decap_8 FILLER_77_251 ();
 sg13g2_decap_8 FILLER_77_258 ();
 sg13g2_decap_8 FILLER_77_265 ();
 sg13g2_fill_1 FILLER_77_272 ();
 sg13g2_decap_8 FILLER_77_288 ();
 sg13g2_decap_8 FILLER_77_295 ();
 sg13g2_decap_8 FILLER_77_302 ();
 sg13g2_fill_2 FILLER_77_309 ();
 sg13g2_fill_1 FILLER_77_326 ();
 sg13g2_decap_8 FILLER_77_331 ();
 sg13g2_decap_8 FILLER_77_338 ();
 sg13g2_decap_8 FILLER_77_345 ();
 sg13g2_decap_8 FILLER_77_352 ();
 sg13g2_decap_8 FILLER_77_359 ();
 sg13g2_decap_8 FILLER_77_366 ();
 sg13g2_decap_8 FILLER_77_373 ();
 sg13g2_decap_8 FILLER_77_380 ();
 sg13g2_fill_2 FILLER_77_387 ();
 sg13g2_fill_1 FILLER_77_389 ();
 sg13g2_decap_8 FILLER_77_399 ();
 sg13g2_decap_8 FILLER_77_406 ();
 sg13g2_decap_8 FILLER_77_413 ();
 sg13g2_fill_2 FILLER_77_420 ();
 sg13g2_decap_8 FILLER_77_427 ();
 sg13g2_decap_8 FILLER_77_434 ();
 sg13g2_decap_8 FILLER_77_441 ();
 sg13g2_fill_2 FILLER_77_448 ();
 sg13g2_fill_2 FILLER_77_454 ();
 sg13g2_fill_1 FILLER_77_456 ();
 sg13g2_decap_8 FILLER_77_470 ();
 sg13g2_fill_2 FILLER_77_477 ();
 sg13g2_fill_2 FILLER_77_483 ();
 sg13g2_fill_2 FILLER_77_489 ();
 sg13g2_decap_8 FILLER_77_496 ();
 sg13g2_decap_8 FILLER_77_503 ();
 sg13g2_decap_8 FILLER_77_510 ();
 sg13g2_decap_8 FILLER_77_517 ();
 sg13g2_decap_8 FILLER_77_524 ();
 sg13g2_decap_8 FILLER_77_531 ();
 sg13g2_decap_8 FILLER_77_538 ();
 sg13g2_fill_2 FILLER_77_545 ();
 sg13g2_fill_1 FILLER_77_547 ();
 sg13g2_decap_8 FILLER_77_551 ();
 sg13g2_decap_8 FILLER_77_558 ();
 sg13g2_decap_8 FILLER_77_565 ();
 sg13g2_decap_4 FILLER_77_572 ();
 sg13g2_fill_2 FILLER_77_576 ();
 sg13g2_decap_8 FILLER_77_583 ();
 sg13g2_decap_8 FILLER_77_590 ();
 sg13g2_decap_8 FILLER_77_597 ();
 sg13g2_decap_8 FILLER_77_604 ();
 sg13g2_decap_8 FILLER_77_611 ();
 sg13g2_decap_8 FILLER_77_618 ();
 sg13g2_decap_4 FILLER_77_625 ();
 sg13g2_decap_8 FILLER_77_633 ();
 sg13g2_fill_2 FILLER_77_640 ();
 sg13g2_decap_8 FILLER_77_647 ();
 sg13g2_decap_8 FILLER_77_654 ();
 sg13g2_fill_2 FILLER_77_661 ();
 sg13g2_fill_1 FILLER_77_663 ();
 sg13g2_decap_8 FILLER_77_675 ();
 sg13g2_decap_8 FILLER_77_682 ();
 sg13g2_decap_4 FILLER_77_689 ();
 sg13g2_fill_1 FILLER_77_693 ();
 sg13g2_decap_4 FILLER_77_699 ();
 sg13g2_decap_8 FILLER_77_734 ();
 sg13g2_decap_4 FILLER_77_741 ();
 sg13g2_fill_2 FILLER_77_745 ();
 sg13g2_fill_1 FILLER_77_757 ();
 sg13g2_fill_2 FILLER_77_761 ();
 sg13g2_fill_1 FILLER_77_773 ();
 sg13g2_decap_8 FILLER_77_797 ();
 sg13g2_decap_8 FILLER_77_804 ();
 sg13g2_decap_8 FILLER_77_811 ();
 sg13g2_decap_8 FILLER_77_830 ();
 sg13g2_decap_8 FILLER_77_837 ();
 sg13g2_decap_8 FILLER_77_844 ();
 sg13g2_decap_8 FILLER_77_859 ();
 sg13g2_decap_8 FILLER_77_866 ();
 sg13g2_fill_1 FILLER_77_878 ();
 sg13g2_decap_8 FILLER_77_883 ();
 sg13g2_decap_8 FILLER_77_890 ();
 sg13g2_decap_8 FILLER_77_897 ();
 sg13g2_fill_2 FILLER_77_904 ();
 sg13g2_fill_1 FILLER_77_906 ();
 sg13g2_decap_4 FILLER_77_916 ();
 sg13g2_decap_8 FILLER_77_925 ();
 sg13g2_decap_8 FILLER_77_932 ();
 sg13g2_decap_8 FILLER_77_939 ();
 sg13g2_decap_8 FILLER_77_946 ();
 sg13g2_decap_8 FILLER_77_953 ();
 sg13g2_decap_8 FILLER_77_960 ();
 sg13g2_fill_2 FILLER_77_967 ();
 sg13g2_fill_1 FILLER_77_969 ();
 sg13g2_decap_8 FILLER_77_985 ();
 sg13g2_decap_4 FILLER_77_992 ();
 sg13g2_fill_1 FILLER_77_1004 ();
 sg13g2_fill_1 FILLER_77_1021 ();
 sg13g2_decap_8 FILLER_77_1032 ();
 sg13g2_decap_8 FILLER_77_1039 ();
 sg13g2_decap_8 FILLER_77_1046 ();
 sg13g2_decap_8 FILLER_77_1053 ();
 sg13g2_decap_8 FILLER_77_1060 ();
 sg13g2_decap_8 FILLER_77_1067 ();
 sg13g2_fill_2 FILLER_77_1074 ();
 sg13g2_fill_2 FILLER_77_1080 ();
 sg13g2_decap_8 FILLER_77_1087 ();
 sg13g2_decap_8 FILLER_77_1094 ();
 sg13g2_decap_8 FILLER_77_1101 ();
 sg13g2_fill_2 FILLER_77_1108 ();
 sg13g2_decap_8 FILLER_77_1114 ();
 sg13g2_decap_8 FILLER_77_1121 ();
 sg13g2_fill_1 FILLER_77_1128 ();
 sg13g2_decap_4 FILLER_77_1133 ();
 sg13g2_fill_1 FILLER_77_1137 ();
 sg13g2_decap_4 FILLER_77_1143 ();
 sg13g2_decap_8 FILLER_77_1156 ();
 sg13g2_decap_8 FILLER_77_1163 ();
 sg13g2_decap_8 FILLER_77_1170 ();
 sg13g2_decap_4 FILLER_77_1177 ();
 sg13g2_fill_1 FILLER_77_1181 ();
 sg13g2_decap_8 FILLER_77_1186 ();
 sg13g2_decap_4 FILLER_77_1193 ();
 sg13g2_decap_8 FILLER_77_1205 ();
 sg13g2_decap_8 FILLER_77_1212 ();
 sg13g2_decap_8 FILLER_77_1219 ();
 sg13g2_fill_1 FILLER_77_1226 ();
 sg13g2_decap_8 FILLER_77_1231 ();
 sg13g2_decap_8 FILLER_77_1238 ();
 sg13g2_decap_8 FILLER_77_1245 ();
 sg13g2_fill_2 FILLER_77_1252 ();
 sg13g2_fill_1 FILLER_77_1254 ();
 sg13g2_fill_2 FILLER_77_1270 ();
 sg13g2_fill_1 FILLER_77_1272 ();
 sg13g2_decap_8 FILLER_77_1280 ();
 sg13g2_decap_8 FILLER_77_1302 ();
 sg13g2_decap_8 FILLER_77_1309 ();
 sg13g2_decap_4 FILLER_77_1316 ();
 sg13g2_decap_8 FILLER_77_1325 ();
 sg13g2_decap_8 FILLER_77_1332 ();
 sg13g2_decap_8 FILLER_77_1339 ();
 sg13g2_decap_4 FILLER_77_1346 ();
 sg13g2_fill_1 FILLER_77_1350 ();
 sg13g2_decap_8 FILLER_77_1355 ();
 sg13g2_fill_1 FILLER_77_1362 ();
 sg13g2_decap_8 FILLER_77_1368 ();
 sg13g2_decap_4 FILLER_77_1375 ();
 sg13g2_fill_1 FILLER_77_1379 ();
 sg13g2_decap_8 FILLER_77_1398 ();
 sg13g2_fill_1 FILLER_77_1405 ();
 sg13g2_decap_4 FILLER_77_1410 ();
 sg13g2_fill_2 FILLER_77_1414 ();
 sg13g2_decap_8 FILLER_77_1420 ();
 sg13g2_decap_4 FILLER_77_1427 ();
 sg13g2_fill_1 FILLER_77_1431 ();
 sg13g2_decap_8 FILLER_77_1437 ();
 sg13g2_decap_4 FILLER_77_1444 ();
 sg13g2_decap_4 FILLER_77_1452 ();
 sg13g2_decap_8 FILLER_77_1461 ();
 sg13g2_decap_8 FILLER_77_1468 ();
 sg13g2_decap_8 FILLER_77_1475 ();
 sg13g2_decap_4 FILLER_77_1482 ();
 sg13g2_fill_1 FILLER_77_1486 ();
 sg13g2_decap_8 FILLER_77_1491 ();
 sg13g2_decap_8 FILLER_77_1498 ();
 sg13g2_decap_8 FILLER_77_1505 ();
 sg13g2_decap_8 FILLER_77_1512 ();
 sg13g2_fill_1 FILLER_77_1519 ();
 sg13g2_fill_1 FILLER_77_1525 ();
 sg13g2_decap_4 FILLER_77_1530 ();
 sg13g2_fill_2 FILLER_77_1534 ();
 sg13g2_decap_8 FILLER_77_1541 ();
 sg13g2_decap_8 FILLER_77_1548 ();
 sg13g2_decap_8 FILLER_77_1555 ();
 sg13g2_fill_2 FILLER_77_1562 ();
 sg13g2_fill_1 FILLER_77_1575 ();
 sg13g2_fill_1 FILLER_77_1586 ();
 sg13g2_decap_8 FILLER_77_1594 ();
 sg13g2_fill_2 FILLER_77_1601 ();
 sg13g2_fill_1 FILLER_77_1603 ();
 sg13g2_decap_8 FILLER_77_1609 ();
 sg13g2_decap_4 FILLER_77_1616 ();
 sg13g2_fill_2 FILLER_77_1629 ();
 sg13g2_decap_8 FILLER_77_1639 ();
 sg13g2_decap_8 FILLER_77_1646 ();
 sg13g2_decap_8 FILLER_77_1653 ();
 sg13g2_decap_4 FILLER_77_1660 ();
 sg13g2_decap_8 FILLER_77_1668 ();
 sg13g2_decap_8 FILLER_77_1683 ();
 sg13g2_decap_8 FILLER_77_1690 ();
 sg13g2_decap_8 FILLER_77_1697 ();
 sg13g2_decap_8 FILLER_77_1704 ();
 sg13g2_decap_8 FILLER_77_1711 ();
 sg13g2_decap_8 FILLER_77_1718 ();
 sg13g2_decap_8 FILLER_77_1725 ();
 sg13g2_decap_8 FILLER_77_1732 ();
 sg13g2_decap_8 FILLER_77_1739 ();
 sg13g2_decap_8 FILLER_77_1746 ();
 sg13g2_decap_8 FILLER_77_1753 ();
 sg13g2_decap_8 FILLER_77_1760 ();
 sg13g2_decap_8 FILLER_77_1767 ();
 sg13g2_decap_8 FILLER_77_1774 ();
 sg13g2_decap_8 FILLER_77_1781 ();
 sg13g2_decap_8 FILLER_77_1788 ();
 sg13g2_decap_8 FILLER_77_1795 ();
 sg13g2_decap_8 FILLER_77_1802 ();
 sg13g2_decap_8 FILLER_77_1809 ();
 sg13g2_decap_8 FILLER_77_1816 ();
 sg13g2_decap_8 FILLER_77_1823 ();
 sg13g2_decap_8 FILLER_77_1830 ();
 sg13g2_decap_8 FILLER_77_1837 ();
 sg13g2_decap_8 FILLER_77_1844 ();
 sg13g2_decap_8 FILLER_77_1851 ();
 sg13g2_decap_8 FILLER_77_1858 ();
 sg13g2_decap_8 FILLER_77_1865 ();
 sg13g2_decap_8 FILLER_77_1872 ();
 sg13g2_decap_8 FILLER_77_1879 ();
 sg13g2_decap_8 FILLER_77_1886 ();
 sg13g2_decap_8 FILLER_77_1893 ();
 sg13g2_decap_8 FILLER_77_1900 ();
 sg13g2_decap_8 FILLER_77_1907 ();
 sg13g2_decap_8 FILLER_77_1914 ();
 sg13g2_decap_8 FILLER_77_1921 ();
 sg13g2_decap_8 FILLER_77_1928 ();
 sg13g2_decap_8 FILLER_77_1935 ();
 sg13g2_decap_8 FILLER_77_1942 ();
 sg13g2_decap_8 FILLER_77_1949 ();
 sg13g2_decap_8 FILLER_77_1956 ();
 sg13g2_decap_8 FILLER_77_1963 ();
 sg13g2_decap_8 FILLER_77_1970 ();
 sg13g2_decap_8 FILLER_77_1977 ();
 sg13g2_decap_8 FILLER_77_1984 ();
 sg13g2_decap_8 FILLER_77_1991 ();
 sg13g2_decap_8 FILLER_77_1998 ();
 sg13g2_decap_8 FILLER_77_2005 ();
 sg13g2_decap_8 FILLER_77_2012 ();
 sg13g2_decap_8 FILLER_77_2019 ();
 sg13g2_decap_8 FILLER_77_2026 ();
 sg13g2_decap_4 FILLER_77_2033 ();
 sg13g2_fill_2 FILLER_77_2037 ();
 sg13g2_decap_8 FILLER_77_2069 ();
 sg13g2_decap_8 FILLER_77_2076 ();
 sg13g2_decap_4 FILLER_77_2083 ();
 sg13g2_decap_8 FILLER_77_2091 ();
 sg13g2_decap_8 FILLER_77_2098 ();
 sg13g2_decap_8 FILLER_77_2105 ();
 sg13g2_decap_8 FILLER_77_2112 ();
 sg13g2_decap_8 FILLER_77_2119 ();
 sg13g2_decap_8 FILLER_77_2126 ();
 sg13g2_decap_8 FILLER_77_2137 ();
 sg13g2_decap_8 FILLER_77_2144 ();
 sg13g2_decap_8 FILLER_77_2151 ();
 sg13g2_decap_8 FILLER_77_2188 ();
 sg13g2_decap_8 FILLER_77_2195 ();
 sg13g2_decap_8 FILLER_77_2202 ();
 sg13g2_decap_8 FILLER_77_2209 ();
 sg13g2_decap_8 FILLER_77_2216 ();
 sg13g2_decap_8 FILLER_77_2223 ();
 sg13g2_decap_8 FILLER_77_2230 ();
 sg13g2_decap_8 FILLER_77_2237 ();
 sg13g2_decap_8 FILLER_77_2244 ();
 sg13g2_decap_8 FILLER_77_2251 ();
 sg13g2_decap_8 FILLER_77_2258 ();
 sg13g2_decap_8 FILLER_77_2265 ();
 sg13g2_decap_8 FILLER_77_2272 ();
 sg13g2_decap_8 FILLER_77_2279 ();
 sg13g2_decap_8 FILLER_77_2286 ();
 sg13g2_decap_8 FILLER_77_2293 ();
 sg13g2_decap_8 FILLER_77_2300 ();
 sg13g2_decap_8 FILLER_77_2307 ();
 sg13g2_decap_8 FILLER_77_2314 ();
 sg13g2_decap_8 FILLER_77_2321 ();
 sg13g2_decap_8 FILLER_77_2328 ();
 sg13g2_decap_8 FILLER_77_2335 ();
 sg13g2_decap_8 FILLER_77_2342 ();
 sg13g2_decap_8 FILLER_77_2349 ();
 sg13g2_decap_8 FILLER_77_2356 ();
 sg13g2_decap_8 FILLER_77_2363 ();
 sg13g2_decap_8 FILLER_77_2370 ();
 sg13g2_decap_8 FILLER_77_2377 ();
 sg13g2_decap_8 FILLER_77_2384 ();
 sg13g2_decap_8 FILLER_77_2391 ();
 sg13g2_decap_8 FILLER_77_2398 ();
 sg13g2_decap_8 FILLER_77_2405 ();
 sg13g2_decap_8 FILLER_77_2412 ();
 sg13g2_decap_8 FILLER_77_2419 ();
 sg13g2_decap_8 FILLER_77_2426 ();
 sg13g2_decap_8 FILLER_77_2433 ();
 sg13g2_decap_8 FILLER_77_2440 ();
 sg13g2_decap_8 FILLER_77_2447 ();
 sg13g2_decap_8 FILLER_77_2454 ();
 sg13g2_decap_8 FILLER_77_2461 ();
 sg13g2_decap_8 FILLER_77_2468 ();
 sg13g2_decap_8 FILLER_77_2475 ();
 sg13g2_decap_8 FILLER_77_2482 ();
 sg13g2_decap_8 FILLER_77_2489 ();
 sg13g2_decap_8 FILLER_77_2496 ();
 sg13g2_decap_8 FILLER_77_2503 ();
 sg13g2_decap_8 FILLER_77_2510 ();
 sg13g2_decap_8 FILLER_77_2517 ();
 sg13g2_decap_8 FILLER_77_2524 ();
 sg13g2_decap_8 FILLER_77_2531 ();
 sg13g2_decap_8 FILLER_77_2538 ();
 sg13g2_decap_8 FILLER_77_2545 ();
 sg13g2_decap_8 FILLER_77_2552 ();
 sg13g2_decap_8 FILLER_77_2559 ();
 sg13g2_decap_8 FILLER_77_2566 ();
 sg13g2_decap_8 FILLER_77_2573 ();
 sg13g2_decap_8 FILLER_77_2580 ();
 sg13g2_decap_8 FILLER_77_2587 ();
 sg13g2_decap_8 FILLER_77_2594 ();
 sg13g2_decap_8 FILLER_77_2601 ();
 sg13g2_decap_8 FILLER_77_2608 ();
 sg13g2_decap_8 FILLER_77_2615 ();
 sg13g2_decap_8 FILLER_77_2622 ();
 sg13g2_decap_8 FILLER_77_2629 ();
 sg13g2_decap_8 FILLER_77_2636 ();
 sg13g2_decap_8 FILLER_77_2643 ();
 sg13g2_decap_8 FILLER_77_2650 ();
 sg13g2_decap_8 FILLER_77_2657 ();
 sg13g2_decap_4 FILLER_77_2664 ();
 sg13g2_fill_2 FILLER_77_2668 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_4 FILLER_78_28 ();
 sg13g2_fill_1 FILLER_78_32 ();
 sg13g2_decap_8 FILLER_78_37 ();
 sg13g2_decap_4 FILLER_78_44 ();
 sg13g2_fill_2 FILLER_78_48 ();
 sg13g2_decap_8 FILLER_78_76 ();
 sg13g2_decap_8 FILLER_78_83 ();
 sg13g2_decap_8 FILLER_78_90 ();
 sg13g2_decap_8 FILLER_78_97 ();
 sg13g2_decap_8 FILLER_78_104 ();
 sg13g2_decap_8 FILLER_78_111 ();
 sg13g2_decap_8 FILLER_78_118 ();
 sg13g2_decap_8 FILLER_78_125 ();
 sg13g2_decap_8 FILLER_78_132 ();
 sg13g2_decap_8 FILLER_78_139 ();
 sg13g2_decap_8 FILLER_78_146 ();
 sg13g2_decap_8 FILLER_78_153 ();
 sg13g2_decap_8 FILLER_78_160 ();
 sg13g2_decap_4 FILLER_78_167 ();
 sg13g2_decap_8 FILLER_78_175 ();
 sg13g2_decap_8 FILLER_78_182 ();
 sg13g2_decap_8 FILLER_78_189 ();
 sg13g2_decap_8 FILLER_78_196 ();
 sg13g2_decap_8 FILLER_78_244 ();
 sg13g2_decap_4 FILLER_78_251 ();
 sg13g2_fill_2 FILLER_78_255 ();
 sg13g2_decap_8 FILLER_78_302 ();
 sg13g2_fill_2 FILLER_78_309 ();
 sg13g2_decap_8 FILLER_78_346 ();
 sg13g2_decap_8 FILLER_78_353 ();
 sg13g2_decap_8 FILLER_78_360 ();
 sg13g2_decap_8 FILLER_78_367 ();
 sg13g2_decap_8 FILLER_78_374 ();
 sg13g2_decap_8 FILLER_78_381 ();
 sg13g2_decap_8 FILLER_78_388 ();
 sg13g2_decap_8 FILLER_78_395 ();
 sg13g2_decap_8 FILLER_78_402 ();
 sg13g2_decap_8 FILLER_78_409 ();
 sg13g2_decap_8 FILLER_78_416 ();
 sg13g2_decap_8 FILLER_78_423 ();
 sg13g2_decap_8 FILLER_78_430 ();
 sg13g2_decap_8 FILLER_78_437 ();
 sg13g2_decap_8 FILLER_78_444 ();
 sg13g2_decap_8 FILLER_78_451 ();
 sg13g2_decap_8 FILLER_78_458 ();
 sg13g2_decap_8 FILLER_78_465 ();
 sg13g2_decap_8 FILLER_78_472 ();
 sg13g2_decap_8 FILLER_78_479 ();
 sg13g2_decap_4 FILLER_78_486 ();
 sg13g2_decap_8 FILLER_78_499 ();
 sg13g2_decap_8 FILLER_78_506 ();
 sg13g2_decap_8 FILLER_78_513 ();
 sg13g2_decap_8 FILLER_78_520 ();
 sg13g2_decap_8 FILLER_78_527 ();
 sg13g2_decap_8 FILLER_78_534 ();
 sg13g2_decap_8 FILLER_78_541 ();
 sg13g2_decap_8 FILLER_78_552 ();
 sg13g2_fill_1 FILLER_78_559 ();
 sg13g2_decap_4 FILLER_78_568 ();
 sg13g2_fill_1 FILLER_78_572 ();
 sg13g2_decap_8 FILLER_78_577 ();
 sg13g2_decap_8 FILLER_78_584 ();
 sg13g2_decap_8 FILLER_78_591 ();
 sg13g2_decap_8 FILLER_78_598 ();
 sg13g2_decap_8 FILLER_78_605 ();
 sg13g2_decap_8 FILLER_78_612 ();
 sg13g2_decap_8 FILLER_78_619 ();
 sg13g2_decap_8 FILLER_78_626 ();
 sg13g2_decap_8 FILLER_78_637 ();
 sg13g2_decap_8 FILLER_78_644 ();
 sg13g2_decap_8 FILLER_78_651 ();
 sg13g2_decap_8 FILLER_78_658 ();
 sg13g2_decap_8 FILLER_78_665 ();
 sg13g2_decap_8 FILLER_78_672 ();
 sg13g2_decap_4 FILLER_78_679 ();
 sg13g2_fill_2 FILLER_78_683 ();
 sg13g2_decap_8 FILLER_78_690 ();
 sg13g2_decap_8 FILLER_78_697 ();
 sg13g2_decap_8 FILLER_78_704 ();
 sg13g2_fill_2 FILLER_78_711 ();
 sg13g2_decap_8 FILLER_78_717 ();
 sg13g2_fill_2 FILLER_78_724 ();
 sg13g2_decap_8 FILLER_78_730 ();
 sg13g2_decap_8 FILLER_78_737 ();
 sg13g2_decap_8 FILLER_78_744 ();
 sg13g2_decap_8 FILLER_78_751 ();
 sg13g2_decap_8 FILLER_78_758 ();
 sg13g2_decap_8 FILLER_78_765 ();
 sg13g2_decap_8 FILLER_78_772 ();
 sg13g2_decap_4 FILLER_78_779 ();
 sg13g2_decap_8 FILLER_78_792 ();
 sg13g2_decap_8 FILLER_78_799 ();
 sg13g2_decap_8 FILLER_78_806 ();
 sg13g2_decap_8 FILLER_78_813 ();
 sg13g2_decap_8 FILLER_78_820 ();
 sg13g2_decap_8 FILLER_78_827 ();
 sg13g2_decap_8 FILLER_78_834 ();
 sg13g2_decap_8 FILLER_78_841 ();
 sg13g2_decap_8 FILLER_78_848 ();
 sg13g2_decap_8 FILLER_78_855 ();
 sg13g2_decap_8 FILLER_78_862 ();
 sg13g2_decap_8 FILLER_78_869 ();
 sg13g2_decap_8 FILLER_78_876 ();
 sg13g2_decap_8 FILLER_78_883 ();
 sg13g2_decap_8 FILLER_78_890 ();
 sg13g2_decap_8 FILLER_78_897 ();
 sg13g2_fill_2 FILLER_78_904 ();
 sg13g2_decap_8 FILLER_78_914 ();
 sg13g2_decap_8 FILLER_78_921 ();
 sg13g2_decap_8 FILLER_78_928 ();
 sg13g2_decap_8 FILLER_78_935 ();
 sg13g2_decap_8 FILLER_78_942 ();
 sg13g2_fill_2 FILLER_78_949 ();
 sg13g2_fill_1 FILLER_78_951 ();
 sg13g2_decap_4 FILLER_78_956 ();
 sg13g2_fill_1 FILLER_78_960 ();
 sg13g2_decap_8 FILLER_78_980 ();
 sg13g2_decap_8 FILLER_78_987 ();
 sg13g2_decap_8 FILLER_78_994 ();
 sg13g2_decap_8 FILLER_78_1001 ();
 sg13g2_decap_8 FILLER_78_1008 ();
 sg13g2_decap_8 FILLER_78_1015 ();
 sg13g2_decap_8 FILLER_78_1022 ();
 sg13g2_decap_8 FILLER_78_1029 ();
 sg13g2_fill_2 FILLER_78_1036 ();
 sg13g2_decap_4 FILLER_78_1042 ();
 sg13g2_decap_8 FILLER_78_1054 ();
 sg13g2_decap_8 FILLER_78_1061 ();
 sg13g2_decap_8 FILLER_78_1068 ();
 sg13g2_decap_8 FILLER_78_1075 ();
 sg13g2_decap_8 FILLER_78_1082 ();
 sg13g2_decap_8 FILLER_78_1089 ();
 sg13g2_decap_8 FILLER_78_1096 ();
 sg13g2_decap_8 FILLER_78_1103 ();
 sg13g2_fill_2 FILLER_78_1110 ();
 sg13g2_decap_8 FILLER_78_1116 ();
 sg13g2_decap_8 FILLER_78_1123 ();
 sg13g2_decap_8 FILLER_78_1130 ();
 sg13g2_decap_8 FILLER_78_1137 ();
 sg13g2_fill_1 FILLER_78_1144 ();
 sg13g2_decap_8 FILLER_78_1149 ();
 sg13g2_decap_8 FILLER_78_1156 ();
 sg13g2_decap_8 FILLER_78_1163 ();
 sg13g2_decap_8 FILLER_78_1170 ();
 sg13g2_decap_8 FILLER_78_1177 ();
 sg13g2_decap_8 FILLER_78_1184 ();
 sg13g2_decap_8 FILLER_78_1191 ();
 sg13g2_decap_8 FILLER_78_1203 ();
 sg13g2_decap_4 FILLER_78_1210 ();
 sg13g2_fill_1 FILLER_78_1214 ();
 sg13g2_decap_8 FILLER_78_1219 ();
 sg13g2_decap_8 FILLER_78_1226 ();
 sg13g2_decap_8 FILLER_78_1233 ();
 sg13g2_decap_8 FILLER_78_1240 ();
 sg13g2_decap_8 FILLER_78_1247 ();
 sg13g2_fill_1 FILLER_78_1254 ();
 sg13g2_decap_8 FILLER_78_1265 ();
 sg13g2_decap_4 FILLER_78_1272 ();
 sg13g2_fill_1 FILLER_78_1286 ();
 sg13g2_decap_8 FILLER_78_1298 ();
 sg13g2_decap_8 FILLER_78_1305 ();
 sg13g2_decap_8 FILLER_78_1312 ();
 sg13g2_decap_8 FILLER_78_1319 ();
 sg13g2_decap_8 FILLER_78_1326 ();
 sg13g2_decap_8 FILLER_78_1333 ();
 sg13g2_decap_8 FILLER_78_1340 ();
 sg13g2_decap_8 FILLER_78_1347 ();
 sg13g2_decap_8 FILLER_78_1354 ();
 sg13g2_decap_8 FILLER_78_1361 ();
 sg13g2_decap_8 FILLER_78_1368 ();
 sg13g2_decap_8 FILLER_78_1375 ();
 sg13g2_decap_8 FILLER_78_1382 ();
 sg13g2_fill_2 FILLER_78_1389 ();
 sg13g2_decap_8 FILLER_78_1395 ();
 sg13g2_decap_8 FILLER_78_1402 ();
 sg13g2_decap_8 FILLER_78_1409 ();
 sg13g2_decap_8 FILLER_78_1416 ();
 sg13g2_decap_8 FILLER_78_1427 ();
 sg13g2_decap_8 FILLER_78_1434 ();
 sg13g2_decap_8 FILLER_78_1441 ();
 sg13g2_decap_8 FILLER_78_1448 ();
 sg13g2_decap_8 FILLER_78_1455 ();
 sg13g2_decap_8 FILLER_78_1462 ();
 sg13g2_decap_8 FILLER_78_1469 ();
 sg13g2_decap_8 FILLER_78_1476 ();
 sg13g2_decap_8 FILLER_78_1483 ();
 sg13g2_fill_1 FILLER_78_1490 ();
 sg13g2_decap_8 FILLER_78_1495 ();
 sg13g2_decap_8 FILLER_78_1502 ();
 sg13g2_decap_8 FILLER_78_1509 ();
 sg13g2_decap_8 FILLER_78_1516 ();
 sg13g2_decap_8 FILLER_78_1523 ();
 sg13g2_decap_8 FILLER_78_1530 ();
 sg13g2_decap_8 FILLER_78_1537 ();
 sg13g2_decap_8 FILLER_78_1544 ();
 sg13g2_decap_8 FILLER_78_1551 ();
 sg13g2_fill_2 FILLER_78_1558 ();
 sg13g2_fill_1 FILLER_78_1560 ();
 sg13g2_decap_8 FILLER_78_1578 ();
 sg13g2_decap_8 FILLER_78_1585 ();
 sg13g2_decap_8 FILLER_78_1592 ();
 sg13g2_decap_8 FILLER_78_1599 ();
 sg13g2_decap_8 FILLER_78_1606 ();
 sg13g2_decap_8 FILLER_78_1613 ();
 sg13g2_decap_8 FILLER_78_1620 ();
 sg13g2_decap_8 FILLER_78_1627 ();
 sg13g2_decap_8 FILLER_78_1634 ();
 sg13g2_decap_8 FILLER_78_1641 ();
 sg13g2_fill_2 FILLER_78_1648 ();
 sg13g2_fill_1 FILLER_78_1650 ();
 sg13g2_decap_8 FILLER_78_1659 ();
 sg13g2_decap_8 FILLER_78_1666 ();
 sg13g2_decap_8 FILLER_78_1673 ();
 sg13g2_fill_2 FILLER_78_1680 ();
 sg13g2_fill_1 FILLER_78_1682 ();
 sg13g2_decap_8 FILLER_78_1696 ();
 sg13g2_decap_8 FILLER_78_1703 ();
 sg13g2_decap_8 FILLER_78_1710 ();
 sg13g2_decap_8 FILLER_78_1717 ();
 sg13g2_decap_8 FILLER_78_1724 ();
 sg13g2_decap_8 FILLER_78_1731 ();
 sg13g2_decap_8 FILLER_78_1738 ();
 sg13g2_decap_8 FILLER_78_1745 ();
 sg13g2_decap_8 FILLER_78_1752 ();
 sg13g2_decap_8 FILLER_78_1759 ();
 sg13g2_decap_8 FILLER_78_1766 ();
 sg13g2_decap_8 FILLER_78_1773 ();
 sg13g2_decap_8 FILLER_78_1780 ();
 sg13g2_decap_8 FILLER_78_1787 ();
 sg13g2_decap_8 FILLER_78_1794 ();
 sg13g2_decap_8 FILLER_78_1801 ();
 sg13g2_decap_8 FILLER_78_1808 ();
 sg13g2_decap_8 FILLER_78_1815 ();
 sg13g2_decap_8 FILLER_78_1822 ();
 sg13g2_decap_8 FILLER_78_1829 ();
 sg13g2_decap_8 FILLER_78_1836 ();
 sg13g2_decap_8 FILLER_78_1843 ();
 sg13g2_decap_8 FILLER_78_1850 ();
 sg13g2_decap_8 FILLER_78_1857 ();
 sg13g2_decap_8 FILLER_78_1864 ();
 sg13g2_decap_8 FILLER_78_1871 ();
 sg13g2_decap_8 FILLER_78_1878 ();
 sg13g2_decap_8 FILLER_78_1885 ();
 sg13g2_decap_8 FILLER_78_1892 ();
 sg13g2_decap_8 FILLER_78_1899 ();
 sg13g2_decap_8 FILLER_78_1906 ();
 sg13g2_decap_8 FILLER_78_1913 ();
 sg13g2_decap_8 FILLER_78_1920 ();
 sg13g2_decap_8 FILLER_78_1927 ();
 sg13g2_decap_8 FILLER_78_1934 ();
 sg13g2_decap_8 FILLER_78_1941 ();
 sg13g2_decap_8 FILLER_78_1948 ();
 sg13g2_decap_8 FILLER_78_1955 ();
 sg13g2_decap_8 FILLER_78_1962 ();
 sg13g2_decap_8 FILLER_78_1969 ();
 sg13g2_decap_8 FILLER_78_1976 ();
 sg13g2_decap_8 FILLER_78_1983 ();
 sg13g2_decap_8 FILLER_78_1990 ();
 sg13g2_decap_8 FILLER_78_1997 ();
 sg13g2_decap_8 FILLER_78_2004 ();
 sg13g2_decap_8 FILLER_78_2011 ();
 sg13g2_decap_8 FILLER_78_2018 ();
 sg13g2_decap_8 FILLER_78_2025 ();
 sg13g2_decap_8 FILLER_78_2032 ();
 sg13g2_decap_8 FILLER_78_2039 ();
 sg13g2_decap_8 FILLER_78_2046 ();
 sg13g2_decap_8 FILLER_78_2053 ();
 sg13g2_decap_8 FILLER_78_2060 ();
 sg13g2_decap_8 FILLER_78_2067 ();
 sg13g2_decap_8 FILLER_78_2074 ();
 sg13g2_decap_8 FILLER_78_2107 ();
 sg13g2_decap_8 FILLER_78_2114 ();
 sg13g2_decap_4 FILLER_78_2121 ();
 sg13g2_fill_1 FILLER_78_2125 ();
 sg13g2_decap_8 FILLER_78_2152 ();
 sg13g2_decap_8 FILLER_78_2159 ();
 sg13g2_decap_8 FILLER_78_2166 ();
 sg13g2_decap_8 FILLER_78_2173 ();
 sg13g2_decap_8 FILLER_78_2180 ();
 sg13g2_decap_8 FILLER_78_2187 ();
 sg13g2_decap_8 FILLER_78_2194 ();
 sg13g2_decap_8 FILLER_78_2201 ();
 sg13g2_decap_8 FILLER_78_2208 ();
 sg13g2_decap_8 FILLER_78_2215 ();
 sg13g2_decap_8 FILLER_78_2222 ();
 sg13g2_decap_8 FILLER_78_2229 ();
 sg13g2_decap_8 FILLER_78_2236 ();
 sg13g2_decap_8 FILLER_78_2243 ();
 sg13g2_decap_8 FILLER_78_2250 ();
 sg13g2_decap_8 FILLER_78_2257 ();
 sg13g2_decap_8 FILLER_78_2264 ();
 sg13g2_decap_8 FILLER_78_2271 ();
 sg13g2_decap_8 FILLER_78_2278 ();
 sg13g2_decap_8 FILLER_78_2285 ();
 sg13g2_decap_8 FILLER_78_2292 ();
 sg13g2_decap_8 FILLER_78_2299 ();
 sg13g2_decap_8 FILLER_78_2306 ();
 sg13g2_decap_8 FILLER_78_2313 ();
 sg13g2_decap_8 FILLER_78_2320 ();
 sg13g2_decap_8 FILLER_78_2327 ();
 sg13g2_decap_8 FILLER_78_2334 ();
 sg13g2_decap_8 FILLER_78_2341 ();
 sg13g2_decap_8 FILLER_78_2348 ();
 sg13g2_decap_8 FILLER_78_2355 ();
 sg13g2_decap_8 FILLER_78_2362 ();
 sg13g2_decap_8 FILLER_78_2369 ();
 sg13g2_decap_8 FILLER_78_2376 ();
 sg13g2_decap_8 FILLER_78_2383 ();
 sg13g2_decap_8 FILLER_78_2390 ();
 sg13g2_decap_8 FILLER_78_2397 ();
 sg13g2_decap_8 FILLER_78_2404 ();
 sg13g2_decap_8 FILLER_78_2411 ();
 sg13g2_decap_8 FILLER_78_2418 ();
 sg13g2_decap_8 FILLER_78_2425 ();
 sg13g2_decap_8 FILLER_78_2432 ();
 sg13g2_decap_8 FILLER_78_2439 ();
 sg13g2_decap_8 FILLER_78_2446 ();
 sg13g2_decap_8 FILLER_78_2453 ();
 sg13g2_decap_8 FILLER_78_2460 ();
 sg13g2_decap_8 FILLER_78_2467 ();
 sg13g2_decap_8 FILLER_78_2474 ();
 sg13g2_decap_8 FILLER_78_2481 ();
 sg13g2_decap_8 FILLER_78_2488 ();
 sg13g2_decap_8 FILLER_78_2495 ();
 sg13g2_decap_8 FILLER_78_2502 ();
 sg13g2_decap_8 FILLER_78_2509 ();
 sg13g2_decap_8 FILLER_78_2516 ();
 sg13g2_decap_8 FILLER_78_2523 ();
 sg13g2_decap_8 FILLER_78_2530 ();
 sg13g2_decap_8 FILLER_78_2537 ();
 sg13g2_decap_8 FILLER_78_2544 ();
 sg13g2_decap_8 FILLER_78_2551 ();
 sg13g2_decap_8 FILLER_78_2558 ();
 sg13g2_decap_8 FILLER_78_2565 ();
 sg13g2_decap_8 FILLER_78_2572 ();
 sg13g2_decap_8 FILLER_78_2579 ();
 sg13g2_decap_8 FILLER_78_2586 ();
 sg13g2_decap_8 FILLER_78_2593 ();
 sg13g2_decap_8 FILLER_78_2600 ();
 sg13g2_decap_8 FILLER_78_2607 ();
 sg13g2_decap_8 FILLER_78_2614 ();
 sg13g2_decap_8 FILLER_78_2621 ();
 sg13g2_decap_8 FILLER_78_2628 ();
 sg13g2_decap_8 FILLER_78_2635 ();
 sg13g2_decap_8 FILLER_78_2642 ();
 sg13g2_decap_8 FILLER_78_2649 ();
 sg13g2_decap_8 FILLER_78_2656 ();
 sg13g2_decap_8 FILLER_78_2663 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_4 FILLER_79_84 ();
 sg13g2_fill_1 FILLER_79_88 ();
 sg13g2_decap_8 FILLER_79_93 ();
 sg13g2_fill_2 FILLER_79_100 ();
 sg13g2_decap_8 FILLER_79_106 ();
 sg13g2_decap_8 FILLER_79_113 ();
 sg13g2_decap_8 FILLER_79_120 ();
 sg13g2_decap_8 FILLER_79_127 ();
 sg13g2_decap_8 FILLER_79_134 ();
 sg13g2_decap_4 FILLER_79_141 ();
 sg13g2_fill_2 FILLER_79_145 ();
 sg13g2_decap_8 FILLER_79_151 ();
 sg13g2_decap_8 FILLER_79_158 ();
 sg13g2_decap_8 FILLER_79_165 ();
 sg13g2_decap_8 FILLER_79_172 ();
 sg13g2_decap_8 FILLER_79_179 ();
 sg13g2_decap_8 FILLER_79_186 ();
 sg13g2_decap_8 FILLER_79_193 ();
 sg13g2_decap_8 FILLER_79_200 ();
 sg13g2_decap_8 FILLER_79_207 ();
 sg13g2_decap_8 FILLER_79_214 ();
 sg13g2_fill_2 FILLER_79_221 ();
 sg13g2_fill_1 FILLER_79_223 ();
 sg13g2_decap_8 FILLER_79_228 ();
 sg13g2_decap_8 FILLER_79_235 ();
 sg13g2_decap_8 FILLER_79_242 ();
 sg13g2_decap_8 FILLER_79_249 ();
 sg13g2_decap_8 FILLER_79_256 ();
 sg13g2_decap_8 FILLER_79_263 ();
 sg13g2_decap_8 FILLER_79_270 ();
 sg13g2_decap_8 FILLER_79_277 ();
 sg13g2_decap_8 FILLER_79_284 ();
 sg13g2_decap_8 FILLER_79_291 ();
 sg13g2_decap_8 FILLER_79_298 ();
 sg13g2_decap_8 FILLER_79_305 ();
 sg13g2_decap_8 FILLER_79_312 ();
 sg13g2_decap_4 FILLER_79_319 ();
 sg13g2_fill_2 FILLER_79_323 ();
 sg13g2_decap_8 FILLER_79_329 ();
 sg13g2_decap_4 FILLER_79_336 ();
 sg13g2_fill_2 FILLER_79_340 ();
 sg13g2_decap_8 FILLER_79_346 ();
 sg13g2_decap_8 FILLER_79_353 ();
 sg13g2_decap_8 FILLER_79_360 ();
 sg13g2_decap_8 FILLER_79_367 ();
 sg13g2_decap_8 FILLER_79_374 ();
 sg13g2_decap_8 FILLER_79_381 ();
 sg13g2_decap_8 FILLER_79_388 ();
 sg13g2_decap_8 FILLER_79_395 ();
 sg13g2_decap_8 FILLER_79_402 ();
 sg13g2_decap_8 FILLER_79_409 ();
 sg13g2_decap_8 FILLER_79_416 ();
 sg13g2_decap_8 FILLER_79_423 ();
 sg13g2_decap_8 FILLER_79_430 ();
 sg13g2_decap_8 FILLER_79_437 ();
 sg13g2_decap_8 FILLER_79_444 ();
 sg13g2_decap_8 FILLER_79_451 ();
 sg13g2_decap_8 FILLER_79_458 ();
 sg13g2_decap_8 FILLER_79_465 ();
 sg13g2_decap_8 FILLER_79_472 ();
 sg13g2_decap_8 FILLER_79_479 ();
 sg13g2_decap_8 FILLER_79_486 ();
 sg13g2_decap_8 FILLER_79_493 ();
 sg13g2_decap_8 FILLER_79_500 ();
 sg13g2_decap_8 FILLER_79_507 ();
 sg13g2_decap_8 FILLER_79_514 ();
 sg13g2_decap_8 FILLER_79_521 ();
 sg13g2_decap_8 FILLER_79_528 ();
 sg13g2_decap_8 FILLER_79_535 ();
 sg13g2_decap_8 FILLER_79_542 ();
 sg13g2_decap_8 FILLER_79_549 ();
 sg13g2_decap_8 FILLER_79_556 ();
 sg13g2_decap_8 FILLER_79_563 ();
 sg13g2_decap_8 FILLER_79_570 ();
 sg13g2_decap_8 FILLER_79_577 ();
 sg13g2_decap_8 FILLER_79_584 ();
 sg13g2_decap_8 FILLER_79_591 ();
 sg13g2_decap_8 FILLER_79_598 ();
 sg13g2_decap_8 FILLER_79_605 ();
 sg13g2_decap_8 FILLER_79_612 ();
 sg13g2_decap_8 FILLER_79_619 ();
 sg13g2_decap_8 FILLER_79_626 ();
 sg13g2_decap_8 FILLER_79_633 ();
 sg13g2_decap_8 FILLER_79_640 ();
 sg13g2_decap_8 FILLER_79_647 ();
 sg13g2_decap_8 FILLER_79_654 ();
 sg13g2_decap_8 FILLER_79_661 ();
 sg13g2_decap_8 FILLER_79_668 ();
 sg13g2_decap_8 FILLER_79_675 ();
 sg13g2_decap_8 FILLER_79_682 ();
 sg13g2_decap_8 FILLER_79_689 ();
 sg13g2_decap_8 FILLER_79_696 ();
 sg13g2_decap_8 FILLER_79_703 ();
 sg13g2_decap_8 FILLER_79_710 ();
 sg13g2_decap_8 FILLER_79_717 ();
 sg13g2_decap_8 FILLER_79_724 ();
 sg13g2_decap_8 FILLER_79_731 ();
 sg13g2_decap_8 FILLER_79_738 ();
 sg13g2_decap_8 FILLER_79_745 ();
 sg13g2_decap_8 FILLER_79_752 ();
 sg13g2_decap_8 FILLER_79_759 ();
 sg13g2_decap_8 FILLER_79_766 ();
 sg13g2_decap_8 FILLER_79_773 ();
 sg13g2_decap_8 FILLER_79_780 ();
 sg13g2_decap_8 FILLER_79_787 ();
 sg13g2_decap_8 FILLER_79_794 ();
 sg13g2_decap_8 FILLER_79_801 ();
 sg13g2_decap_8 FILLER_79_808 ();
 sg13g2_decap_8 FILLER_79_815 ();
 sg13g2_decap_8 FILLER_79_822 ();
 sg13g2_decap_8 FILLER_79_829 ();
 sg13g2_decap_8 FILLER_79_836 ();
 sg13g2_decap_8 FILLER_79_843 ();
 sg13g2_decap_8 FILLER_79_850 ();
 sg13g2_decap_8 FILLER_79_857 ();
 sg13g2_decap_8 FILLER_79_864 ();
 sg13g2_decap_8 FILLER_79_871 ();
 sg13g2_decap_8 FILLER_79_878 ();
 sg13g2_decap_8 FILLER_79_885 ();
 sg13g2_decap_8 FILLER_79_892 ();
 sg13g2_decap_8 FILLER_79_899 ();
 sg13g2_decap_8 FILLER_79_906 ();
 sg13g2_decap_8 FILLER_79_913 ();
 sg13g2_decap_8 FILLER_79_920 ();
 sg13g2_decap_8 FILLER_79_927 ();
 sg13g2_decap_8 FILLER_79_934 ();
 sg13g2_decap_8 FILLER_79_941 ();
 sg13g2_decap_8 FILLER_79_948 ();
 sg13g2_decap_8 FILLER_79_955 ();
 sg13g2_decap_8 FILLER_79_962 ();
 sg13g2_decap_8 FILLER_79_969 ();
 sg13g2_decap_8 FILLER_79_976 ();
 sg13g2_decap_8 FILLER_79_983 ();
 sg13g2_decap_8 FILLER_79_990 ();
 sg13g2_decap_8 FILLER_79_997 ();
 sg13g2_decap_8 FILLER_79_1004 ();
 sg13g2_decap_8 FILLER_79_1011 ();
 sg13g2_decap_8 FILLER_79_1018 ();
 sg13g2_decap_8 FILLER_79_1025 ();
 sg13g2_decap_8 FILLER_79_1032 ();
 sg13g2_decap_8 FILLER_79_1039 ();
 sg13g2_decap_8 FILLER_79_1046 ();
 sg13g2_decap_8 FILLER_79_1053 ();
 sg13g2_decap_8 FILLER_79_1060 ();
 sg13g2_decap_8 FILLER_79_1067 ();
 sg13g2_decap_8 FILLER_79_1074 ();
 sg13g2_decap_8 FILLER_79_1081 ();
 sg13g2_decap_8 FILLER_79_1088 ();
 sg13g2_decap_8 FILLER_79_1095 ();
 sg13g2_decap_8 FILLER_79_1102 ();
 sg13g2_decap_8 FILLER_79_1109 ();
 sg13g2_decap_8 FILLER_79_1116 ();
 sg13g2_decap_8 FILLER_79_1123 ();
 sg13g2_decap_8 FILLER_79_1130 ();
 sg13g2_decap_8 FILLER_79_1137 ();
 sg13g2_decap_8 FILLER_79_1144 ();
 sg13g2_decap_8 FILLER_79_1151 ();
 sg13g2_decap_8 FILLER_79_1158 ();
 sg13g2_decap_8 FILLER_79_1165 ();
 sg13g2_decap_8 FILLER_79_1172 ();
 sg13g2_decap_8 FILLER_79_1179 ();
 sg13g2_decap_8 FILLER_79_1186 ();
 sg13g2_decap_8 FILLER_79_1193 ();
 sg13g2_decap_8 FILLER_79_1200 ();
 sg13g2_decap_8 FILLER_79_1207 ();
 sg13g2_decap_8 FILLER_79_1214 ();
 sg13g2_decap_8 FILLER_79_1221 ();
 sg13g2_decap_8 FILLER_79_1228 ();
 sg13g2_decap_8 FILLER_79_1235 ();
 sg13g2_decap_8 FILLER_79_1242 ();
 sg13g2_decap_8 FILLER_79_1249 ();
 sg13g2_fill_2 FILLER_79_1256 ();
 sg13g2_decap_8 FILLER_79_1261 ();
 sg13g2_decap_8 FILLER_79_1268 ();
 sg13g2_decap_8 FILLER_79_1275 ();
 sg13g2_decap_4 FILLER_79_1282 ();
 sg13g2_fill_1 FILLER_79_1286 ();
 sg13g2_decap_8 FILLER_79_1299 ();
 sg13g2_decap_8 FILLER_79_1306 ();
 sg13g2_decap_8 FILLER_79_1313 ();
 sg13g2_decap_8 FILLER_79_1320 ();
 sg13g2_decap_8 FILLER_79_1327 ();
 sg13g2_decap_8 FILLER_79_1334 ();
 sg13g2_decap_8 FILLER_79_1341 ();
 sg13g2_decap_8 FILLER_79_1348 ();
 sg13g2_decap_8 FILLER_79_1355 ();
 sg13g2_decap_8 FILLER_79_1362 ();
 sg13g2_decap_8 FILLER_79_1369 ();
 sg13g2_decap_8 FILLER_79_1376 ();
 sg13g2_decap_8 FILLER_79_1383 ();
 sg13g2_decap_8 FILLER_79_1390 ();
 sg13g2_decap_8 FILLER_79_1397 ();
 sg13g2_decap_8 FILLER_79_1404 ();
 sg13g2_decap_8 FILLER_79_1411 ();
 sg13g2_decap_8 FILLER_79_1418 ();
 sg13g2_decap_8 FILLER_79_1425 ();
 sg13g2_decap_8 FILLER_79_1432 ();
 sg13g2_decap_8 FILLER_79_1439 ();
 sg13g2_decap_8 FILLER_79_1446 ();
 sg13g2_decap_8 FILLER_79_1453 ();
 sg13g2_decap_8 FILLER_79_1460 ();
 sg13g2_decap_8 FILLER_79_1467 ();
 sg13g2_decap_8 FILLER_79_1474 ();
 sg13g2_decap_8 FILLER_79_1481 ();
 sg13g2_decap_8 FILLER_79_1488 ();
 sg13g2_decap_8 FILLER_79_1495 ();
 sg13g2_decap_8 FILLER_79_1502 ();
 sg13g2_decap_8 FILLER_79_1509 ();
 sg13g2_decap_8 FILLER_79_1516 ();
 sg13g2_decap_8 FILLER_79_1523 ();
 sg13g2_decap_8 FILLER_79_1530 ();
 sg13g2_decap_8 FILLER_79_1537 ();
 sg13g2_decap_8 FILLER_79_1544 ();
 sg13g2_decap_8 FILLER_79_1551 ();
 sg13g2_decap_4 FILLER_79_1558 ();
 sg13g2_fill_2 FILLER_79_1562 ();
 sg13g2_decap_8 FILLER_79_1570 ();
 sg13g2_decap_8 FILLER_79_1577 ();
 sg13g2_decap_8 FILLER_79_1584 ();
 sg13g2_decap_8 FILLER_79_1591 ();
 sg13g2_decap_8 FILLER_79_1598 ();
 sg13g2_decap_8 FILLER_79_1605 ();
 sg13g2_decap_8 FILLER_79_1612 ();
 sg13g2_decap_8 FILLER_79_1619 ();
 sg13g2_decap_8 FILLER_79_1626 ();
 sg13g2_decap_8 FILLER_79_1633 ();
 sg13g2_decap_8 FILLER_79_1640 ();
 sg13g2_decap_8 FILLER_79_1647 ();
 sg13g2_decap_8 FILLER_79_1654 ();
 sg13g2_decap_8 FILLER_79_1661 ();
 sg13g2_decap_8 FILLER_79_1668 ();
 sg13g2_decap_8 FILLER_79_1675 ();
 sg13g2_decap_8 FILLER_79_1682 ();
 sg13g2_decap_8 FILLER_79_1689 ();
 sg13g2_decap_8 FILLER_79_1696 ();
 sg13g2_decap_8 FILLER_79_1703 ();
 sg13g2_decap_8 FILLER_79_1710 ();
 sg13g2_decap_8 FILLER_79_1717 ();
 sg13g2_decap_8 FILLER_79_1724 ();
 sg13g2_decap_8 FILLER_79_1731 ();
 sg13g2_decap_8 FILLER_79_1738 ();
 sg13g2_decap_8 FILLER_79_1745 ();
 sg13g2_decap_8 FILLER_79_1752 ();
 sg13g2_decap_8 FILLER_79_1759 ();
 sg13g2_decap_8 FILLER_79_1766 ();
 sg13g2_decap_8 FILLER_79_1773 ();
 sg13g2_decap_8 FILLER_79_1780 ();
 sg13g2_decap_8 FILLER_79_1787 ();
 sg13g2_decap_8 FILLER_79_1794 ();
 sg13g2_decap_8 FILLER_79_1801 ();
 sg13g2_decap_8 FILLER_79_1808 ();
 sg13g2_decap_8 FILLER_79_1815 ();
 sg13g2_decap_8 FILLER_79_1822 ();
 sg13g2_decap_8 FILLER_79_1829 ();
 sg13g2_decap_8 FILLER_79_1836 ();
 sg13g2_decap_8 FILLER_79_1843 ();
 sg13g2_decap_8 FILLER_79_1850 ();
 sg13g2_decap_8 FILLER_79_1857 ();
 sg13g2_decap_8 FILLER_79_1864 ();
 sg13g2_decap_8 FILLER_79_1871 ();
 sg13g2_decap_8 FILLER_79_1878 ();
 sg13g2_decap_8 FILLER_79_1885 ();
 sg13g2_decap_8 FILLER_79_1892 ();
 sg13g2_decap_8 FILLER_79_1899 ();
 sg13g2_decap_8 FILLER_79_1906 ();
 sg13g2_decap_8 FILLER_79_1913 ();
 sg13g2_decap_8 FILLER_79_1920 ();
 sg13g2_decap_8 FILLER_79_1927 ();
 sg13g2_decap_8 FILLER_79_1934 ();
 sg13g2_decap_8 FILLER_79_1941 ();
 sg13g2_decap_8 FILLER_79_1948 ();
 sg13g2_decap_8 FILLER_79_1955 ();
 sg13g2_decap_8 FILLER_79_1962 ();
 sg13g2_decap_8 FILLER_79_1969 ();
 sg13g2_decap_8 FILLER_79_1976 ();
 sg13g2_decap_8 FILLER_79_1983 ();
 sg13g2_decap_8 FILLER_79_1990 ();
 sg13g2_decap_8 FILLER_79_1997 ();
 sg13g2_decap_8 FILLER_79_2004 ();
 sg13g2_decap_8 FILLER_79_2011 ();
 sg13g2_decap_8 FILLER_79_2018 ();
 sg13g2_decap_8 FILLER_79_2025 ();
 sg13g2_decap_8 FILLER_79_2032 ();
 sg13g2_decap_8 FILLER_79_2039 ();
 sg13g2_decap_8 FILLER_79_2046 ();
 sg13g2_decap_8 FILLER_79_2053 ();
 sg13g2_decap_8 FILLER_79_2060 ();
 sg13g2_decap_8 FILLER_79_2067 ();
 sg13g2_decap_8 FILLER_79_2074 ();
 sg13g2_decap_8 FILLER_79_2081 ();
 sg13g2_decap_8 FILLER_79_2088 ();
 sg13g2_decap_8 FILLER_79_2095 ();
 sg13g2_decap_8 FILLER_79_2102 ();
 sg13g2_decap_8 FILLER_79_2109 ();
 sg13g2_decap_8 FILLER_79_2116 ();
 sg13g2_decap_8 FILLER_79_2123 ();
 sg13g2_decap_8 FILLER_79_2130 ();
 sg13g2_decap_8 FILLER_79_2137 ();
 sg13g2_decap_8 FILLER_79_2144 ();
 sg13g2_decap_8 FILLER_79_2151 ();
 sg13g2_decap_8 FILLER_79_2158 ();
 sg13g2_decap_8 FILLER_79_2165 ();
 sg13g2_decap_8 FILLER_79_2172 ();
 sg13g2_decap_8 FILLER_79_2179 ();
 sg13g2_decap_8 FILLER_79_2186 ();
 sg13g2_decap_8 FILLER_79_2193 ();
 sg13g2_decap_8 FILLER_79_2200 ();
 sg13g2_decap_8 FILLER_79_2207 ();
 sg13g2_decap_8 FILLER_79_2214 ();
 sg13g2_decap_8 FILLER_79_2221 ();
 sg13g2_decap_8 FILLER_79_2228 ();
 sg13g2_decap_8 FILLER_79_2235 ();
 sg13g2_decap_8 FILLER_79_2242 ();
 sg13g2_decap_8 FILLER_79_2249 ();
 sg13g2_decap_8 FILLER_79_2256 ();
 sg13g2_decap_8 FILLER_79_2263 ();
 sg13g2_decap_8 FILLER_79_2270 ();
 sg13g2_decap_8 FILLER_79_2277 ();
 sg13g2_decap_8 FILLER_79_2284 ();
 sg13g2_decap_8 FILLER_79_2291 ();
 sg13g2_decap_8 FILLER_79_2298 ();
 sg13g2_decap_8 FILLER_79_2305 ();
 sg13g2_decap_8 FILLER_79_2312 ();
 sg13g2_decap_8 FILLER_79_2319 ();
 sg13g2_decap_8 FILLER_79_2326 ();
 sg13g2_decap_8 FILLER_79_2333 ();
 sg13g2_decap_8 FILLER_79_2340 ();
 sg13g2_decap_8 FILLER_79_2347 ();
 sg13g2_decap_8 FILLER_79_2354 ();
 sg13g2_decap_8 FILLER_79_2361 ();
 sg13g2_decap_8 FILLER_79_2368 ();
 sg13g2_decap_8 FILLER_79_2375 ();
 sg13g2_decap_8 FILLER_79_2382 ();
 sg13g2_decap_8 FILLER_79_2389 ();
 sg13g2_decap_8 FILLER_79_2396 ();
 sg13g2_decap_8 FILLER_79_2403 ();
 sg13g2_decap_8 FILLER_79_2410 ();
 sg13g2_decap_8 FILLER_79_2417 ();
 sg13g2_decap_8 FILLER_79_2424 ();
 sg13g2_decap_8 FILLER_79_2431 ();
 sg13g2_decap_8 FILLER_79_2438 ();
 sg13g2_decap_8 FILLER_79_2445 ();
 sg13g2_decap_8 FILLER_79_2452 ();
 sg13g2_decap_8 FILLER_79_2459 ();
 sg13g2_decap_8 FILLER_79_2466 ();
 sg13g2_decap_8 FILLER_79_2473 ();
 sg13g2_decap_8 FILLER_79_2480 ();
 sg13g2_decap_8 FILLER_79_2487 ();
 sg13g2_decap_8 FILLER_79_2494 ();
 sg13g2_decap_8 FILLER_79_2501 ();
 sg13g2_decap_8 FILLER_79_2508 ();
 sg13g2_decap_8 FILLER_79_2515 ();
 sg13g2_decap_8 FILLER_79_2522 ();
 sg13g2_decap_8 FILLER_79_2529 ();
 sg13g2_decap_8 FILLER_79_2536 ();
 sg13g2_decap_8 FILLER_79_2543 ();
 sg13g2_decap_8 FILLER_79_2550 ();
 sg13g2_decap_8 FILLER_79_2557 ();
 sg13g2_decap_8 FILLER_79_2564 ();
 sg13g2_decap_8 FILLER_79_2571 ();
 sg13g2_decap_8 FILLER_79_2578 ();
 sg13g2_decap_8 FILLER_79_2585 ();
 sg13g2_decap_8 FILLER_79_2592 ();
 sg13g2_decap_8 FILLER_79_2599 ();
 sg13g2_decap_8 FILLER_79_2606 ();
 sg13g2_decap_8 FILLER_79_2613 ();
 sg13g2_decap_8 FILLER_79_2620 ();
 sg13g2_decap_8 FILLER_79_2627 ();
 sg13g2_decap_8 FILLER_79_2634 ();
 sg13g2_decap_8 FILLER_79_2641 ();
 sg13g2_decap_8 FILLER_79_2648 ();
 sg13g2_decap_8 FILLER_79_2655 ();
 sg13g2_decap_8 FILLER_79_2662 ();
 sg13g2_fill_1 FILLER_79_2669 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_fill_1 FILLER_80_70 ();
 sg13g2_decap_4 FILLER_80_87 ();
 sg13g2_fill_1 FILLER_80_111 ();
 sg13g2_fill_2 FILLER_80_124 ();
 sg13g2_decap_4 FILLER_80_134 ();
 sg13g2_fill_1 FILLER_80_146 ();
 sg13g2_fill_1 FILLER_80_151 ();
 sg13g2_decap_8 FILLER_80_156 ();
 sg13g2_fill_1 FILLER_80_163 ();
 sg13g2_decap_8 FILLER_80_168 ();
 sg13g2_fill_1 FILLER_80_175 ();
 sg13g2_decap_8 FILLER_80_192 ();
 sg13g2_decap_8 FILLER_80_199 ();
 sg13g2_decap_8 FILLER_80_206 ();
 sg13g2_decap_8 FILLER_80_217 ();
 sg13g2_decap_4 FILLER_80_224 ();
 sg13g2_fill_2 FILLER_80_228 ();
 sg13g2_decap_8 FILLER_80_238 ();
 sg13g2_fill_2 FILLER_80_245 ();
 sg13g2_fill_1 FILLER_80_247 ();
 sg13g2_decap_8 FILLER_80_252 ();
 sg13g2_decap_8 FILLER_80_267 ();
 sg13g2_decap_8 FILLER_80_278 ();
 sg13g2_decap_8 FILLER_80_285 ();
 sg13g2_fill_1 FILLER_80_292 ();
 sg13g2_decap_8 FILLER_80_297 ();
 sg13g2_decap_8 FILLER_80_304 ();
 sg13g2_decap_8 FILLER_80_311 ();
 sg13g2_decap_8 FILLER_80_318 ();
 sg13g2_decap_8 FILLER_80_325 ();
 sg13g2_decap_4 FILLER_80_332 ();
 sg13g2_decap_8 FILLER_80_340 ();
 sg13g2_decap_8 FILLER_80_347 ();
 sg13g2_decap_8 FILLER_80_354 ();
 sg13g2_decap_8 FILLER_80_361 ();
 sg13g2_decap_8 FILLER_80_368 ();
 sg13g2_decap_8 FILLER_80_375 ();
 sg13g2_decap_8 FILLER_80_382 ();
 sg13g2_decap_8 FILLER_80_389 ();
 sg13g2_decap_8 FILLER_80_401 ();
 sg13g2_decap_8 FILLER_80_408 ();
 sg13g2_decap_8 FILLER_80_415 ();
 sg13g2_decap_8 FILLER_80_422 ();
 sg13g2_decap_8 FILLER_80_429 ();
 sg13g2_decap_8 FILLER_80_436 ();
 sg13g2_decap_8 FILLER_80_443 ();
 sg13g2_decap_8 FILLER_80_450 ();
 sg13g2_decap_8 FILLER_80_457 ();
 sg13g2_decap_8 FILLER_80_464 ();
 sg13g2_decap_8 FILLER_80_471 ();
 sg13g2_decap_8 FILLER_80_478 ();
 sg13g2_decap_8 FILLER_80_485 ();
 sg13g2_decap_8 FILLER_80_492 ();
 sg13g2_decap_8 FILLER_80_499 ();
 sg13g2_decap_8 FILLER_80_506 ();
 sg13g2_decap_8 FILLER_80_513 ();
 sg13g2_decap_8 FILLER_80_520 ();
 sg13g2_decap_8 FILLER_80_527 ();
 sg13g2_decap_8 FILLER_80_534 ();
 sg13g2_decap_8 FILLER_80_541 ();
 sg13g2_decap_8 FILLER_80_548 ();
 sg13g2_decap_8 FILLER_80_555 ();
 sg13g2_decap_8 FILLER_80_562 ();
 sg13g2_decap_8 FILLER_80_569 ();
 sg13g2_decap_8 FILLER_80_576 ();
 sg13g2_decap_8 FILLER_80_583 ();
 sg13g2_decap_8 FILLER_80_590 ();
 sg13g2_decap_8 FILLER_80_597 ();
 sg13g2_decap_8 FILLER_80_604 ();
 sg13g2_decap_8 FILLER_80_611 ();
 sg13g2_decap_8 FILLER_80_618 ();
 sg13g2_decap_8 FILLER_80_625 ();
 sg13g2_decap_8 FILLER_80_632 ();
 sg13g2_decap_8 FILLER_80_639 ();
 sg13g2_decap_8 FILLER_80_646 ();
 sg13g2_decap_8 FILLER_80_653 ();
 sg13g2_decap_8 FILLER_80_660 ();
 sg13g2_decap_8 FILLER_80_667 ();
 sg13g2_decap_8 FILLER_80_674 ();
 sg13g2_decap_8 FILLER_80_681 ();
 sg13g2_decap_8 FILLER_80_688 ();
 sg13g2_decap_8 FILLER_80_695 ();
 sg13g2_decap_8 FILLER_80_702 ();
 sg13g2_decap_8 FILLER_80_709 ();
 sg13g2_decap_8 FILLER_80_716 ();
 sg13g2_decap_8 FILLER_80_723 ();
 sg13g2_decap_8 FILLER_80_730 ();
 sg13g2_decap_8 FILLER_80_737 ();
 sg13g2_decap_8 FILLER_80_744 ();
 sg13g2_decap_8 FILLER_80_751 ();
 sg13g2_decap_8 FILLER_80_758 ();
 sg13g2_decap_8 FILLER_80_765 ();
 sg13g2_decap_8 FILLER_80_772 ();
 sg13g2_decap_8 FILLER_80_779 ();
 sg13g2_decap_8 FILLER_80_786 ();
 sg13g2_decap_8 FILLER_80_793 ();
 sg13g2_decap_8 FILLER_80_800 ();
 sg13g2_decap_8 FILLER_80_807 ();
 sg13g2_decap_8 FILLER_80_814 ();
 sg13g2_decap_8 FILLER_80_821 ();
 sg13g2_decap_8 FILLER_80_828 ();
 sg13g2_decap_8 FILLER_80_835 ();
 sg13g2_decap_8 FILLER_80_842 ();
 sg13g2_decap_8 FILLER_80_849 ();
 sg13g2_decap_8 FILLER_80_856 ();
 sg13g2_decap_8 FILLER_80_863 ();
 sg13g2_decap_8 FILLER_80_870 ();
 sg13g2_decap_8 FILLER_80_877 ();
 sg13g2_decap_8 FILLER_80_884 ();
 sg13g2_decap_8 FILLER_80_891 ();
 sg13g2_decap_8 FILLER_80_898 ();
 sg13g2_decap_8 FILLER_80_905 ();
 sg13g2_decap_8 FILLER_80_912 ();
 sg13g2_decap_8 FILLER_80_919 ();
 sg13g2_decap_8 FILLER_80_926 ();
 sg13g2_decap_8 FILLER_80_933 ();
 sg13g2_decap_8 FILLER_80_940 ();
 sg13g2_decap_8 FILLER_80_947 ();
 sg13g2_decap_8 FILLER_80_954 ();
 sg13g2_decap_8 FILLER_80_961 ();
 sg13g2_decap_8 FILLER_80_968 ();
 sg13g2_decap_8 FILLER_80_975 ();
 sg13g2_decap_8 FILLER_80_982 ();
 sg13g2_decap_8 FILLER_80_989 ();
 sg13g2_decap_8 FILLER_80_996 ();
 sg13g2_decap_8 FILLER_80_1003 ();
 sg13g2_decap_8 FILLER_80_1010 ();
 sg13g2_decap_8 FILLER_80_1017 ();
 sg13g2_decap_8 FILLER_80_1024 ();
 sg13g2_decap_8 FILLER_80_1031 ();
 sg13g2_decap_8 FILLER_80_1038 ();
 sg13g2_decap_8 FILLER_80_1045 ();
 sg13g2_decap_8 FILLER_80_1052 ();
 sg13g2_decap_8 FILLER_80_1059 ();
 sg13g2_decap_8 FILLER_80_1066 ();
 sg13g2_decap_8 FILLER_80_1073 ();
 sg13g2_decap_8 FILLER_80_1080 ();
 sg13g2_decap_8 FILLER_80_1087 ();
 sg13g2_decap_8 FILLER_80_1094 ();
 sg13g2_decap_8 FILLER_80_1101 ();
 sg13g2_decap_8 FILLER_80_1108 ();
 sg13g2_decap_8 FILLER_80_1115 ();
 sg13g2_decap_8 FILLER_80_1122 ();
 sg13g2_decap_8 FILLER_80_1129 ();
 sg13g2_decap_8 FILLER_80_1136 ();
 sg13g2_decap_8 FILLER_80_1143 ();
 sg13g2_decap_8 FILLER_80_1150 ();
 sg13g2_decap_8 FILLER_80_1157 ();
 sg13g2_decap_8 FILLER_80_1164 ();
 sg13g2_decap_8 FILLER_80_1171 ();
 sg13g2_decap_8 FILLER_80_1178 ();
 sg13g2_decap_8 FILLER_80_1185 ();
 sg13g2_decap_8 FILLER_80_1192 ();
 sg13g2_decap_8 FILLER_80_1199 ();
 sg13g2_decap_8 FILLER_80_1206 ();
 sg13g2_decap_8 FILLER_80_1213 ();
 sg13g2_decap_8 FILLER_80_1220 ();
 sg13g2_decap_8 FILLER_80_1227 ();
 sg13g2_decap_8 FILLER_80_1234 ();
 sg13g2_decap_8 FILLER_80_1241 ();
 sg13g2_decap_8 FILLER_80_1248 ();
 sg13g2_decap_8 FILLER_80_1255 ();
 sg13g2_decap_8 FILLER_80_1262 ();
 sg13g2_decap_8 FILLER_80_1269 ();
 sg13g2_decap_8 FILLER_80_1276 ();
 sg13g2_decap_8 FILLER_80_1283 ();
 sg13g2_decap_8 FILLER_80_1290 ();
 sg13g2_decap_8 FILLER_80_1297 ();
 sg13g2_decap_8 FILLER_80_1304 ();
 sg13g2_decap_8 FILLER_80_1311 ();
 sg13g2_decap_8 FILLER_80_1318 ();
 sg13g2_decap_8 FILLER_80_1325 ();
 sg13g2_decap_8 FILLER_80_1332 ();
 sg13g2_decap_8 FILLER_80_1339 ();
 sg13g2_decap_8 FILLER_80_1346 ();
 sg13g2_decap_8 FILLER_80_1353 ();
 sg13g2_decap_8 FILLER_80_1360 ();
 sg13g2_decap_8 FILLER_80_1367 ();
 sg13g2_decap_8 FILLER_80_1374 ();
 sg13g2_decap_8 FILLER_80_1381 ();
 sg13g2_decap_8 FILLER_80_1388 ();
 sg13g2_decap_8 FILLER_80_1395 ();
 sg13g2_decap_8 FILLER_80_1402 ();
 sg13g2_decap_8 FILLER_80_1409 ();
 sg13g2_decap_8 FILLER_80_1416 ();
 sg13g2_decap_8 FILLER_80_1423 ();
 sg13g2_decap_8 FILLER_80_1430 ();
 sg13g2_decap_8 FILLER_80_1437 ();
 sg13g2_decap_8 FILLER_80_1444 ();
 sg13g2_decap_8 FILLER_80_1451 ();
 sg13g2_decap_8 FILLER_80_1458 ();
 sg13g2_decap_8 FILLER_80_1465 ();
 sg13g2_decap_8 FILLER_80_1472 ();
 sg13g2_decap_8 FILLER_80_1479 ();
 sg13g2_decap_8 FILLER_80_1486 ();
 sg13g2_decap_8 FILLER_80_1493 ();
 sg13g2_decap_8 FILLER_80_1500 ();
 sg13g2_decap_8 FILLER_80_1507 ();
 sg13g2_decap_8 FILLER_80_1514 ();
 sg13g2_decap_8 FILLER_80_1521 ();
 sg13g2_decap_8 FILLER_80_1528 ();
 sg13g2_decap_8 FILLER_80_1535 ();
 sg13g2_decap_8 FILLER_80_1542 ();
 sg13g2_decap_8 FILLER_80_1549 ();
 sg13g2_decap_8 FILLER_80_1556 ();
 sg13g2_decap_8 FILLER_80_1563 ();
 sg13g2_decap_8 FILLER_80_1570 ();
 sg13g2_decap_8 FILLER_80_1577 ();
 sg13g2_decap_8 FILLER_80_1584 ();
 sg13g2_decap_8 FILLER_80_1591 ();
 sg13g2_decap_8 FILLER_80_1598 ();
 sg13g2_decap_8 FILLER_80_1605 ();
 sg13g2_decap_8 FILLER_80_1612 ();
 sg13g2_decap_8 FILLER_80_1619 ();
 sg13g2_decap_8 FILLER_80_1626 ();
 sg13g2_decap_8 FILLER_80_1633 ();
 sg13g2_decap_8 FILLER_80_1640 ();
 sg13g2_decap_8 FILLER_80_1647 ();
 sg13g2_decap_8 FILLER_80_1654 ();
 sg13g2_decap_8 FILLER_80_1661 ();
 sg13g2_decap_8 FILLER_80_1668 ();
 sg13g2_decap_8 FILLER_80_1675 ();
 sg13g2_decap_8 FILLER_80_1682 ();
 sg13g2_decap_8 FILLER_80_1689 ();
 sg13g2_decap_8 FILLER_80_1696 ();
 sg13g2_decap_8 FILLER_80_1703 ();
 sg13g2_decap_8 FILLER_80_1710 ();
 sg13g2_decap_8 FILLER_80_1717 ();
 sg13g2_decap_8 FILLER_80_1724 ();
 sg13g2_decap_8 FILLER_80_1731 ();
 sg13g2_decap_8 FILLER_80_1738 ();
 sg13g2_decap_8 FILLER_80_1745 ();
 sg13g2_decap_8 FILLER_80_1752 ();
 sg13g2_decap_8 FILLER_80_1759 ();
 sg13g2_decap_8 FILLER_80_1766 ();
 sg13g2_decap_8 FILLER_80_1773 ();
 sg13g2_decap_8 FILLER_80_1780 ();
 sg13g2_decap_8 FILLER_80_1787 ();
 sg13g2_decap_8 FILLER_80_1794 ();
 sg13g2_decap_8 FILLER_80_1801 ();
 sg13g2_decap_8 FILLER_80_1808 ();
 sg13g2_decap_8 FILLER_80_1815 ();
 sg13g2_decap_8 FILLER_80_1822 ();
 sg13g2_decap_8 FILLER_80_1829 ();
 sg13g2_decap_8 FILLER_80_1836 ();
 sg13g2_decap_8 FILLER_80_1843 ();
 sg13g2_decap_8 FILLER_80_1850 ();
 sg13g2_decap_8 FILLER_80_1857 ();
 sg13g2_decap_8 FILLER_80_1864 ();
 sg13g2_decap_8 FILLER_80_1871 ();
 sg13g2_decap_8 FILLER_80_1878 ();
 sg13g2_decap_8 FILLER_80_1885 ();
 sg13g2_decap_8 FILLER_80_1892 ();
 sg13g2_decap_8 FILLER_80_1899 ();
 sg13g2_decap_8 FILLER_80_1906 ();
 sg13g2_decap_8 FILLER_80_1913 ();
 sg13g2_decap_8 FILLER_80_1920 ();
 sg13g2_decap_8 FILLER_80_1927 ();
 sg13g2_decap_8 FILLER_80_1934 ();
 sg13g2_decap_8 FILLER_80_1941 ();
 sg13g2_decap_8 FILLER_80_1948 ();
 sg13g2_decap_8 FILLER_80_1955 ();
 sg13g2_decap_8 FILLER_80_1962 ();
 sg13g2_decap_8 FILLER_80_1969 ();
 sg13g2_decap_8 FILLER_80_1976 ();
 sg13g2_decap_8 FILLER_80_1983 ();
 sg13g2_decap_8 FILLER_80_1990 ();
 sg13g2_decap_8 FILLER_80_1997 ();
 sg13g2_decap_8 FILLER_80_2004 ();
 sg13g2_decap_8 FILLER_80_2011 ();
 sg13g2_decap_8 FILLER_80_2018 ();
 sg13g2_decap_8 FILLER_80_2025 ();
 sg13g2_decap_8 FILLER_80_2032 ();
 sg13g2_decap_8 FILLER_80_2039 ();
 sg13g2_decap_8 FILLER_80_2046 ();
 sg13g2_decap_8 FILLER_80_2053 ();
 sg13g2_decap_8 FILLER_80_2060 ();
 sg13g2_decap_8 FILLER_80_2067 ();
 sg13g2_decap_8 FILLER_80_2074 ();
 sg13g2_decap_8 FILLER_80_2081 ();
 sg13g2_decap_8 FILLER_80_2088 ();
 sg13g2_decap_8 FILLER_80_2095 ();
 sg13g2_decap_8 FILLER_80_2102 ();
 sg13g2_decap_8 FILLER_80_2109 ();
 sg13g2_decap_8 FILLER_80_2116 ();
 sg13g2_decap_8 FILLER_80_2123 ();
 sg13g2_decap_8 FILLER_80_2130 ();
 sg13g2_decap_8 FILLER_80_2137 ();
 sg13g2_decap_8 FILLER_80_2144 ();
 sg13g2_decap_8 FILLER_80_2151 ();
 sg13g2_decap_8 FILLER_80_2158 ();
 sg13g2_decap_8 FILLER_80_2165 ();
 sg13g2_decap_8 FILLER_80_2172 ();
 sg13g2_decap_8 FILLER_80_2179 ();
 sg13g2_decap_8 FILLER_80_2186 ();
 sg13g2_decap_8 FILLER_80_2193 ();
 sg13g2_decap_8 FILLER_80_2200 ();
 sg13g2_decap_8 FILLER_80_2207 ();
 sg13g2_decap_8 FILLER_80_2214 ();
 sg13g2_decap_8 FILLER_80_2221 ();
 sg13g2_decap_8 FILLER_80_2228 ();
 sg13g2_decap_8 FILLER_80_2235 ();
 sg13g2_decap_8 FILLER_80_2242 ();
 sg13g2_decap_8 FILLER_80_2249 ();
 sg13g2_decap_8 FILLER_80_2256 ();
 sg13g2_decap_8 FILLER_80_2263 ();
 sg13g2_decap_8 FILLER_80_2270 ();
 sg13g2_decap_8 FILLER_80_2277 ();
 sg13g2_decap_8 FILLER_80_2284 ();
 sg13g2_decap_8 FILLER_80_2291 ();
 sg13g2_decap_8 FILLER_80_2298 ();
 sg13g2_decap_8 FILLER_80_2305 ();
 sg13g2_decap_8 FILLER_80_2312 ();
 sg13g2_decap_8 FILLER_80_2319 ();
 sg13g2_decap_8 FILLER_80_2326 ();
 sg13g2_decap_8 FILLER_80_2333 ();
 sg13g2_decap_8 FILLER_80_2340 ();
 sg13g2_decap_8 FILLER_80_2347 ();
 sg13g2_decap_8 FILLER_80_2354 ();
 sg13g2_decap_8 FILLER_80_2361 ();
 sg13g2_decap_8 FILLER_80_2368 ();
 sg13g2_decap_8 FILLER_80_2375 ();
 sg13g2_decap_8 FILLER_80_2382 ();
 sg13g2_decap_8 FILLER_80_2389 ();
 sg13g2_decap_8 FILLER_80_2396 ();
 sg13g2_decap_8 FILLER_80_2403 ();
 sg13g2_decap_8 FILLER_80_2410 ();
 sg13g2_decap_8 FILLER_80_2417 ();
 sg13g2_decap_8 FILLER_80_2424 ();
 sg13g2_decap_8 FILLER_80_2431 ();
 sg13g2_decap_8 FILLER_80_2438 ();
 sg13g2_decap_8 FILLER_80_2445 ();
 sg13g2_decap_8 FILLER_80_2452 ();
 sg13g2_decap_8 FILLER_80_2459 ();
 sg13g2_decap_8 FILLER_80_2466 ();
 sg13g2_decap_8 FILLER_80_2473 ();
 sg13g2_decap_8 FILLER_80_2480 ();
 sg13g2_decap_8 FILLER_80_2487 ();
 sg13g2_decap_8 FILLER_80_2494 ();
 sg13g2_decap_8 FILLER_80_2501 ();
 sg13g2_decap_8 FILLER_80_2508 ();
 sg13g2_decap_8 FILLER_80_2515 ();
 sg13g2_decap_8 FILLER_80_2522 ();
 sg13g2_decap_8 FILLER_80_2529 ();
 sg13g2_decap_8 FILLER_80_2536 ();
 sg13g2_decap_8 FILLER_80_2543 ();
 sg13g2_decap_8 FILLER_80_2550 ();
 sg13g2_decap_8 FILLER_80_2557 ();
 sg13g2_decap_8 FILLER_80_2564 ();
 sg13g2_decap_8 FILLER_80_2571 ();
 sg13g2_decap_8 FILLER_80_2578 ();
 sg13g2_decap_8 FILLER_80_2585 ();
 sg13g2_decap_8 FILLER_80_2592 ();
 sg13g2_decap_8 FILLER_80_2599 ();
 sg13g2_decap_8 FILLER_80_2606 ();
 sg13g2_decap_8 FILLER_80_2613 ();
 sg13g2_decap_8 FILLER_80_2620 ();
 sg13g2_decap_8 FILLER_80_2627 ();
 sg13g2_decap_8 FILLER_80_2634 ();
 sg13g2_decap_8 FILLER_80_2641 ();
 sg13g2_decap_8 FILLER_80_2648 ();
 sg13g2_decap_8 FILLER_80_2655 ();
 sg13g2_decap_8 FILLER_80_2662 ();
 sg13g2_fill_1 FILLER_80_2669 ();
endmodule
